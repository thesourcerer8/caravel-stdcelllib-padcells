magic
tech sky130A
magscale 1 2
timestamp 1608118436
<< locali >>
rect 219081 685899 219115 695453
rect 154313 676243 154347 685797
rect 218989 666587 219023 676141
rect 299857 666587 299891 684437
rect 219265 647275 219299 656829
rect 219357 616879 219391 626501
rect 219081 608719 219115 611405
rect 219265 601579 219299 608549
rect 299673 601715 299707 608549
rect 219173 589339 219207 598893
rect 299857 589339 299891 598893
rect 154313 579751 154347 589237
rect 218897 569959 218931 579581
rect 218897 550647 218931 553401
rect 154405 521679 154439 531233
rect 154405 502367 154439 511921
rect 219081 505087 219115 510561
rect 299673 485775 299707 492609
rect 299673 466395 299707 473297
rect 154221 444431 154255 453985
rect 218989 444431 219023 453985
rect 299489 440283 299523 449837
rect 299581 427771 299615 436781
rect 299673 405739 299707 415361
rect 154589 402951 154623 403053
rect 164157 402951 164191 403053
rect 251189 402951 251223 403121
rect 260757 403019 260791 403121
rect 105955 402781 106013 402815
rect 105771 402713 106105 402747
rect 244841 401591 244875 401965
rect 248337 401591 248371 401829
rect 253949 401591 253983 402101
rect 254133 402067 254167 402713
rect 254777 402611 254811 402781
rect 255973 402679 256007 402917
rect 254225 402135 254259 402577
rect 254041 401931 254075 402033
rect 257905 401931 257939 402713
rect 261309 402679 261343 402917
rect 257997 401931 258031 402169
rect 259503 402033 259653 402067
rect 272349 401931 272383 402033
rect 244197 399279 244231 400129
rect 253949 399279 253983 400129
rect 263517 399279 263551 400129
rect 279801 399449 280077 399483
rect 279801 399279 279835 399449
rect 279927 399381 279985 399415
rect 280169 399279 280203 399449
rect 282837 399415 282871 399517
rect 289829 399415 289863 399517
rect 299397 399211 299431 399517
rect 338129 399483 338163 399585
rect 347697 399415 347731 399585
rect 357449 399483 357483 399585
rect 367017 399415 367051 399585
rect 376769 399483 376803 399585
rect 386337 399415 386371 399585
rect 331171 399381 331229 399415
rect 350491 399381 350549 399415
rect 369811 399381 369869 399415
rect 309149 399075 309183 399177
rect 318717 399075 318751 399245
rect 386981 398191 387015 399381
rect 235641 337739 235675 337977
rect 235733 337807 235767 338045
rect 235917 337875 235951 338045
rect 232053 337059 232087 337297
rect 57989 336039 58023 336141
rect 62773 335971 62807 336141
rect 104909 336107 104943 336345
rect 114477 336243 114511 336345
rect 115891 336209 115983 336243
rect 115949 336175 115983 336209
rect 132509 336107 132543 336209
rect 142077 336107 142111 336209
rect 143549 336107 143583 336209
rect 211203 336141 211445 336175
rect 96537 336039 96571 336073
rect 96479 336005 96571 336039
rect 176611 336005 176795 336039
rect 67649 335835 67683 335937
rect 77217 335835 77251 335937
rect 77309 335835 77343 335937
rect 81633 335835 81667 335937
rect 86969 335835 87003 335937
rect 96537 335835 96571 335937
rect 96629 335835 96663 335937
rect 106289 335937 106473 335971
rect 106289 335903 106323 335937
rect 115949 335835 115983 335937
rect 129105 335903 129139 336005
rect 176761 335971 176795 336005
rect 129047 335869 129139 335903
rect 132509 335835 132543 335937
rect 143583 335937 143675 335971
rect 142077 335835 142111 335937
rect 143641 335903 143675 335937
rect 179429 335835 179463 335937
rect 188997 335835 189031 335937
rect 189089 335835 189123 335937
rect 196081 335835 196115 335937
rect 198749 335835 198783 335937
rect 209731 335937 209789 335971
rect 208317 335835 208351 335937
rect 229569 328491 229603 334169
rect 230581 329511 230615 337025
rect 231869 336107 231903 336549
rect 234997 336243 235031 337365
rect 236009 337263 236043 337841
rect 240701 328491 240735 338045
rect 241529 337399 241563 337637
rect 241805 337331 241839 337705
rect 243093 330667 243127 338045
rect 260849 337467 260883 337909
rect 263517 337671 263551 337909
rect 245577 335019 245611 335733
rect 246221 334815 246255 335801
rect 248705 328491 248739 336073
rect 251557 330871 251591 335665
rect 251741 335359 251775 336957
rect 260665 336787 260699 337161
rect 261217 336651 261251 337229
rect 262965 336787 262999 337569
rect 263149 336991 263183 337365
rect 263241 336855 263275 337637
rect 263793 337127 263827 337569
rect 263643 337093 263827 337127
rect 263701 336787 263735 336889
rect 266093 336787 266127 337229
rect 256433 331755 256467 335257
rect 267473 328491 267507 338045
rect 231501 318835 231535 328389
rect 229477 309247 229511 318733
rect 233525 317475 233559 327029
rect 237573 317475 237607 327029
rect 267933 325703 267967 337773
rect 270509 336719 270543 337501
rect 270693 336787 270727 337501
rect 275293 337467 275327 337637
rect 277409 337603 277443 337705
rect 277961 337671 277995 337841
rect 280169 337739 280203 337909
rect 277685 337399 277719 337501
rect 277869 337467 277903 337637
rect 277627 337365 277719 337399
rect 271061 331211 271095 337161
rect 274649 337127 274683 337297
rect 277685 337263 277719 337297
rect 277685 337229 278145 337263
rect 274833 331143 274867 337093
rect 276305 336787 276339 337161
rect 276397 329307 276431 336889
rect 277501 336855 277535 337229
rect 278973 335155 279007 337229
rect 280169 335223 280203 337297
rect 280445 335291 280479 337841
rect 280813 336787 280847 337637
rect 281457 336923 281491 337229
rect 282469 335155 282503 337161
rect 282837 337059 282871 337773
rect 282929 337331 282963 337705
rect 282745 336787 282779 337025
rect 283113 336991 283147 337297
rect 283055 336957 283147 336991
rect 283021 336719 283055 336821
rect 283389 332095 283423 332401
rect 283665 328559 283699 337909
rect 287345 337841 288023 337875
rect 287345 337807 287379 337841
rect 284033 336923 284067 337501
rect 287437 337399 287471 337773
rect 287621 337773 287931 337807
rect 287621 337739 287655 337773
rect 287529 337399 287563 337569
rect 287713 337127 287747 337705
rect 287805 337059 287839 337501
rect 287897 337127 287931 337773
rect 287989 337059 288023 337841
rect 290933 337671 290967 337909
rect 291025 337263 291059 337909
rect 284401 328899 284435 335733
rect 279893 326519 279927 326757
rect 238953 317475 238987 319481
rect 284585 318835 284619 328389
rect 287621 327131 287655 335665
rect 289829 331823 289863 331925
rect 249165 309179 249199 318733
rect 229477 299523 229511 309077
rect 233525 305643 233559 309077
rect 238953 299523 238987 309077
rect 251741 298163 251775 307717
rect 260205 299387 260239 307717
rect 283021 302923 283055 309009
rect 283757 299591 283791 317373
rect 284677 302175 284711 309077
rect 288173 307819 288207 317373
rect 237573 288439 237607 298061
rect 243461 280211 243495 289765
rect 251649 287079 251683 292485
rect 229569 270555 229603 280109
rect 241161 260899 241195 270453
rect 229569 251243 229603 260797
rect 243461 256751 243495 278681
rect 259929 267767 259963 278681
rect 277869 277423 277903 289561
rect 283757 288439 283791 298061
rect 288173 288439 288207 298061
rect 253949 258111 253983 260865
rect 237573 244171 237607 248353
rect 243461 240227 243495 255221
rect 260113 249747 260147 258009
rect 260205 248455 260239 258009
rect 275293 248455 275327 249781
rect 258549 240159 258583 244409
rect 237481 227783 237515 231965
rect 243461 219487 243495 237337
rect 254041 230299 254075 238697
rect 260297 230503 260331 240057
rect 251833 222207 251867 224961
rect 277961 220847 277995 225165
rect 237665 214591 237699 219317
rect 238953 205343 238987 218841
rect 243461 202895 243495 219317
rect 270969 211191 271003 220745
rect 277869 209831 277903 219385
rect 275293 205615 275327 209729
rect 260205 191879 260239 201433
rect 243369 186303 243403 191777
rect 243461 174403 243495 182053
rect 237573 166991 237607 172465
rect 238217 162911 238251 172465
rect 256525 169779 256559 173961
rect 258641 171207 258675 180761
rect 260297 178755 260331 183481
rect 270969 182223 271003 191777
rect 275293 190519 275327 190621
rect 270785 171139 270819 180761
rect 275201 171139 275235 180761
rect 241161 153255 241195 162809
rect 258641 161483 258675 171037
rect 259377 161551 259411 171037
rect 243461 153323 243495 157369
rect 237573 147611 237607 153153
rect 238217 143599 238251 153153
rect 238953 147203 238987 153153
rect 237573 134011 237607 143429
rect 238125 122859 238159 133841
rect 243461 124219 243495 142069
rect 251649 132515 251683 137105
rect 254041 132515 254075 142069
rect 256433 139451 256467 149005
rect 258641 142171 258675 151725
rect 259285 142171 259319 160021
rect 260205 153323 260239 162809
rect 275201 161483 275235 170969
rect 276489 135303 276523 144857
rect 238033 113135 238067 121397
rect 238769 115379 238803 121397
rect 241069 114563 241103 124117
rect 243553 108987 243587 118881
rect 253949 111843 253983 122757
rect 256525 113203 256559 122757
rect 258549 121499 258583 131053
rect 260297 124287 260331 133841
rect 275385 124219 275419 133841
rect 278145 128299 278179 135201
rect 260113 114563 260147 124117
rect 260297 114563 260331 124117
rect 272441 111843 272475 121397
rect 237573 85595 237607 95149
rect 238125 92531 238159 102085
rect 248981 97835 249015 106165
rect 251741 100759 251775 110381
rect 258641 102187 258675 111741
rect 272349 102187 272383 111673
rect 276489 107627 276523 119357
rect 278329 104907 278363 114461
rect 253857 91103 253891 95217
rect 229569 77367 229603 80121
rect 229569 67643 229603 77197
rect 237573 73219 237607 82773
rect 243553 77299 243587 86921
rect 248797 82127 248831 86921
rect 248981 78455 249015 86853
rect 249165 77299 249199 86921
rect 258549 84235 258583 97257
rect 260113 92531 260147 102085
rect 251741 74579 251775 84133
rect 253949 75871 253983 80121
rect 259285 74579 259319 84133
rect 260297 75939 260331 86513
rect 272349 74579 272383 97257
rect 275293 84235 275327 93789
rect 238953 64923 238987 74477
rect 229569 48331 229603 57885
rect 238217 55267 238251 64821
rect 240517 57987 240551 67541
rect 258549 64991 258583 74477
rect 241161 55267 241195 64821
rect 238217 46971 238251 51085
rect 238953 45611 238987 55165
rect 229569 29019 229603 38573
rect 237573 35955 237607 45509
rect 238309 36023 238343 45509
rect 241253 35955 241287 45509
rect 238125 26299 238159 35853
rect 243461 27659 243495 48229
rect 258641 45611 258675 63461
rect 275293 51051 275327 56525
rect 260113 46971 260147 48365
rect 260297 46971 260331 48365
rect 278053 37315 278087 46869
rect 243461 22083 243495 27489
rect 256617 26299 256651 35853
rect 259285 26299 259319 35853
rect 238861 16643 238895 21437
rect 253949 16643 253983 18037
rect 259929 18003 259963 19465
rect 237573 9299 237607 16541
rect 260205 8347 260239 17833
rect 274925 16643 274959 26197
rect 276489 9707 276523 19261
rect 278237 9707 278271 27489
rect 244289 5219 244323 5457
rect 224141 4607 224175 4981
rect 224233 4811 224267 4981
rect 74549 3111 74583 3961
rect 84025 3111 84059 3961
rect 93869 2975 93903 3961
rect 93961 2907 93995 4029
rect 103345 2907 103379 4029
rect 103437 2975 103471 3961
rect 231133 3383 231167 3553
rect 232329 3451 232363 4029
rect 232421 3723 232455 4029
rect 233065 2975 233099 3689
rect 248981 3519 249015 3893
rect 275385 3723 275419 8245
rect 433349 3859 433383 3961
rect 571073 3247 571107 3553
rect 571993 3383 572027 3485
<< viali >>
rect 219081 695453 219115 695487
rect 219081 685865 219115 685899
rect 154313 685797 154347 685831
rect 154313 676209 154347 676243
rect 299857 684437 299891 684471
rect 218989 676141 219023 676175
rect 218989 666553 219023 666587
rect 299857 666553 299891 666587
rect 219265 656829 219299 656863
rect 219265 647241 219299 647275
rect 219357 626501 219391 626535
rect 219357 616845 219391 616879
rect 219081 611405 219115 611439
rect 219081 608685 219115 608719
rect 219265 608549 219299 608583
rect 299673 608549 299707 608583
rect 299673 601681 299707 601715
rect 219265 601545 219299 601579
rect 219173 598893 219207 598927
rect 219173 589305 219207 589339
rect 299857 598893 299891 598927
rect 299857 589305 299891 589339
rect 154313 589237 154347 589271
rect 154313 579717 154347 579751
rect 218897 579581 218931 579615
rect 218897 569925 218931 569959
rect 218897 553401 218931 553435
rect 218897 550613 218931 550647
rect 154405 531233 154439 531267
rect 154405 521645 154439 521679
rect 154405 511921 154439 511955
rect 219081 510561 219115 510595
rect 219081 505053 219115 505087
rect 154405 502333 154439 502367
rect 299673 492609 299707 492643
rect 299673 485741 299707 485775
rect 299673 473297 299707 473331
rect 299673 466361 299707 466395
rect 154221 453985 154255 454019
rect 154221 444397 154255 444431
rect 218989 453985 219023 454019
rect 218989 444397 219023 444431
rect 299489 449837 299523 449871
rect 299489 440249 299523 440283
rect 299581 436781 299615 436815
rect 299581 427737 299615 427771
rect 299673 415361 299707 415395
rect 299673 405705 299707 405739
rect 251189 403121 251223 403155
rect 154589 403053 154623 403087
rect 154589 402917 154623 402951
rect 164157 403053 164191 403087
rect 164157 402917 164191 402951
rect 260757 403121 260791 403155
rect 260757 402985 260791 403019
rect 251189 402917 251223 402951
rect 255973 402917 256007 402951
rect 105921 402781 105955 402815
rect 106013 402781 106047 402815
rect 254777 402781 254811 402815
rect 105737 402713 105771 402747
rect 106105 402713 106139 402747
rect 254133 402713 254167 402747
rect 253949 402101 253983 402135
rect 244841 401965 244875 401999
rect 244841 401557 244875 401591
rect 248337 401829 248371 401863
rect 248337 401557 248371 401591
rect 261309 402917 261343 402951
rect 255973 402645 256007 402679
rect 257905 402713 257939 402747
rect 254225 402577 254259 402611
rect 254777 402577 254811 402611
rect 254225 402101 254259 402135
rect 254041 402033 254075 402067
rect 254133 402033 254167 402067
rect 254041 401897 254075 401931
rect 261309 402645 261343 402679
rect 257905 401897 257939 401931
rect 257997 402169 258031 402203
rect 259469 402033 259503 402067
rect 259653 402033 259687 402067
rect 272349 402033 272383 402067
rect 257997 401897 258031 401931
rect 272349 401897 272383 401931
rect 253949 401557 253983 401591
rect 244197 400129 244231 400163
rect 244197 399245 244231 399279
rect 253949 400129 253983 400163
rect 253949 399245 253983 399279
rect 263517 400129 263551 400163
rect 338129 399585 338163 399619
rect 282837 399517 282871 399551
rect 263517 399245 263551 399279
rect 280077 399449 280111 399483
rect 280169 399449 280203 399483
rect 279893 399381 279927 399415
rect 279985 399381 280019 399415
rect 279801 399245 279835 399279
rect 282837 399381 282871 399415
rect 289829 399517 289863 399551
rect 289829 399381 289863 399415
rect 299397 399517 299431 399551
rect 280169 399245 280203 399279
rect 338129 399449 338163 399483
rect 347697 399585 347731 399619
rect 357449 399585 357483 399619
rect 357449 399449 357483 399483
rect 367017 399585 367051 399619
rect 376769 399585 376803 399619
rect 376769 399449 376803 399483
rect 386337 399585 386371 399619
rect 331137 399381 331171 399415
rect 331229 399381 331263 399415
rect 347697 399381 347731 399415
rect 350457 399381 350491 399415
rect 350549 399381 350583 399415
rect 367017 399381 367051 399415
rect 369777 399381 369811 399415
rect 369869 399381 369903 399415
rect 386337 399381 386371 399415
rect 386981 399381 387015 399415
rect 318717 399245 318751 399279
rect 299397 399177 299431 399211
rect 309149 399177 309183 399211
rect 309149 399041 309183 399075
rect 318717 399041 318751 399075
rect 386981 398157 387015 398191
rect 235733 338045 235767 338079
rect 235641 337977 235675 338011
rect 235917 338045 235951 338079
rect 240701 338045 240735 338079
rect 235917 337841 235951 337875
rect 236009 337841 236043 337875
rect 235733 337773 235767 337807
rect 235641 337705 235675 337739
rect 234997 337365 235031 337399
rect 232053 337297 232087 337331
rect 230581 337025 230615 337059
rect 232053 337025 232087 337059
rect 104909 336345 104943 336379
rect 57989 336141 58023 336175
rect 57989 336005 58023 336039
rect 62773 336141 62807 336175
rect 114477 336345 114511 336379
rect 114477 336209 114511 336243
rect 115857 336209 115891 336243
rect 115949 336141 115983 336175
rect 132509 336209 132543 336243
rect 96537 336073 96571 336107
rect 104909 336073 104943 336107
rect 132509 336073 132543 336107
rect 142077 336209 142111 336243
rect 142077 336073 142111 336107
rect 143549 336209 143583 336243
rect 211169 336141 211203 336175
rect 211445 336141 211479 336175
rect 143549 336073 143583 336107
rect 96445 336005 96479 336039
rect 129105 336005 129139 336039
rect 176577 336005 176611 336039
rect 62773 335937 62807 335971
rect 67649 335937 67683 335971
rect 67649 335801 67683 335835
rect 77217 335937 77251 335971
rect 77217 335801 77251 335835
rect 77309 335937 77343 335971
rect 77309 335801 77343 335835
rect 81633 335937 81667 335971
rect 81633 335801 81667 335835
rect 86969 335937 87003 335971
rect 86969 335801 87003 335835
rect 96537 335937 96571 335971
rect 96537 335801 96571 335835
rect 96629 335937 96663 335971
rect 106473 335937 106507 335971
rect 115949 335937 115983 335971
rect 106289 335869 106323 335903
rect 96629 335801 96663 335835
rect 129013 335869 129047 335903
rect 132509 335937 132543 335971
rect 115949 335801 115983 335835
rect 132509 335801 132543 335835
rect 142077 335937 142111 335971
rect 143549 335937 143583 335971
rect 176761 335937 176795 335971
rect 179429 335937 179463 335971
rect 143641 335869 143675 335903
rect 142077 335801 142111 335835
rect 179429 335801 179463 335835
rect 188997 335937 189031 335971
rect 188997 335801 189031 335835
rect 189089 335937 189123 335971
rect 189089 335801 189123 335835
rect 196081 335937 196115 335971
rect 196081 335801 196115 335835
rect 198749 335937 198783 335971
rect 198749 335801 198783 335835
rect 208317 335937 208351 335971
rect 209697 335937 209731 335971
rect 209789 335937 209823 335971
rect 208317 335801 208351 335835
rect 229569 334169 229603 334203
rect 231869 336549 231903 336583
rect 236009 337229 236043 337263
rect 234997 336209 235031 336243
rect 231869 336073 231903 336107
rect 230581 329477 230615 329511
rect 229569 328457 229603 328491
rect 243093 338045 243127 338079
rect 241805 337705 241839 337739
rect 241529 337637 241563 337671
rect 241529 337365 241563 337399
rect 241805 337297 241839 337331
rect 267473 338045 267507 338079
rect 260849 337909 260883 337943
rect 263517 337909 263551 337943
rect 263241 337637 263275 337671
rect 263517 337637 263551 337671
rect 260849 337433 260883 337467
rect 262965 337569 262999 337603
rect 261217 337229 261251 337263
rect 260665 337161 260699 337195
rect 251741 336957 251775 336991
rect 248705 336073 248739 336107
rect 246221 335801 246255 335835
rect 245577 335733 245611 335767
rect 245577 334985 245611 335019
rect 246221 334781 246255 334815
rect 243093 330633 243127 330667
rect 240701 328457 240735 328491
rect 251557 335665 251591 335699
rect 260665 336753 260699 336787
rect 263149 337365 263183 337399
rect 263149 336957 263183 336991
rect 263793 337569 263827 337603
rect 263609 337093 263643 337127
rect 266093 337229 266127 337263
rect 263241 336821 263275 336855
rect 263701 336889 263735 336923
rect 262965 336753 262999 336787
rect 263701 336753 263735 336787
rect 266093 336753 266127 336787
rect 261217 336617 261251 336651
rect 251741 335325 251775 335359
rect 256433 335257 256467 335291
rect 256433 331721 256467 331755
rect 251557 330837 251591 330871
rect 248705 328457 248739 328491
rect 280169 337909 280203 337943
rect 277961 337841 277995 337875
rect 267473 328457 267507 328491
rect 267933 337773 267967 337807
rect 231501 328389 231535 328423
rect 231501 318801 231535 318835
rect 233525 327029 233559 327063
rect 229477 318733 229511 318767
rect 233525 317441 233559 317475
rect 237573 327029 237607 327063
rect 277409 337705 277443 337739
rect 275293 337637 275327 337671
rect 270509 337501 270543 337535
rect 270693 337501 270727 337535
rect 283665 337909 283699 337943
rect 280169 337705 280203 337739
rect 280445 337841 280479 337875
rect 277409 337569 277443 337603
rect 277869 337637 277903 337671
rect 277961 337637 277995 337671
rect 275293 337433 275327 337467
rect 277685 337501 277719 337535
rect 277869 337433 277903 337467
rect 277593 337365 277627 337399
rect 274649 337297 274683 337331
rect 270693 336753 270727 336787
rect 271061 337161 271095 337195
rect 270509 336685 270543 336719
rect 277685 337297 277719 337331
rect 280169 337297 280203 337331
rect 277501 337229 277535 337263
rect 278145 337229 278179 337263
rect 278973 337229 279007 337263
rect 276305 337161 276339 337195
rect 274649 337093 274683 337127
rect 274833 337093 274867 337127
rect 271061 331177 271095 331211
rect 276305 336753 276339 336787
rect 276397 336889 276431 336923
rect 274833 331109 274867 331143
rect 277501 336821 277535 336855
rect 282837 337773 282871 337807
rect 280813 337637 280847 337671
rect 281457 337229 281491 337263
rect 281457 336889 281491 336923
rect 282469 337161 282503 337195
rect 280813 336753 280847 336787
rect 280445 335257 280479 335291
rect 280169 335189 280203 335223
rect 278973 335121 279007 335155
rect 282929 337705 282963 337739
rect 282929 337297 282963 337331
rect 283113 337297 283147 337331
rect 282745 337025 282779 337059
rect 282837 337025 282871 337059
rect 283021 336957 283055 336991
rect 282745 336753 282779 336787
rect 283021 336821 283055 336855
rect 283021 336685 283055 336719
rect 282469 335121 282503 335155
rect 283389 332401 283423 332435
rect 283389 332061 283423 332095
rect 276397 329273 276431 329307
rect 290933 337909 290967 337943
rect 287345 337773 287379 337807
rect 287437 337773 287471 337807
rect 284033 337501 284067 337535
rect 287621 337705 287655 337739
rect 287713 337705 287747 337739
rect 287437 337365 287471 337399
rect 287529 337569 287563 337603
rect 287529 337365 287563 337399
rect 287713 337093 287747 337127
rect 287805 337501 287839 337535
rect 287897 337093 287931 337127
rect 287805 337025 287839 337059
rect 290933 337637 290967 337671
rect 291025 337909 291059 337943
rect 291025 337229 291059 337263
rect 287989 337025 288023 337059
rect 284033 336889 284067 336923
rect 284401 335733 284435 335767
rect 284401 328865 284435 328899
rect 287621 335665 287655 335699
rect 283665 328525 283699 328559
rect 284585 328389 284619 328423
rect 279893 326757 279927 326791
rect 279893 326485 279927 326519
rect 267933 325669 267967 325703
rect 237573 317441 237607 317475
rect 238953 319481 238987 319515
rect 289829 331925 289863 331959
rect 289829 331789 289863 331823
rect 287621 327097 287655 327131
rect 284585 318801 284619 318835
rect 238953 317441 238987 317475
rect 249165 318733 249199 318767
rect 229477 309213 229511 309247
rect 249165 309145 249199 309179
rect 283757 317373 283791 317407
rect 229477 309077 229511 309111
rect 233525 309077 233559 309111
rect 233525 305609 233559 305643
rect 238953 309077 238987 309111
rect 229477 299489 229511 299523
rect 283021 309009 283055 309043
rect 238953 299489 238987 299523
rect 251741 307717 251775 307751
rect 260205 307717 260239 307751
rect 283021 302889 283055 302923
rect 288173 317373 288207 317407
rect 284677 309077 284711 309111
rect 288173 307785 288207 307819
rect 284677 302141 284711 302175
rect 283757 299557 283791 299591
rect 260205 299353 260239 299387
rect 251741 298129 251775 298163
rect 237573 298061 237607 298095
rect 283757 298061 283791 298095
rect 251649 292485 251683 292519
rect 237573 288405 237607 288439
rect 243461 289765 243495 289799
rect 251649 287045 251683 287079
rect 277869 289561 277903 289595
rect 243461 280177 243495 280211
rect 229569 280109 229603 280143
rect 229569 270521 229603 270555
rect 243461 278681 243495 278715
rect 241161 270453 241195 270487
rect 241161 260865 241195 260899
rect 229569 260797 229603 260831
rect 259929 278681 259963 278715
rect 283757 288405 283791 288439
rect 288173 298061 288207 298095
rect 288173 288405 288207 288439
rect 277869 277389 277903 277423
rect 259929 267733 259963 267767
rect 253949 260865 253983 260899
rect 253949 258077 253983 258111
rect 243461 256717 243495 256751
rect 260113 258009 260147 258043
rect 229569 251209 229603 251243
rect 243461 255221 243495 255255
rect 237573 248353 237607 248387
rect 237573 244137 237607 244171
rect 260113 249713 260147 249747
rect 260205 258009 260239 258043
rect 260205 248421 260239 248455
rect 275293 249781 275327 249815
rect 275293 248421 275327 248455
rect 243461 240193 243495 240227
rect 258549 244409 258583 244443
rect 258549 240125 258583 240159
rect 260297 240057 260331 240091
rect 254041 238697 254075 238731
rect 243461 237337 243495 237371
rect 237481 231965 237515 231999
rect 237481 227749 237515 227783
rect 260297 230469 260331 230503
rect 254041 230265 254075 230299
rect 277961 225165 277995 225199
rect 251833 224961 251867 224995
rect 251833 222173 251867 222207
rect 277961 220813 277995 220847
rect 243461 219453 243495 219487
rect 270969 220745 271003 220779
rect 237665 219317 237699 219351
rect 243461 219317 243495 219351
rect 237665 214557 237699 214591
rect 238953 218841 238987 218875
rect 238953 205309 238987 205343
rect 270969 211157 271003 211191
rect 277869 219385 277903 219419
rect 277869 209797 277903 209831
rect 275293 209729 275327 209763
rect 275293 205581 275327 205615
rect 243461 202861 243495 202895
rect 260205 201433 260239 201467
rect 260205 191845 260239 191879
rect 243369 191777 243403 191811
rect 243369 186269 243403 186303
rect 270969 191777 271003 191811
rect 260297 183481 260331 183515
rect 243461 182053 243495 182087
rect 243461 174369 243495 174403
rect 258641 180761 258675 180795
rect 256525 173961 256559 173995
rect 237573 172465 237607 172499
rect 237573 166957 237607 166991
rect 238217 172465 238251 172499
rect 275293 190621 275327 190655
rect 275293 190485 275327 190519
rect 270969 182189 271003 182223
rect 260297 178721 260331 178755
rect 270785 180761 270819 180795
rect 258641 171173 258675 171207
rect 270785 171105 270819 171139
rect 275201 180761 275235 180795
rect 275201 171105 275235 171139
rect 256525 169745 256559 169779
rect 258641 171037 258675 171071
rect 238217 162877 238251 162911
rect 241161 162809 241195 162843
rect 259377 171037 259411 171071
rect 275201 170969 275235 171003
rect 259377 161517 259411 161551
rect 260205 162809 260239 162843
rect 258641 161449 258675 161483
rect 259285 160021 259319 160055
rect 243461 157369 243495 157403
rect 243461 153289 243495 153323
rect 241161 153221 241195 153255
rect 237573 153153 237607 153187
rect 237573 147577 237607 147611
rect 238217 153153 238251 153187
rect 238953 153153 238987 153187
rect 258641 151725 258675 151759
rect 238953 147169 238987 147203
rect 256433 149005 256467 149039
rect 238217 143565 238251 143599
rect 237573 143429 237607 143463
rect 237573 133977 237607 134011
rect 243461 142069 243495 142103
rect 238125 133841 238159 133875
rect 254041 142069 254075 142103
rect 251649 137105 251683 137139
rect 251649 132481 251683 132515
rect 258641 142137 258675 142171
rect 275201 161449 275235 161483
rect 260205 153289 260239 153323
rect 259285 142137 259319 142171
rect 276489 144857 276523 144891
rect 256433 139417 256467 139451
rect 276489 135269 276523 135303
rect 278145 135201 278179 135235
rect 254041 132481 254075 132515
rect 260297 133841 260331 133875
rect 243461 124185 243495 124219
rect 258549 131053 258583 131087
rect 238125 122825 238159 122859
rect 241069 124117 241103 124151
rect 238033 121397 238067 121431
rect 238769 121397 238803 121431
rect 238769 115345 238803 115379
rect 253949 122757 253983 122791
rect 241069 114529 241103 114563
rect 243553 118881 243587 118915
rect 238033 113101 238067 113135
rect 256525 122757 256559 122791
rect 260297 124253 260331 124287
rect 275385 133841 275419 133875
rect 278145 128265 278179 128299
rect 275385 124185 275419 124219
rect 258549 121465 258583 121499
rect 260113 124117 260147 124151
rect 260113 114529 260147 114563
rect 260297 124117 260331 124151
rect 260297 114529 260331 114563
rect 272441 121397 272475 121431
rect 256525 113169 256559 113203
rect 253949 111809 253983 111843
rect 272441 111809 272475 111843
rect 276489 119357 276523 119391
rect 258641 111741 258675 111775
rect 243553 108953 243587 108987
rect 251741 110381 251775 110415
rect 248981 106165 249015 106199
rect 238125 102085 238159 102119
rect 237573 95149 237607 95183
rect 258641 102153 258675 102187
rect 272349 111673 272383 111707
rect 276489 107593 276523 107627
rect 278329 114461 278363 114495
rect 278329 104873 278363 104907
rect 272349 102153 272383 102187
rect 251741 100725 251775 100759
rect 260113 102085 260147 102119
rect 248981 97801 249015 97835
rect 258549 97257 258583 97291
rect 238125 92497 238159 92531
rect 253857 95217 253891 95251
rect 253857 91069 253891 91103
rect 237573 85561 237607 85595
rect 243553 86921 243587 86955
rect 237573 82773 237607 82807
rect 229569 80121 229603 80155
rect 229569 77333 229603 77367
rect 229569 77197 229603 77231
rect 248797 86921 248831 86955
rect 249165 86921 249199 86955
rect 248797 82093 248831 82127
rect 248981 86853 249015 86887
rect 248981 78421 249015 78455
rect 243553 77265 243587 77299
rect 260113 92497 260147 92531
rect 272349 97257 272383 97291
rect 258549 84201 258583 84235
rect 260297 86513 260331 86547
rect 249165 77265 249199 77299
rect 251741 84133 251775 84167
rect 259285 84133 259319 84167
rect 253949 80121 253983 80155
rect 253949 75837 253983 75871
rect 251741 74545 251775 74579
rect 260297 75905 260331 75939
rect 259285 74545 259319 74579
rect 275293 93789 275327 93823
rect 275293 84201 275327 84235
rect 272349 74545 272383 74579
rect 237573 73185 237607 73219
rect 238953 74477 238987 74511
rect 229569 67609 229603 67643
rect 258549 74477 258583 74511
rect 238953 64889 238987 64923
rect 240517 67541 240551 67575
rect 238217 64821 238251 64855
rect 229569 57885 229603 57919
rect 258549 64957 258583 64991
rect 240517 57953 240551 57987
rect 241161 64821 241195 64855
rect 238217 55233 238251 55267
rect 241161 55233 241195 55267
rect 258641 63461 258675 63495
rect 238953 55165 238987 55199
rect 229569 48297 229603 48331
rect 238217 51085 238251 51119
rect 238217 46937 238251 46971
rect 238953 45577 238987 45611
rect 243461 48229 243495 48263
rect 237573 45509 237607 45543
rect 229569 38573 229603 38607
rect 238309 45509 238343 45543
rect 238309 35989 238343 36023
rect 241253 45509 241287 45543
rect 237573 35921 237607 35955
rect 241253 35921 241287 35955
rect 229569 28985 229603 29019
rect 238125 35853 238159 35887
rect 275293 56525 275327 56559
rect 275293 51017 275327 51051
rect 260113 48365 260147 48399
rect 260113 46937 260147 46971
rect 260297 48365 260331 48399
rect 260297 46937 260331 46971
rect 258641 45577 258675 45611
rect 278053 46869 278087 46903
rect 278053 37281 278087 37315
rect 243461 27625 243495 27659
rect 256617 35853 256651 35887
rect 238125 26265 238159 26299
rect 243461 27489 243495 27523
rect 256617 26265 256651 26299
rect 259285 35853 259319 35887
rect 259285 26265 259319 26299
rect 278237 27489 278271 27523
rect 243461 22049 243495 22083
rect 274925 26197 274959 26231
rect 238861 21437 238895 21471
rect 259929 19465 259963 19499
rect 238861 16609 238895 16643
rect 253949 18037 253983 18071
rect 259929 17969 259963 18003
rect 253949 16609 253983 16643
rect 260205 17833 260239 17867
rect 237573 16541 237607 16575
rect 237573 9265 237607 9299
rect 274925 16609 274959 16643
rect 276489 19261 276523 19295
rect 276489 9673 276523 9707
rect 278237 9673 278271 9707
rect 260205 8313 260239 8347
rect 275385 8245 275419 8279
rect 244289 5457 244323 5491
rect 244289 5185 244323 5219
rect 224141 4981 224175 5015
rect 224233 4981 224267 5015
rect 224233 4777 224267 4811
rect 224141 4573 224175 4607
rect 93961 4029 93995 4063
rect 74549 3961 74583 3995
rect 74549 3077 74583 3111
rect 84025 3961 84059 3995
rect 84025 3077 84059 3111
rect 93869 3961 93903 3995
rect 93869 2941 93903 2975
rect 93961 2873 93995 2907
rect 103345 4029 103379 4063
rect 232329 4029 232363 4063
rect 103437 3961 103471 3995
rect 231133 3553 231167 3587
rect 232421 4029 232455 4063
rect 248981 3893 249015 3927
rect 232421 3689 232455 3723
rect 233065 3689 233099 3723
rect 232329 3417 232363 3451
rect 231133 3349 231167 3383
rect 103437 2941 103471 2975
rect 433349 3961 433383 3995
rect 433349 3825 433383 3859
rect 275385 3689 275419 3723
rect 248981 3485 249015 3519
rect 571073 3553 571107 3587
rect 571993 3485 572027 3519
rect 571993 3349 572027 3383
rect 571073 3213 571107 3247
rect 233065 2941 233099 2975
rect 103345 2873 103379 2907
<< metal1 >>
rect 257890 700952 257896 701004
rect 257948 700992 257954 701004
rect 397454 700992 397460 701004
rect 257948 700964 397460 700992
rect 257948 700952 257954 700964
rect 397454 700952 397460 700964
rect 397512 700952 397518 701004
rect 259362 700884 259368 700936
rect 259420 700924 259426 700936
rect 413646 700924 413652 700936
rect 259420 700896 413652 700924
rect 259420 700884 259426 700896
rect 413646 700884 413652 700896
rect 413704 700884 413710 700936
rect 257982 700816 257988 700868
rect 258040 700856 258046 700868
rect 429838 700856 429844 700868
rect 258040 700828 429844 700856
rect 258040 700816 258046 700828
rect 429838 700816 429844 700828
rect 429896 700816 429902 700868
rect 72970 700748 72976 700800
rect 73028 700788 73034 700800
rect 265066 700788 265072 700800
rect 73028 700760 265072 700788
rect 73028 700748 73034 700760
rect 265066 700748 265072 700760
rect 265124 700748 265130 700800
rect 256510 700680 256516 700732
rect 256568 700720 256574 700732
rect 462314 700720 462320 700732
rect 256568 700692 462320 700720
rect 256568 700680 256574 700692
rect 462314 700680 462320 700692
rect 462372 700680 462378 700732
rect 256602 700612 256608 700664
rect 256660 700652 256666 700664
rect 478506 700652 478512 700664
rect 256660 700624 478512 700652
rect 256660 700612 256666 700624
rect 478506 700612 478512 700624
rect 478564 700612 478570 700664
rect 256418 700544 256424 700596
rect 256476 700584 256482 700596
rect 494790 700584 494796 700596
rect 256476 700556 494796 700584
rect 256476 700544 256482 700556
rect 494790 700544 494796 700556
rect 494848 700544 494854 700596
rect 8110 700476 8116 700528
rect 8168 700516 8174 700528
rect 266538 700516 266544 700528
rect 8168 700488 266544 700516
rect 8168 700476 8174 700488
rect 266538 700476 266544 700488
rect 266596 700476 266602 700528
rect 255222 700408 255228 700460
rect 255280 700448 255286 700460
rect 527174 700448 527180 700460
rect 255280 700420 527180 700448
rect 255280 700408 255286 700420
rect 527174 700408 527180 700420
rect 527232 700408 527238 700460
rect 40494 700340 40500 700392
rect 40552 700380 40558 700392
rect 41322 700380 41328 700392
rect 40552 700352 41328 700380
rect 40552 700340 40558 700352
rect 41322 700340 41328 700352
rect 41380 700340 41386 700392
rect 255130 700340 255136 700392
rect 255188 700380 255194 700392
rect 543458 700380 543464 700392
rect 255188 700352 543464 700380
rect 255188 700340 255194 700352
rect 543458 700340 543464 700352
rect 543516 700340 543522 700392
rect 253842 700272 253848 700324
rect 253900 700312 253906 700324
rect 559650 700312 559656 700324
rect 253900 700284 559656 700312
rect 253900 700272 253906 700284
rect 559650 700272 559656 700284
rect 559708 700272 559714 700324
rect 137830 700204 137836 700256
rect 137888 700244 137894 700256
rect 263778 700244 263784 700256
rect 137888 700216 263784 700244
rect 137888 700204 137894 700216
rect 263778 700204 263784 700216
rect 263836 700204 263842 700256
rect 259270 700136 259276 700188
rect 259328 700176 259334 700188
rect 364978 700176 364984 700188
rect 259328 700148 364984 700176
rect 259328 700136 259334 700148
rect 364978 700136 364984 700148
rect 365036 700136 365042 700188
rect 260650 700068 260656 700120
rect 260708 700108 260714 700120
rect 348786 700108 348792 700120
rect 260708 700080 348792 700108
rect 260708 700068 260714 700080
rect 348786 700068 348792 700080
rect 348844 700068 348850 700120
rect 259178 700000 259184 700052
rect 259236 700040 259242 700052
rect 332502 700040 332508 700052
rect 259236 700012 332508 700040
rect 259236 700000 259242 700012
rect 332502 700000 332508 700012
rect 332560 700000 332566 700052
rect 202782 699932 202788 699984
rect 202840 699972 202846 699984
rect 262214 699972 262220 699984
rect 202840 699944 262220 699972
rect 202840 699932 202846 699944
rect 262214 699932 262220 699944
rect 262272 699932 262278 699984
rect 262122 699864 262128 699916
rect 262180 699904 262186 699916
rect 283834 699904 283840 699916
rect 262180 699876 283840 699904
rect 262180 699864 262186 699876
rect 283834 699864 283840 699876
rect 283892 699864 283898 699916
rect 24302 699660 24308 699712
rect 24360 699700 24366 699712
rect 24762 699700 24768 699712
rect 24360 699672 24768 699700
rect 24360 699660 24366 699672
rect 24762 699660 24768 699672
rect 24820 699660 24826 699712
rect 89162 699660 89168 699712
rect 89220 699700 89226 699712
rect 89622 699700 89628 699712
rect 89220 699672 89628 699700
rect 89220 699660 89226 699672
rect 89622 699660 89628 699672
rect 89680 699660 89686 699712
rect 105446 699660 105452 699712
rect 105504 699700 105510 699712
rect 106182 699700 106188 699712
rect 105504 699672 106188 699700
rect 105504 699660 105510 699672
rect 106182 699660 106188 699672
rect 106240 699660 106246 699712
rect 170306 699660 170312 699712
rect 170364 699700 170370 699712
rect 171042 699700 171048 699712
rect 170364 699672 171048 699700
rect 170364 699660 170370 699672
rect 171042 699660 171048 699672
rect 171100 699660 171106 699712
rect 235166 699660 235172 699712
rect 235224 699700 235230 699712
rect 235902 699700 235908 699712
rect 235224 699672 235908 699700
rect 235224 699660 235230 699672
rect 235902 699660 235908 699672
rect 235960 699660 235966 699712
rect 260742 699660 260748 699712
rect 260800 699700 260806 699712
rect 267642 699700 267648 699712
rect 260800 699672 267648 699700
rect 260800 699660 260806 699672
rect 267642 699660 267648 699672
rect 267700 699660 267706 699712
rect 253750 696940 253756 696992
rect 253808 696980 253814 696992
rect 580166 696980 580172 696992
rect 253808 696952 580172 696980
rect 253808 696940 253814 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 154114 695512 154120 695564
rect 154172 695552 154178 695564
rect 154206 695552 154212 695564
rect 154172 695524 154212 695552
rect 154172 695512 154178 695524
rect 154206 695512 154212 695524
rect 154264 695512 154270 695564
rect 219069 695487 219127 695493
rect 219069 695453 219081 695487
rect 219115 695484 219127 695487
rect 219158 695484 219164 695496
rect 219115 695456 219164 695484
rect 219115 695453 219127 695456
rect 219069 695447 219127 695453
rect 219158 695444 219164 695456
rect 219216 695444 219222 695496
rect 154206 688576 154212 688628
rect 154264 688616 154270 688628
rect 154390 688616 154396 688628
rect 154264 688588 154396 688616
rect 154264 688576 154270 688588
rect 154390 688576 154396 688588
rect 154448 688576 154454 688628
rect 299658 688576 299664 688628
rect 299716 688616 299722 688628
rect 300118 688616 300124 688628
rect 299716 688588 300124 688616
rect 299716 688576 299722 688588
rect 300118 688576 300124 688588
rect 300176 688576 300182 688628
rect 299492 685936 301268 685964
rect 219066 685896 219072 685908
rect 219027 685868 219072 685896
rect 219066 685856 219072 685868
rect 219124 685856 219130 685908
rect 253658 685856 253664 685908
rect 253716 685896 253722 685908
rect 299492 685896 299520 685936
rect 253716 685868 299520 685896
rect 301240 685896 301268 685936
rect 580166 685896 580172 685908
rect 301240 685868 580172 685896
rect 253716 685856 253722 685868
rect 580166 685856 580172 685868
rect 580224 685856 580230 685908
rect 154301 685831 154359 685837
rect 154301 685797 154313 685831
rect 154347 685828 154359 685831
rect 154390 685828 154396 685840
rect 154347 685800 154396 685828
rect 154347 685797 154359 685800
rect 154301 685791 154359 685797
rect 154390 685788 154396 685800
rect 154448 685788 154454 685840
rect 299566 684428 299572 684480
rect 299624 684468 299630 684480
rect 299845 684471 299903 684477
rect 299845 684468 299857 684471
rect 299624 684440 299857 684468
rect 299624 684428 299630 684440
rect 299845 684437 299857 684440
rect 299891 684437 299903 684471
rect 299845 684431 299903 684437
rect 154298 676240 154304 676252
rect 154259 676212 154304 676240
rect 154298 676200 154304 676212
rect 154356 676200 154362 676252
rect 218974 676172 218980 676184
rect 218935 676144 218980 676172
rect 218974 676132 218980 676144
rect 219032 676132 219038 676184
rect 154298 673480 154304 673532
rect 154356 673520 154362 673532
rect 154482 673520 154488 673532
rect 154356 673492 154488 673520
rect 154356 673480 154362 673492
rect 154482 673480 154488 673492
rect 154540 673480 154546 673532
rect 252462 673480 252468 673532
rect 252520 673520 252526 673532
rect 580166 673520 580172 673532
rect 252520 673492 580172 673520
rect 252520 673480 252526 673492
rect 580166 673480 580172 673492
rect 580224 673480 580230 673532
rect 218977 666587 219035 666593
rect 218977 666553 218989 666587
rect 219023 666584 219035 666587
rect 219066 666584 219072 666596
rect 219023 666556 219072 666584
rect 219023 666553 219035 666556
rect 218977 666547 219035 666553
rect 219066 666544 219072 666556
rect 219124 666544 219130 666596
rect 299845 666587 299903 666593
rect 299845 666553 299857 666587
rect 299891 666584 299903 666587
rect 299934 666584 299940 666596
rect 299891 666556 299940 666584
rect 299891 666553 299903 666556
rect 299845 666547 299903 666553
rect 299934 666544 299940 666556
rect 299992 666544 299998 666596
rect 219158 659608 219164 659660
rect 219216 659648 219222 659660
rect 219342 659648 219348 659660
rect 219216 659620 219348 659648
rect 219216 659608 219222 659620
rect 219342 659608 219348 659620
rect 219400 659608 219406 659660
rect 219253 656863 219311 656869
rect 219253 656829 219265 656863
rect 219299 656860 219311 656863
rect 219342 656860 219348 656872
rect 219299 656832 219348 656860
rect 219299 656829 219311 656832
rect 219253 656823 219311 656829
rect 219342 656820 219348 656832
rect 219400 656820 219406 656872
rect 154298 654100 154304 654152
rect 154356 654140 154362 654152
rect 154482 654140 154488 654152
rect 154356 654112 154488 654140
rect 154356 654100 154362 654112
rect 154482 654100 154488 654112
rect 154540 654100 154546 654152
rect 3326 652740 3332 652792
rect 3384 652780 3390 652792
rect 267826 652780 267832 652792
rect 3384 652752 267832 652780
rect 3384 652740 3390 652752
rect 267826 652740 267832 652752
rect 267884 652740 267890 652792
rect 252370 650020 252376 650072
rect 252428 650060 252434 650072
rect 580166 650060 580172 650072
rect 252428 650032 580172 650060
rect 252428 650020 252434 650032
rect 580166 650020 580172 650032
rect 580224 650020 580230 650072
rect 219250 647272 219256 647284
rect 219211 647244 219256 647272
rect 219250 647232 219256 647244
rect 219308 647232 219314 647284
rect 299658 647232 299664 647284
rect 299716 647272 299722 647284
rect 299750 647272 299756 647284
rect 299716 647244 299756 647272
rect 299716 647232 299722 647244
rect 299750 647232 299756 647244
rect 299808 647232 299814 647284
rect 219250 640404 219256 640416
rect 219084 640376 219256 640404
rect 219084 640280 219112 640376
rect 219250 640364 219256 640376
rect 219308 640364 219314 640416
rect 299658 640364 299664 640416
rect 299716 640404 299722 640416
rect 299750 640404 299756 640416
rect 299716 640376 299756 640404
rect 299716 640364 299722 640376
rect 299750 640364 299756 640376
rect 299808 640364 299814 640416
rect 219066 640228 219072 640280
rect 219124 640228 219130 640280
rect 252278 638936 252284 638988
rect 252336 638976 252342 638988
rect 580166 638976 580172 638988
rect 252336 638948 580172 638976
rect 252336 638936 252342 638948
rect 580166 638936 580172 638948
rect 580224 638936 580230 638988
rect 219066 637508 219072 637560
rect 219124 637548 219130 637560
rect 219158 637548 219164 637560
rect 219124 637520 219164 637548
rect 219124 637508 219130 637520
rect 219158 637508 219164 637520
rect 219216 637508 219222 637560
rect 154298 634788 154304 634840
rect 154356 634828 154362 634840
rect 154482 634828 154488 634840
rect 154356 634800 154488 634828
rect 154356 634788 154362 634800
rect 154482 634788 154488 634800
rect 154540 634788 154546 634840
rect 299566 630640 299572 630692
rect 299624 630680 299630 630692
rect 299750 630680 299756 630692
rect 299624 630652 299756 630680
rect 299624 630640 299630 630652
rect 299750 630640 299756 630652
rect 299808 630640 299814 630692
rect 251082 626560 251088 626612
rect 251140 626600 251146 626612
rect 580166 626600 580172 626612
rect 251140 626572 580172 626600
rect 251140 626560 251146 626572
rect 580166 626560 580172 626572
rect 580224 626560 580230 626612
rect 219342 626532 219348 626544
rect 219303 626504 219348 626532
rect 219342 626492 219348 626504
rect 219400 626492 219406 626544
rect 219342 616876 219348 616888
rect 219303 616848 219348 616876
rect 219342 616836 219348 616848
rect 219400 616836 219406 616888
rect 154298 615476 154304 615528
rect 154356 615516 154362 615528
rect 154482 615516 154488 615528
rect 154356 615488 154488 615516
rect 154356 615476 154362 615488
rect 154482 615476 154488 615488
rect 154540 615476 154546 615528
rect 219069 611439 219127 611445
rect 219069 611405 219081 611439
rect 219115 611436 219127 611439
rect 219342 611436 219348 611448
rect 219115 611408 219348 611436
rect 219115 611405 219127 611408
rect 219069 611399 219127 611405
rect 219342 611396 219348 611408
rect 219400 611396 219406 611448
rect 299566 611328 299572 611380
rect 299624 611368 299630 611380
rect 299750 611368 299756 611380
rect 299624 611340 299756 611368
rect 299624 611328 299630 611340
rect 299750 611328 299756 611340
rect 299808 611328 299814 611380
rect 219066 608716 219072 608728
rect 219027 608688 219072 608716
rect 219066 608676 219072 608688
rect 219124 608676 219130 608728
rect 219066 608540 219072 608592
rect 219124 608580 219130 608592
rect 219253 608583 219311 608589
rect 219253 608580 219265 608583
rect 219124 608552 219265 608580
rect 219124 608540 219130 608552
rect 219253 608549 219265 608552
rect 219299 608549 219311 608583
rect 299658 608580 299664 608592
rect 299619 608552 299664 608580
rect 219253 608543 219311 608549
rect 299658 608540 299664 608552
rect 299716 608540 299722 608592
rect 249702 603100 249708 603152
rect 249760 603140 249766 603152
rect 580166 603140 580172 603152
rect 249760 603112 580172 603140
rect 249760 603100 249766 603112
rect 580166 603100 580172 603112
rect 580224 603100 580230 603152
rect 299661 601715 299719 601721
rect 299661 601681 299673 601715
rect 299707 601712 299719 601715
rect 299842 601712 299848 601724
rect 299707 601684 299848 601712
rect 299707 601681 299719 601684
rect 299661 601675 299719 601681
rect 299842 601672 299848 601684
rect 299900 601672 299906 601724
rect 219250 601576 219256 601588
rect 219211 601548 219256 601576
rect 219250 601536 219256 601548
rect 219308 601536 219314 601588
rect 219161 598927 219219 598933
rect 219161 598893 219173 598927
rect 219207 598924 219219 598927
rect 219250 598924 219256 598936
rect 219207 598896 219256 598924
rect 219207 598893 219219 598896
rect 219161 598887 219219 598893
rect 219250 598884 219256 598896
rect 219308 598884 219314 598936
rect 299842 598924 299848 598936
rect 299803 598896 299848 598924
rect 299842 598884 299848 598896
rect 299900 598884 299906 598936
rect 154298 596164 154304 596216
rect 154356 596204 154362 596216
rect 154482 596204 154488 596216
rect 154356 596176 154488 596204
rect 154356 596164 154362 596176
rect 154482 596164 154488 596176
rect 154540 596164 154546 596216
rect 3050 594804 3056 594856
rect 3108 594844 3114 594856
rect 269298 594844 269304 594856
rect 3108 594816 269304 594844
rect 3108 594804 3114 594816
rect 269298 594804 269304 594816
rect 269356 594804 269362 594856
rect 250990 592016 250996 592068
rect 251048 592056 251054 592068
rect 580166 592056 580172 592068
rect 251048 592028 580172 592056
rect 251048 592016 251054 592028
rect 580166 592016 580172 592028
rect 580224 592016 580230 592068
rect 219158 589336 219164 589348
rect 219119 589308 219164 589336
rect 219158 589296 219164 589308
rect 219216 589296 219222 589348
rect 299845 589339 299903 589345
rect 299845 589305 299857 589339
rect 299891 589336 299903 589339
rect 299934 589336 299940 589348
rect 299891 589308 299940 589336
rect 299891 589305 299903 589308
rect 299845 589299 299903 589305
rect 299934 589296 299940 589308
rect 299992 589296 299998 589348
rect 154298 589268 154304 589280
rect 154259 589240 154304 589268
rect 154298 589228 154304 589240
rect 154356 589228 154362 589280
rect 299934 582468 299940 582480
rect 299860 582440 299940 582468
rect 218974 582360 218980 582412
rect 219032 582400 219038 582412
rect 219158 582400 219164 582412
rect 219032 582372 219164 582400
rect 219032 582360 219038 582372
rect 219158 582360 219164 582372
rect 219216 582360 219222 582412
rect 299860 582344 299888 582440
rect 299934 582428 299940 582440
rect 299992 582428 299998 582480
rect 299842 582292 299848 582344
rect 299900 582292 299906 582344
rect 154298 579748 154304 579760
rect 154259 579720 154304 579748
rect 154298 579708 154304 579720
rect 154356 579708 154362 579760
rect 249610 579640 249616 579692
rect 249668 579680 249674 579692
rect 580166 579680 580172 579692
rect 249668 579652 580172 579680
rect 249668 579640 249674 579652
rect 580166 579640 580172 579652
rect 580224 579640 580230 579692
rect 154206 579572 154212 579624
rect 154264 579612 154270 579624
rect 154390 579612 154396 579624
rect 154264 579584 154396 579612
rect 154264 579572 154270 579584
rect 154390 579572 154396 579584
rect 154448 579572 154454 579624
rect 218885 579615 218943 579621
rect 218885 579581 218897 579615
rect 218931 579612 218943 579615
rect 218974 579612 218980 579624
rect 218931 579584 218980 579612
rect 218931 579581 218943 579584
rect 218885 579575 218943 579581
rect 218974 579572 218980 579584
rect 219032 579572 219038 579624
rect 218882 569956 218888 569968
rect 218843 569928 218888 569956
rect 218882 569916 218888 569928
rect 218940 569916 218946 569968
rect 299566 563116 299572 563168
rect 299624 563116 299630 563168
rect 218882 563048 218888 563100
rect 218940 563048 218946 563100
rect 154206 562912 154212 562964
rect 154264 562952 154270 562964
rect 154390 562952 154396 562964
rect 154264 562924 154396 562952
rect 154264 562912 154270 562924
rect 154390 562912 154396 562924
rect 154448 562912 154454 562964
rect 218900 562952 218928 563048
rect 299584 563032 299612 563116
rect 299566 562980 299572 563032
rect 299624 562980 299630 563032
rect 218974 562952 218980 562964
rect 218900 562924 218980 562952
rect 218974 562912 218980 562924
rect 219032 562912 219038 562964
rect 248322 556180 248328 556232
rect 248380 556220 248386 556232
rect 580166 556220 580172 556232
rect 248380 556192 580172 556220
rect 248380 556180 248386 556192
rect 580166 556180 580172 556192
rect 580224 556180 580230 556232
rect 299566 553500 299572 553512
rect 299492 553472 299572 553500
rect 218882 553432 218888 553444
rect 218843 553404 218888 553432
rect 218882 553392 218888 553404
rect 218940 553392 218946 553444
rect 299492 553376 299520 553472
rect 299566 553460 299572 553472
rect 299624 553460 299630 553512
rect 299474 553324 299480 553376
rect 299532 553324 299538 553376
rect 2958 552032 2964 552084
rect 3016 552072 3022 552084
rect 262858 552072 262864 552084
rect 3016 552044 262864 552072
rect 3016 552032 3022 552044
rect 262858 552032 262864 552044
rect 262916 552032 262922 552084
rect 218882 550644 218888 550656
rect 218843 550616 218888 550644
rect 218882 550604 218888 550616
rect 218940 550604 218946 550656
rect 249518 545096 249524 545148
rect 249576 545136 249582 545148
rect 580166 545136 580172 545148
rect 249576 545108 580172 545136
rect 249576 545096 249582 545108
rect 580166 545096 580172 545108
rect 580224 545096 580230 545148
rect 218882 543736 218888 543788
rect 218940 543736 218946 543788
rect 218900 543640 218928 543736
rect 299290 543668 299296 543720
rect 299348 543708 299354 543720
rect 299474 543708 299480 543720
rect 299348 543680 299480 543708
rect 299348 543668 299354 543680
rect 299474 543668 299480 543680
rect 299532 543668 299538 543720
rect 218974 543640 218980 543652
rect 218900 543612 218980 543640
rect 218974 543600 218980 543612
rect 219032 543600 219038 543652
rect 3142 538228 3148 538280
rect 3200 538268 3206 538280
rect 270770 538268 270776 538280
rect 3200 538240 270776 538268
rect 3200 538228 3206 538240
rect 270770 538228 270776 538240
rect 270828 538228 270834 538280
rect 248230 532720 248236 532772
rect 248288 532760 248294 532772
rect 580166 532760 580172 532772
rect 248288 532732 580172 532760
rect 248288 532720 248294 532732
rect 580166 532720 580172 532732
rect 580224 532720 580230 532772
rect 299566 531292 299572 531344
rect 299624 531332 299630 531344
rect 299750 531332 299756 531344
rect 299624 531304 299756 531332
rect 299624 531292 299630 531304
rect 299750 531292 299756 531304
rect 299808 531292 299814 531344
rect 154390 531264 154396 531276
rect 154351 531236 154396 531264
rect 154390 531224 154396 531236
rect 154448 531224 154454 531276
rect 299750 524424 299756 524476
rect 299808 524424 299814 524476
rect 299768 524396 299796 524424
rect 299842 524396 299848 524408
rect 299768 524368 299848 524396
rect 299842 524356 299848 524368
rect 299900 524356 299906 524408
rect 218974 524288 218980 524340
rect 219032 524328 219038 524340
rect 219158 524328 219164 524340
rect 219032 524300 219164 524328
rect 219032 524288 219038 524300
rect 219158 524288 219164 524300
rect 219216 524288 219222 524340
rect 154393 521679 154451 521685
rect 154393 521645 154405 521679
rect 154439 521676 154451 521679
rect 154482 521676 154488 521688
rect 154439 521648 154488 521676
rect 154439 521645 154451 521648
rect 154393 521639 154451 521645
rect 154482 521636 154488 521648
rect 154540 521636 154546 521688
rect 218790 514632 218796 514684
rect 218848 514672 218854 514684
rect 219066 514672 219072 514684
rect 218848 514644 219072 514672
rect 218848 514632 218854 514644
rect 219066 514632 219072 514644
rect 219124 514632 219130 514684
rect 299658 511980 299664 512032
rect 299716 512020 299722 512032
rect 299934 512020 299940 512032
rect 299716 511992 299940 512020
rect 299716 511980 299722 511992
rect 299934 511980 299940 511992
rect 299992 511980 299998 512032
rect 154390 511952 154396 511964
rect 154351 511924 154396 511952
rect 154390 511912 154396 511924
rect 154448 511912 154454 511964
rect 219066 510592 219072 510604
rect 219027 510564 219072 510592
rect 219066 510552 219072 510564
rect 219124 510552 219130 510604
rect 246942 509260 246948 509312
rect 247000 509300 247006 509312
rect 580166 509300 580172 509312
rect 247000 509272 580172 509300
rect 247000 509260 247006 509272
rect 580166 509260 580172 509272
rect 580224 509260 580230 509312
rect 219066 505084 219072 505096
rect 219027 505056 219072 505084
rect 219066 505044 219072 505056
rect 219124 505044 219130 505096
rect 154393 502367 154451 502373
rect 154393 502333 154405 502367
rect 154439 502364 154451 502367
rect 154482 502364 154488 502376
rect 154439 502336 154488 502364
rect 154439 502333 154451 502336
rect 154393 502327 154451 502333
rect 154482 502324 154488 502336
rect 154540 502324 154546 502376
rect 299750 502324 299756 502376
rect 299808 502364 299814 502376
rect 299934 502364 299940 502376
rect 299808 502336 299940 502364
rect 299808 502324 299814 502336
rect 299934 502324 299940 502336
rect 299992 502324 299998 502376
rect 248138 498176 248144 498228
rect 248196 498216 248202 498228
rect 580166 498216 580172 498228
rect 248196 498188 580172 498216
rect 248196 498176 248202 498188
rect 580166 498176 580172 498188
rect 580224 498176 580230 498228
rect 3326 495456 3332 495508
rect 3384 495496 3390 495508
rect 264238 495496 264244 495508
rect 3384 495468 264244 495496
rect 3384 495456 3390 495468
rect 264238 495456 264244 495468
rect 264296 495456 264302 495508
rect 219066 492668 219072 492720
rect 219124 492708 219130 492720
rect 219158 492708 219164 492720
rect 219124 492680 219164 492708
rect 219124 492668 219130 492680
rect 219158 492668 219164 492680
rect 219216 492668 219222 492720
rect 154206 492600 154212 492652
rect 154264 492640 154270 492652
rect 154390 492640 154396 492652
rect 154264 492612 154396 492640
rect 154264 492600 154270 492612
rect 154390 492600 154396 492612
rect 154448 492600 154454 492652
rect 299658 492640 299664 492652
rect 299619 492612 299664 492640
rect 299658 492600 299664 492612
rect 299716 492600 299722 492652
rect 219158 485800 219164 485852
rect 219216 485800 219222 485852
rect 246850 485800 246856 485852
rect 246908 485840 246914 485852
rect 580166 485840 580172 485852
rect 246908 485812 580172 485840
rect 246908 485800 246914 485812
rect 580166 485800 580172 485812
rect 580224 485800 580230 485852
rect 219176 485704 219204 485800
rect 299658 485772 299664 485784
rect 299619 485744 299664 485772
rect 299658 485732 299664 485744
rect 299716 485732 299722 485784
rect 219250 485704 219256 485716
rect 219176 485676 219256 485704
rect 219250 485664 219256 485676
rect 219308 485664 219314 485716
rect 3142 480224 3148 480276
rect 3200 480264 3206 480276
rect 272518 480264 272524 480276
rect 3200 480236 272524 480264
rect 3200 480224 3206 480236
rect 272518 480224 272524 480236
rect 272576 480224 272582 480276
rect 299566 476076 299572 476128
rect 299624 476116 299630 476128
rect 299750 476116 299756 476128
rect 299624 476088 299756 476116
rect 299624 476076 299630 476088
rect 299750 476076 299756 476088
rect 299808 476076 299814 476128
rect 299658 473328 299664 473340
rect 299619 473300 299664 473328
rect 299658 473288 299664 473300
rect 299716 473288 299722 473340
rect 154298 466420 154304 466472
rect 154356 466460 154362 466472
rect 154482 466460 154488 466472
rect 154356 466432 154488 466460
rect 154356 466420 154362 466432
rect 154482 466420 154488 466432
rect 154540 466420 154546 466472
rect 218974 466420 218980 466472
rect 219032 466420 219038 466472
rect 218992 466324 219020 466420
rect 299658 466392 299664 466404
rect 299619 466364 299664 466392
rect 299658 466352 299664 466364
rect 299716 466352 299722 466404
rect 219342 466324 219348 466336
rect 218992 466296 219348 466324
rect 219342 466284 219348 466296
rect 219400 466284 219406 466336
rect 245562 462340 245568 462392
rect 245620 462380 245626 462392
rect 580166 462380 580172 462392
rect 245620 462352 580172 462380
rect 245620 462340 245626 462352
rect 580166 462340 580172 462352
rect 580224 462340 580230 462392
rect 299382 460844 299388 460896
rect 299440 460884 299446 460896
rect 299750 460884 299756 460896
rect 299440 460856 299756 460884
rect 299440 460844 299446 460856
rect 299750 460844 299756 460856
rect 299808 460844 299814 460896
rect 154209 454019 154267 454025
rect 154209 453985 154221 454019
rect 154255 454016 154267 454019
rect 154298 454016 154304 454028
rect 154255 453988 154304 454016
rect 154255 453985 154267 453988
rect 154209 453979 154267 453985
rect 154298 453976 154304 453988
rect 154356 453976 154362 454028
rect 218977 454019 219035 454025
rect 218977 453985 218989 454019
rect 219023 454016 219035 454019
rect 219066 454016 219072 454028
rect 219023 453988 219072 454016
rect 219023 453985 219035 453988
rect 218977 453979 219035 453985
rect 219066 453976 219072 453988
rect 219124 453976 219130 454028
rect 299400 451336 299888 451364
rect 245470 451256 245476 451308
rect 245528 451296 245534 451308
rect 299400 451296 299428 451336
rect 245528 451268 299428 451296
rect 299860 451296 299888 451336
rect 580166 451296 580172 451308
rect 299860 451268 580172 451296
rect 245528 451256 245534 451268
rect 580166 451256 580172 451268
rect 580224 451256 580230 451308
rect 299474 449868 299480 449880
rect 299435 449840 299480 449868
rect 299474 449828 299480 449840
rect 299532 449828 299538 449880
rect 154206 444428 154212 444440
rect 154167 444400 154212 444428
rect 154206 444388 154212 444400
rect 154264 444388 154270 444440
rect 218974 444428 218980 444440
rect 218935 444400 218980 444428
rect 218974 444388 218980 444400
rect 219032 444388 219038 444440
rect 299477 440283 299535 440289
rect 299477 440249 299489 440283
rect 299523 440280 299535 440283
rect 299566 440280 299572 440292
rect 299523 440252 299572 440280
rect 299523 440249 299535 440252
rect 299477 440243 299535 440249
rect 299566 440240 299572 440252
rect 299624 440240 299630 440292
rect 245378 438880 245384 438932
rect 245436 438920 245442 438932
rect 580166 438920 580172 438932
rect 245436 438892 580172 438920
rect 245436 438880 245442 438892
rect 580166 438880 580172 438892
rect 580224 438880 580230 438932
rect 2958 437452 2964 437504
rect 3016 437492 3022 437504
rect 265618 437492 265624 437504
rect 3016 437464 265624 437492
rect 3016 437452 3022 437464
rect 265618 437452 265624 437464
rect 265676 437452 265682 437504
rect 299566 436812 299572 436824
rect 299527 436784 299572 436812
rect 299566 436772 299572 436784
rect 299624 436772 299630 436824
rect 218974 434664 218980 434716
rect 219032 434704 219038 434716
rect 219066 434704 219072 434716
rect 219032 434676 219072 434704
rect 219032 434664 219038 434676
rect 219066 434664 219072 434676
rect 219124 434664 219130 434716
rect 154298 427796 154304 427848
rect 154356 427796 154362 427848
rect 154316 427768 154344 427796
rect 154390 427768 154396 427780
rect 154316 427740 154396 427768
rect 154390 427728 154396 427740
rect 154448 427728 154454 427780
rect 299566 427768 299572 427780
rect 299527 427740 299572 427768
rect 299566 427728 299572 427740
rect 299624 427728 299630 427780
rect 154114 425008 154120 425060
rect 154172 425048 154178 425060
rect 154390 425048 154396 425060
rect 154172 425020 154396 425048
rect 154172 425008 154178 425020
rect 154390 425008 154396 425020
rect 154448 425008 154454 425060
rect 3326 423648 3332 423700
rect 3384 423688 3390 423700
rect 273898 423688 273904 423700
rect 3384 423660 273904 423688
rect 3384 423648 3390 423660
rect 273898 423648 273904 423660
rect 273956 423648 273962 423700
rect 244182 415420 244188 415472
rect 244240 415460 244246 415472
rect 580166 415460 580172 415472
rect 244240 415432 580172 415460
rect 244240 415420 244246 415432
rect 580166 415420 580172 415432
rect 580224 415420 580230 415472
rect 299661 415395 299719 415401
rect 299661 415361 299673 415395
rect 299707 415392 299719 415395
rect 299750 415392 299756 415404
rect 299707 415364 299756 415392
rect 299707 415361 299719 415364
rect 299661 415355 299719 415361
rect 299750 415352 299756 415364
rect 299808 415352 299814 415404
rect 154482 408484 154488 408536
rect 154540 408484 154546 408536
rect 154500 408400 154528 408484
rect 154482 408348 154488 408400
rect 154540 408348 154546 408400
rect 299658 405736 299664 405748
rect 299619 405708 299664 405736
rect 299658 405696 299664 405708
rect 299716 405696 299722 405748
rect 243814 404336 243820 404388
rect 243872 404376 243878 404388
rect 580166 404376 580172 404388
rect 243872 404348 580172 404376
rect 243872 404336 243878 404348
rect 580166 404336 580172 404348
rect 580224 404336 580230 404388
rect 106182 403152 106188 403164
rect 106108 403124 106188 403152
rect 106108 403016 106136 403124
rect 106182 403112 106188 403124
rect 106240 403112 106246 403164
rect 251177 403155 251235 403161
rect 251177 403121 251189 403155
rect 251223 403152 251235 403155
rect 260745 403155 260803 403161
rect 260745 403152 260757 403155
rect 251223 403124 260757 403152
rect 251223 403121 251235 403124
rect 251177 403115 251235 403121
rect 260745 403121 260757 403124
rect 260791 403121 260803 403155
rect 260745 403115 260803 403121
rect 154577 403087 154635 403093
rect 154577 403053 154589 403087
rect 154623 403084 154635 403087
rect 164145 403087 164203 403093
rect 164145 403084 164157 403087
rect 154623 403056 164157 403084
rect 154623 403053 154635 403056
rect 154577 403047 154635 403053
rect 164145 403053 164157 403056
rect 164191 403053 164203 403087
rect 164145 403047 164203 403053
rect 260745 403019 260803 403025
rect 106108 402988 106228 403016
rect 106200 402948 106228 402988
rect 260745 402985 260757 403019
rect 260791 403016 260803 403019
rect 264882 403016 264888 403028
rect 260791 402988 264888 403016
rect 260791 402985 260803 402988
rect 260745 402979 260803 402985
rect 264882 402976 264888 402988
rect 264940 402976 264946 403028
rect 154577 402951 154635 402957
rect 154577 402948 154589 402951
rect 106200 402920 154589 402948
rect 154577 402917 154589 402920
rect 154623 402917 154635 402951
rect 154577 402911 154635 402917
rect 164145 402951 164203 402957
rect 164145 402917 164157 402951
rect 164191 402948 164203 402951
rect 251177 402951 251235 402957
rect 251177 402948 251189 402951
rect 164191 402920 251189 402948
rect 164191 402917 164203 402920
rect 164145 402911 164203 402917
rect 251177 402917 251189 402920
rect 251223 402917 251235 402951
rect 251177 402911 251235 402917
rect 255961 402951 256019 402957
rect 255961 402917 255973 402951
rect 256007 402948 256019 402951
rect 261297 402951 261355 402957
rect 261297 402948 261309 402951
rect 256007 402920 261309 402948
rect 256007 402917 256019 402920
rect 255961 402911 256019 402917
rect 261297 402917 261309 402920
rect 261343 402917 261355 402951
rect 261297 402911 261355 402917
rect 264238 402908 264244 402960
rect 264296 402948 264302 402960
rect 273806 402948 273812 402960
rect 264296 402920 273812 402948
rect 264296 402908 264302 402920
rect 273806 402908 273812 402920
rect 273864 402908 273870 402960
rect 273898 402908 273904 402960
rect 273956 402948 273962 402960
rect 274910 402948 274916 402960
rect 273956 402920 274916 402948
rect 273956 402908 273962 402920
rect 274910 402908 274916 402920
rect 274968 402908 274974 402960
rect 89622 402840 89628 402892
rect 89680 402880 89686 402892
rect 89680 402852 254900 402880
rect 89680 402840 89686 402852
rect 41322 402772 41328 402824
rect 41380 402812 41386 402824
rect 105909 402815 105967 402821
rect 105909 402812 105921 402815
rect 41380 402784 105921 402812
rect 41380 402772 41386 402784
rect 105909 402781 105921 402784
rect 105955 402781 105967 402815
rect 105909 402775 105967 402781
rect 106001 402815 106059 402821
rect 106001 402781 106013 402815
rect 106047 402812 106059 402815
rect 254765 402815 254823 402821
rect 254765 402812 254777 402815
rect 106047 402784 254777 402812
rect 106047 402781 106059 402784
rect 106001 402775 106059 402781
rect 254765 402781 254777 402784
rect 254811 402781 254823 402815
rect 254872 402812 254900 402852
rect 255406 402840 255412 402892
rect 255464 402880 255470 402892
rect 256418 402880 256424 402892
rect 255464 402852 256424 402880
rect 255464 402840 255470 402852
rect 256418 402840 256424 402852
rect 256476 402840 256482 402892
rect 256970 402840 256976 402892
rect 257028 402880 257034 402892
rect 257982 402880 257988 402892
rect 257028 402852 257988 402880
rect 257028 402840 257034 402852
rect 257982 402840 257988 402852
rect 258040 402840 258046 402892
rect 258534 402840 258540 402892
rect 258592 402880 258598 402892
rect 259270 402880 259276 402892
rect 258592 402852 259276 402880
rect 258592 402840 258598 402852
rect 259270 402840 259276 402852
rect 259328 402840 259334 402892
rect 259638 402840 259644 402892
rect 259696 402880 259702 402892
rect 260650 402880 260656 402892
rect 259696 402852 260656 402880
rect 259696 402840 259702 402852
rect 260650 402840 260656 402852
rect 260708 402840 260714 402892
rect 261202 402840 261208 402892
rect 261260 402880 261266 402892
rect 262122 402880 262128 402892
rect 261260 402852 262128 402880
rect 261260 402840 261266 402852
rect 262122 402840 262128 402852
rect 262180 402840 262186 402892
rect 265618 402840 265624 402892
rect 265676 402880 265682 402892
rect 275370 402880 275376 402892
rect 265676 402852 275376 402880
rect 265676 402840 265682 402852
rect 275370 402840 275376 402852
rect 275428 402840 275434 402892
rect 265894 402812 265900 402824
rect 254872 402784 265900 402812
rect 254765 402775 254823 402781
rect 265894 402772 265900 402784
rect 265952 402772 265958 402824
rect 24762 402704 24768 402756
rect 24820 402744 24826 402756
rect 105725 402747 105783 402753
rect 105725 402744 105737 402747
rect 24820 402716 105737 402744
rect 24820 402704 24826 402716
rect 105725 402713 105737 402716
rect 105771 402713 105783 402747
rect 105725 402707 105783 402713
rect 106093 402747 106151 402753
rect 106093 402713 106105 402747
rect 106139 402744 106151 402747
rect 254121 402747 254179 402753
rect 254121 402744 254133 402747
rect 106139 402716 254133 402744
rect 106139 402713 106151 402716
rect 106093 402707 106151 402713
rect 254121 402713 254133 402716
rect 254167 402713 254179 402747
rect 254121 402707 254179 402713
rect 254394 402704 254400 402756
rect 254452 402744 254458 402756
rect 255222 402744 255228 402756
rect 254452 402716 255228 402744
rect 254452 402704 254458 402716
rect 255222 402704 255228 402716
rect 255280 402704 255286 402756
rect 257893 402747 257951 402753
rect 257893 402713 257905 402747
rect 257939 402744 257951 402747
rect 262766 402744 262772 402756
rect 257939 402716 262772 402744
rect 257939 402713 257951 402716
rect 257893 402707 257951 402713
rect 262766 402704 262772 402716
rect 262824 402704 262830 402756
rect 3418 402636 3424 402688
rect 3476 402676 3482 402688
rect 255961 402679 256019 402685
rect 255961 402676 255973 402679
rect 3476 402648 255973 402676
rect 3476 402636 3482 402648
rect 255961 402645 255973 402648
rect 256007 402645 256019 402679
rect 255961 402639 256019 402645
rect 261297 402679 261355 402685
rect 261297 402645 261309 402679
rect 261343 402676 261355 402679
rect 268010 402676 268016 402688
rect 261343 402648 268016 402676
rect 261343 402645 261355 402648
rect 261297 402639 261355 402645
rect 268010 402636 268016 402648
rect 268068 402636 268074 402688
rect 3602 402568 3608 402620
rect 3660 402608 3666 402620
rect 254213 402611 254271 402617
rect 254213 402608 254225 402611
rect 3660 402580 254225 402608
rect 3660 402568 3666 402580
rect 254213 402577 254225 402580
rect 254259 402577 254271 402611
rect 254213 402571 254271 402577
rect 254765 402611 254823 402617
rect 254765 402577 254777 402611
rect 254811 402608 254823 402611
rect 266446 402608 266452 402620
rect 254811 402580 266452 402608
rect 254811 402577 254823 402580
rect 254765 402571 254823 402577
rect 266446 402568 266452 402580
rect 266504 402568 266510 402620
rect 3510 402500 3516 402552
rect 3568 402540 3574 402552
rect 269114 402540 269120 402552
rect 3568 402512 269120 402540
rect 3568 402500 3574 402512
rect 269114 402500 269120 402512
rect 269172 402500 269178 402552
rect 3878 402432 3884 402484
rect 3936 402472 3942 402484
rect 271230 402472 271236 402484
rect 3936 402444 271236 402472
rect 3936 402432 3942 402444
rect 271230 402432 271236 402444
rect 271288 402432 271294 402484
rect 3694 402364 3700 402416
rect 3752 402404 3758 402416
rect 270678 402404 270684 402416
rect 3752 402376 270684 402404
rect 3752 402364 3758 402376
rect 270678 402364 270684 402376
rect 270736 402364 270742 402416
rect 4062 402296 4068 402348
rect 4120 402336 4126 402348
rect 272794 402336 272800 402348
rect 4120 402308 272800 402336
rect 4120 402296 4126 402308
rect 272794 402296 272800 402308
rect 272852 402296 272858 402348
rect 3234 402228 3240 402280
rect 3292 402268 3298 402280
rect 274358 402268 274364 402280
rect 3292 402240 274364 402268
rect 3292 402228 3298 402240
rect 274358 402228 274364 402240
rect 274416 402228 274422 402280
rect 154482 402160 154488 402212
rect 154540 402200 154546 402212
rect 257985 402203 258043 402209
rect 257985 402200 257997 402203
rect 154540 402172 257997 402200
rect 154540 402160 154546 402172
rect 257985 402169 257997 402172
rect 258031 402169 258043 402203
rect 257985 402163 258043 402169
rect 258074 402160 258080 402212
rect 258132 402200 258138 402212
rect 259362 402200 259368 402212
rect 258132 402172 259368 402200
rect 258132 402160 258138 402172
rect 259362 402160 259368 402172
rect 259420 402160 259426 402212
rect 269574 402200 269580 402212
rect 259472 402172 269580 402200
rect 171042 402092 171048 402144
rect 171100 402132 171106 402144
rect 253937 402135 253995 402141
rect 253937 402132 253949 402135
rect 171100 402104 253949 402132
rect 171100 402092 171106 402104
rect 253937 402101 253949 402104
rect 253983 402101 253995 402135
rect 253937 402095 253995 402101
rect 254213 402135 254271 402141
rect 254213 402101 254225 402135
rect 254259 402132 254271 402135
rect 259472 402132 259500 402172
rect 269574 402160 269580 402172
rect 269632 402160 269638 402212
rect 261754 402132 261760 402144
rect 254259 402104 259500 402132
rect 259564 402104 261760 402132
rect 254259 402101 254271 402104
rect 254213 402095 254271 402101
rect 219342 402024 219348 402076
rect 219400 402064 219406 402076
rect 254029 402067 254087 402073
rect 254029 402064 254041 402067
rect 219400 402036 254041 402064
rect 219400 402024 219406 402036
rect 254029 402033 254041 402036
rect 254075 402033 254087 402067
rect 254029 402027 254087 402033
rect 254121 402067 254179 402073
rect 254121 402033 254133 402067
rect 254167 402064 254179 402067
rect 259457 402067 259515 402073
rect 259457 402064 259469 402067
rect 254167 402036 259469 402064
rect 254167 402033 254179 402036
rect 254121 402027 254179 402033
rect 259457 402033 259469 402036
rect 259503 402033 259515 402067
rect 259457 402027 259515 402033
rect 242250 401956 242256 402008
rect 242308 401996 242314 402008
rect 244829 401999 244887 402005
rect 244829 401996 244841 401999
rect 242308 401968 244841 401996
rect 242308 401956 242314 401968
rect 244829 401965 244841 401968
rect 244875 401965 244887 401999
rect 244829 401959 244887 401965
rect 244918 401956 244924 402008
rect 244976 401996 244982 402008
rect 245562 401996 245568 402008
rect 244976 401968 245568 401996
rect 244976 401956 244982 401968
rect 245562 401956 245568 401968
rect 245620 401956 245626 402008
rect 247034 401956 247040 402008
rect 247092 401996 247098 402008
rect 248138 401996 248144 402008
rect 247092 401968 248144 401996
rect 247092 401956 247098 401968
rect 248138 401956 248144 401968
rect 248196 401956 248202 402008
rect 248598 401956 248604 402008
rect 248656 401996 248662 402008
rect 249518 401996 249524 402008
rect 248656 401968 249524 401996
rect 248656 401956 248662 401968
rect 249518 401956 249524 401968
rect 249576 401956 249582 402008
rect 250162 401956 250168 402008
rect 250220 401996 250226 402008
rect 250990 401996 250996 402008
rect 250220 401968 250996 401996
rect 250220 401956 250226 401968
rect 250990 401956 250996 401968
rect 251048 401956 251054 402008
rect 251174 401956 251180 402008
rect 251232 401996 251238 402008
rect 252370 401996 252376 402008
rect 251232 401968 252376 401996
rect 251232 401956 251238 401968
rect 252370 401956 252376 401968
rect 252428 401956 252434 402008
rect 252738 401956 252744 402008
rect 252796 401996 252802 402008
rect 253750 401996 253756 402008
rect 252796 401968 253756 401996
rect 252796 401956 252802 401968
rect 253750 401956 253756 401968
rect 253808 401956 253814 402008
rect 259564 401996 259592 402104
rect 261754 402092 261760 402104
rect 261812 402092 261818 402144
rect 262858 402092 262864 402144
rect 262916 402132 262922 402144
rect 272242 402132 272248 402144
rect 262916 402104 272248 402132
rect 262916 402092 262922 402104
rect 272242 402092 272248 402104
rect 272300 402092 272306 402144
rect 259641 402067 259699 402073
rect 259641 402033 259653 402067
rect 259687 402064 259699 402067
rect 267550 402064 267556 402076
rect 259687 402036 267556 402064
rect 259687 402033 259699 402036
rect 259641 402027 259699 402033
rect 267550 402024 267556 402036
rect 267608 402024 267614 402076
rect 272337 402067 272395 402073
rect 272337 402033 272349 402067
rect 272383 402064 272395 402067
rect 277026 402064 277032 402076
rect 272383 402036 277032 402064
rect 272383 402033 272395 402036
rect 272337 402027 272395 402033
rect 277026 402024 277032 402036
rect 277084 402024 277090 402076
rect 253952 401968 259592 401996
rect 235902 401888 235908 401940
rect 235960 401928 235966 401940
rect 253952 401928 253980 401968
rect 260190 401956 260196 402008
rect 260248 401996 260254 402008
rect 299658 401996 299664 402008
rect 260248 401968 299664 401996
rect 260248 401956 260254 401968
rect 299658 401956 299664 401968
rect 299716 401956 299722 402008
rect 235960 401900 253980 401928
rect 254029 401931 254087 401937
rect 235960 401888 235966 401900
rect 254029 401897 254041 401931
rect 254075 401928 254087 401931
rect 257893 401931 257951 401937
rect 257893 401928 257905 401931
rect 254075 401900 257905 401928
rect 254075 401897 254087 401900
rect 254029 401891 254087 401897
rect 257893 401897 257905 401900
rect 257939 401897 257951 401931
rect 257893 401891 257951 401897
rect 257985 401931 258043 401937
rect 257985 401897 257997 401931
rect 258031 401928 258043 401931
rect 264330 401928 264336 401940
rect 258031 401900 264336 401928
rect 258031 401897 258043 401900
rect 257985 401891 258043 401897
rect 264330 401888 264336 401900
rect 264388 401888 264394 401940
rect 264974 401888 264980 401940
rect 265032 401928 265038 401940
rect 272337 401931 272395 401937
rect 272337 401928 272349 401931
rect 265032 401900 272349 401928
rect 265032 401888 265038 401900
rect 272337 401897 272349 401900
rect 272383 401897 272395 401931
rect 272337 401891 272395 401897
rect 272518 401888 272524 401940
rect 272576 401928 272582 401940
rect 273254 401928 273260 401940
rect 272576 401900 273260 401928
rect 272576 401888 272582 401900
rect 273254 401888 273260 401900
rect 273312 401888 273318 401940
rect 243262 401820 243268 401872
rect 243320 401860 243326 401872
rect 244182 401860 244188 401872
rect 243320 401832 244188 401860
rect 243320 401820 243326 401832
rect 244182 401820 244188 401832
rect 244240 401820 244246 401872
rect 244366 401820 244372 401872
rect 244424 401860 244430 401872
rect 245378 401860 245384 401872
rect 244424 401832 245384 401860
rect 244424 401820 244430 401832
rect 245378 401820 245384 401832
rect 245436 401820 245442 401872
rect 245930 401820 245936 401872
rect 245988 401860 245994 401872
rect 246850 401860 246856 401872
rect 245988 401832 246856 401860
rect 245988 401820 245994 401832
rect 246850 401820 246856 401832
rect 246908 401820 246914 401872
rect 247494 401820 247500 401872
rect 247552 401860 247558 401872
rect 248230 401860 248236 401872
rect 247552 401832 248236 401860
rect 247552 401820 247558 401832
rect 248230 401820 248236 401832
rect 248288 401820 248294 401872
rect 248325 401863 248383 401869
rect 248325 401829 248337 401863
rect 248371 401860 248383 401863
rect 489178 401860 489184 401872
rect 248371 401832 489184 401860
rect 248371 401829 248383 401832
rect 248325 401823 248383 401829
rect 489178 401820 489184 401832
rect 489236 401820 489242 401872
rect 3326 401752 3332 401804
rect 3384 401792 3390 401804
rect 278590 401792 278596 401804
rect 3384 401764 278596 401792
rect 3384 401752 3390 401764
rect 278590 401752 278596 401764
rect 278648 401752 278654 401804
rect 3970 401684 3976 401736
rect 4028 401724 4034 401736
rect 280154 401724 280160 401736
rect 4028 401696 280160 401724
rect 4028 401684 4034 401696
rect 280154 401684 280160 401696
rect 280212 401684 280218 401736
rect 3786 401616 3792 401668
rect 3844 401656 3850 401668
rect 281718 401656 281724 401668
rect 3844 401628 281724 401656
rect 3844 401616 3850 401628
rect 281718 401616 281724 401628
rect 281776 401616 281782 401668
rect 244829 401591 244887 401597
rect 244829 401557 244841 401591
rect 244875 401588 244887 401591
rect 248325 401591 248383 401597
rect 248325 401588 248337 401591
rect 244875 401560 248337 401588
rect 244875 401557 244887 401560
rect 244829 401551 244887 401557
rect 248325 401557 248337 401560
rect 248371 401557 248383 401591
rect 248325 401551 248383 401557
rect 253937 401591 253995 401597
rect 253937 401557 253949 401591
rect 253983 401588 253995 401591
rect 262950 401588 262956 401600
rect 253983 401560 262956 401588
rect 253983 401557 253995 401560
rect 253937 401551 253995 401557
rect 262950 401548 262956 401560
rect 263008 401548 263014 401600
rect 10962 401412 10968 401464
rect 11020 401452 11026 401464
rect 275922 401452 275928 401464
rect 11020 401424 275928 401452
rect 11020 401412 11026 401424
rect 275922 401412 275928 401424
rect 275980 401412 275986 401464
rect 14550 401344 14556 401396
rect 14608 401384 14614 401396
rect 277486 401384 277492 401396
rect 14608 401356 277492 401384
rect 14608 401344 14614 401356
rect 277486 401344 277492 401356
rect 277544 401344 277550 401396
rect 227162 401276 227168 401328
rect 227220 401316 227226 401328
rect 279050 401316 279056 401328
rect 227220 401288 279056 401316
rect 227220 401276 227226 401288
rect 279050 401276 279056 401288
rect 279108 401276 279114 401328
rect 225782 401208 225788 401260
rect 225840 401248 225846 401260
rect 280706 401248 280712 401260
rect 225840 401220 280712 401248
rect 225840 401208 225846 401220
rect 280706 401208 280712 401220
rect 280764 401208 280770 401260
rect 227070 401140 227076 401192
rect 227128 401180 227134 401192
rect 284386 401180 284392 401192
rect 227128 401152 284392 401180
rect 227128 401140 227134 401152
rect 284386 401140 284392 401152
rect 284444 401140 284450 401192
rect 233326 401072 233332 401124
rect 233384 401112 233390 401124
rect 291930 401112 291936 401124
rect 233384 401084 291936 401112
rect 233384 401072 233390 401084
rect 291930 401072 291936 401084
rect 291988 401072 291994 401124
rect 222838 401004 222844 401056
rect 222896 401044 222902 401056
rect 283834 401044 283840 401056
rect 222896 401016 283840 401044
rect 222896 401004 222902 401016
rect 283834 401004 283840 401016
rect 283892 401004 283898 401056
rect 225598 400936 225604 400988
rect 225656 400976 225662 400988
rect 287514 400976 287520 400988
rect 225656 400948 287520 400976
rect 225656 400936 225662 400948
rect 287514 400936 287520 400948
rect 287572 400936 287578 400988
rect 234890 400868 234896 400920
rect 234948 400908 234954 400920
rect 297450 400908 297456 400920
rect 234948 400880 297456 400908
rect 234948 400868 234954 400880
rect 297450 400868 297456 400880
rect 297508 400868 297514 400920
rect 231762 400800 231768 400852
rect 231820 400840 231826 400852
rect 294598 400840 294604 400852
rect 231820 400812 294604 400840
rect 231820 400800 231826 400812
rect 294598 400800 294604 400812
rect 294656 400800 294662 400852
rect 238018 400732 238024 400784
rect 238076 400772 238082 400784
rect 301590 400772 301596 400784
rect 238076 400744 301596 400772
rect 238076 400732 238082 400744
rect 301590 400732 301596 400744
rect 301648 400732 301654 400784
rect 211798 400664 211804 400716
rect 211856 400704 211862 400716
rect 279602 400704 279608 400716
rect 211856 400676 279608 400704
rect 211856 400664 211862 400676
rect 279602 400664 279608 400676
rect 279660 400664 279666 400716
rect 215938 400596 215944 400648
rect 215996 400636 216002 400648
rect 286962 400636 286968 400648
rect 215996 400608 286968 400636
rect 215996 400596 216002 400608
rect 286962 400596 286968 400608
rect 287020 400596 287026 400648
rect 209038 400528 209044 400580
rect 209096 400568 209102 400580
rect 281166 400568 281172 400580
rect 209096 400540 281172 400568
rect 209096 400528 209102 400540
rect 281166 400528 281172 400540
rect 281224 400528 281230 400580
rect 235442 400460 235448 400512
rect 235500 400500 235506 400512
rect 308398 400500 308404 400512
rect 235500 400472 308404 400500
rect 235500 400460 235506 400472
rect 308398 400460 308404 400472
rect 308456 400460 308462 400512
rect 230658 400392 230664 400444
rect 230716 400432 230722 400444
rect 304258 400432 304264 400444
rect 230716 400404 304264 400432
rect 230716 400392 230722 400404
rect 304258 400392 304264 400404
rect 304316 400392 304322 400444
rect 233878 400324 233884 400376
rect 233936 400364 233942 400376
rect 496078 400364 496084 400376
rect 233936 400336 496084 400364
rect 233936 400324 233942 400336
rect 496078 400324 496084 400336
rect 496136 400324 496142 400376
rect 241698 400256 241704 400308
rect 241756 400296 241762 400308
rect 290550 400296 290556 400308
rect 241756 400268 290556 400296
rect 241756 400256 241762 400268
rect 290550 400256 290556 400268
rect 290608 400256 290614 400308
rect 241238 400188 241244 400240
rect 241296 400228 241302 400240
rect 290458 400228 290464 400240
rect 241296 400200 290464 400228
rect 241296 400188 241302 400200
rect 290458 400188 290464 400200
rect 290516 400188 290522 400240
rect 238570 400120 238576 400172
rect 238628 400160 238634 400172
rect 244185 400163 244243 400169
rect 244185 400160 244197 400163
rect 238628 400132 244197 400160
rect 238628 400120 238634 400132
rect 244185 400129 244197 400132
rect 244231 400129 244243 400163
rect 244185 400123 244243 400129
rect 253937 400163 253995 400169
rect 253937 400129 253949 400163
rect 253983 400160 253995 400163
rect 263505 400163 263563 400169
rect 263505 400160 263517 400163
rect 253983 400132 263517 400160
rect 253983 400129 253995 400132
rect 253937 400123 253995 400129
rect 263505 400129 263517 400132
rect 263551 400129 263563 400163
rect 263505 400123 263563 400129
rect 226978 400052 226984 400104
rect 227036 400092 227042 400104
rect 276474 400092 276480 400104
rect 227036 400064 276480 400092
rect 227036 400052 227042 400064
rect 276474 400052 276480 400064
rect 276532 400052 276538 400104
rect 242618 399984 242624 400036
rect 242676 400024 242682 400036
rect 290642 400024 290648 400036
rect 242676 399996 290648 400024
rect 242676 399984 242682 399996
rect 290642 399984 290648 399996
rect 290700 399984 290706 400036
rect 236730 399916 236736 399968
rect 236788 399956 236794 399968
rect 298830 399956 298836 399968
rect 236788 399928 298836 399956
rect 236788 399916 236794 399928
rect 298830 399916 298836 399928
rect 298888 399916 298894 399968
rect 239858 399848 239864 399900
rect 239916 399888 239922 399900
rect 302970 399888 302976 399900
rect 239916 399860 302976 399888
rect 239916 399848 239922 399860
rect 302970 399848 302976 399860
rect 303028 399848 303034 399900
rect 213178 399780 213184 399832
rect 213236 399820 213242 399832
rect 277670 399820 277676 399832
rect 213236 399792 277676 399820
rect 213236 399780 213242 399792
rect 277670 399780 277676 399792
rect 277728 399780 277734 399832
rect 218698 399712 218704 399764
rect 218756 399752 218762 399764
rect 285030 399752 285036 399764
rect 218756 399724 285036 399752
rect 218756 399712 218762 399724
rect 285030 399712 285036 399724
rect 285088 399712 285094 399764
rect 232498 399644 232504 399696
rect 232556 399684 232562 399696
rect 305638 399684 305644 399696
rect 232556 399656 305644 399684
rect 232556 399644 232562 399656
rect 305638 399644 305644 399656
rect 305696 399644 305702 399696
rect 214558 399576 214564 399628
rect 214616 399616 214622 399628
rect 288342 399616 288348 399628
rect 214616 399588 288348 399616
rect 214616 399576 214622 399588
rect 288342 399576 288348 399588
rect 288400 399576 288406 399628
rect 338117 399619 338175 399625
rect 338117 399585 338129 399619
rect 338163 399616 338175 399619
rect 347685 399619 347743 399625
rect 347685 399616 347697 399619
rect 338163 399588 347697 399616
rect 338163 399585 338175 399588
rect 338117 399579 338175 399585
rect 347685 399585 347697 399588
rect 347731 399585 347743 399619
rect 347685 399579 347743 399585
rect 357437 399619 357495 399625
rect 357437 399585 357449 399619
rect 357483 399616 357495 399619
rect 367005 399619 367063 399625
rect 367005 399616 367017 399619
rect 357483 399588 367017 399616
rect 357483 399585 357495 399588
rect 357437 399579 357495 399585
rect 367005 399585 367017 399588
rect 367051 399585 367063 399619
rect 367005 399579 367063 399585
rect 376757 399619 376815 399625
rect 376757 399585 376769 399619
rect 376803 399616 376815 399619
rect 386325 399619 386383 399625
rect 386325 399616 386337 399619
rect 376803 399588 386337 399616
rect 376803 399585 376815 399588
rect 376757 399579 376815 399585
rect 386325 399585 386337 399588
rect 386371 399585 386383 399619
rect 386325 399579 386383 399585
rect 207658 399508 207664 399560
rect 207716 399548 207722 399560
rect 282454 399548 282460 399560
rect 207716 399520 282460 399548
rect 207716 399508 207722 399520
rect 282454 399508 282460 399520
rect 282512 399508 282518 399560
rect 282825 399551 282883 399557
rect 282825 399517 282837 399551
rect 282871 399548 282883 399551
rect 285582 399548 285588 399560
rect 282871 399520 285588 399548
rect 282871 399517 282883 399520
rect 282825 399511 282883 399517
rect 285582 399508 285588 399520
rect 285640 399508 285646 399560
rect 289817 399551 289875 399557
rect 289817 399517 289829 399551
rect 289863 399548 289875 399551
rect 299385 399551 299443 399557
rect 299385 399548 299397 399551
rect 289863 399520 299397 399548
rect 289863 399517 289875 399520
rect 289817 399511 289875 399517
rect 299385 399517 299397 399520
rect 299431 399517 299443 399551
rect 299385 399511 299443 399517
rect 3418 399440 3424 399492
rect 3476 399480 3482 399492
rect 264974 399480 264980 399492
rect 3476 399452 264980 399480
rect 3476 399440 3482 399452
rect 264974 399440 264980 399452
rect 265032 399440 265038 399492
rect 280065 399483 280123 399489
rect 280065 399449 280077 399483
rect 280111 399480 280123 399483
rect 280157 399483 280215 399489
rect 280157 399480 280169 399483
rect 280111 399452 280169 399480
rect 280111 399449 280123 399452
rect 280065 399443 280123 399449
rect 280157 399449 280169 399452
rect 280203 399449 280215 399483
rect 338117 399483 338175 399489
rect 338117 399480 338129 399483
rect 280157 399443 280215 399449
rect 332428 399452 338129 399480
rect 204898 399372 204904 399424
rect 204956 399412 204962 399424
rect 279881 399415 279939 399421
rect 279881 399412 279893 399415
rect 204956 399384 279893 399412
rect 204956 399372 204962 399384
rect 279881 399381 279893 399384
rect 279927 399381 279939 399415
rect 279881 399375 279939 399381
rect 279973 399415 280031 399421
rect 279973 399381 279985 399415
rect 280019 399412 280031 399415
rect 282825 399415 282883 399421
rect 282825 399412 282837 399415
rect 280019 399384 282837 399412
rect 280019 399381 280031 399384
rect 279973 399375 280031 399381
rect 282825 399381 282837 399384
rect 282871 399381 282883 399415
rect 289817 399415 289875 399421
rect 289817 399412 289829 399415
rect 282825 399375 282883 399381
rect 285876 399384 289829 399412
rect 180058 399304 180064 399356
rect 180116 399344 180122 399356
rect 281902 399344 281908 399356
rect 180116 399316 281908 399344
rect 180116 399304 180122 399316
rect 281902 399304 281908 399316
rect 281960 399304 281966 399356
rect 244185 399279 244243 399285
rect 244185 399245 244197 399279
rect 244231 399276 244243 399279
rect 253937 399279 253995 399285
rect 253937 399276 253949 399279
rect 244231 399248 253949 399276
rect 244231 399245 244243 399248
rect 244185 399239 244243 399245
rect 253937 399245 253949 399248
rect 253983 399245 253995 399279
rect 253937 399239 253995 399245
rect 263505 399279 263563 399285
rect 263505 399245 263517 399279
rect 263551 399276 263563 399279
rect 279789 399279 279847 399285
rect 279789 399276 279801 399279
rect 263551 399248 279801 399276
rect 263551 399245 263563 399248
rect 263505 399239 263563 399245
rect 279789 399245 279801 399248
rect 279835 399245 279847 399279
rect 279789 399239 279847 399245
rect 280157 399279 280215 399285
rect 280157 399245 280169 399279
rect 280203 399276 280215 399279
rect 285876 399276 285904 399384
rect 289817 399381 289829 399384
rect 289863 399381 289875 399415
rect 331125 399415 331183 399421
rect 331125 399412 331137 399415
rect 289817 399375 289875 399381
rect 321480 399384 331137 399412
rect 288710 399304 288716 399356
rect 288768 399304 288774 399356
rect 280203 399248 285904 399276
rect 280203 399245 280215 399248
rect 280157 399239 280215 399245
rect 13078 399168 13084 399220
rect 13136 399208 13142 399220
rect 288728 399208 288756 399304
rect 318705 399279 318763 399285
rect 318705 399245 318717 399279
rect 318751 399276 318763 399279
rect 321480 399276 321508 399384
rect 331125 399381 331137 399384
rect 331171 399381 331183 399415
rect 331125 399375 331183 399381
rect 331217 399415 331275 399421
rect 331217 399381 331229 399415
rect 331263 399412 331275 399415
rect 332428 399412 332456 399452
rect 338117 399449 338129 399452
rect 338163 399449 338175 399483
rect 357437 399483 357495 399489
rect 357437 399480 357449 399483
rect 338117 399443 338175 399449
rect 351748 399452 357449 399480
rect 331263 399384 332456 399412
rect 347685 399415 347743 399421
rect 331263 399381 331275 399384
rect 331217 399375 331275 399381
rect 347685 399381 347697 399415
rect 347731 399412 347743 399415
rect 350445 399415 350503 399421
rect 350445 399412 350457 399415
rect 347731 399384 350457 399412
rect 347731 399381 347743 399384
rect 347685 399375 347743 399381
rect 350445 399381 350457 399384
rect 350491 399381 350503 399415
rect 350445 399375 350503 399381
rect 350537 399415 350595 399421
rect 350537 399381 350549 399415
rect 350583 399412 350595 399415
rect 351748 399412 351776 399452
rect 357437 399449 357449 399452
rect 357483 399449 357495 399483
rect 376757 399483 376815 399489
rect 376757 399480 376769 399483
rect 357437 399443 357495 399449
rect 371068 399452 376769 399480
rect 350583 399384 351776 399412
rect 367005 399415 367063 399421
rect 350583 399381 350595 399384
rect 350537 399375 350595 399381
rect 367005 399381 367017 399415
rect 367051 399412 367063 399415
rect 369765 399415 369823 399421
rect 369765 399412 369777 399415
rect 367051 399384 369777 399412
rect 367051 399381 367063 399384
rect 367005 399375 367063 399381
rect 369765 399381 369777 399384
rect 369811 399381 369823 399415
rect 369765 399375 369823 399381
rect 369857 399415 369915 399421
rect 369857 399381 369869 399415
rect 369903 399412 369915 399415
rect 371068 399412 371096 399452
rect 376757 399449 376769 399452
rect 376803 399449 376815 399483
rect 376757 399443 376815 399449
rect 369903 399384 371096 399412
rect 386325 399415 386383 399421
rect 369903 399381 369915 399384
rect 369857 399375 369915 399381
rect 386325 399381 386337 399415
rect 386371 399412 386383 399415
rect 386969 399415 387027 399421
rect 386969 399412 386981 399415
rect 386371 399384 386981 399412
rect 386371 399381 386383 399384
rect 386325 399375 386383 399381
rect 386969 399381 386981 399384
rect 387015 399381 387027 399415
rect 386969 399375 387027 399381
rect 318751 399248 321508 399276
rect 318751 399245 318763 399248
rect 318705 399239 318763 399245
rect 13136 399180 288756 399208
rect 299385 399211 299443 399217
rect 13136 399168 13142 399180
rect 299385 399177 299397 399211
rect 299431 399208 299443 399211
rect 309137 399211 309195 399217
rect 309137 399208 309149 399211
rect 299431 399180 309149 399208
rect 299431 399177 299443 399180
rect 299385 399171 299443 399177
rect 309137 399177 309149 399180
rect 309183 399177 309195 399211
rect 309137 399171 309195 399177
rect 309137 399075 309195 399081
rect 309137 399041 309149 399075
rect 309183 399072 309195 399075
rect 318705 399075 318763 399081
rect 318705 399072 318717 399075
rect 309183 399044 318717 399072
rect 309183 399041 309195 399044
rect 309137 399035 309195 399041
rect 318705 399041 318717 399044
rect 318751 399041 318763 399075
rect 318705 399035 318763 399041
rect 386969 398191 387027 398197
rect 386969 398157 386981 398191
rect 387015 398188 387027 398191
rect 393958 398188 393964 398200
rect 387015 398160 393964 398188
rect 387015 398157 387027 398160
rect 386969 398151 387027 398157
rect 393958 398148 393964 398160
rect 394016 398148 394022 398200
rect 3142 395972 3148 396024
rect 3200 396012 3206 396024
rect 10962 396012 10968 396024
rect 3200 395984 10968 396012
rect 3200 395972 3206 395984
rect 10962 395972 10968 395984
rect 11020 395972 11026 396024
rect 290642 393252 290648 393304
rect 290700 393292 290706 393304
rect 579798 393292 579804 393304
rect 290700 393264 579804 393292
rect 290700 393252 290706 393264
rect 579798 393252 579804 393264
rect 579856 393252 579862 393304
rect 290550 369792 290556 369844
rect 290608 369832 290614 369844
rect 580166 369832 580172 369844
rect 290608 369804 580172 369832
rect 290608 369792 290614 369804
rect 580166 369792 580172 369804
rect 580224 369792 580230 369844
rect 2958 367004 2964 367056
rect 3016 367044 3022 367056
rect 226978 367044 226984 367056
rect 3016 367016 226984 367044
rect 3016 367004 3022 367016
rect 226978 367004 226984 367016
rect 227036 367004 227042 367056
rect 489178 358708 489184 358760
rect 489236 358748 489242 358760
rect 580074 358748 580080 358760
rect 489236 358720 580080 358748
rect 489236 358708 489242 358720
rect 580074 358708 580080 358720
rect 580132 358708 580138 358760
rect 290458 346332 290464 346384
rect 290516 346372 290522 346384
rect 579798 346372 579804 346384
rect 290516 346344 579804 346372
rect 290516 346332 290522 346344
rect 579798 346332 579804 346344
rect 579856 346332 579862 346384
rect 277854 338104 277860 338156
rect 277912 338144 277918 338156
rect 278130 338144 278136 338156
rect 277912 338116 278136 338144
rect 277912 338104 277918 338116
rect 278130 338104 278136 338116
rect 278188 338104 278194 338156
rect 3418 338036 3424 338088
rect 3476 338076 3482 338088
rect 14550 338076 14556 338088
rect 3476 338048 14556 338076
rect 3476 338036 3482 338048
rect 14550 338036 14556 338048
rect 14608 338036 14614 338088
rect 125502 338036 125508 338088
rect 125560 338076 125566 338088
rect 235721 338079 235779 338085
rect 235721 338076 235733 338079
rect 125560 338048 235733 338076
rect 125560 338036 125566 338048
rect 235721 338045 235733 338048
rect 235767 338045 235779 338079
rect 235721 338039 235779 338045
rect 235905 338079 235963 338085
rect 235905 338045 235917 338079
rect 235951 338076 235963 338079
rect 240226 338076 240232 338088
rect 235951 338048 240232 338076
rect 235951 338045 235963 338048
rect 235905 338039 235963 338045
rect 240226 338036 240232 338048
rect 240284 338036 240290 338088
rect 240689 338079 240747 338085
rect 240689 338045 240701 338079
rect 240735 338076 240747 338079
rect 240870 338076 240876 338088
rect 240735 338048 240876 338076
rect 240735 338045 240747 338048
rect 240689 338039 240747 338045
rect 240870 338036 240876 338048
rect 240928 338036 240934 338088
rect 243078 338076 243084 338088
rect 243039 338048 243084 338076
rect 243078 338036 243084 338048
rect 243136 338036 243142 338088
rect 267461 338079 267519 338085
rect 267461 338045 267473 338079
rect 267507 338076 267519 338079
rect 267550 338076 267556 338088
rect 267507 338048 267556 338076
rect 267507 338045 267519 338048
rect 267461 338039 267519 338045
rect 267550 338036 267556 338048
rect 267608 338036 267614 338088
rect 274910 338036 274916 338088
rect 274968 338076 274974 338088
rect 278774 338076 278780 338088
rect 274968 338048 278780 338076
rect 274968 338036 274974 338048
rect 278774 338036 278780 338048
rect 278832 338036 278838 338088
rect 279694 338036 279700 338088
rect 279752 338076 279758 338088
rect 289998 338076 290004 338088
rect 279752 338048 290004 338076
rect 279752 338036 279758 338048
rect 289998 338036 290004 338048
rect 290056 338036 290062 338088
rect 107562 337968 107568 338020
rect 107620 338008 107626 338020
rect 235629 338011 235687 338017
rect 235629 338008 235641 338011
rect 107620 337980 235641 338008
rect 107620 337968 107626 337980
rect 235629 337977 235641 337980
rect 235675 337977 235687 338011
rect 241698 338008 241704 338020
rect 235629 337971 235687 337977
rect 235920 337980 241704 338008
rect 115842 337900 115848 337952
rect 115900 337940 115906 337952
rect 235920 337940 235948 337980
rect 241698 337968 241704 337980
rect 241756 337968 241762 338020
rect 277486 337968 277492 338020
rect 277544 338008 277550 338020
rect 278498 338008 278504 338020
rect 277544 337980 278504 338008
rect 277544 337968 277550 337980
rect 278498 337968 278504 337980
rect 278556 337968 278562 338020
rect 284846 337968 284852 338020
rect 284904 338008 284910 338020
rect 294690 338008 294696 338020
rect 284904 337980 294696 338008
rect 284904 337968 284910 337980
rect 294690 337968 294696 337980
rect 294748 337968 294754 338020
rect 115900 337912 235948 337940
rect 115900 337900 115906 337912
rect 253198 337900 253204 337952
rect 253256 337940 253262 337952
rect 254210 337940 254216 337952
rect 253256 337912 254216 337940
rect 253256 337900 253262 337912
rect 254210 337900 254216 337912
rect 254268 337900 254274 337952
rect 260837 337943 260895 337949
rect 260837 337909 260849 337943
rect 260883 337940 260895 337943
rect 263505 337943 263563 337949
rect 263505 337940 263517 337943
rect 260883 337912 263517 337940
rect 260883 337909 260895 337912
rect 260837 337903 260895 337909
rect 263505 337909 263517 337912
rect 263551 337909 263563 337943
rect 263505 337903 263563 337909
rect 263594 337900 263600 337952
rect 263652 337940 263658 337952
rect 267734 337940 267740 337952
rect 263652 337912 267740 337940
rect 263652 337900 263658 337912
rect 267734 337900 267740 337912
rect 267792 337900 267798 337952
rect 271966 337900 271972 337952
rect 272024 337940 272030 337952
rect 272024 337912 278084 337940
rect 272024 337900 272030 337912
rect 100662 337832 100668 337884
rect 100720 337872 100726 337884
rect 235905 337875 235963 337881
rect 235905 337872 235917 337875
rect 100720 337844 235917 337872
rect 100720 337832 100726 337844
rect 235905 337841 235917 337844
rect 235951 337841 235963 337875
rect 235905 337835 235963 337841
rect 235997 337875 236055 337881
rect 235997 337841 236009 337875
rect 236043 337872 236055 337875
rect 245102 337872 245108 337884
rect 236043 337844 245108 337872
rect 236043 337841 236055 337844
rect 235997 337835 236055 337841
rect 245102 337832 245108 337844
rect 245160 337832 245166 337884
rect 257154 337832 257160 337884
rect 257212 337872 257218 337884
rect 263410 337872 263416 337884
rect 257212 337844 263416 337872
rect 257212 337832 257218 337844
rect 263410 337832 263416 337844
rect 263468 337832 263474 337884
rect 277949 337875 278007 337881
rect 277949 337872 277961 337875
rect 275296 337844 277961 337872
rect 39298 337764 39304 337816
rect 39356 337804 39362 337816
rect 233602 337804 233608 337816
rect 39356 337776 233608 337804
rect 39356 337764 39362 337776
rect 233602 337764 233608 337776
rect 233660 337764 233666 337816
rect 235721 337807 235779 337813
rect 235721 337773 235733 337807
rect 235767 337804 235779 337807
rect 242802 337804 242808 337816
rect 235767 337776 242808 337804
rect 235767 337773 235779 337776
rect 235721 337767 235779 337773
rect 242802 337764 242808 337776
rect 242860 337764 242866 337816
rect 262398 337764 262404 337816
rect 262456 337804 262462 337816
rect 265526 337804 265532 337816
rect 262456 337776 265532 337804
rect 262456 337764 262462 337776
rect 265526 337764 265532 337776
rect 265584 337764 265590 337816
rect 266354 337764 266360 337816
rect 266412 337804 266418 337816
rect 266998 337804 267004 337816
rect 266412 337776 267004 337804
rect 266412 337764 266418 337776
rect 266998 337764 267004 337776
rect 267056 337764 267062 337816
rect 267918 337804 267924 337816
rect 267879 337776 267924 337804
rect 267918 337764 267924 337776
rect 267976 337764 267982 337816
rect 273898 337764 273904 337816
rect 273956 337804 273962 337816
rect 274542 337804 274548 337816
rect 273956 337776 274548 337804
rect 273956 337764 273962 337776
rect 274542 337764 274548 337776
rect 274600 337764 274606 337816
rect 32398 337696 32404 337748
rect 32456 337736 32462 337748
rect 231946 337736 231952 337748
rect 32456 337708 231952 337736
rect 32456 337696 32462 337708
rect 231946 337696 231952 337708
rect 232004 337696 232010 337748
rect 235629 337739 235687 337745
rect 235629 337705 235641 337739
rect 235675 337736 235687 337739
rect 240962 337736 240968 337748
rect 235675 337708 240968 337736
rect 235675 337705 235687 337708
rect 235629 337699 235687 337705
rect 240962 337696 240968 337708
rect 241020 337696 241026 337748
rect 241793 337739 241851 337745
rect 241793 337705 241805 337739
rect 241839 337736 241851 337739
rect 246942 337736 246948 337748
rect 241839 337708 246948 337736
rect 241839 337705 241851 337708
rect 241793 337699 241851 337705
rect 246942 337696 246948 337708
rect 247000 337696 247006 337748
rect 257522 337696 257528 337748
rect 257580 337736 257586 337748
rect 262214 337736 262220 337748
rect 257580 337708 262220 337736
rect 257580 337696 257586 337708
rect 262214 337696 262220 337708
rect 262272 337696 262278 337748
rect 262306 337696 262312 337748
rect 262364 337736 262370 337748
rect 275296 337736 275324 337844
rect 277949 337841 277961 337844
rect 277995 337841 278007 337875
rect 278056 337872 278084 337912
rect 279234 337900 279240 337952
rect 279292 337940 279298 337952
rect 280157 337943 280215 337949
rect 280157 337940 280169 337943
rect 279292 337912 280169 337940
rect 279292 337900 279298 337912
rect 280157 337909 280169 337912
rect 280203 337909 280215 337943
rect 280157 337903 280215 337909
rect 283558 337900 283564 337952
rect 283616 337940 283622 337952
rect 283653 337943 283711 337949
rect 283653 337940 283665 337943
rect 283616 337912 283665 337940
rect 283616 337900 283622 337912
rect 283653 337909 283665 337912
rect 283699 337909 283711 337943
rect 283653 337903 283711 337909
rect 285950 337900 285956 337952
rect 286008 337940 286014 337952
rect 290921 337943 290979 337949
rect 290921 337940 290933 337943
rect 286008 337912 290933 337940
rect 286008 337900 286014 337912
rect 290921 337909 290933 337912
rect 290967 337909 290979 337943
rect 290921 337903 290979 337909
rect 291013 337943 291071 337949
rect 291013 337909 291025 337943
rect 291059 337940 291071 337943
rect 297358 337940 297364 337952
rect 291059 337912 297364 337940
rect 291059 337909 291071 337912
rect 291013 337903 291071 337909
rect 297358 337900 297364 337912
rect 297416 337900 297422 337952
rect 280433 337875 280491 337881
rect 280433 337872 280445 337875
rect 278056 337844 280445 337872
rect 277949 337835 278007 337841
rect 280433 337841 280445 337844
rect 280479 337841 280491 337875
rect 280433 337835 280491 337841
rect 282638 337832 282644 337884
rect 282696 337872 282702 337884
rect 298738 337872 298744 337884
rect 282696 337844 298744 337872
rect 282696 337832 282702 337844
rect 298738 337832 298744 337844
rect 298796 337832 298802 337884
rect 276014 337764 276020 337816
rect 276072 337804 276078 337816
rect 282825 337807 282883 337813
rect 282825 337804 282837 337807
rect 276072 337776 282837 337804
rect 276072 337764 276078 337776
rect 282825 337773 282837 337776
rect 282871 337773 282883 337807
rect 282825 337767 282883 337773
rect 283006 337764 283012 337816
rect 283064 337804 283070 337816
rect 287333 337807 287391 337813
rect 287333 337804 287345 337807
rect 283064 337776 287345 337804
rect 283064 337764 283070 337776
rect 287333 337773 287345 337776
rect 287379 337773 287391 337807
rect 287333 337767 287391 337773
rect 287425 337807 287483 337813
rect 287425 337773 287437 337807
rect 287471 337804 287483 337807
rect 301498 337804 301504 337816
rect 287471 337776 301504 337804
rect 287471 337773 287483 337776
rect 287425 337767 287483 337773
rect 301498 337764 301504 337776
rect 301556 337764 301562 337816
rect 262364 337708 275324 337736
rect 277397 337739 277455 337745
rect 262364 337696 262370 337708
rect 277397 337705 277409 337739
rect 277443 337736 277455 337739
rect 279602 337736 279608 337748
rect 277443 337708 279608 337736
rect 277443 337705 277455 337708
rect 277397 337699 277455 337705
rect 279602 337696 279608 337708
rect 279660 337696 279666 337748
rect 280157 337739 280215 337745
rect 280157 337705 280169 337739
rect 280203 337736 280215 337739
rect 282917 337739 282975 337745
rect 280203 337708 280936 337736
rect 280203 337705 280215 337708
rect 280157 337699 280215 337705
rect 35158 337628 35164 337680
rect 35216 337668 35222 337680
rect 232866 337668 232872 337680
rect 35216 337640 232872 337668
rect 35216 337628 35222 337640
rect 232866 337628 232872 337640
rect 232924 337628 232930 337680
rect 241517 337671 241575 337677
rect 241517 337637 241529 337671
rect 241563 337668 241575 337671
rect 246574 337668 246580 337680
rect 241563 337640 246580 337668
rect 241563 337637 241575 337640
rect 241517 337631 241575 337637
rect 246574 337628 246580 337640
rect 246632 337628 246638 337680
rect 257246 337628 257252 337680
rect 257304 337668 257310 337680
rect 263229 337671 263287 337677
rect 263229 337668 263241 337671
rect 257304 337640 263241 337668
rect 257304 337628 257310 337640
rect 263229 337637 263241 337640
rect 263275 337637 263287 337671
rect 263229 337631 263287 337637
rect 263505 337671 263563 337677
rect 263505 337637 263517 337671
rect 263551 337668 263563 337671
rect 275186 337668 275192 337680
rect 263551 337640 275192 337668
rect 263551 337637 263563 337640
rect 263505 337631 263563 337637
rect 275186 337628 275192 337640
rect 275244 337628 275250 337680
rect 275281 337671 275339 337677
rect 275281 337637 275293 337671
rect 275327 337668 275339 337671
rect 277857 337671 277915 337677
rect 277857 337668 277869 337671
rect 275327 337640 277869 337668
rect 275327 337637 275339 337640
rect 275281 337631 275339 337637
rect 277857 337637 277869 337640
rect 277903 337637 277915 337671
rect 277857 337631 277915 337637
rect 277949 337671 278007 337677
rect 277949 337637 277961 337671
rect 277995 337668 278007 337671
rect 280801 337671 280859 337677
rect 280801 337668 280813 337671
rect 277995 337640 280813 337668
rect 277995 337637 278007 337640
rect 277949 337631 278007 337637
rect 280801 337637 280813 337640
rect 280847 337637 280859 337671
rect 280908 337668 280936 337708
rect 282917 337705 282929 337739
rect 282963 337736 282975 337739
rect 287609 337739 287667 337745
rect 287609 337736 287621 337739
rect 282963 337708 287621 337736
rect 282963 337705 282975 337708
rect 282917 337699 282975 337705
rect 287609 337705 287621 337708
rect 287655 337705 287667 337739
rect 287609 337699 287667 337705
rect 287701 337739 287759 337745
rect 287701 337705 287713 337739
rect 287747 337736 287759 337739
rect 302878 337736 302884 337748
rect 287747 337708 302884 337736
rect 287747 337705 287759 337708
rect 287701 337699 287759 337705
rect 302878 337696 302884 337708
rect 302936 337696 302942 337748
rect 283558 337668 283564 337680
rect 280908 337640 283564 337668
rect 280801 337631 280859 337637
rect 283558 337628 283564 337640
rect 283616 337628 283622 337680
rect 286318 337628 286324 337680
rect 286376 337668 286382 337680
rect 286594 337668 286600 337680
rect 286376 337640 286600 337668
rect 286376 337628 286382 337640
rect 286594 337628 286600 337640
rect 286652 337628 286658 337680
rect 287422 337628 287428 337680
rect 287480 337668 287486 337680
rect 290826 337668 290832 337680
rect 287480 337640 290832 337668
rect 287480 337628 287486 337640
rect 290826 337628 290832 337640
rect 290884 337628 290890 337680
rect 290921 337671 290979 337677
rect 290921 337637 290933 337671
rect 290967 337668 290979 337671
rect 320818 337668 320824 337680
rect 290967 337640 320824 337668
rect 290967 337637 290979 337640
rect 290921 337631 290979 337637
rect 320818 337628 320824 337640
rect 320876 337628 320882 337680
rect 28258 337560 28264 337612
rect 28316 337600 28322 337612
rect 232038 337600 232044 337612
rect 28316 337572 232044 337600
rect 28316 337560 28322 337572
rect 232038 337560 232044 337572
rect 232096 337560 232102 337612
rect 258258 337560 258264 337612
rect 258316 337600 258322 337612
rect 262953 337603 263011 337609
rect 262953 337600 262965 337603
rect 258316 337572 262965 337600
rect 258316 337560 258322 337572
rect 262953 337569 262965 337572
rect 262999 337569 263011 337603
rect 262953 337563 263011 337569
rect 263781 337603 263839 337609
rect 263781 337569 263793 337603
rect 263827 337600 263839 337603
rect 277397 337603 277455 337609
rect 277397 337600 277409 337603
rect 263827 337572 277409 337600
rect 263827 337569 263839 337572
rect 263781 337563 263839 337569
rect 277397 337569 277409 337572
rect 277443 337569 277455 337603
rect 277397 337563 277455 337569
rect 277486 337560 277492 337612
rect 277544 337600 277550 337612
rect 278682 337600 278688 337612
rect 277544 337572 278688 337600
rect 277544 337560 277550 337572
rect 278682 337560 278688 337572
rect 278740 337560 278746 337612
rect 281166 337560 281172 337612
rect 281224 337600 281230 337612
rect 287517 337603 287575 337609
rect 287517 337600 287529 337603
rect 281224 337572 287529 337600
rect 281224 337560 281230 337572
rect 287517 337569 287529 337572
rect 287563 337569 287575 337603
rect 316678 337600 316684 337612
rect 287517 337563 287575 337569
rect 287624 337572 316684 337600
rect 15838 337492 15844 337544
rect 15896 337532 15902 337544
rect 231026 337532 231032 337544
rect 15896 337504 231032 337532
rect 15896 337492 15902 337504
rect 231026 337492 231032 337504
rect 231084 337492 231090 337544
rect 241146 337492 241152 337544
rect 241204 337532 241210 337544
rect 242986 337532 242992 337544
rect 241204 337504 242992 337532
rect 241204 337492 241210 337504
rect 242986 337492 242992 337504
rect 243044 337492 243050 337544
rect 260926 337492 260932 337544
rect 260984 337532 260990 337544
rect 270497 337535 270555 337541
rect 270497 337532 270509 337535
rect 260984 337504 270509 337532
rect 260984 337492 260990 337504
rect 270497 337501 270509 337504
rect 270543 337501 270555 337535
rect 270497 337495 270555 337501
rect 270681 337535 270739 337541
rect 270681 337501 270693 337535
rect 270727 337532 270739 337535
rect 271138 337532 271144 337544
rect 270727 337504 271144 337532
rect 270727 337501 270739 337504
rect 270681 337495 270739 337501
rect 271138 337492 271144 337504
rect 271196 337492 271202 337544
rect 277673 337535 277731 337541
rect 277673 337501 277685 337535
rect 277719 337532 277731 337535
rect 280706 337532 280712 337544
rect 277719 337504 280712 337532
rect 277719 337501 277731 337504
rect 277673 337495 277731 337501
rect 280706 337492 280712 337504
rect 280764 337492 280770 337544
rect 284021 337535 284079 337541
rect 284021 337501 284033 337535
rect 284067 337532 284079 337535
rect 287624 337532 287652 337572
rect 316678 337560 316684 337572
rect 316736 337560 316742 337612
rect 284067 337504 287652 337532
rect 287793 337535 287851 337541
rect 284067 337501 284079 337504
rect 284021 337495 284079 337501
rect 287793 337501 287805 337535
rect 287839 337532 287851 337535
rect 319438 337532 319444 337544
rect 287839 337504 319444 337532
rect 287839 337501 287851 337504
rect 287793 337495 287851 337501
rect 319438 337492 319444 337504
rect 319496 337492 319502 337544
rect 14458 337424 14464 337476
rect 14516 337464 14522 337476
rect 230934 337464 230940 337476
rect 14516 337436 230940 337464
rect 14516 337424 14522 337436
rect 230934 337424 230940 337436
rect 230992 337424 230998 337476
rect 242894 337424 242900 337476
rect 242952 337464 242958 337476
rect 253290 337464 253296 337476
rect 242952 337436 253296 337464
rect 242952 337424 242958 337436
rect 253290 337424 253296 337436
rect 253348 337424 253354 337476
rect 259638 337424 259644 337476
rect 259696 337464 259702 337476
rect 260837 337467 260895 337473
rect 260837 337464 260849 337467
rect 259696 337436 260849 337464
rect 259696 337424 259702 337436
rect 260837 337433 260849 337436
rect 260883 337433 260895 337467
rect 260837 337427 260895 337433
rect 265618 337424 265624 337476
rect 265676 337464 265682 337476
rect 275281 337467 275339 337473
rect 275281 337464 275293 337467
rect 265676 337436 275293 337464
rect 265676 337424 265682 337436
rect 275281 337433 275293 337436
rect 275327 337433 275339 337467
rect 275281 337427 275339 337433
rect 277857 337467 277915 337473
rect 277857 337433 277869 337467
rect 277903 337464 277915 337467
rect 346394 337464 346400 337476
rect 277903 337436 346400 337464
rect 277903 337433 277915 337436
rect 277857 337427 277915 337433
rect 346394 337424 346400 337436
rect 346452 337424 346458 337476
rect 10318 337356 10324 337408
rect 10376 337396 10382 337408
rect 230474 337396 230480 337408
rect 10376 337368 230480 337396
rect 10376 337356 10382 337368
rect 230474 337356 230480 337368
rect 230532 337356 230538 337408
rect 234985 337399 235043 337405
rect 234985 337365 234997 337399
rect 235031 337396 235043 337399
rect 241517 337399 241575 337405
rect 241517 337396 241529 337399
rect 235031 337368 241529 337396
rect 235031 337365 235043 337368
rect 234985 337359 235043 337365
rect 241517 337365 241529 337368
rect 241563 337365 241575 337399
rect 241517 337359 241575 337365
rect 245562 337356 245568 337408
rect 245620 337396 245626 337408
rect 251266 337396 251272 337408
rect 245620 337368 251272 337396
rect 245620 337356 245626 337368
rect 251266 337356 251272 337368
rect 251324 337356 251330 337408
rect 260190 337356 260196 337408
rect 260248 337396 260254 337408
rect 263137 337399 263195 337405
rect 263137 337396 263149 337399
rect 260248 337368 263149 337396
rect 260248 337356 260254 337368
rect 263137 337365 263149 337368
rect 263183 337365 263195 337399
rect 277581 337399 277639 337405
rect 277581 337396 277593 337399
rect 263137 337359 263195 337365
rect 263704 337368 277593 337396
rect 232041 337331 232099 337337
rect 232041 337297 232053 337331
rect 232087 337328 232099 337331
rect 241793 337331 241851 337337
rect 241793 337328 241805 337331
rect 232087 337300 241805 337328
rect 232087 337297 232099 337300
rect 232041 337291 232099 337297
rect 241793 337297 241805 337300
rect 241839 337297 241851 337331
rect 241793 337291 241851 337297
rect 260558 337288 260564 337340
rect 260616 337328 260622 337340
rect 260616 337300 262260 337328
rect 260616 337288 260622 337300
rect 225690 337220 225696 337272
rect 225748 337260 225754 337272
rect 235997 337263 236055 337269
rect 235997 337260 236009 337263
rect 225748 337232 236009 337260
rect 225748 337220 225754 337232
rect 235997 337229 236009 337232
rect 236043 337229 236055 337263
rect 235997 337223 236055 337229
rect 257430 337220 257436 337272
rect 257488 337260 257494 337272
rect 261205 337263 261263 337269
rect 261205 337260 261217 337263
rect 257488 337232 261217 337260
rect 257488 337220 257494 337232
rect 261205 337229 261217 337232
rect 261251 337229 261263 337263
rect 261205 337223 261263 337229
rect 261478 337220 261484 337272
rect 261536 337260 261542 337272
rect 261662 337260 261668 337272
rect 261536 337232 261668 337260
rect 261536 337220 261542 337232
rect 261662 337220 261668 337232
rect 261720 337220 261726 337272
rect 228358 337152 228364 337204
rect 228416 337192 228422 337204
rect 228416 337164 239444 337192
rect 228416 337152 228422 337164
rect 231946 337084 231952 337136
rect 232004 337124 232010 337136
rect 234890 337124 234896 337136
rect 232004 337096 234896 337124
rect 232004 337084 232010 337096
rect 234890 337084 234896 337096
rect 234948 337084 234954 337136
rect 239416 337124 239444 337164
rect 251266 337152 251272 337204
rect 251324 337192 251330 337204
rect 254854 337192 254860 337204
rect 251324 337164 254860 337192
rect 251324 337152 251330 337164
rect 254854 337152 254860 337164
rect 254912 337152 254918 337204
rect 260466 337152 260472 337204
rect 260524 337192 260530 337204
rect 260653 337195 260711 337201
rect 260653 337192 260665 337195
rect 260524 337164 260665 337192
rect 260524 337152 260530 337164
rect 260653 337161 260665 337164
rect 260699 337161 260711 337195
rect 260653 337155 260711 337161
rect 262122 337152 262128 337204
rect 262180 337152 262186 337204
rect 246758 337124 246764 337136
rect 239416 337096 246764 337124
rect 246758 337084 246764 337096
rect 246816 337084 246822 337136
rect 256694 337084 256700 337136
rect 256752 337124 256758 337136
rect 258442 337124 258448 337136
rect 256752 337096 258448 337124
rect 256752 337084 256758 337096
rect 258442 337084 258448 337096
rect 258500 337084 258506 337136
rect 258626 337084 258632 337136
rect 258684 337124 258690 337136
rect 260926 337124 260932 337136
rect 258684 337096 260932 337124
rect 258684 337084 258690 337096
rect 260926 337084 260932 337096
rect 260984 337084 260990 337136
rect 261294 337084 261300 337136
rect 261352 337124 261358 337136
rect 261662 337124 261668 337136
rect 261352 337096 261668 337124
rect 261352 337084 261358 337096
rect 261662 337084 261668 337096
rect 261720 337084 261726 337136
rect 230569 337059 230627 337065
rect 230569 337025 230581 337059
rect 230615 337056 230627 337059
rect 232041 337059 232099 337065
rect 232041 337056 232053 337059
rect 230615 337028 232053 337056
rect 230615 337025 230627 337028
rect 230569 337019 230627 337025
rect 232041 337025 232053 337028
rect 232087 337025 232099 337059
rect 232041 337019 232099 337025
rect 247678 337016 247684 337068
rect 247736 337056 247742 337068
rect 255038 337056 255044 337068
rect 247736 337028 255044 337056
rect 247736 337016 247742 337028
rect 255038 337016 255044 337028
rect 255096 337016 255102 337068
rect 256878 337016 256884 337068
rect 256936 337056 256942 337068
rect 258074 337056 258080 337068
rect 256936 337028 258080 337056
rect 256936 337016 256942 337028
rect 258074 337016 258080 337028
rect 258132 337016 258138 337068
rect 260098 337016 260104 337068
rect 260156 337056 260162 337068
rect 260558 337056 260564 337068
rect 260156 337028 260564 337056
rect 260156 337016 260162 337028
rect 260558 337016 260564 337028
rect 260616 337016 260622 337068
rect 260834 337016 260840 337068
rect 260892 337056 260898 337068
rect 261846 337056 261852 337068
rect 260892 337028 261852 337056
rect 260892 337016 260898 337028
rect 261846 337016 261852 337028
rect 261904 337016 261910 337068
rect 230382 336948 230388 337000
rect 230440 336988 230446 337000
rect 236822 336988 236828 337000
rect 230440 336960 236828 336988
rect 230440 336948 230446 336960
rect 236822 336948 236828 336960
rect 236880 336948 236886 337000
rect 248506 336948 248512 337000
rect 248564 336988 248570 337000
rect 251358 336988 251364 337000
rect 248564 336960 251364 336988
rect 248564 336948 248570 336960
rect 251358 336948 251364 336960
rect 251416 336948 251422 337000
rect 251729 336991 251787 336997
rect 251729 336957 251741 336991
rect 251775 336988 251787 336991
rect 253566 336988 253572 337000
rect 251775 336960 253572 336988
rect 251775 336957 251787 336960
rect 251729 336951 251787 336957
rect 253566 336948 253572 336960
rect 253624 336948 253630 337000
rect 257062 336948 257068 337000
rect 257120 336988 257126 337000
rect 257798 336988 257804 337000
rect 257120 336960 257804 336988
rect 257120 336948 257126 336960
rect 257798 336948 257804 336960
rect 257856 336948 257862 337000
rect 258350 336948 258356 337000
rect 258408 336988 258414 337000
rect 259178 336988 259184 337000
rect 258408 336960 259184 336988
rect 258408 336948 258414 336960
rect 259178 336948 259184 336960
rect 259236 336948 259242 337000
rect 261018 336948 261024 337000
rect 261076 336988 261082 337000
rect 261938 336988 261944 337000
rect 261076 336960 261944 336988
rect 261076 336948 261082 336960
rect 261938 336948 261944 336960
rect 261996 336948 262002 337000
rect 233234 336880 233240 336932
rect 233292 336920 233298 336932
rect 234430 336920 234436 336932
rect 233292 336892 234436 336920
rect 233292 336880 233298 336892
rect 234430 336880 234436 336892
rect 234488 336880 234494 336932
rect 249610 336880 249616 336932
rect 249668 336920 249674 336932
rect 252830 336920 252836 336932
rect 249668 336892 252836 336920
rect 249668 336880 249674 336892
rect 252830 336880 252836 336892
rect 252888 336880 252894 336932
rect 257154 336880 257160 336932
rect 257212 336920 257218 336932
rect 257890 336920 257896 336932
rect 257212 336892 257896 336920
rect 257212 336880 257218 336892
rect 257890 336880 257896 336892
rect 257948 336880 257954 336932
rect 258258 336880 258264 336932
rect 258316 336920 258322 336932
rect 259270 336920 259276 336932
rect 258316 336892 259276 336920
rect 258316 336880 258322 336892
rect 259270 336880 259276 336892
rect 259328 336880 259334 336932
rect 259822 336880 259828 336932
rect 259880 336920 259886 336932
rect 260650 336920 260656 336932
rect 259880 336892 260656 336920
rect 259880 336880 259886 336892
rect 260650 336880 260656 336892
rect 260708 336880 260714 336932
rect 261202 336880 261208 336932
rect 261260 336920 261266 336932
rect 262030 336920 262036 336932
rect 261260 336892 262036 336920
rect 261260 336880 261266 336892
rect 262030 336880 262036 336892
rect 262088 336880 262094 336932
rect 252278 336812 252284 336864
rect 252336 336852 252342 336864
rect 253750 336852 253756 336864
rect 252336 336824 253756 336852
rect 252336 336812 252342 336824
rect 253750 336812 253756 336824
rect 253808 336812 253814 336864
rect 254854 336812 254860 336864
rect 254912 336852 254918 336864
rect 255774 336852 255780 336864
rect 254912 336824 255780 336852
rect 254912 336812 254918 336824
rect 255774 336812 255780 336824
rect 255832 336812 255838 336864
rect 257062 336812 257068 336864
rect 257120 336852 257126 336864
rect 257614 336852 257620 336864
rect 257120 336824 257620 336852
rect 257120 336812 257126 336824
rect 257614 336812 257620 336824
rect 257672 336812 257678 336864
rect 258350 336812 258356 336864
rect 258408 336852 258414 336864
rect 259086 336852 259092 336864
rect 258408 336824 259092 336852
rect 258408 336812 258414 336824
rect 259086 336812 259092 336824
rect 259144 336812 259150 336864
rect 260834 336812 260840 336864
rect 260892 336852 260898 336864
rect 261570 336852 261576 336864
rect 260892 336824 261576 336852
rect 260892 336812 260898 336824
rect 261570 336812 261576 336824
rect 261628 336812 261634 336864
rect 261938 336812 261944 336864
rect 261996 336852 262002 336864
rect 262140 336852 262168 337152
rect 262232 337124 262260 337300
rect 263597 337127 263655 337133
rect 263597 337124 263609 337127
rect 262232 337096 263609 337124
rect 263597 337093 263609 337096
rect 263643 337093 263655 337127
rect 263597 337087 263655 337093
rect 262766 337016 262772 337068
rect 262824 337056 262830 337068
rect 262950 337056 262956 337068
rect 262824 337028 262956 337056
rect 262824 337016 262830 337028
rect 262950 337016 262956 337028
rect 263008 337016 263014 337068
rect 262398 336948 262404 337000
rect 262456 336988 262462 337000
rect 263042 336988 263048 337000
rect 262456 336960 263048 336988
rect 262456 336948 262462 336960
rect 263042 336948 263048 336960
rect 263100 336948 263106 337000
rect 263137 336991 263195 336997
rect 263137 336957 263149 336991
rect 263183 336988 263195 336991
rect 263704 336988 263732 337368
rect 277581 337365 277593 337368
rect 277627 337365 277639 337399
rect 277581 337359 277639 337365
rect 277762 337356 277768 337408
rect 277820 337396 277826 337408
rect 278314 337396 278320 337408
rect 277820 337368 278320 337396
rect 277820 337356 277826 337368
rect 278314 337356 278320 337368
rect 278372 337356 278378 337408
rect 281902 337356 281908 337408
rect 281960 337396 281966 337408
rect 287425 337399 287483 337405
rect 287425 337396 287437 337399
rect 281960 337368 287437 337396
rect 281960 337356 281966 337368
rect 287425 337365 287437 337368
rect 287471 337365 287483 337399
rect 287425 337359 287483 337365
rect 287517 337399 287575 337405
rect 287517 337365 287529 337399
rect 287563 337396 287575 337399
rect 489178 337396 489184 337408
rect 287563 337368 489184 337396
rect 287563 337365 287575 337368
rect 287517 337359 287575 337365
rect 489178 337356 489184 337368
rect 489236 337356 489242 337408
rect 263962 337288 263968 337340
rect 264020 337328 264026 337340
rect 271322 337328 271328 337340
rect 264020 337300 271328 337328
rect 264020 337288 264026 337300
rect 271322 337288 271328 337300
rect 271380 337288 271386 337340
rect 273438 337288 273444 337340
rect 273496 337328 273502 337340
rect 274542 337328 274548 337340
rect 273496 337300 274548 337328
rect 273496 337288 273502 337300
rect 274542 337288 274548 337300
rect 274600 337288 274606 337340
rect 274637 337331 274695 337337
rect 274637 337297 274649 337331
rect 274683 337328 274695 337331
rect 277673 337331 277731 337337
rect 277673 337328 277685 337331
rect 274683 337300 277685 337328
rect 274683 337297 274695 337300
rect 274637 337291 274695 337297
rect 277673 337297 277685 337300
rect 277719 337297 277731 337331
rect 277673 337291 277731 337297
rect 277854 337288 277860 337340
rect 277912 337328 277918 337340
rect 278590 337328 278596 337340
rect 277912 337300 278596 337328
rect 277912 337288 277918 337300
rect 278590 337288 278596 337300
rect 278648 337288 278654 337340
rect 280157 337331 280215 337337
rect 280157 337328 280169 337331
rect 278700 337300 280169 337328
rect 265250 337220 265256 337272
rect 265308 337260 265314 337272
rect 266081 337263 266139 337269
rect 266081 337260 266093 337263
rect 265308 337232 266093 337260
rect 265308 337220 265314 337232
rect 266081 337229 266093 337232
rect 266127 337229 266139 337263
rect 266081 337223 266139 337229
rect 271230 337220 271236 337272
rect 271288 337260 271294 337272
rect 277489 337263 277547 337269
rect 277489 337260 277501 337263
rect 271288 337232 277501 337260
rect 271288 337220 271294 337232
rect 277489 337229 277501 337232
rect 277535 337229 277547 337263
rect 277489 337223 277547 337229
rect 278133 337263 278191 337269
rect 278133 337229 278145 337263
rect 278179 337260 278191 337263
rect 278700 337260 278728 337300
rect 280157 337297 280169 337300
rect 280203 337297 280215 337331
rect 280157 337291 280215 337297
rect 282917 337331 282975 337337
rect 282917 337297 282929 337331
rect 282963 337297 282975 337331
rect 282917 337291 282975 337297
rect 283101 337331 283159 337337
rect 283101 337297 283113 337331
rect 283147 337328 283159 337331
rect 289906 337328 289912 337340
rect 283147 337300 289912 337328
rect 283147 337297 283159 337300
rect 283101 337291 283159 337297
rect 278179 337232 278728 337260
rect 278179 337229 278191 337232
rect 278133 337223 278191 337229
rect 278774 337220 278780 337272
rect 278832 337260 278838 337272
rect 278961 337263 279019 337269
rect 278961 337260 278973 337263
rect 278832 337232 278973 337260
rect 278832 337220 278838 337232
rect 278961 337229 278973 337232
rect 279007 337229 279019 337263
rect 278961 337223 279019 337229
rect 280062 337220 280068 337272
rect 280120 337260 280126 337272
rect 281445 337263 281503 337269
rect 281445 337260 281457 337263
rect 280120 337232 281457 337260
rect 280120 337220 280126 337232
rect 281445 337229 281457 337232
rect 281491 337229 281503 337263
rect 281445 337223 281503 337229
rect 282270 337220 282276 337272
rect 282328 337260 282334 337272
rect 282932 337260 282960 337291
rect 289906 337288 289912 337300
rect 289964 337288 289970 337340
rect 282328 337232 282960 337260
rect 282328 337220 282334 337232
rect 283006 337220 283012 337272
rect 283064 337260 283070 337272
rect 284202 337260 284208 337272
rect 283064 337232 284208 337260
rect 283064 337220 283070 337232
rect 284202 337220 284208 337232
rect 284260 337220 284266 337272
rect 284294 337220 284300 337272
rect 284352 337260 284358 337272
rect 291013 337263 291071 337269
rect 291013 337260 291025 337263
rect 284352 337232 291025 337260
rect 284352 337220 284358 337232
rect 291013 337229 291025 337232
rect 291059 337229 291071 337263
rect 291013 337223 291071 337229
rect 271049 337195 271107 337201
rect 271049 337192 271061 337195
rect 263183 336960 263732 336988
rect 263796 337164 271061 337192
rect 263183 336957 263195 336960
rect 263137 336951 263195 336957
rect 262766 336880 262772 336932
rect 262824 336920 262830 336932
rect 263502 336920 263508 336932
rect 262824 336892 263508 336920
rect 262824 336880 262830 336892
rect 263502 336880 263508 336892
rect 263560 336880 263566 336932
rect 263689 336923 263747 336929
rect 263689 336889 263701 336923
rect 263735 336920 263747 336923
rect 263796 336920 263824 337164
rect 271049 337161 271061 337164
rect 271095 337161 271107 337195
rect 271049 337155 271107 337161
rect 272518 337152 272524 337204
rect 272576 337192 272582 337204
rect 273070 337192 273076 337204
rect 272576 337164 273076 337192
rect 272576 337152 272582 337164
rect 273070 337152 273076 337164
rect 273128 337152 273134 337204
rect 276293 337195 276351 337201
rect 276293 337161 276305 337195
rect 276339 337192 276351 337195
rect 282457 337195 282515 337201
rect 282457 337192 282469 337195
rect 276339 337164 282469 337192
rect 276339 337161 276351 337164
rect 276293 337155 276351 337161
rect 282457 337161 282469 337164
rect 282503 337161 282515 337195
rect 282457 337155 282515 337161
rect 282546 337152 282552 337204
rect 282604 337192 282610 337204
rect 282822 337192 282828 337204
rect 282604 337164 282828 337192
rect 282604 337152 282610 337164
rect 282822 337152 282828 337164
rect 282880 337152 282886 337204
rect 282914 337152 282920 337204
rect 282972 337192 282978 337204
rect 283466 337192 283472 337204
rect 282972 337164 283472 337192
rect 282972 337152 282978 337164
rect 283466 337152 283472 337164
rect 283524 337152 283530 337204
rect 286042 337152 286048 337204
rect 286100 337192 286106 337204
rect 286962 337192 286968 337204
rect 286100 337164 286968 337192
rect 286100 337152 286106 337164
rect 286962 337152 286968 337164
rect 287020 337152 287026 337204
rect 287422 337152 287428 337204
rect 287480 337192 287486 337204
rect 288342 337192 288348 337204
rect 287480 337164 288348 337192
rect 287480 337152 287486 337164
rect 288342 337152 288348 337164
rect 288400 337152 288406 337204
rect 264974 337084 264980 337136
rect 265032 337124 265038 337136
rect 265894 337124 265900 337136
rect 265032 337096 265900 337124
rect 265032 337084 265038 337096
rect 265894 337084 265900 337096
rect 265952 337084 265958 337136
rect 270494 337084 270500 337136
rect 270552 337124 270558 337136
rect 274637 337127 274695 337133
rect 274637 337124 274649 337127
rect 270552 337096 274649 337124
rect 270552 337084 270558 337096
rect 274637 337093 274649 337096
rect 274683 337093 274695 337127
rect 274818 337124 274824 337136
rect 274779 337096 274824 337124
rect 274637 337087 274695 337093
rect 274818 337084 274824 337096
rect 274876 337084 274882 337136
rect 279234 337084 279240 337136
rect 279292 337124 279298 337136
rect 279878 337124 279884 337136
rect 279292 337096 279884 337124
rect 279292 337084 279298 337096
rect 279878 337084 279884 337096
rect 279936 337084 279942 337136
rect 280798 337084 280804 337136
rect 280856 337124 280862 337136
rect 287701 337127 287759 337133
rect 287701 337124 287713 337127
rect 280856 337096 287713 337124
rect 280856 337084 280862 337096
rect 287701 337093 287713 337096
rect 287747 337093 287759 337127
rect 287701 337087 287759 337093
rect 287885 337127 287943 337133
rect 287885 337093 287897 337127
rect 287931 337124 287943 337127
rect 291838 337124 291844 337136
rect 287931 337096 291844 337124
rect 287931 337093 287943 337096
rect 287885 337087 287943 337093
rect 291838 337084 291844 337096
rect 291896 337084 291902 337136
rect 265158 337016 265164 337068
rect 265216 337056 265222 337068
rect 265986 337056 265992 337068
rect 265216 337028 265992 337056
rect 265216 337016 265222 337028
rect 265986 337016 265992 337028
rect 266044 337016 266050 337068
rect 266722 337016 266728 337068
rect 266780 337056 266786 337068
rect 266780 337028 267780 337056
rect 266780 337016 266786 337028
rect 264974 336988 264980 337000
rect 263735 336892 263824 336920
rect 263888 336960 264980 336988
rect 263735 336889 263747 336892
rect 263689 336883 263747 336889
rect 261996 336824 262168 336852
rect 261996 336812 262002 336824
rect 262674 336812 262680 336864
rect 262732 336852 262738 336864
rect 263134 336852 263140 336864
rect 262732 336824 263140 336852
rect 262732 336812 262738 336824
rect 263134 336812 263140 336824
rect 263192 336812 263198 336864
rect 263229 336855 263287 336861
rect 263229 336821 263241 336855
rect 263275 336852 263287 336855
rect 263888 336852 263916 336960
rect 264974 336948 264980 336960
rect 265032 336948 265038 337000
rect 265250 336948 265256 337000
rect 265308 336988 265314 337000
rect 266078 336988 266084 337000
rect 265308 336960 266084 336988
rect 265308 336948 265314 336960
rect 266078 336948 266084 336960
rect 266136 336948 266142 337000
rect 266354 336948 266360 337000
rect 266412 336988 266418 337000
rect 267642 336988 267648 337000
rect 266412 336960 267648 336988
rect 266412 336948 266418 336960
rect 267642 336948 267648 336960
rect 267700 336948 267706 337000
rect 265434 336880 265440 336932
rect 265492 336920 265498 336932
rect 266262 336920 266268 336932
rect 265492 336892 266268 336920
rect 265492 336880 265498 336892
rect 266262 336880 266268 336892
rect 266320 336880 266326 336932
rect 266722 336880 266728 336932
rect 266780 336920 266786 336932
rect 267182 336920 267188 336932
rect 266780 336892 267188 336920
rect 266780 336880 266786 336892
rect 267182 336880 267188 336892
rect 267240 336880 267246 336932
rect 267752 336920 267780 337028
rect 272334 337016 272340 337068
rect 272392 337056 272398 337068
rect 273070 337056 273076 337068
rect 272392 337028 273076 337056
rect 272392 337016 272398 337028
rect 273070 337016 273076 337028
rect 273128 337016 273134 337068
rect 273346 337016 273352 337068
rect 273404 337056 273410 337068
rect 274358 337056 274364 337068
rect 273404 337028 274364 337056
rect 273404 337016 273410 337028
rect 274358 337016 274364 337028
rect 274416 337016 274422 337068
rect 274726 337016 274732 337068
rect 274784 337056 274790 337068
rect 275646 337056 275652 337068
rect 274784 337028 275652 337056
rect 274784 337016 274790 337028
rect 275646 337016 275652 337028
rect 275704 337016 275710 337068
rect 278130 337016 278136 337068
rect 278188 337016 278194 337068
rect 278222 337016 278228 337068
rect 278280 337056 278286 337068
rect 278774 337056 278780 337068
rect 278280 337028 278780 337056
rect 278280 337016 278286 337028
rect 278774 337016 278780 337028
rect 278832 337016 278838 337068
rect 279142 337016 279148 337068
rect 279200 337056 279206 337068
rect 280062 337056 280068 337068
rect 279200 337028 280068 337056
rect 279200 337016 279206 337028
rect 280062 337016 280068 337028
rect 280120 337016 280126 337068
rect 280430 337016 280436 337068
rect 280488 337056 280494 337068
rect 282733 337059 282791 337065
rect 282733 337056 282745 337059
rect 280488 337028 282745 337056
rect 280488 337016 280494 337028
rect 282733 337025 282745 337028
rect 282779 337025 282791 337059
rect 282733 337019 282791 337025
rect 282825 337059 282883 337065
rect 282825 337025 282837 337059
rect 282871 337056 282883 337059
rect 283466 337056 283472 337068
rect 282871 337028 283472 337056
rect 282871 337025 282883 337028
rect 282825 337019 282883 337025
rect 283466 337016 283472 337028
rect 283524 337016 283530 337068
rect 283742 337016 283748 337068
rect 283800 337056 283806 337068
rect 284018 337056 284024 337068
rect 283800 337028 284024 337056
rect 283800 337016 283806 337028
rect 284018 337016 284024 337028
rect 284076 337016 284082 337068
rect 287793 337059 287851 337065
rect 287793 337056 287805 337059
rect 284220 337028 287805 337056
rect 267918 336948 267924 337000
rect 267976 336988 267982 337000
rect 268654 336988 268660 337000
rect 267976 336960 268660 336988
rect 267976 336948 267982 336960
rect 268654 336948 268660 336960
rect 268712 336948 268718 337000
rect 273438 336948 273444 337000
rect 273496 336988 273502 337000
rect 274450 336988 274456 337000
rect 273496 336960 274456 336988
rect 273496 336948 273502 336960
rect 274450 336948 274456 336960
rect 274508 336948 274514 337000
rect 276106 336948 276112 337000
rect 276164 336988 276170 337000
rect 277026 336988 277032 337000
rect 276164 336960 277032 336988
rect 276164 336948 276170 336960
rect 277026 336948 277032 336960
rect 277084 336948 277090 337000
rect 278148 336988 278176 337016
rect 278590 336988 278596 337000
rect 278148 336960 278596 336988
rect 278590 336948 278596 336960
rect 278648 336948 278654 337000
rect 279050 336948 279056 337000
rect 279108 336988 279114 337000
rect 279694 336988 279700 337000
rect 279108 336960 279700 336988
rect 279108 336948 279114 336960
rect 279694 336948 279700 336960
rect 279752 336948 279758 337000
rect 280338 336948 280344 337000
rect 280396 336988 280402 337000
rect 280890 336988 280896 337000
rect 280396 336960 280896 336988
rect 280396 336948 280402 336960
rect 280890 336948 280896 336960
rect 280948 336948 280954 337000
rect 281534 336948 281540 337000
rect 281592 336988 281598 337000
rect 283009 336991 283067 336997
rect 283009 336988 283021 336991
rect 281592 336960 283021 336988
rect 281592 336948 281598 336960
rect 283009 336957 283021 336960
rect 283055 336957 283067 336991
rect 283009 336951 283067 336957
rect 283190 336948 283196 337000
rect 283248 336988 283254 337000
rect 284110 336988 284116 337000
rect 283248 336960 284116 336988
rect 283248 336948 283254 336960
rect 284110 336948 284116 336960
rect 284168 336948 284174 337000
rect 267660 336892 267780 336920
rect 267660 336864 267688 336892
rect 268286 336880 268292 336932
rect 268344 336920 268350 336932
rect 268838 336920 268844 336932
rect 268344 336892 268844 336920
rect 268344 336880 268350 336892
rect 268838 336880 268844 336892
rect 268896 336880 268902 336932
rect 270586 336880 270592 336932
rect 270644 336920 270650 336932
rect 271230 336920 271236 336932
rect 270644 336892 271236 336920
rect 270644 336880 270650 336892
rect 271230 336880 271236 336892
rect 271288 336880 271294 336932
rect 272334 336880 272340 336932
rect 272392 336920 272398 336932
rect 272702 336920 272708 336932
rect 272392 336892 272708 336920
rect 272392 336880 272398 336892
rect 272702 336880 272708 336892
rect 272760 336880 272766 336932
rect 273254 336880 273260 336932
rect 273312 336920 273318 336932
rect 274082 336920 274088 336932
rect 273312 336892 274088 336920
rect 273312 336880 273318 336892
rect 274082 336880 274088 336892
rect 274140 336880 274146 336932
rect 274818 336880 274824 336932
rect 274876 336920 274882 336932
rect 275370 336920 275376 336932
rect 274876 336892 275376 336920
rect 274876 336880 274882 336892
rect 275370 336880 275376 336892
rect 275428 336880 275434 336932
rect 276385 336923 276443 336929
rect 276385 336889 276397 336923
rect 276431 336920 276443 336923
rect 276934 336920 276940 336932
rect 276431 336892 276940 336920
rect 276431 336889 276443 336892
rect 276385 336883 276443 336889
rect 276934 336880 276940 336892
rect 276992 336880 276998 336932
rect 279326 336880 279332 336932
rect 279384 336920 279390 336932
rect 279878 336920 279884 336932
rect 279384 336892 279884 336920
rect 279384 336880 279390 336892
rect 279878 336880 279884 336892
rect 279936 336880 279942 336932
rect 280614 336880 280620 336932
rect 280672 336920 280678 336932
rect 281166 336920 281172 336932
rect 280672 336892 281172 336920
rect 280672 336880 280678 336892
rect 281166 336880 281172 336892
rect 281224 336880 281230 336932
rect 281445 336923 281503 336929
rect 281445 336889 281457 336923
rect 281491 336920 281503 336923
rect 284021 336923 284079 336929
rect 284021 336920 284033 336923
rect 281491 336892 284033 336920
rect 281491 336889 281503 336892
rect 281445 336883 281503 336889
rect 284021 336889 284033 336892
rect 284067 336889 284079 336923
rect 284021 336883 284079 336889
rect 263275 336824 263916 336852
rect 263275 336821 263287 336824
rect 263229 336815 263287 336821
rect 263962 336812 263968 336864
rect 264020 336852 264026 336864
rect 264882 336852 264888 336864
rect 264020 336824 264888 336852
rect 264020 336812 264026 336824
rect 264882 336812 264888 336824
rect 264940 336812 264946 336864
rect 265618 336812 265624 336864
rect 265676 336852 265682 336864
rect 266170 336852 266176 336864
rect 265676 336824 266176 336852
rect 265676 336812 265682 336824
rect 266170 336812 266176 336824
rect 266228 336812 266234 336864
rect 266906 336812 266912 336864
rect 266964 336852 266970 336864
rect 267366 336852 267372 336864
rect 266964 336824 267372 336852
rect 266964 336812 266970 336824
rect 267366 336812 267372 336824
rect 267424 336812 267430 336864
rect 267642 336812 267648 336864
rect 267700 336812 267706 336864
rect 271874 336812 271880 336864
rect 271932 336852 271938 336864
rect 272150 336852 272156 336864
rect 271932 336824 272156 336852
rect 271932 336812 271938 336824
rect 272150 336812 272156 336824
rect 272208 336812 272214 336864
rect 273346 336812 273352 336864
rect 273404 336852 273410 336864
rect 273806 336852 273812 336864
rect 273404 336824 273812 336852
rect 273404 336812 273410 336824
rect 273806 336812 273812 336824
rect 273864 336812 273870 336864
rect 274910 336812 274916 336864
rect 274968 336852 274974 336864
rect 275462 336852 275468 336864
rect 274968 336824 275468 336852
rect 274968 336812 274974 336824
rect 275462 336812 275468 336824
rect 275520 336812 275526 336864
rect 276014 336812 276020 336864
rect 276072 336852 276078 336864
rect 276474 336852 276480 336864
rect 276072 336824 276480 336852
rect 276072 336812 276078 336824
rect 276474 336812 276480 336824
rect 276532 336812 276538 336864
rect 277302 336852 277308 336864
rect 276768 336824 277308 336852
rect 233234 336744 233240 336796
rect 233292 336784 233298 336796
rect 235258 336784 235264 336796
rect 233292 336756 235264 336784
rect 233292 336744 233298 336756
rect 235258 336744 235264 336756
rect 235316 336744 235322 336796
rect 240226 336744 240232 336796
rect 240284 336784 240290 336796
rect 241606 336784 241612 336796
rect 240284 336756 241612 336784
rect 240284 336744 240290 336756
rect 241606 336744 241612 336756
rect 241664 336744 241670 336796
rect 245286 336744 245292 336796
rect 245344 336784 245350 336796
rect 245838 336784 245844 336796
rect 245344 336756 245844 336784
rect 245344 336744 245350 336756
rect 245838 336744 245844 336756
rect 245896 336744 245902 336796
rect 247034 336744 247040 336796
rect 247092 336784 247098 336796
rect 248414 336784 248420 336796
rect 247092 336756 248420 336784
rect 247092 336744 247098 336756
rect 248414 336744 248420 336756
rect 248472 336744 248478 336796
rect 251910 336744 251916 336796
rect 251968 336784 251974 336796
rect 253474 336784 253480 336796
rect 251968 336756 253480 336784
rect 251968 336744 251974 336756
rect 253474 336744 253480 336756
rect 253532 336744 253538 336796
rect 254762 336744 254768 336796
rect 254820 336784 254826 336796
rect 255406 336784 255412 336796
rect 254820 336756 255412 336784
rect 254820 336744 254826 336756
rect 255406 336744 255412 336756
rect 255464 336744 255470 336796
rect 256510 336744 256516 336796
rect 256568 336784 256574 336796
rect 257338 336784 257344 336796
rect 256568 336756 257344 336784
rect 256568 336744 256574 336756
rect 257338 336744 257344 336756
rect 257396 336744 257402 336796
rect 257522 336744 257528 336796
rect 257580 336784 257586 336796
rect 257982 336784 257988 336796
rect 257580 336756 257988 336784
rect 257580 336744 257586 336756
rect 257982 336744 257988 336756
rect 258040 336744 258046 336796
rect 258534 336744 258540 336796
rect 258592 336784 258598 336796
rect 258902 336784 258908 336796
rect 258592 336756 258908 336784
rect 258592 336744 258598 336756
rect 258902 336744 258908 336756
rect 258960 336744 258966 336796
rect 260006 336744 260012 336796
rect 260064 336784 260070 336796
rect 260466 336784 260472 336796
rect 260064 336756 260472 336784
rect 260064 336744 260070 336756
rect 260466 336744 260472 336756
rect 260524 336744 260530 336796
rect 260650 336784 260656 336796
rect 260611 336756 260656 336784
rect 260650 336744 260656 336756
rect 260708 336744 260714 336796
rect 260926 336744 260932 336796
rect 260984 336784 260990 336796
rect 260984 336756 261248 336784
rect 260984 336744 260990 336756
rect 261220 336716 261248 336756
rect 261294 336744 261300 336796
rect 261352 336784 261358 336796
rect 261754 336784 261760 336796
rect 261352 336756 261760 336784
rect 261352 336744 261358 336756
rect 261754 336744 261760 336756
rect 261812 336744 261818 336796
rect 262214 336744 262220 336796
rect 262272 336784 262278 336796
rect 262272 336756 262444 336784
rect 262272 336744 262278 336756
rect 261570 336716 261576 336728
rect 261220 336688 261576 336716
rect 261570 336676 261576 336688
rect 261628 336676 261634 336728
rect 261202 336648 261208 336660
rect 261163 336620 261208 336648
rect 261202 336608 261208 336620
rect 261260 336608 261266 336660
rect 262416 336648 262444 336756
rect 262490 336744 262496 336796
rect 262548 336784 262554 336796
rect 262858 336784 262864 336796
rect 262548 336756 262864 336784
rect 262548 336744 262554 336756
rect 262858 336744 262864 336756
rect 262916 336744 262922 336796
rect 262953 336787 263011 336793
rect 262953 336753 262965 336787
rect 262999 336784 263011 336787
rect 263689 336787 263747 336793
rect 263689 336784 263701 336787
rect 262999 336756 263701 336784
rect 262999 336753 263011 336756
rect 262953 336747 263011 336753
rect 263689 336753 263701 336756
rect 263735 336753 263747 336787
rect 263689 336747 263747 336753
rect 263778 336744 263784 336796
rect 263836 336784 263842 336796
rect 264146 336784 264152 336796
rect 263836 336756 264152 336784
rect 263836 336744 263842 336756
rect 264146 336744 264152 336756
rect 264204 336744 264210 336796
rect 264330 336744 264336 336796
rect 264388 336784 264394 336796
rect 264606 336784 264612 336796
rect 264388 336756 264612 336784
rect 264388 336744 264394 336756
rect 264606 336744 264612 336756
rect 264664 336744 264670 336796
rect 265710 336744 265716 336796
rect 265768 336784 265774 336796
rect 265894 336784 265900 336796
rect 265768 336756 265900 336784
rect 265768 336744 265774 336756
rect 265894 336744 265900 336756
rect 265952 336744 265958 336796
rect 266078 336784 266084 336796
rect 266039 336756 266084 336784
rect 266078 336744 266084 336756
rect 266136 336744 266142 336796
rect 266630 336744 266636 336796
rect 266688 336784 266694 336796
rect 267090 336784 267096 336796
rect 266688 336756 267096 336784
rect 266688 336744 266694 336756
rect 267090 336744 267096 336756
rect 267148 336744 267154 336796
rect 267182 336744 267188 336796
rect 267240 336784 267246 336796
rect 267458 336784 267464 336796
rect 267240 336756 267464 336784
rect 267240 336744 267246 336756
rect 267458 336744 267464 336756
rect 267516 336744 267522 336796
rect 268286 336744 268292 336796
rect 268344 336784 268350 336796
rect 268562 336784 268568 336796
rect 268344 336756 268568 336784
rect 268344 336744 268350 336756
rect 268562 336744 268568 336756
rect 268620 336744 268626 336796
rect 268654 336744 268660 336796
rect 268712 336784 268718 336796
rect 268930 336784 268936 336796
rect 268712 336756 268936 336784
rect 268712 336744 268718 336756
rect 268930 336744 268936 336756
rect 268988 336744 268994 336796
rect 269482 336744 269488 336796
rect 269540 336784 269546 336796
rect 269758 336784 269764 336796
rect 269540 336756 269764 336784
rect 269540 336744 269546 336756
rect 269758 336744 269764 336756
rect 269816 336744 269822 336796
rect 270034 336744 270040 336796
rect 270092 336784 270098 336796
rect 270218 336784 270224 336796
rect 270092 336756 270224 336784
rect 270092 336744 270098 336756
rect 270218 336744 270224 336756
rect 270276 336744 270282 336796
rect 270678 336784 270684 336796
rect 270639 336756 270684 336784
rect 270678 336744 270684 336756
rect 270736 336744 270742 336796
rect 271046 336744 271052 336796
rect 271104 336784 271110 336796
rect 271506 336784 271512 336796
rect 271104 336756 271512 336784
rect 271104 336744 271110 336756
rect 271506 336744 271512 336756
rect 271564 336744 271570 336796
rect 271966 336744 271972 336796
rect 272024 336784 272030 336796
rect 272242 336784 272248 336796
rect 272024 336756 272248 336784
rect 272024 336744 272030 336756
rect 272242 336744 272248 336756
rect 272300 336744 272306 336796
rect 272426 336744 272432 336796
rect 272484 336784 272490 336796
rect 272702 336784 272708 336796
rect 272484 336756 272708 336784
rect 272484 336744 272490 336756
rect 272702 336744 272708 336756
rect 272760 336744 272766 336796
rect 272886 336744 272892 336796
rect 272944 336784 272950 336796
rect 273162 336784 273168 336796
rect 272944 336756 273168 336784
rect 272944 336744 272950 336756
rect 273162 336744 273168 336756
rect 273220 336744 273226 336796
rect 273622 336744 273628 336796
rect 273680 336784 273686 336796
rect 274174 336784 274180 336796
rect 273680 336756 274180 336784
rect 273680 336744 273686 336756
rect 274174 336744 274180 336756
rect 274232 336744 274238 336796
rect 275002 336744 275008 336796
rect 275060 336784 275066 336796
rect 275370 336784 275376 336796
rect 275060 336756 275376 336784
rect 275060 336744 275066 336756
rect 275370 336744 275376 336756
rect 275428 336744 275434 336796
rect 276293 336787 276351 336793
rect 276293 336784 276305 336787
rect 275480 336756 276305 336784
rect 270497 336719 270555 336725
rect 270497 336685 270509 336719
rect 270543 336716 270555 336719
rect 275480 336716 275508 336756
rect 276293 336753 276305 336756
rect 276339 336753 276351 336787
rect 276293 336747 276351 336753
rect 276382 336744 276388 336796
rect 276440 336784 276446 336796
rect 276658 336784 276664 336796
rect 276440 336756 276664 336784
rect 276440 336744 276446 336756
rect 276658 336744 276664 336756
rect 276716 336744 276722 336796
rect 270543 336688 275508 336716
rect 270543 336685 270555 336688
rect 270497 336679 270555 336685
rect 276106 336676 276112 336728
rect 276164 336716 276170 336728
rect 276768 336716 276796 336824
rect 277302 336812 277308 336824
rect 277360 336812 277366 336864
rect 277489 336855 277547 336861
rect 277489 336821 277501 336855
rect 277535 336852 277547 336855
rect 283009 336855 283067 336861
rect 283009 336852 283021 336855
rect 277535 336824 283021 336852
rect 277535 336821 277547 336824
rect 277489 336815 277547 336821
rect 283009 336821 283021 336824
rect 283055 336821 283067 336855
rect 283009 336815 283067 336821
rect 276934 336744 276940 336796
rect 276992 336784 276998 336796
rect 277210 336784 277216 336796
rect 276992 336756 277216 336784
rect 276992 336744 276998 336756
rect 277210 336744 277216 336756
rect 277268 336744 277274 336796
rect 277578 336744 277584 336796
rect 277636 336784 277642 336796
rect 277762 336784 277768 336796
rect 277636 336756 277768 336784
rect 277636 336744 277642 336756
rect 277762 336744 277768 336756
rect 277820 336744 277826 336796
rect 277946 336744 277952 336796
rect 278004 336784 278010 336796
rect 278222 336784 278228 336796
rect 278004 336756 278228 336784
rect 278004 336744 278010 336756
rect 278222 336744 278228 336756
rect 278280 336744 278286 336796
rect 278498 336744 278504 336796
rect 278556 336784 278562 336796
rect 278556 336756 279464 336784
rect 278556 336744 278562 336756
rect 276164 336688 276796 336716
rect 276164 336676 276170 336688
rect 262858 336648 262864 336660
rect 262416 336620 262864 336648
rect 262858 336608 262864 336620
rect 262916 336608 262922 336660
rect 279436 336648 279464 336756
rect 279510 336744 279516 336796
rect 279568 336784 279574 336796
rect 279970 336784 279976 336796
rect 279568 336756 279976 336784
rect 279568 336744 279574 336756
rect 279970 336744 279976 336756
rect 280028 336744 280034 336796
rect 280154 336744 280160 336796
rect 280212 336784 280218 336796
rect 280430 336784 280436 336796
rect 280212 336756 280436 336784
rect 280212 336744 280218 336756
rect 280430 336744 280436 336756
rect 280488 336744 280494 336796
rect 280522 336744 280528 336796
rect 280580 336784 280586 336796
rect 280798 336784 280804 336796
rect 280580 336756 280660 336784
rect 280759 336756 280804 336784
rect 280580 336744 280586 336756
rect 280632 336716 280660 336756
rect 280798 336744 280804 336756
rect 280856 336744 280862 336796
rect 280982 336744 280988 336796
rect 281040 336784 281046 336796
rect 281442 336784 281448 336796
rect 281040 336756 281448 336784
rect 281040 336744 281046 336756
rect 281442 336744 281448 336756
rect 281500 336744 281506 336796
rect 281626 336744 281632 336796
rect 281684 336784 281690 336796
rect 281684 336756 282040 336784
rect 281684 336744 281690 336756
rect 280890 336716 280896 336728
rect 280632 336688 280896 336716
rect 280890 336676 280896 336688
rect 280948 336676 280954 336728
rect 282012 336716 282040 336756
rect 282086 336744 282092 336796
rect 282144 336784 282150 336796
rect 282638 336784 282644 336796
rect 282144 336756 282644 336784
rect 282144 336744 282150 336756
rect 282638 336744 282644 336756
rect 282696 336744 282702 336796
rect 282733 336787 282791 336793
rect 282733 336753 282745 336787
rect 282779 336784 282791 336787
rect 284220 336784 284248 337028
rect 287793 337025 287805 337028
rect 287839 337025 287851 337059
rect 287793 337019 287851 337025
rect 287977 337059 288035 337065
rect 287977 337025 287989 337059
rect 288023 337056 288035 337059
rect 290458 337056 290464 337068
rect 288023 337028 290464 337056
rect 288023 337025 288035 337028
rect 287977 337019 288035 337025
rect 290458 337016 290464 337028
rect 290516 337016 290522 337068
rect 284478 336948 284484 337000
rect 284536 336988 284542 337000
rect 285490 336988 285496 337000
rect 284536 336960 285496 336988
rect 284536 336948 284542 336960
rect 285490 336948 285496 336960
rect 285548 336948 285554 337000
rect 286226 336948 286232 337000
rect 286284 336988 286290 337000
rect 286870 336988 286876 337000
rect 286284 336960 286876 336988
rect 286284 336948 286290 336960
rect 286870 336948 286876 336960
rect 286928 336948 286934 337000
rect 288526 336948 288532 337000
rect 288584 336988 288590 337000
rect 290734 336988 290740 337000
rect 288584 336960 290740 336988
rect 288584 336948 288590 336960
rect 290734 336948 290740 336960
rect 290792 336948 290798 337000
rect 285674 336880 285680 336932
rect 285732 336920 285738 336932
rect 286318 336920 286324 336932
rect 285732 336892 286324 336920
rect 285732 336880 285738 336892
rect 286318 336880 286324 336892
rect 286376 336880 286382 336932
rect 288618 336880 288624 336932
rect 288676 336920 288682 336932
rect 290550 336920 290556 336932
rect 288676 336892 290556 336920
rect 288676 336880 288682 336892
rect 290550 336880 290556 336892
rect 290608 336880 290614 336932
rect 285950 336812 285956 336864
rect 286008 336852 286014 336864
rect 286410 336852 286416 336864
rect 286008 336824 286416 336852
rect 286008 336812 286014 336824
rect 286410 336812 286416 336824
rect 286468 336812 286474 336864
rect 287514 336812 287520 336864
rect 287572 336852 287578 336864
rect 288066 336852 288072 336864
rect 287572 336824 288072 336852
rect 287572 336812 287578 336824
rect 288066 336812 288072 336824
rect 288124 336812 288130 336864
rect 288894 336812 288900 336864
rect 288952 336852 288958 336864
rect 290642 336852 290648 336864
rect 288952 336824 290648 336852
rect 288952 336812 288958 336824
rect 290642 336812 290648 336824
rect 290700 336812 290706 336864
rect 282779 336756 284248 336784
rect 282779 336753 282791 336756
rect 282733 336747 282791 336753
rect 284294 336744 284300 336796
rect 284352 336784 284358 336796
rect 284570 336784 284576 336796
rect 284352 336756 284576 336784
rect 284352 336744 284358 336756
rect 284570 336744 284576 336756
rect 284628 336744 284634 336796
rect 286042 336744 286048 336796
rect 286100 336784 286106 336796
rect 286502 336784 286508 336796
rect 286100 336756 286508 336784
rect 286100 336744 286106 336756
rect 286502 336744 286508 336756
rect 286560 336744 286566 336796
rect 286686 336744 286692 336796
rect 286744 336784 286750 336796
rect 286870 336784 286876 336796
rect 286744 336756 286876 336784
rect 286744 336744 286750 336756
rect 286870 336744 286876 336756
rect 286928 336744 286934 336796
rect 287698 336744 287704 336796
rect 287756 336784 287762 336796
rect 287974 336784 287980 336796
rect 287756 336756 287980 336784
rect 287756 336744 287762 336756
rect 287974 336744 287980 336756
rect 288032 336744 288038 336796
rect 289078 336744 289084 336796
rect 289136 336784 289142 336796
rect 289446 336784 289452 336796
rect 289136 336756 289452 336784
rect 289136 336744 289142 336756
rect 289446 336744 289452 336756
rect 289504 336744 289510 336796
rect 289814 336744 289820 336796
rect 289872 336784 289878 336796
rect 291102 336784 291108 336796
rect 289872 336756 291108 336784
rect 289872 336744 289878 336756
rect 291102 336744 291108 336756
rect 291160 336744 291166 336796
rect 282822 336716 282828 336728
rect 282012 336688 282828 336716
rect 282822 336676 282828 336688
rect 282880 336676 282886 336728
rect 283009 336719 283067 336725
rect 283009 336685 283021 336719
rect 283055 336716 283067 336719
rect 283282 336716 283288 336728
rect 283055 336688 283288 336716
rect 283055 336685 283067 336688
rect 283009 336679 283067 336685
rect 283282 336676 283288 336688
rect 283340 336676 283346 336728
rect 280154 336648 280160 336660
rect 279436 336620 280160 336648
rect 280154 336608 280160 336620
rect 280212 336608 280218 336660
rect 280706 336608 280712 336660
rect 280764 336648 280770 336660
rect 293954 336648 293960 336660
rect 280764 336620 293960 336648
rect 280764 336608 280770 336620
rect 293954 336608 293960 336620
rect 294012 336608 294018 336660
rect 231857 336583 231915 336589
rect 231857 336549 231869 336583
rect 231903 336580 231915 336583
rect 239030 336580 239036 336592
rect 231903 336552 239036 336580
rect 231903 336549 231915 336552
rect 231857 336543 231915 336549
rect 239030 336540 239036 336552
rect 239088 336540 239094 336592
rect 279602 336540 279608 336592
rect 279660 336580 279666 336592
rect 296714 336580 296720 336592
rect 279660 336552 296720 336580
rect 279660 336540 279666 336552
rect 296714 336540 296720 336552
rect 296772 336540 296778 336592
rect 227622 336472 227628 336524
rect 227680 336512 227686 336524
rect 242894 336512 242900 336524
rect 227680 336484 242900 336512
rect 227680 336472 227686 336484
rect 242894 336472 242900 336484
rect 242952 336472 242958 336524
rect 261662 336472 261668 336524
rect 261720 336512 261726 336524
rect 304994 336512 305000 336524
rect 261720 336484 305000 336512
rect 261720 336472 261726 336484
rect 304994 336472 305000 336484
rect 305052 336472 305058 336524
rect 220722 336404 220728 336456
rect 220780 336444 220786 336456
rect 252646 336444 252652 336456
rect 220780 336416 252652 336444
rect 220780 336404 220786 336416
rect 252646 336404 252652 336416
rect 252704 336404 252710 336456
rect 265526 336404 265532 336456
rect 265584 336444 265590 336456
rect 314654 336444 314660 336456
rect 265584 336416 314660 336444
rect 265584 336404 265590 336416
rect 314654 336404 314660 336416
rect 314712 336404 314718 336456
rect 104897 336379 104955 336385
rect 104897 336345 104909 336379
rect 104943 336376 104955 336379
rect 114465 336379 114523 336385
rect 114465 336376 114477 336379
rect 104943 336348 114477 336376
rect 104943 336345 104955 336348
rect 104897 336339 104955 336345
rect 114465 336345 114477 336348
rect 114511 336345 114523 336379
rect 114465 336339 114523 336345
rect 216582 336336 216588 336388
rect 216640 336376 216646 336388
rect 252094 336376 252100 336388
rect 216640 336348 252100 336376
rect 216640 336336 216646 336348
rect 252094 336336 252100 336348
rect 252152 336336 252158 336388
rect 267734 336336 267740 336388
rect 267792 336376 267798 336388
rect 327074 336376 327080 336388
rect 267792 336348 327080 336376
rect 267792 336336 267798 336348
rect 327074 336336 327080 336348
rect 327132 336336 327138 336388
rect 209682 336268 209688 336320
rect 209740 336308 209746 336320
rect 248506 336308 248512 336320
rect 209740 336280 248512 336308
rect 209740 336268 209746 336280
rect 248506 336268 248512 336280
rect 248564 336268 248570 336320
rect 265342 336268 265348 336320
rect 265400 336308 265406 336320
rect 265526 336308 265532 336320
rect 265400 336280 265532 336308
rect 265400 336268 265406 336280
rect 265526 336268 265532 336280
rect 265584 336268 265590 336320
rect 266998 336268 267004 336320
rect 267056 336308 267062 336320
rect 353294 336308 353300 336320
rect 267056 336280 353300 336308
rect 267056 336268 267062 336280
rect 353294 336268 353300 336280
rect 353352 336268 353358 336320
rect 114465 336243 114523 336249
rect 114465 336209 114477 336243
rect 114511 336240 114523 336243
rect 115845 336243 115903 336249
rect 115845 336240 115857 336243
rect 114511 336212 115857 336240
rect 114511 336209 114523 336212
rect 114465 336203 114523 336209
rect 115845 336209 115857 336212
rect 115891 336209 115903 336243
rect 115845 336203 115903 336209
rect 132497 336243 132555 336249
rect 132497 336209 132509 336243
rect 132543 336240 132555 336243
rect 142065 336243 142123 336249
rect 142065 336240 142077 336243
rect 132543 336212 142077 336240
rect 132543 336209 132555 336212
rect 132497 336203 132555 336209
rect 142065 336209 142077 336212
rect 142111 336209 142123 336243
rect 142065 336203 142123 336209
rect 143537 336243 143595 336249
rect 143537 336209 143549 336243
rect 143583 336240 143595 336243
rect 143583 336212 153148 336240
rect 143583 336209 143595 336212
rect 143537 336203 143595 336209
rect 57977 336175 58035 336181
rect 57977 336141 57989 336175
rect 58023 336172 58035 336175
rect 62761 336175 62819 336181
rect 62761 336172 62773 336175
rect 58023 336144 62773 336172
rect 58023 336141 58035 336144
rect 57977 336135 58035 336141
rect 62761 336141 62773 336144
rect 62807 336141 62819 336175
rect 62761 336135 62819 336141
rect 115937 336175 115995 336181
rect 115937 336141 115949 336175
rect 115983 336172 115995 336175
rect 115983 336144 128860 336172
rect 115983 336141 115995 336144
rect 115937 336135 115995 336141
rect 96525 336107 96583 336113
rect 96525 336073 96537 336107
rect 96571 336104 96583 336107
rect 104897 336107 104955 336113
rect 104897 336104 104909 336107
rect 96571 336076 104909 336104
rect 96571 336073 96583 336076
rect 96525 336067 96583 336073
rect 104897 336073 104909 336076
rect 104943 336073 104955 336107
rect 128832 336104 128860 336144
rect 132497 336107 132555 336113
rect 132497 336104 132509 336107
rect 128832 336076 132509 336104
rect 104897 336067 104955 336073
rect 132497 336073 132509 336076
rect 132543 336073 132555 336107
rect 132497 336067 132555 336073
rect 142065 336107 142123 336113
rect 142065 336073 142077 336107
rect 142111 336104 142123 336107
rect 143537 336107 143595 336113
rect 143537 336104 143549 336107
rect 142111 336076 143549 336104
rect 142111 336073 142123 336076
rect 142065 336067 142123 336073
rect 143537 336073 143549 336076
rect 143583 336073 143595 336107
rect 153120 336104 153148 336212
rect 162762 336200 162768 336252
rect 162820 336240 162826 336252
rect 234985 336243 235043 336249
rect 234985 336240 234997 336243
rect 162820 336212 234997 336240
rect 162820 336200 162826 336212
rect 234985 336209 234997 336212
rect 235031 336209 235043 336243
rect 234985 336203 235043 336209
rect 275278 336200 275284 336252
rect 275336 336240 275342 336252
rect 440234 336240 440240 336252
rect 275336 336212 440240 336240
rect 275336 336200 275342 336212
rect 440234 336200 440240 336212
rect 440292 336200 440298 336252
rect 176562 336132 176568 336184
rect 176620 336172 176626 336184
rect 211157 336175 211215 336181
rect 211157 336172 211169 336175
rect 176620 336144 211169 336172
rect 176620 336132 176626 336144
rect 211157 336141 211169 336144
rect 211203 336141 211215 336175
rect 211157 336135 211215 336141
rect 211433 336175 211491 336181
rect 211433 336141 211445 336175
rect 211479 336172 211491 336175
rect 248046 336172 248052 336184
rect 211479 336144 248052 336172
rect 211479 336141 211491 336144
rect 211433 336135 211491 336141
rect 248046 336132 248052 336144
rect 248104 336132 248110 336184
rect 289998 336132 290004 336184
rect 290056 336172 290062 336184
rect 483014 336172 483020 336184
rect 290056 336144 483020 336172
rect 290056 336132 290062 336144
rect 483014 336132 483020 336144
rect 483072 336132 483078 336184
rect 153194 336104 153200 336116
rect 153120 336076 153200 336104
rect 143537 336067 143595 336073
rect 153194 336064 153200 336076
rect 153252 336064 153258 336116
rect 153286 336064 153292 336116
rect 153344 336104 153350 336116
rect 211246 336104 211252 336116
rect 153344 336076 211252 336104
rect 153344 336064 153350 336076
rect 211246 336064 211252 336076
rect 211304 336064 211310 336116
rect 211338 336064 211344 336116
rect 211396 336104 211402 336116
rect 231857 336107 231915 336113
rect 231857 336104 231869 336107
rect 211396 336076 231869 336104
rect 211396 336064 211402 336076
rect 231857 336073 231869 336076
rect 231903 336073 231915 336107
rect 231857 336067 231915 336073
rect 236270 336064 236276 336116
rect 236328 336104 236334 336116
rect 236546 336104 236552 336116
rect 236328 336076 236552 336104
rect 236328 336064 236334 336076
rect 236546 336064 236552 336076
rect 236604 336064 236610 336116
rect 248690 336104 248696 336116
rect 248651 336076 248696 336104
rect 248690 336064 248696 336076
rect 248748 336064 248754 336116
rect 284018 336064 284024 336116
rect 284076 336104 284082 336116
rect 521654 336104 521660 336116
rect 284076 336076 521660 336104
rect 284076 336064 284082 336076
rect 521654 336064 521660 336076
rect 521712 336064 521718 336116
rect 52362 335996 52368 336048
rect 52420 336036 52426 336048
rect 57977 336039 58035 336045
rect 57977 336036 57989 336039
rect 52420 336008 57989 336036
rect 52420 335996 52426 336008
rect 57977 336005 57989 336008
rect 58023 336005 58035 336039
rect 57977 335999 58035 336005
rect 77220 336008 77340 336036
rect 77220 335977 77248 336008
rect 77312 335977 77340 336008
rect 89622 335996 89628 336048
rect 89680 336036 89686 336048
rect 96433 336039 96491 336045
rect 96433 336036 96445 336039
rect 89680 336008 96445 336036
rect 89680 335996 89686 336008
rect 96433 336005 96445 336008
rect 96479 336005 96491 336039
rect 129093 336039 129151 336045
rect 96433 335999 96491 336005
rect 96540 336008 96660 336036
rect 96540 335977 96568 336008
rect 96632 335977 96660 336008
rect 109236 336008 115980 336036
rect 62761 335971 62819 335977
rect 62761 335937 62773 335971
rect 62807 335968 62819 335971
rect 67637 335971 67695 335977
rect 67637 335968 67649 335971
rect 62807 335940 67649 335968
rect 62807 335937 62819 335940
rect 62761 335931 62819 335937
rect 67637 335937 67649 335940
rect 67683 335937 67695 335971
rect 67637 335931 67695 335937
rect 77205 335971 77263 335977
rect 77205 335937 77217 335971
rect 77251 335937 77263 335971
rect 77205 335931 77263 335937
rect 77297 335971 77355 335977
rect 77297 335937 77309 335971
rect 77343 335937 77355 335971
rect 77297 335931 77355 335937
rect 81621 335971 81679 335977
rect 81621 335937 81633 335971
rect 81667 335968 81679 335971
rect 86957 335971 87015 335977
rect 86957 335968 86969 335971
rect 81667 335940 86969 335968
rect 81667 335937 81679 335940
rect 81621 335931 81679 335937
rect 86957 335937 86969 335940
rect 87003 335937 87015 335971
rect 86957 335931 87015 335937
rect 96525 335971 96583 335977
rect 96525 335937 96537 335971
rect 96571 335937 96583 335971
rect 96525 335931 96583 335937
rect 96617 335971 96675 335977
rect 96617 335937 96629 335971
rect 96663 335937 96675 335971
rect 106461 335971 106519 335977
rect 96617 335931 96675 335937
rect 106200 335940 106320 335968
rect 67637 335835 67695 335841
rect 67637 335801 67649 335835
rect 67683 335832 67695 335835
rect 77205 335835 77263 335841
rect 77205 335832 77217 335835
rect 67683 335804 77217 335832
rect 67683 335801 67695 335804
rect 67637 335795 67695 335801
rect 77205 335801 77217 335804
rect 77251 335801 77263 335835
rect 77205 335795 77263 335801
rect 77297 335835 77355 335841
rect 77297 335801 77309 335835
rect 77343 335832 77355 335835
rect 81621 335835 81679 335841
rect 81621 335832 81633 335835
rect 77343 335804 81633 335832
rect 77343 335801 77355 335804
rect 77297 335795 77355 335801
rect 81621 335801 81633 335804
rect 81667 335801 81679 335835
rect 81621 335795 81679 335801
rect 86957 335835 87015 335841
rect 86957 335801 86969 335835
rect 87003 335832 87015 335835
rect 96525 335835 96583 335841
rect 96525 335832 96537 335835
rect 87003 335804 96537 335832
rect 87003 335801 87015 335804
rect 86957 335795 87015 335801
rect 96525 335801 96537 335804
rect 96571 335801 96583 335835
rect 96525 335795 96583 335801
rect 96617 335835 96675 335841
rect 96617 335801 96629 335835
rect 96663 335832 96675 335835
rect 106200 335832 106228 335940
rect 106292 335909 106320 335940
rect 106461 335937 106473 335971
rect 106507 335968 106519 335971
rect 109236 335968 109264 336008
rect 115952 335977 115980 336008
rect 129093 336005 129105 336039
rect 129139 336036 129151 336039
rect 129139 336008 132540 336036
rect 129139 336005 129151 336008
rect 129093 335999 129151 336005
rect 132512 335977 132540 336008
rect 153102 335996 153108 336048
rect 153160 336036 153166 336048
rect 176565 336039 176623 336045
rect 176565 336036 176577 336039
rect 153160 336008 153240 336036
rect 153160 335996 153166 336008
rect 106507 335940 109264 335968
rect 115937 335971 115995 335977
rect 106507 335937 106519 335940
rect 106461 335931 106519 335937
rect 115937 335937 115949 335971
rect 115983 335937 115995 335971
rect 115937 335931 115995 335937
rect 132497 335971 132555 335977
rect 132497 335937 132509 335971
rect 132543 335937 132555 335971
rect 132497 335931 132555 335937
rect 142065 335971 142123 335977
rect 142065 335937 142077 335971
rect 142111 335968 142123 335971
rect 143537 335971 143595 335977
rect 143537 335968 143549 335971
rect 142111 335940 143549 335968
rect 142111 335937 142123 335940
rect 142065 335931 142123 335937
rect 143537 335937 143549 335940
rect 143583 335937 143595 335971
rect 153212 335968 153240 336008
rect 153304 336008 176577 336036
rect 153304 335968 153332 336008
rect 176565 336005 176577 336008
rect 176611 336005 176623 336039
rect 176565 335999 176623 336005
rect 189000 336008 189120 336036
rect 189000 335977 189028 336008
rect 189092 335977 189120 336008
rect 232038 335996 232044 336048
rect 232096 336036 232102 336048
rect 232682 336036 232688 336048
rect 232096 336008 232688 336036
rect 232096 335996 232102 336008
rect 232682 335996 232688 336008
rect 232740 335996 232746 336048
rect 287054 335996 287060 336048
rect 287112 336036 287118 336048
rect 554774 336036 554780 336048
rect 287112 336008 554780 336036
rect 287112 335996 287118 336008
rect 554774 335996 554780 336008
rect 554832 335996 554838 336048
rect 153212 335940 153332 335968
rect 176749 335971 176807 335977
rect 143537 335931 143595 335937
rect 176749 335937 176761 335971
rect 176795 335968 176807 335971
rect 179417 335971 179475 335977
rect 179417 335968 179429 335971
rect 176795 335940 179429 335968
rect 176795 335937 176807 335940
rect 176749 335931 176807 335937
rect 179417 335937 179429 335940
rect 179463 335937 179475 335971
rect 179417 335931 179475 335937
rect 188985 335971 189043 335977
rect 188985 335937 188997 335971
rect 189031 335937 189043 335971
rect 188985 335931 189043 335937
rect 189077 335971 189135 335977
rect 189077 335937 189089 335971
rect 189123 335937 189135 335971
rect 189077 335931 189135 335937
rect 196069 335971 196127 335977
rect 196069 335937 196081 335971
rect 196115 335968 196127 335971
rect 198737 335971 198795 335977
rect 198737 335968 198749 335971
rect 196115 335940 198749 335968
rect 196115 335937 196127 335940
rect 196069 335931 196127 335937
rect 198737 335937 198749 335940
rect 198783 335937 198795 335971
rect 198737 335931 198795 335937
rect 208305 335971 208363 335977
rect 208305 335937 208317 335971
rect 208351 335968 208363 335971
rect 209685 335971 209743 335977
rect 209685 335968 209697 335971
rect 208351 335940 209697 335968
rect 208351 335937 208363 335940
rect 208305 335931 208363 335937
rect 209685 335937 209697 335940
rect 209731 335937 209743 335971
rect 209685 335931 209743 335937
rect 209777 335971 209835 335977
rect 209777 335937 209789 335971
rect 209823 335968 209835 335971
rect 209823 335940 218008 335968
rect 209823 335937 209835 335940
rect 209777 335931 209835 335937
rect 106277 335903 106335 335909
rect 106277 335869 106289 335903
rect 106323 335869 106335 335903
rect 129001 335903 129059 335909
rect 129001 335900 129013 335903
rect 106277 335863 106335 335869
rect 119172 335872 129013 335900
rect 96663 335804 106228 335832
rect 115937 335835 115995 335841
rect 96663 335801 96675 335804
rect 96617 335795 96675 335801
rect 115937 335801 115949 335835
rect 115983 335832 115995 335835
rect 119172 335832 119200 335872
rect 129001 335869 129013 335872
rect 129047 335869 129059 335903
rect 129001 335863 129059 335869
rect 143629 335903 143687 335909
rect 143629 335869 143641 335903
rect 143675 335900 143687 335903
rect 153102 335900 153108 335912
rect 143675 335872 153108 335900
rect 143675 335869 143687 335872
rect 143629 335863 143687 335869
rect 153102 335860 153108 335872
rect 153160 335860 153166 335912
rect 217980 335900 218008 335940
rect 232222 335928 232228 335980
rect 232280 335968 232286 335980
rect 232774 335968 232780 335980
rect 232280 335940 232780 335968
rect 232280 335928 232286 335940
rect 232774 335928 232780 335940
rect 232832 335928 232838 335980
rect 233234 335900 233240 335912
rect 217980 335872 233240 335900
rect 233234 335860 233240 335872
rect 233292 335860 233298 335912
rect 244642 335860 244648 335912
rect 244700 335900 244706 335912
rect 245102 335900 245108 335912
rect 244700 335872 245108 335900
rect 244700 335860 244706 335872
rect 245102 335860 245108 335872
rect 245160 335860 245166 335912
rect 251358 335860 251364 335912
rect 251416 335900 251422 335912
rect 251726 335900 251732 335912
rect 251416 335872 251732 335900
rect 251416 335860 251422 335872
rect 251726 335860 251732 335872
rect 251784 335860 251790 335912
rect 115983 335804 119200 335832
rect 132497 335835 132555 335841
rect 115983 335801 115995 335804
rect 115937 335795 115995 335801
rect 132497 335801 132509 335835
rect 132543 335832 132555 335835
rect 142065 335835 142123 335841
rect 142065 335832 142077 335835
rect 132543 335804 142077 335832
rect 132543 335801 132555 335804
rect 132497 335795 132555 335801
rect 142065 335801 142077 335804
rect 142111 335801 142123 335835
rect 142065 335795 142123 335801
rect 179417 335835 179475 335841
rect 179417 335801 179429 335835
rect 179463 335832 179475 335835
rect 188985 335835 189043 335841
rect 188985 335832 188997 335835
rect 179463 335804 188997 335832
rect 179463 335801 179475 335804
rect 179417 335795 179475 335801
rect 188985 335801 188997 335804
rect 189031 335801 189043 335835
rect 188985 335795 189043 335801
rect 189077 335835 189135 335841
rect 189077 335801 189089 335835
rect 189123 335832 189135 335835
rect 196069 335835 196127 335841
rect 196069 335832 196081 335835
rect 189123 335804 196081 335832
rect 189123 335801 189135 335804
rect 189077 335795 189135 335801
rect 196069 335801 196081 335804
rect 196115 335801 196127 335835
rect 196069 335795 196127 335801
rect 198737 335835 198795 335841
rect 198737 335801 198749 335835
rect 198783 335832 198795 335835
rect 208305 335835 208363 335841
rect 208305 335832 208317 335835
rect 198783 335804 208317 335832
rect 198783 335801 198795 335804
rect 198737 335795 198795 335801
rect 208305 335801 208317 335804
rect 208351 335801 208363 335835
rect 208305 335795 208363 335801
rect 233510 335792 233516 335844
rect 233568 335832 233574 335844
rect 233694 335832 233700 335844
rect 233568 335804 233700 335832
rect 233568 335792 233574 335804
rect 233694 335792 233700 335804
rect 233752 335792 233758 335844
rect 240502 335792 240508 335844
rect 240560 335832 240566 335844
rect 241422 335832 241428 335844
rect 240560 335804 241428 335832
rect 240560 335792 240566 335804
rect 241422 335792 241428 335804
rect 241480 335792 241486 335844
rect 244274 335792 244280 335844
rect 244332 335832 244338 335844
rect 244734 335832 244740 335844
rect 244332 335804 244740 335832
rect 244332 335792 244338 335804
rect 244734 335792 244740 335804
rect 244792 335792 244798 335844
rect 246206 335832 246212 335844
rect 246167 335804 246212 335832
rect 246206 335792 246212 335804
rect 246264 335792 246270 335844
rect 248506 335792 248512 335844
rect 248564 335832 248570 335844
rect 249518 335832 249524 335844
rect 248564 335804 249524 335832
rect 248564 335792 248570 335804
rect 249518 335792 249524 335804
rect 249576 335792 249582 335844
rect 236454 335724 236460 335776
rect 236512 335764 236518 335776
rect 236730 335764 236736 335776
rect 236512 335736 236736 335764
rect 236512 335724 236518 335736
rect 236730 335724 236736 335736
rect 236788 335724 236794 335776
rect 237742 335724 237748 335776
rect 237800 335764 237806 335776
rect 238478 335764 238484 335776
rect 237800 335736 238484 335764
rect 237800 335724 237806 335736
rect 238478 335724 238484 335736
rect 238536 335724 238542 335776
rect 245562 335764 245568 335776
rect 245523 335736 245568 335764
rect 245562 335724 245568 335736
rect 245620 335724 245626 335776
rect 250346 335724 250352 335776
rect 250404 335764 250410 335776
rect 251082 335764 251088 335776
rect 250404 335736 251088 335764
rect 250404 335724 250410 335736
rect 251082 335724 251088 335736
rect 251140 335724 251146 335776
rect 251450 335724 251456 335776
rect 251508 335764 251514 335776
rect 252186 335764 252192 335776
rect 251508 335736 252192 335764
rect 251508 335724 251514 335736
rect 252186 335724 252192 335736
rect 252244 335724 252250 335776
rect 284389 335767 284447 335773
rect 284389 335733 284401 335767
rect 284435 335764 284447 335767
rect 284938 335764 284944 335776
rect 284435 335736 284944 335764
rect 284435 335733 284447 335736
rect 284389 335727 284447 335733
rect 284938 335724 284944 335736
rect 284996 335724 285002 335776
rect 230198 335696 230204 335708
rect 229388 335668 230204 335696
rect 229388 335640 229416 335668
rect 230198 335656 230204 335668
rect 230256 335656 230262 335708
rect 236362 335656 236368 335708
rect 236420 335696 236426 335708
rect 236638 335696 236644 335708
rect 236420 335668 236644 335696
rect 236420 335656 236426 335668
rect 236638 335656 236644 335668
rect 236696 335656 236702 335708
rect 240318 335656 240324 335708
rect 240376 335696 240382 335708
rect 241054 335696 241060 335708
rect 240376 335668 241060 335696
rect 240376 335656 240382 335668
rect 241054 335656 241060 335668
rect 241112 335656 241118 335708
rect 244458 335656 244464 335708
rect 244516 335656 244522 335708
rect 245746 335656 245752 335708
rect 245804 335656 245810 335708
rect 246022 335656 246028 335708
rect 246080 335696 246086 335708
rect 246666 335696 246672 335708
rect 246080 335668 246672 335696
rect 246080 335656 246086 335668
rect 246666 335656 246672 335668
rect 246724 335656 246730 335708
rect 248414 335656 248420 335708
rect 248472 335696 248478 335708
rect 248782 335696 248788 335708
rect 248472 335668 248788 335696
rect 248472 335656 248478 335668
rect 248782 335656 248788 335668
rect 248840 335656 248846 335708
rect 248966 335656 248972 335708
rect 249024 335696 249030 335708
rect 249334 335696 249340 335708
rect 249024 335668 249340 335696
rect 249024 335656 249030 335668
rect 249334 335656 249340 335668
rect 249392 335656 249398 335708
rect 250162 335656 250168 335708
rect 250220 335696 250226 335708
rect 250714 335696 250720 335708
rect 250220 335668 250720 335696
rect 250220 335656 250226 335668
rect 250714 335656 250720 335668
rect 250772 335656 250778 335708
rect 251542 335696 251548 335708
rect 251503 335668 251548 335696
rect 251542 335656 251548 335668
rect 251600 335656 251606 335708
rect 251634 335656 251640 335708
rect 251692 335696 251698 335708
rect 252094 335696 252100 335708
rect 251692 335668 252100 335696
rect 251692 335656 251698 335668
rect 252094 335656 252100 335668
rect 252152 335656 252158 335708
rect 252278 335656 252284 335708
rect 252336 335656 252342 335708
rect 254026 335656 254032 335708
rect 254084 335696 254090 335708
rect 254394 335696 254400 335708
rect 254084 335668 254400 335696
rect 254084 335656 254090 335668
rect 254394 335656 254400 335668
rect 254452 335656 254458 335708
rect 269298 335656 269304 335708
rect 269356 335696 269362 335708
rect 269850 335696 269856 335708
rect 269356 335668 269856 335696
rect 269356 335656 269362 335668
rect 269850 335656 269856 335668
rect 269908 335656 269914 335708
rect 287606 335696 287612 335708
rect 287567 335668 287612 335696
rect 287606 335656 287612 335668
rect 287664 335656 287670 335708
rect 229370 335588 229376 335640
rect 229428 335588 229434 335640
rect 230658 335588 230664 335640
rect 230716 335628 230722 335640
rect 231394 335628 231400 335640
rect 230716 335600 231400 335628
rect 230716 335588 230722 335600
rect 231394 335588 231400 335600
rect 231452 335588 231458 335640
rect 236086 335588 236092 335640
rect 236144 335628 236150 335640
rect 236822 335628 236828 335640
rect 236144 335600 236828 335628
rect 236144 335588 236150 335600
rect 236822 335588 236828 335600
rect 236880 335588 236886 335640
rect 237742 335588 237748 335640
rect 237800 335628 237806 335640
rect 238110 335628 238116 335640
rect 237800 335600 238116 335628
rect 237800 335588 237806 335600
rect 238110 335588 238116 335600
rect 238168 335588 238174 335640
rect 238846 335588 238852 335640
rect 238904 335628 238910 335640
rect 239766 335628 239772 335640
rect 238904 335600 239772 335628
rect 238904 335588 238910 335600
rect 239766 335588 239772 335600
rect 239824 335588 239830 335640
rect 240686 335588 240692 335640
rect 240744 335628 240750 335640
rect 240962 335628 240968 335640
rect 240744 335600 240968 335628
rect 240744 335588 240750 335600
rect 240962 335588 240968 335600
rect 241020 335588 241026 335640
rect 241514 335588 241520 335640
rect 241572 335628 241578 335640
rect 241882 335628 241888 335640
rect 241572 335600 241888 335628
rect 241572 335588 241578 335600
rect 241882 335588 241888 335600
rect 241940 335588 241946 335640
rect 242158 335588 242164 335640
rect 242216 335628 242222 335640
rect 242434 335628 242440 335640
rect 242216 335600 242440 335628
rect 242216 335588 242222 335600
rect 242434 335588 242440 335600
rect 242492 335588 242498 335640
rect 242526 335588 242532 335640
rect 242584 335628 242590 335640
rect 242710 335628 242716 335640
rect 242584 335600 242716 335628
rect 242584 335588 242590 335600
rect 242710 335588 242716 335600
rect 242768 335588 242774 335640
rect 240410 335520 240416 335572
rect 240468 335560 240474 335572
rect 240778 335560 240784 335572
rect 240468 335532 240784 335560
rect 240468 335520 240474 335532
rect 240778 335520 240784 335532
rect 240836 335520 240842 335572
rect 233326 335452 233332 335504
rect 233384 335492 233390 335504
rect 234154 335492 234160 335504
rect 233384 335464 234160 335492
rect 233384 335452 233390 335464
rect 234154 335452 234160 335464
rect 234212 335452 234218 335504
rect 235994 335452 236000 335504
rect 236052 335492 236058 335504
rect 236454 335492 236460 335504
rect 236052 335464 236460 335492
rect 236052 335452 236058 335464
rect 236454 335452 236460 335464
rect 236512 335452 236518 335504
rect 244476 335424 244504 335656
rect 244642 335588 244648 335640
rect 244700 335628 244706 335640
rect 244918 335628 244924 335640
rect 244700 335600 244924 335628
rect 244700 335588 244706 335600
rect 244918 335588 244924 335600
rect 244976 335588 244982 335640
rect 245010 335588 245016 335640
rect 245068 335628 245074 335640
rect 245562 335628 245568 335640
rect 245068 335600 245568 335628
rect 245068 335588 245074 335600
rect 245562 335588 245568 335600
rect 245620 335588 245626 335640
rect 245764 335560 245792 335656
rect 247402 335588 247408 335640
rect 247460 335628 247466 335640
rect 247586 335628 247592 335640
rect 247460 335600 247592 335628
rect 247460 335588 247466 335600
rect 247586 335588 247592 335600
rect 247644 335588 247650 335640
rect 249242 335588 249248 335640
rect 249300 335628 249306 335640
rect 249610 335628 249616 335640
rect 249300 335600 249616 335628
rect 249300 335588 249306 335600
rect 249610 335588 249616 335600
rect 249668 335588 249674 335640
rect 245764 335532 246436 335560
rect 246408 335504 246436 335532
rect 245930 335452 245936 335504
rect 245988 335492 245994 335504
rect 246206 335492 246212 335504
rect 245988 335464 246212 335492
rect 245988 335452 245994 335464
rect 246206 335452 246212 335464
rect 246264 335452 246270 335504
rect 246390 335452 246396 335504
rect 246448 335452 246454 335504
rect 249794 335452 249800 335504
rect 249852 335492 249858 335504
rect 250070 335492 250076 335504
rect 249852 335464 250076 335492
rect 249852 335452 249858 335464
rect 250070 335452 250076 335464
rect 250128 335452 250134 335504
rect 251910 335452 251916 335504
rect 251968 335492 251974 335504
rect 252296 335492 252324 335656
rect 252922 335588 252928 335640
rect 252980 335628 252986 335640
rect 253842 335628 253848 335640
rect 252980 335600 253848 335628
rect 252980 335588 252986 335600
rect 253842 335588 253848 335600
rect 253900 335588 253906 335640
rect 255498 335588 255504 335640
rect 255556 335628 255562 335640
rect 256234 335628 256240 335640
rect 255556 335600 256240 335628
rect 255556 335588 255562 335600
rect 256234 335588 256240 335600
rect 256292 335588 256298 335640
rect 254118 335520 254124 335572
rect 254176 335520 254182 335572
rect 256050 335560 256056 335572
rect 255608 335532 256056 335560
rect 251968 335464 252324 335492
rect 251968 335452 251974 335464
rect 244292 335396 244504 335424
rect 244292 335368 244320 335396
rect 244274 335316 244280 335368
rect 244332 335316 244338 335368
rect 244366 335316 244372 335368
rect 244424 335356 244430 335368
rect 245194 335356 245200 335368
rect 244424 335328 245200 335356
rect 244424 335316 244430 335328
rect 245194 335316 245200 335328
rect 245252 335316 245258 335368
rect 248874 335316 248880 335368
rect 248932 335356 248938 335368
rect 249702 335356 249708 335368
rect 248932 335328 249708 335356
rect 248932 335316 248938 335328
rect 249702 335316 249708 335328
rect 249760 335316 249766 335368
rect 249794 335316 249800 335368
rect 249852 335356 249858 335368
rect 250438 335356 250444 335368
rect 249852 335328 250444 335356
rect 249852 335316 249858 335328
rect 250438 335316 250444 335328
rect 250496 335316 250502 335368
rect 251726 335356 251732 335368
rect 251687 335328 251732 335356
rect 251726 335316 251732 335328
rect 251784 335316 251790 335368
rect 249886 335248 249892 335300
rect 249944 335288 249950 335300
rect 250622 335288 250628 335300
rect 249944 335260 250628 335288
rect 249944 335248 249950 335260
rect 250622 335248 250628 335260
rect 250680 335248 250686 335300
rect 254136 335220 254164 335520
rect 254302 335316 254308 335368
rect 254360 335356 254366 335368
rect 254670 335356 254676 335368
rect 254360 335328 254676 335356
rect 254360 335316 254366 335328
rect 254670 335316 254676 335328
rect 254728 335316 254734 335368
rect 254486 335220 254492 335232
rect 254136 335192 254492 335220
rect 254486 335180 254492 335192
rect 254544 335180 254550 335232
rect 255608 335220 255636 335532
rect 256050 335520 256056 335532
rect 256108 335520 256114 335572
rect 277670 335520 277676 335572
rect 277728 335520 277734 335572
rect 256786 335452 256792 335504
rect 256844 335492 256850 335504
rect 257798 335492 257804 335504
rect 256844 335464 257804 335492
rect 256844 335452 256850 335464
rect 257798 335452 257804 335464
rect 257856 335452 257862 335504
rect 269574 335452 269580 335504
rect 269632 335492 269638 335504
rect 269942 335492 269948 335504
rect 269632 335464 269948 335492
rect 269632 335452 269638 335464
rect 269942 335452 269948 335464
rect 270000 335452 270006 335504
rect 272150 335452 272156 335504
rect 272208 335492 272214 335504
rect 272518 335492 272524 335504
rect 272208 335464 272524 335492
rect 272208 335452 272214 335464
rect 272518 335452 272524 335464
rect 272576 335452 272582 335504
rect 269390 335384 269396 335436
rect 269448 335424 269454 335436
rect 270126 335424 270132 335436
rect 269448 335396 270132 335424
rect 269448 335384 269454 335396
rect 270126 335384 270132 335396
rect 270184 335384 270190 335436
rect 277688 335368 277716 335520
rect 279510 335452 279516 335504
rect 279568 335492 279574 335504
rect 279786 335492 279792 335504
rect 279568 335464 279792 335492
rect 279568 335452 279574 335464
rect 279786 335452 279792 335464
rect 279844 335452 279850 335504
rect 255682 335316 255688 335368
rect 255740 335356 255746 335368
rect 256050 335356 256056 335368
rect 255740 335328 256056 335356
rect 255740 335316 255746 335328
rect 256050 335316 256056 335328
rect 256108 335316 256114 335368
rect 269574 335316 269580 335368
rect 269632 335356 269638 335368
rect 270310 335356 270316 335368
rect 269632 335328 270316 335356
rect 269632 335316 269638 335328
rect 270310 335316 270316 335328
rect 270368 335316 270374 335368
rect 277670 335316 277676 335368
rect 277728 335316 277734 335368
rect 280154 335316 280160 335368
rect 280212 335356 280218 335368
rect 280522 335356 280528 335368
rect 280212 335328 280528 335356
rect 280212 335316 280218 335328
rect 280522 335316 280528 335328
rect 280580 335316 280586 335368
rect 256418 335288 256424 335300
rect 256379 335260 256424 335288
rect 256418 335248 256424 335260
rect 256476 335248 256482 335300
rect 280430 335288 280436 335300
rect 280391 335260 280436 335288
rect 280430 335248 280436 335260
rect 280488 335248 280494 335300
rect 255682 335220 255688 335232
rect 255608 335192 255688 335220
rect 255682 335180 255688 335192
rect 255740 335180 255746 335232
rect 278866 335180 278872 335232
rect 278924 335220 278930 335232
rect 279326 335220 279332 335232
rect 278924 335192 279332 335220
rect 278924 335180 278930 335192
rect 279326 335180 279332 335192
rect 279384 335180 279390 335232
rect 280154 335220 280160 335232
rect 280115 335192 280160 335220
rect 280154 335180 280160 335192
rect 280212 335180 280218 335232
rect 229002 335112 229008 335164
rect 229060 335152 229066 335164
rect 253382 335152 253388 335164
rect 229060 335124 253388 335152
rect 229060 335112 229066 335124
rect 253382 335112 253388 335124
rect 253440 335112 253446 335164
rect 278958 335152 278964 335164
rect 278919 335124 278964 335152
rect 278958 335112 278964 335124
rect 279016 335112 279022 335164
rect 282457 335155 282515 335161
rect 282457 335121 282469 335155
rect 282503 335152 282515 335155
rect 282503 335124 282684 335152
rect 282503 335121 282515 335124
rect 282457 335115 282515 335121
rect 223482 335044 223488 335096
rect 223540 335084 223546 335096
rect 249518 335084 249524 335096
rect 223540 335056 249524 335084
rect 223540 335044 223546 335056
rect 249518 335044 249524 335056
rect 249576 335044 249582 335096
rect 281626 335044 281632 335096
rect 281684 335084 281690 335096
rect 282546 335084 282552 335096
rect 281684 335056 282552 335084
rect 281684 335044 281690 335056
rect 282546 335044 282552 335056
rect 282604 335044 282610 335096
rect 282656 335084 282684 335124
rect 300854 335084 300860 335096
rect 282656 335056 300860 335084
rect 300854 335044 300860 335056
rect 300912 335044 300918 335096
rect 208302 334976 208308 335028
rect 208360 335016 208366 335028
rect 245565 335019 245623 335025
rect 245565 335016 245577 335019
rect 208360 334988 245577 335016
rect 208360 334976 208366 334988
rect 245565 334985 245577 334988
rect 245611 334985 245623 335019
rect 245565 334979 245623 334985
rect 262122 334976 262128 335028
rect 262180 335016 262186 335028
rect 311894 335016 311900 335028
rect 262180 334988 311900 335016
rect 262180 334976 262186 334988
rect 311894 334976 311900 334988
rect 311952 334976 311958 335028
rect 212442 334908 212448 334960
rect 212500 334948 212506 334960
rect 251358 334948 251364 334960
rect 212500 334920 251364 334948
rect 212500 334908 212506 334920
rect 251358 334908 251364 334920
rect 251416 334908 251422 334960
rect 262306 334908 262312 334960
rect 262364 334948 262370 334960
rect 316034 334948 316040 334960
rect 262364 334920 316040 334948
rect 262364 334908 262370 334920
rect 316034 334908 316040 334920
rect 316092 334908 316098 334960
rect 169662 334840 169668 334892
rect 169720 334880 169726 334892
rect 247310 334880 247316 334892
rect 169720 334852 247316 334880
rect 169720 334840 169726 334852
rect 247310 334840 247316 334852
rect 247368 334840 247374 334892
rect 264422 334840 264428 334892
rect 264480 334880 264486 334892
rect 333974 334880 333980 334892
rect 264480 334852 333980 334880
rect 264480 334840 264486 334852
rect 333974 334840 333980 334852
rect 334032 334840 334038 334892
rect 160002 334772 160008 334824
rect 160060 334812 160066 334824
rect 246209 334815 246267 334821
rect 246209 334812 246221 334815
rect 160060 334784 246221 334812
rect 160060 334772 160066 334784
rect 246209 334781 246221 334784
rect 246255 334781 246267 334815
rect 246209 334775 246267 334781
rect 259914 334772 259920 334824
rect 259972 334812 259978 334824
rect 260190 334812 260196 334824
rect 259972 334784 260196 334812
rect 259972 334772 259978 334784
rect 260190 334772 260196 334784
rect 260248 334772 260254 334824
rect 274542 334772 274548 334824
rect 274600 334812 274606 334824
rect 422294 334812 422300 334824
rect 274600 334784 422300 334812
rect 274600 334772 274606 334784
rect 422294 334772 422300 334784
rect 422352 334772 422358 334824
rect 126882 334704 126888 334756
rect 126940 334744 126946 334756
rect 241146 334744 241152 334756
rect 126940 334716 241152 334744
rect 126940 334704 126946 334716
rect 241146 334704 241152 334716
rect 241204 334704 241210 334756
rect 289906 334704 289912 334756
rect 289964 334744 289970 334756
rect 500954 334744 500960 334756
rect 289964 334716 500960 334744
rect 289964 334704 289970 334716
rect 500954 334704 500960 334716
rect 501012 334704 501018 334756
rect 117222 334636 117228 334688
rect 117280 334676 117286 334688
rect 241974 334676 241980 334688
rect 117280 334648 241980 334676
rect 117280 334636 117286 334648
rect 241974 334636 241980 334648
rect 242032 334636 242038 334688
rect 285490 334636 285496 334688
rect 285548 334676 285554 334688
rect 528554 334676 528560 334688
rect 285548 334648 528560 334676
rect 285548 334636 285554 334648
rect 528554 334636 528560 334648
rect 528612 334636 528618 334688
rect 56502 334568 56508 334620
rect 56560 334608 56566 334620
rect 235626 334608 235632 334620
rect 56560 334580 235632 334608
rect 56560 334568 56566 334580
rect 235626 334568 235632 334580
rect 235684 334568 235690 334620
rect 289262 334568 289268 334620
rect 289320 334608 289326 334620
rect 574738 334608 574744 334620
rect 289320 334580 574744 334608
rect 289320 334568 289326 334580
rect 574738 334568 574744 334580
rect 574796 334568 574802 334620
rect 276198 334500 276204 334552
rect 276256 334540 276262 334552
rect 277118 334540 277124 334552
rect 276256 334512 277124 334540
rect 276256 334500 276262 334512
rect 277118 334500 277124 334512
rect 277176 334500 277182 334552
rect 229557 334203 229615 334209
rect 229557 334169 229569 334203
rect 229603 334200 229615 334203
rect 230290 334200 230296 334212
rect 229603 334172 230296 334200
rect 229603 334169 229615 334172
rect 229557 334163 229615 334169
rect 230290 334160 230296 334172
rect 230348 334160 230354 334212
rect 232130 334064 232136 334076
rect 232056 334036 232136 334064
rect 231670 333888 231676 333940
rect 231728 333888 231734 333940
rect 231688 333804 231716 333888
rect 232056 333872 232084 334036
rect 232130 334024 232136 334036
rect 232188 334024 232194 334076
rect 259454 334024 259460 334076
rect 259512 334064 259518 334076
rect 260374 334064 260380 334076
rect 259512 334036 260380 334064
rect 259512 334024 259518 334036
rect 260374 334024 260380 334036
rect 260432 334024 260438 334076
rect 232038 333820 232044 333872
rect 232096 333820 232102 333872
rect 231670 333752 231676 333804
rect 231728 333752 231734 333804
rect 239214 333752 239220 333804
rect 239272 333792 239278 333804
rect 239582 333792 239588 333804
rect 239272 333764 239588 333792
rect 239272 333752 239278 333764
rect 239582 333752 239588 333764
rect 239640 333752 239646 333804
rect 233602 333684 233608 333736
rect 233660 333724 233666 333736
rect 233878 333724 233884 333736
rect 233660 333696 233884 333724
rect 233660 333684 233666 333696
rect 233878 333684 233884 333696
rect 233936 333684 233942 333736
rect 236270 333684 236276 333736
rect 236328 333724 236334 333736
rect 236914 333724 236920 333736
rect 236328 333696 236920 333724
rect 236328 333684 236334 333696
rect 236914 333684 236920 333696
rect 236972 333684 236978 333736
rect 260558 333684 260564 333736
rect 260616 333724 260622 333736
rect 292574 333724 292580 333736
rect 260616 333696 292580 333724
rect 260616 333684 260622 333696
rect 292574 333684 292580 333696
rect 292632 333684 292638 333736
rect 219342 333616 219348 333668
rect 219400 333656 219406 333668
rect 252370 333656 252376 333668
rect 219400 333628 252376 333656
rect 219400 333616 219406 333628
rect 252370 333616 252376 333628
rect 252428 333616 252434 333668
rect 261478 333616 261484 333668
rect 261536 333656 261542 333668
rect 307754 333656 307760 333668
rect 261536 333628 307760 333656
rect 261536 333616 261542 333628
rect 307754 333616 307760 333628
rect 307812 333616 307818 333668
rect 184842 333548 184848 333600
rect 184900 333588 184906 333600
rect 248414 333588 248420 333600
rect 184900 333560 248420 333588
rect 184900 333548 184906 333560
rect 248414 333548 248420 333560
rect 248472 333548 248478 333600
rect 262950 333548 262956 333600
rect 263008 333588 263014 333600
rect 318794 333588 318800 333600
rect 263008 333560 318800 333588
rect 263008 333548 263014 333560
rect 318794 333548 318800 333560
rect 318852 333548 318858 333600
rect 173802 333480 173808 333532
rect 173860 333520 173866 333532
rect 247770 333520 247776 333532
rect 173860 333492 247776 333520
rect 173860 333480 173866 333492
rect 247770 333480 247776 333492
rect 247828 333480 247834 333532
rect 261202 333480 261208 333532
rect 261260 333520 261266 333532
rect 261478 333520 261484 333532
rect 261260 333492 261484 333520
rect 261260 333480 261266 333492
rect 261478 333480 261484 333492
rect 261536 333480 261542 333532
rect 266078 333480 266084 333532
rect 266136 333520 266142 333532
rect 342254 333520 342260 333532
rect 266136 333492 342260 333520
rect 266136 333480 266142 333492
rect 342254 333480 342260 333492
rect 342312 333480 342318 333532
rect 155862 333412 155868 333464
rect 155920 333452 155926 333464
rect 245286 333452 245292 333464
rect 155920 333424 245292 333452
rect 155920 333412 155926 333424
rect 245286 333412 245292 333424
rect 245344 333412 245350 333464
rect 271598 333412 271604 333464
rect 271656 333452 271662 333464
rect 404354 333452 404360 333464
rect 271656 333424 404360 333452
rect 271656 333412 271662 333424
rect 404354 333412 404360 333424
rect 404412 333412 404418 333464
rect 129642 333344 129648 333396
rect 129700 333384 129706 333396
rect 243170 333384 243176 333396
rect 129700 333356 243176 333384
rect 129700 333344 129706 333356
rect 243170 333344 243176 333356
rect 243228 333344 243234 333396
rect 278590 333344 278596 333396
rect 278648 333384 278654 333396
rect 465074 333384 465080 333396
rect 278648 333356 465080 333384
rect 278648 333344 278654 333356
rect 465074 333344 465080 333356
rect 465132 333344 465138 333396
rect 114462 333276 114468 333328
rect 114520 333316 114526 333328
rect 240226 333316 240232 333328
rect 114520 333288 240232 333316
rect 114520 333276 114526 333288
rect 240226 333276 240232 333288
rect 240284 333276 240290 333328
rect 241054 333276 241060 333328
rect 241112 333316 241118 333328
rect 241330 333316 241336 333328
rect 241112 333288 241336 333316
rect 241112 333276 241118 333288
rect 241330 333276 241336 333288
rect 241388 333276 241394 333328
rect 262858 333276 262864 333328
rect 262916 333316 262922 333328
rect 263410 333316 263416 333328
rect 262916 333288 263416 333316
rect 262916 333276 262922 333288
rect 263410 333276 263416 333288
rect 263468 333276 263474 333328
rect 283374 333276 283380 333328
rect 283432 333316 283438 333328
rect 518894 333316 518900 333328
rect 283432 333288 518900 333316
rect 283432 333276 283438 333288
rect 518894 333276 518900 333288
rect 518952 333276 518958 333328
rect 49602 333208 49608 333260
rect 49660 333248 49666 333260
rect 234982 333248 234988 333260
rect 49660 333220 234988 333248
rect 49660 333208 49666 333220
rect 234982 333208 234988 333220
rect 235040 333208 235046 333260
rect 238938 333208 238944 333260
rect 238996 333248 239002 333260
rect 239122 333248 239128 333260
rect 238996 333220 239128 333248
rect 238996 333208 239002 333220
rect 239122 333208 239128 333220
rect 239180 333208 239186 333260
rect 284018 333208 284024 333260
rect 284076 333248 284082 333260
rect 284938 333248 284944 333260
rect 284076 333220 284944 333248
rect 284076 333208 284082 333220
rect 284938 333208 284944 333220
rect 284996 333208 285002 333260
rect 286594 333208 286600 333260
rect 286652 333248 286658 333260
rect 546494 333248 546500 333260
rect 286652 333220 546500 333248
rect 286652 333208 286658 333220
rect 546494 333208 546500 333220
rect 546552 333208 546558 333260
rect 231578 333140 231584 333192
rect 231636 333180 231642 333192
rect 231762 333180 231768 333192
rect 231636 333152 231768 333180
rect 231636 333140 231642 333152
rect 231762 333140 231768 333152
rect 231820 333140 231826 333192
rect 232222 333140 232228 333192
rect 232280 333180 232286 333192
rect 233050 333180 233056 333192
rect 232280 333152 233056 333180
rect 232280 333140 232286 333152
rect 233050 333140 233056 333152
rect 233108 333140 233114 333192
rect 233878 333140 233884 333192
rect 233936 333180 233942 333192
rect 237558 333180 237564 333192
rect 233936 333152 237564 333180
rect 233936 333140 233942 333152
rect 237558 333140 237564 333152
rect 237616 333140 237622 333192
rect 278038 333180 278044 333192
rect 277964 333152 278044 333180
rect 277964 333124 277992 333152
rect 278038 333140 278044 333152
rect 278096 333140 278102 333192
rect 287422 333140 287428 333192
rect 287480 333180 287486 333192
rect 288158 333180 288164 333192
rect 287480 333152 288164 333180
rect 287480 333140 287486 333152
rect 288158 333140 288164 333152
rect 288216 333140 288222 333192
rect 234614 333072 234620 333124
rect 234672 333112 234678 333124
rect 234982 333112 234988 333124
rect 234672 333084 234988 333112
rect 234672 333072 234678 333084
rect 234982 333072 234988 333084
rect 235040 333072 235046 333124
rect 277946 333072 277952 333124
rect 278004 333072 278010 333124
rect 278038 333004 278044 333056
rect 278096 333044 278102 333056
rect 278406 333044 278412 333056
rect 278096 333016 278412 333044
rect 278096 333004 278102 333016
rect 278406 333004 278412 333016
rect 278464 333004 278470 333056
rect 235166 332936 235172 332988
rect 235224 332976 235230 332988
rect 235442 332976 235448 332988
rect 235224 332948 235448 332976
rect 235224 332936 235230 332948
rect 235442 332936 235448 332948
rect 235500 332936 235506 332988
rect 285858 332868 285864 332920
rect 285916 332908 285922 332920
rect 286778 332908 286784 332920
rect 285916 332880 286784 332908
rect 285916 332868 285922 332880
rect 286778 332868 286784 332880
rect 286836 332868 286842 332920
rect 234062 332392 234068 332444
rect 234120 332432 234126 332444
rect 234338 332432 234344 332444
rect 234120 332404 234344 332432
rect 234120 332392 234126 332404
rect 234338 332392 234344 332404
rect 234396 332392 234402 332444
rect 278774 332392 278780 332444
rect 278832 332432 278838 332444
rect 283377 332435 283435 332441
rect 283377 332432 283389 332435
rect 278832 332404 283389 332432
rect 278832 332392 278838 332404
rect 283377 332401 283389 332404
rect 283423 332401 283435 332435
rect 283377 332395 283435 332401
rect 260650 332324 260656 332376
rect 260708 332364 260714 332376
rect 296806 332364 296812 332376
rect 260708 332336 296812 332364
rect 260708 332324 260714 332336
rect 296806 332324 296812 332336
rect 296864 332324 296870 332376
rect 230382 332256 230388 332308
rect 230440 332296 230446 332308
rect 251726 332296 251732 332308
rect 230440 332268 251732 332296
rect 230440 332256 230446 332268
rect 251726 332256 251732 332268
rect 251784 332256 251790 332308
rect 261938 332256 261944 332308
rect 261996 332296 262002 332308
rect 313274 332296 313280 332308
rect 261996 332268 313280 332296
rect 261996 332256 262002 332268
rect 313274 332256 313280 332268
rect 313332 332256 313338 332308
rect 224862 332188 224868 332240
rect 224920 332228 224926 332240
rect 253014 332228 253020 332240
rect 224920 332200 253020 332228
rect 224920 332188 224926 332200
rect 253014 332188 253020 332200
rect 253072 332188 253078 332240
rect 271322 332188 271328 332240
rect 271380 332228 271386 332240
rect 331214 332228 331220 332240
rect 271380 332200 331220 332228
rect 271380 332188 271386 332200
rect 331214 332188 331220 332200
rect 331272 332188 331278 332240
rect 180702 332120 180708 332172
rect 180760 332160 180766 332172
rect 247034 332160 247040 332172
rect 180760 332132 247040 332160
rect 180760 332120 180766 332132
rect 247034 332120 247040 332132
rect 247092 332120 247098 332172
rect 267642 332120 267648 332172
rect 267700 332160 267706 332172
rect 356054 332160 356060 332172
rect 267700 332132 356060 332160
rect 267700 332120 267706 332132
rect 356054 332120 356060 332132
rect 356112 332120 356118 332172
rect 142062 332052 142068 332104
rect 142120 332092 142126 332104
rect 244274 332092 244280 332104
rect 142120 332064 244280 332092
rect 142120 332052 142126 332064
rect 244274 332052 244280 332064
rect 244332 332052 244338 332104
rect 283377 332095 283435 332101
rect 283377 332061 283389 332095
rect 283423 332092 283435 332095
rect 397454 332092 397460 332104
rect 283423 332064 397460 332092
rect 283423 332061 283435 332064
rect 283377 332055 283435 332061
rect 397454 332052 397460 332064
rect 397512 332052 397518 332104
rect 139302 331984 139308 332036
rect 139360 332024 139366 332036
rect 139360 331996 233924 332024
rect 139360 331984 139366 331996
rect 48222 331916 48228 331968
rect 48280 331956 48286 331968
rect 231946 331956 231952 331968
rect 48280 331928 231952 331956
rect 48280 331916 48286 331928
rect 231946 331916 231952 331928
rect 232004 331916 232010 331968
rect 233896 331956 233924 331996
rect 243354 331984 243360 332036
rect 243412 332024 243418 332036
rect 243630 332024 243636 332036
rect 243412 331996 243636 332024
rect 243412 331984 243418 331996
rect 243630 331984 243636 331996
rect 243688 331984 243694 332036
rect 273898 331984 273904 332036
rect 273956 332024 273962 332036
rect 433334 332024 433340 332036
rect 273956 331996 433340 332024
rect 273956 331984 273962 331996
rect 433334 331984 433340 331996
rect 433392 331984 433398 332036
rect 244182 331956 244188 331968
rect 233896 331928 244188 331956
rect 244182 331916 244188 331928
rect 244240 331916 244246 331968
rect 289170 331916 289176 331968
rect 289228 331956 289234 331968
rect 289722 331956 289728 331968
rect 289228 331928 289728 331956
rect 289228 331916 289234 331928
rect 289722 331916 289728 331928
rect 289780 331916 289786 331968
rect 289817 331959 289875 331965
rect 289817 331925 289829 331959
rect 289863 331956 289875 331959
rect 536834 331956 536840 331968
rect 289863 331928 536840 331956
rect 289863 331925 289875 331928
rect 289817 331919 289875 331925
rect 536834 331916 536840 331928
rect 536892 331916 536898 331968
rect 17218 331848 17224 331900
rect 17276 331888 17282 331900
rect 231302 331888 231308 331900
rect 17276 331860 231308 331888
rect 17276 331848 17282 331860
rect 231302 331848 231308 331860
rect 231360 331848 231366 331900
rect 244734 331848 244740 331900
rect 244792 331888 244798 331900
rect 245470 331888 245476 331900
rect 244792 331860 245476 331888
rect 244792 331848 244798 331860
rect 245470 331848 245476 331860
rect 245528 331848 245534 331900
rect 287790 331848 287796 331900
rect 287848 331888 287854 331900
rect 560938 331888 560944 331900
rect 287848 331860 560944 331888
rect 287848 331848 287854 331860
rect 560938 331848 560944 331860
rect 560996 331848 561002 331900
rect 285214 331780 285220 331832
rect 285272 331820 285278 331832
rect 289817 331823 289875 331829
rect 289817 331820 289829 331823
rect 285272 331792 289829 331820
rect 285272 331780 285278 331792
rect 289817 331789 289829 331792
rect 289863 331789 289875 331823
rect 289817 331783 289875 331789
rect 256421 331755 256479 331761
rect 256421 331721 256433 331755
rect 256467 331752 256479 331755
rect 256602 331752 256608 331764
rect 256467 331724 256608 331752
rect 256467 331721 256479 331724
rect 256421 331715 256479 331721
rect 256602 331712 256608 331724
rect 256660 331712 256666 331764
rect 243262 331304 243268 331356
rect 243320 331344 243326 331356
rect 243814 331344 243820 331356
rect 243320 331316 243820 331344
rect 243320 331304 243326 331316
rect 243814 331304 243820 331316
rect 243872 331304 243878 331356
rect 237006 331236 237012 331288
rect 237064 331276 237070 331288
rect 237282 331276 237288 331288
rect 237064 331248 237288 331276
rect 237064 331236 237070 331248
rect 237282 331236 237288 331248
rect 237340 331236 237346 331288
rect 239398 331236 239404 331288
rect 239456 331236 239462 331288
rect 240502 331236 240508 331288
rect 240560 331236 240566 331288
rect 268010 331236 268016 331288
rect 268068 331236 268074 331288
rect 239416 331208 239444 331236
rect 239582 331208 239588 331220
rect 239416 331180 239588 331208
rect 239582 331168 239588 331180
rect 239640 331168 239646 331220
rect 240520 331152 240548 331236
rect 268028 331208 268056 331236
rect 268470 331208 268476 331220
rect 268028 331180 268476 331208
rect 268470 331168 268476 331180
rect 268528 331168 268534 331220
rect 271049 331211 271107 331217
rect 271049 331177 271061 331211
rect 271095 331208 271107 331211
rect 272518 331208 272524 331220
rect 271095 331180 272524 331208
rect 271095 331177 271107 331180
rect 271049 331171 271107 331177
rect 272518 331168 272524 331180
rect 272576 331168 272582 331220
rect 240502 331100 240508 331152
rect 240560 331100 240566 331152
rect 274821 331143 274879 331149
rect 274821 331109 274833 331143
rect 274867 331140 274879 331143
rect 275738 331140 275744 331152
rect 274867 331112 275744 331140
rect 274867 331109 274879 331112
rect 274821 331103 274879 331109
rect 275738 331100 275744 331112
rect 275796 331100 275802 331152
rect 283190 331100 283196 331152
rect 283248 331140 283254 331152
rect 283834 331140 283840 331152
rect 283248 331112 283840 331140
rect 283248 331100 283254 331112
rect 283834 331100 283840 331112
rect 283892 331100 283898 331152
rect 262490 330896 262496 330948
rect 262548 330936 262554 330948
rect 320174 330936 320180 330948
rect 262548 330908 320180 330936
rect 262548 330896 262554 330908
rect 320174 330896 320180 330908
rect 320232 330896 320238 330948
rect 211062 330828 211068 330880
rect 211120 330868 211126 330880
rect 251545 330871 251603 330877
rect 251545 330868 251557 330871
rect 211120 330840 251557 330868
rect 211120 330828 211126 330840
rect 251545 330837 251557 330840
rect 251591 330837 251603 330871
rect 251545 330831 251603 330837
rect 263686 330828 263692 330880
rect 263744 330868 263750 330880
rect 328454 330868 328460 330880
rect 263744 330840 328460 330868
rect 263744 330828 263750 330840
rect 328454 330828 328460 330840
rect 328512 330828 328518 330880
rect 165522 330760 165528 330812
rect 165580 330800 165586 330812
rect 246850 330800 246856 330812
rect 165580 330772 246856 330800
rect 165580 330760 165586 330772
rect 246850 330760 246856 330772
rect 246908 330760 246914 330812
rect 269206 330760 269212 330812
rect 269264 330800 269270 330812
rect 382274 330800 382280 330812
rect 269264 330772 382280 330800
rect 269264 330760 269270 330772
rect 382274 330760 382280 330772
rect 382332 330760 382338 330812
rect 144822 330692 144828 330744
rect 144880 330732 144886 330744
rect 244458 330732 244464 330744
rect 144880 330704 244464 330732
rect 144880 330692 144886 330704
rect 244458 330692 244464 330704
rect 244516 330692 244522 330744
rect 273070 330692 273076 330744
rect 273128 330732 273134 330744
rect 411254 330732 411260 330744
rect 273128 330704 411260 330732
rect 273128 330692 273134 330704
rect 411254 330692 411260 330704
rect 411312 330692 411318 330744
rect 128262 330624 128268 330676
rect 128320 330664 128326 330676
rect 243081 330667 243139 330673
rect 243081 330664 243093 330667
rect 128320 330636 243093 330664
rect 128320 330624 128326 330636
rect 243081 330633 243093 330636
rect 243127 330633 243139 330667
rect 243081 330627 243139 330633
rect 276658 330624 276664 330676
rect 276716 330664 276722 330676
rect 451274 330664 451280 330676
rect 276716 330636 451280 330664
rect 276716 330624 276722 330636
rect 451274 330624 451280 330636
rect 451332 330624 451338 330676
rect 121362 330556 121368 330608
rect 121420 330596 121426 330608
rect 242342 330596 242348 330608
rect 121420 330568 242348 330596
rect 121420 330556 121426 330568
rect 242342 330556 242348 330568
rect 242400 330556 242406 330608
rect 270512 330568 284340 330596
rect 71682 330488 71688 330540
rect 71740 330528 71746 330540
rect 237190 330528 237196 330540
rect 71740 330500 237196 330528
rect 71740 330488 71746 330500
rect 237190 330488 237196 330500
rect 237248 330488 237254 330540
rect 259730 330420 259736 330472
rect 259788 330460 259794 330472
rect 270512 330460 270540 330568
rect 284312 330528 284340 330568
rect 285582 330556 285588 330608
rect 285640 330596 285646 330608
rect 539594 330596 539600 330608
rect 285640 330568 539600 330596
rect 285640 330556 285646 330568
rect 539594 330556 539600 330568
rect 539652 330556 539658 330608
rect 288434 330528 288440 330540
rect 284312 330500 288440 330528
rect 288434 330488 288440 330500
rect 288492 330488 288498 330540
rect 289630 330488 289636 330540
rect 289688 330528 289694 330540
rect 573358 330528 573364 330540
rect 289688 330500 573364 330528
rect 289688 330488 289694 330500
rect 573358 330488 573364 330500
rect 573416 330488 573422 330540
rect 259788 330432 270540 330460
rect 259788 330420 259794 330432
rect 279142 330012 279148 330064
rect 279200 330052 279206 330064
rect 279878 330052 279884 330064
rect 279200 330024 279884 330052
rect 279200 330012 279206 330024
rect 279878 330012 279884 330024
rect 279936 330012 279942 330064
rect 238110 329740 238116 329792
rect 238168 329780 238174 329792
rect 238386 329780 238392 329792
rect 238168 329752 238392 329780
rect 238168 329740 238174 329752
rect 238386 329740 238392 329752
rect 238444 329740 238450 329792
rect 226978 329468 226984 329520
rect 227036 329508 227042 329520
rect 230569 329511 230627 329517
rect 230569 329508 230581 329511
rect 227036 329480 230581 329508
rect 227036 329468 227042 329480
rect 230569 329477 230581 329480
rect 230615 329477 230627 329511
rect 230569 329471 230627 329477
rect 262030 329468 262036 329520
rect 262088 329508 262094 329520
rect 303614 329508 303620 329520
rect 262088 329480 303620 329508
rect 262088 329468 262094 329480
rect 303614 329468 303620 329480
rect 303672 329468 303678 329520
rect 264882 329400 264888 329452
rect 264940 329440 264946 329452
rect 338114 329440 338120 329452
rect 264940 329412 338120 329440
rect 264940 329400 264946 329412
rect 338114 329400 338120 329412
rect 338172 329400 338178 329452
rect 206922 329332 206928 329384
rect 206980 329372 206986 329384
rect 251174 329372 251180 329384
rect 206980 329344 251180 329372
rect 206980 329332 206986 329344
rect 251174 329332 251180 329344
rect 251232 329332 251238 329384
rect 267826 329332 267832 329384
rect 267884 329372 267890 329384
rect 367094 329372 367100 329384
rect 267884 329344 367100 329372
rect 267884 329332 267890 329344
rect 367094 329332 367100 329344
rect 367152 329332 367158 329384
rect 153102 329264 153108 329316
rect 153160 329304 153166 329316
rect 246022 329304 246028 329316
rect 153160 329276 246028 329304
rect 153160 329264 153166 329276
rect 246022 329264 246028 329276
rect 246080 329264 246086 329316
rect 276382 329304 276388 329316
rect 276343 329276 276388 329304
rect 276382 329264 276388 329276
rect 276440 329264 276446 329316
rect 280154 329264 280160 329316
rect 280212 329304 280218 329316
rect 393314 329304 393320 329316
rect 280212 329276 393320 329304
rect 280212 329264 280218 329276
rect 393314 329264 393320 329276
rect 393372 329264 393378 329316
rect 151722 329196 151728 329248
rect 151780 329236 151786 329248
rect 244734 329236 244740 329248
rect 151780 329208 244740 329236
rect 151780 329196 151786 329208
rect 244734 329196 244740 329208
rect 244792 329196 244798 329248
rect 272334 329196 272340 329248
rect 272392 329236 272398 329248
rect 415394 329236 415400 329248
rect 272392 329208 415400 329236
rect 272392 329196 272398 329208
rect 415394 329196 415400 329208
rect 415452 329196 415458 329248
rect 78582 329128 78588 329180
rect 78640 329168 78646 329180
rect 237926 329168 237932 329180
rect 78640 329140 237932 329168
rect 78640 329128 78646 329140
rect 237926 329128 237932 329140
rect 237984 329128 237990 329180
rect 268010 329128 268016 329180
rect 268068 329168 268074 329180
rect 269022 329168 269028 329180
rect 268068 329140 269028 329168
rect 268068 329128 268074 329140
rect 269022 329128 269028 329140
rect 269080 329128 269086 329180
rect 279050 329128 279056 329180
rect 279108 329168 279114 329180
rect 467834 329168 467840 329180
rect 279108 329140 467840 329168
rect 279108 329128 279114 329140
rect 467834 329128 467840 329140
rect 467892 329128 467898 329180
rect 34422 329060 34428 329112
rect 34480 329100 34486 329112
rect 233234 329100 233240 329112
rect 34480 329072 233240 329100
rect 34480 329060 34486 329072
rect 233234 329060 233240 329072
rect 233292 329060 233298 329112
rect 286870 329060 286876 329112
rect 286928 329100 286934 329112
rect 550634 329100 550640 329112
rect 286928 329072 550640 329100
rect 286928 329060 286934 329072
rect 550634 329060 550640 329072
rect 550692 329060 550698 329112
rect 249058 328992 249064 329044
rect 249116 329032 249122 329044
rect 249426 329032 249432 329044
rect 249116 329004 249432 329032
rect 249116 328992 249122 329004
rect 249426 328992 249432 329004
rect 249484 328992 249490 329044
rect 284386 328896 284392 328908
rect 284347 328868 284392 328896
rect 284386 328856 284392 328868
rect 284444 328856 284450 328908
rect 283650 328556 283656 328568
rect 283611 328528 283656 328556
rect 283650 328516 283656 328528
rect 283708 328516 283714 328568
rect 229554 328488 229560 328500
rect 229515 328460 229560 328488
rect 229554 328448 229560 328460
rect 229612 328448 229618 328500
rect 240686 328488 240692 328500
rect 240647 328460 240692 328488
rect 240686 328448 240692 328460
rect 240744 328448 240750 328500
rect 248693 328491 248751 328497
rect 248693 328457 248705 328491
rect 248739 328488 248751 328491
rect 249150 328488 249156 328500
rect 248739 328460 249156 328488
rect 248739 328457 248751 328460
rect 248693 328451 248751 328457
rect 249150 328448 249156 328460
rect 249208 328448 249214 328500
rect 267458 328488 267464 328500
rect 267419 328460 267464 328488
rect 267458 328448 267464 328460
rect 267516 328448 267522 328500
rect 231489 328423 231547 328429
rect 231489 328389 231501 328423
rect 231535 328420 231547 328423
rect 231578 328420 231584 328432
rect 231535 328392 231584 328420
rect 231535 328389 231547 328392
rect 231489 328383 231547 328389
rect 231578 328380 231584 328392
rect 231636 328380 231642 328432
rect 258534 328380 258540 328432
rect 258592 328420 258598 328432
rect 258626 328420 258632 328432
rect 258592 328392 258632 328420
rect 258592 328380 258598 328392
rect 258626 328380 258632 328392
rect 258684 328380 258690 328432
rect 284570 328420 284576 328432
rect 284531 328392 284576 328420
rect 284570 328380 284576 328392
rect 284628 328380 284634 328432
rect 261846 328040 261852 328092
rect 261904 328080 261910 328092
rect 299474 328080 299480 328092
rect 261904 328052 299480 328080
rect 261904 328040 261910 328052
rect 299474 328040 299480 328052
rect 299532 328040 299538 328092
rect 222102 327972 222108 328024
rect 222160 328012 222166 328024
rect 252738 328012 252744 328024
rect 222160 327984 252744 328012
rect 222160 327972 222166 327984
rect 252738 327972 252744 327984
rect 252796 327972 252802 328024
rect 283282 327972 283288 328024
rect 283340 328012 283346 328024
rect 400306 328012 400312 328024
rect 283340 327984 400312 328012
rect 283340 327972 283346 327984
rect 400306 327972 400312 327984
rect 400364 327972 400370 328024
rect 168282 327904 168288 327956
rect 168340 327944 168346 327956
rect 247126 327944 247132 327956
rect 168340 327916 247132 327944
rect 168340 327904 168346 327916
rect 247126 327904 247132 327916
rect 247184 327904 247190 327956
rect 273346 327904 273352 327956
rect 273404 327944 273410 327956
rect 425146 327944 425152 327956
rect 273404 327916 425152 327944
rect 273404 327904 273410 327916
rect 425146 327904 425152 327916
rect 425204 327904 425210 327956
rect 150342 327836 150348 327888
rect 150400 327876 150406 327888
rect 244366 327876 244372 327888
rect 150400 327848 244372 327876
rect 150400 327836 150406 327848
rect 244366 327836 244372 327848
rect 244424 327836 244430 327888
rect 277394 327836 277400 327888
rect 277452 327876 277458 327888
rect 462314 327876 462320 327888
rect 277452 327848 462320 327876
rect 277452 327836 277458 327848
rect 462314 327836 462320 327848
rect 462372 327836 462378 327888
rect 82722 327768 82728 327820
rect 82780 327808 82786 327820
rect 238294 327808 238300 327820
rect 82780 327780 238300 327808
rect 82780 327768 82786 327780
rect 238294 327768 238300 327780
rect 238352 327768 238358 327820
rect 282822 327768 282828 327820
rect 282880 327808 282886 327820
rect 502334 327808 502340 327820
rect 282880 327780 502340 327808
rect 282880 327768 282886 327780
rect 502334 327768 502340 327780
rect 502392 327768 502398 327820
rect 38562 327700 38568 327752
rect 38620 327740 38626 327752
rect 233510 327740 233516 327752
rect 38620 327712 233516 327740
rect 38620 327700 38626 327712
rect 233510 327700 233516 327712
rect 233568 327700 233574 327752
rect 290826 327700 290832 327752
rect 290884 327740 290890 327752
rect 557534 327740 557540 327752
rect 290884 327712 557540 327740
rect 290884 327700 290890 327712
rect 557534 327700 557540 327712
rect 557592 327700 557598 327752
rect 287609 327131 287667 327137
rect 287609 327097 287621 327131
rect 287655 327128 287667 327131
rect 288158 327128 288164 327140
rect 287655 327100 288164 327128
rect 287655 327097 287667 327100
rect 287609 327091 287667 327097
rect 288158 327088 288164 327100
rect 288216 327088 288222 327140
rect 233513 327063 233571 327069
rect 233513 327029 233525 327063
rect 233559 327060 233571 327063
rect 233602 327060 233608 327072
rect 233559 327032 233608 327060
rect 233559 327029 233571 327032
rect 233513 327023 233571 327029
rect 233602 327020 233608 327032
rect 233660 327020 233666 327072
rect 237561 327063 237619 327069
rect 237561 327029 237573 327063
rect 237607 327060 237619 327063
rect 237650 327060 237656 327072
rect 237607 327032 237656 327060
rect 237607 327029 237619 327032
rect 237561 327023 237619 327029
rect 237650 327020 237656 327032
rect 237708 327020 237714 327072
rect 274634 326748 274640 326800
rect 274692 326788 274698 326800
rect 279881 326791 279939 326797
rect 279881 326788 279893 326791
rect 274692 326760 279893 326788
rect 274692 326748 274698 326760
rect 279881 326757 279893 326760
rect 279927 326757 279939 326791
rect 279881 326751 279939 326757
rect 263226 326680 263232 326732
rect 263284 326720 263290 326732
rect 322934 326720 322940 326732
rect 263284 326692 322940 326720
rect 263284 326680 263290 326692
rect 322934 326680 322940 326692
rect 322992 326680 322998 326732
rect 226242 326612 226248 326664
rect 226300 326652 226306 326664
rect 253106 326652 253112 326664
rect 226300 326624 253112 326652
rect 226300 326612 226306 326624
rect 253106 326612 253112 326624
rect 253164 326612 253170 326664
rect 266630 326612 266636 326664
rect 266688 326652 266694 326664
rect 360194 326652 360200 326664
rect 266688 326624 360200 326652
rect 266688 326612 266694 326624
rect 360194 326612 360200 326624
rect 360252 326612 360258 326664
rect 171042 326544 171048 326596
rect 171100 326584 171106 326596
rect 247586 326584 247592 326596
rect 171100 326556 247592 326584
rect 171100 326544 171106 326556
rect 247586 326544 247592 326556
rect 247644 326544 247650 326596
rect 274726 326544 274732 326596
rect 274784 326584 274790 326596
rect 274784 326556 279832 326584
rect 274784 326544 274790 326556
rect 157242 326476 157248 326528
rect 157300 326516 157306 326528
rect 246666 326516 246672 326528
rect 157300 326488 246672 326516
rect 157300 326476 157306 326488
rect 246666 326476 246672 326488
rect 246724 326476 246730 326528
rect 96522 326408 96528 326460
rect 96580 326448 96586 326460
rect 238846 326448 238852 326460
rect 96580 326420 238852 326448
rect 96580 326408 96586 326420
rect 238846 326408 238852 326420
rect 238904 326408 238910 326460
rect 272518 326408 272524 326460
rect 272576 326408 272582 326460
rect 279602 326408 279608 326460
rect 279660 326448 279666 326460
rect 279804 326448 279832 326556
rect 280430 326544 280436 326596
rect 280488 326584 280494 326596
rect 408494 326584 408500 326596
rect 280488 326556 408500 326584
rect 280488 326544 280494 326556
rect 408494 326544 408500 326556
rect 408552 326544 408558 326596
rect 279881 326519 279939 326525
rect 279881 326485 279893 326519
rect 279927 326516 279939 326519
rect 433426 326516 433432 326528
rect 279927 326488 433432 326516
rect 279927 326485 279939 326488
rect 279881 326479 279939 326485
rect 433426 326476 433432 326488
rect 433484 326476 433490 326528
rect 443086 326448 443092 326460
rect 279660 326420 279740 326448
rect 279804 326420 443092 326448
rect 279660 326408 279666 326420
rect 53742 326340 53748 326392
rect 53800 326380 53806 326392
rect 235350 326380 235356 326392
rect 53800 326352 235356 326380
rect 53800 326340 53806 326352
rect 235350 326340 235356 326352
rect 235408 326340 235414 326392
rect 251266 326340 251272 326392
rect 251324 326380 251330 326392
rect 251726 326380 251732 326392
rect 251324 326352 251732 326380
rect 251324 326340 251330 326352
rect 251726 326340 251732 326352
rect 251784 326340 251790 326392
rect 252094 326340 252100 326392
rect 252152 326380 252158 326392
rect 252278 326380 252284 326392
rect 252152 326352 252284 326380
rect 252152 326340 252158 326352
rect 252278 326340 252284 326352
rect 252336 326340 252342 326392
rect 265894 326340 265900 326392
rect 265952 326380 265958 326392
rect 266078 326380 266084 326392
rect 265952 326352 266084 326380
rect 265952 326340 265958 326352
rect 266078 326340 266084 326352
rect 266136 326340 266142 326392
rect 272536 326256 272564 326408
rect 273254 326340 273260 326392
rect 273312 326380 273318 326392
rect 273714 326380 273720 326392
rect 273312 326352 273720 326380
rect 273312 326340 273318 326352
rect 273714 326340 273720 326352
rect 273772 326340 273778 326392
rect 273806 326340 273812 326392
rect 273864 326380 273870 326392
rect 274358 326380 274364 326392
rect 273864 326352 274364 326380
rect 273864 326340 273870 326352
rect 274358 326340 274364 326352
rect 274416 326340 274422 326392
rect 276290 326340 276296 326392
rect 276348 326380 276354 326392
rect 276934 326380 276940 326392
rect 276348 326352 276940 326380
rect 276348 326340 276354 326352
rect 276934 326340 276940 326352
rect 276992 326340 276998 326392
rect 279712 326256 279740 326420
rect 443086 326408 443092 326420
rect 443144 326408 443150 326460
rect 280338 326340 280344 326392
rect 280396 326380 280402 326392
rect 280982 326380 280988 326392
rect 280396 326352 280988 326380
rect 280396 326340 280402 326352
rect 280982 326340 280988 326352
rect 281040 326340 281046 326392
rect 281074 326340 281080 326392
rect 281132 326380 281138 326392
rect 281258 326380 281264 326392
rect 281132 326352 281264 326380
rect 281132 326340 281138 326352
rect 281258 326340 281264 326352
rect 281316 326340 281322 326392
rect 286686 326340 286692 326392
rect 286744 326380 286750 326392
rect 286962 326380 286968 326392
rect 286744 326352 286968 326380
rect 286744 326340 286750 326352
rect 286962 326340 286968 326352
rect 287020 326340 287026 326392
rect 288894 326340 288900 326392
rect 288952 326380 288958 326392
rect 289170 326380 289176 326392
rect 288952 326352 289176 326380
rect 288952 326340 288958 326352
rect 289170 326340 289176 326352
rect 289228 326340 289234 326392
rect 564434 326380 564440 326392
rect 289280 326352 564440 326380
rect 287422 326272 287428 326324
rect 287480 326312 287486 326324
rect 289280 326312 289308 326352
rect 564434 326340 564440 326352
rect 564492 326340 564498 326392
rect 287480 326284 289308 326312
rect 287480 326272 287486 326284
rect 265894 326204 265900 326256
rect 265952 326244 265958 326256
rect 266262 326244 266268 326256
rect 265952 326216 266268 326244
rect 265952 326204 265958 326216
rect 266262 326204 266268 326216
rect 266320 326204 266326 326256
rect 272518 326204 272524 326256
rect 272576 326204 272582 326256
rect 279694 326204 279700 326256
rect 279752 326204 279758 326256
rect 267921 325703 267979 325709
rect 267921 325669 267933 325703
rect 267967 325700 267979 325703
rect 269022 325700 269028 325712
rect 267967 325672 269028 325700
rect 267967 325669 267979 325672
rect 267921 325663 267979 325669
rect 269022 325660 269028 325672
rect 269080 325660 269086 325712
rect 269114 325660 269120 325712
rect 269172 325700 269178 325712
rect 269206 325700 269212 325712
rect 269172 325672 269212 325700
rect 269172 325660 269178 325672
rect 269206 325660 269212 325672
rect 269264 325660 269270 325712
rect 263778 325184 263784 325236
rect 263836 325224 263842 325236
rect 331306 325224 331312 325236
rect 263836 325196 331312 325224
rect 263836 325184 263842 325196
rect 331306 325184 331312 325196
rect 331364 325184 331370 325236
rect 213822 325116 213828 325168
rect 213880 325156 213886 325168
rect 251542 325156 251548 325168
rect 213880 325128 251548 325156
rect 213880 325116 213886 325128
rect 251542 325116 251548 325128
rect 251600 325116 251606 325168
rect 271230 325116 271236 325168
rect 271288 325156 271294 325168
rect 394694 325156 394700 325168
rect 271288 325128 394700 325156
rect 271288 325116 271294 325128
rect 394694 325116 394700 325128
rect 394752 325116 394758 325168
rect 141970 325048 141976 325100
rect 142028 325088 142034 325100
rect 244826 325088 244832 325100
rect 142028 325060 244832 325088
rect 142028 325048 142034 325060
rect 244826 325048 244832 325060
rect 244884 325048 244890 325100
rect 273622 325048 273628 325100
rect 273680 325088 273686 325100
rect 429194 325088 429200 325100
rect 273680 325060 429200 325088
rect 273680 325048 273686 325060
rect 429194 325048 429200 325060
rect 429252 325048 429258 325100
rect 92382 324980 92388 325032
rect 92440 325020 92446 325032
rect 239582 325020 239588 325032
rect 92440 324992 239588 325020
rect 92440 324980 92446 324992
rect 239582 324980 239588 324992
rect 239640 324980 239646 325032
rect 277854 324980 277860 325032
rect 277912 325020 277918 325032
rect 471974 325020 471980 325032
rect 277912 324992 471980 325020
rect 277912 324980 277918 324992
rect 471974 324980 471980 324992
rect 472032 324980 472038 325032
rect 42058 324912 42064 324964
rect 42116 324952 42122 324964
rect 233326 324952 233332 324964
rect 42116 324924 233332 324952
rect 42116 324912 42122 324924
rect 233326 324912 233332 324924
rect 233384 324912 233390 324964
rect 290734 324912 290740 324964
rect 290792 324952 290798 324964
rect 568574 324952 568580 324964
rect 290792 324924 568580 324952
rect 290792 324912 290798 324924
rect 568574 324912 568580 324924
rect 568632 324912 568638 324964
rect 284846 324232 284852 324284
rect 284904 324272 284910 324284
rect 285398 324272 285404 324284
rect 284904 324244 285404 324272
rect 284904 324232 284910 324244
rect 285398 324232 285404 324244
rect 285456 324232 285462 324284
rect 265158 323824 265164 323876
rect 265216 323864 265222 323876
rect 349154 323864 349160 323876
rect 265216 323836 349160 323864
rect 265216 323824 265222 323836
rect 349154 323824 349160 323836
rect 349212 323824 349218 323876
rect 217962 323756 217968 323808
rect 218020 323796 218026 323808
rect 251450 323796 251456 323808
rect 218020 323768 251456 323796
rect 218020 323756 218026 323768
rect 251450 323756 251456 323768
rect 251508 323756 251514 323808
rect 270954 323756 270960 323808
rect 271012 323796 271018 323808
rect 398834 323796 398840 323808
rect 271012 323768 398840 323796
rect 271012 323756 271018 323768
rect 398834 323756 398840 323768
rect 398892 323756 398898 323808
rect 159910 323688 159916 323740
rect 159968 323728 159974 323740
rect 245930 323728 245936 323740
rect 159968 323700 245936 323728
rect 159968 323688 159974 323700
rect 245930 323688 245936 323700
rect 245988 323688 245994 323740
rect 278958 323688 278964 323740
rect 279016 323728 279022 323740
rect 436094 323728 436100 323740
rect 279016 323700 436100 323728
rect 279016 323688 279022 323700
rect 436094 323688 436100 323700
rect 436152 323688 436158 323740
rect 99282 323620 99288 323672
rect 99340 323660 99346 323672
rect 240226 323660 240232 323672
rect 99340 323632 240232 323660
rect 99340 323620 99346 323632
rect 240226 323620 240232 323632
rect 240284 323620 240290 323672
rect 281810 323620 281816 323672
rect 281868 323660 281874 323672
rect 509234 323660 509240 323672
rect 281868 323632 509240 323660
rect 281868 323620 281874 323632
rect 509234 323620 509240 323632
rect 509292 323620 509298 323672
rect 46198 323552 46204 323604
rect 46256 323592 46262 323604
rect 234522 323592 234528 323604
rect 46256 323564 234528 323592
rect 46256 323552 46262 323564
rect 234522 323552 234528 323564
rect 234580 323552 234586 323604
rect 259362 323552 259368 323604
rect 259420 323592 259426 323604
rect 285674 323592 285680 323604
rect 259420 323564 285680 323592
rect 259420 323552 259426 323564
rect 285674 323552 285680 323564
rect 285732 323552 285738 323604
rect 290642 323552 290648 323604
rect 290700 323592 290706 323604
rect 571334 323592 571340 323604
rect 290700 323564 571340 323592
rect 290700 323552 290706 323564
rect 571334 323552 571340 323564
rect 571392 323552 571398 323604
rect 259178 323416 259184 323468
rect 259236 323456 259242 323468
rect 259362 323456 259368 323468
rect 259236 323428 259368 323456
rect 259236 323416 259242 323428
rect 259362 323416 259368 323428
rect 259420 323416 259426 323468
rect 260834 322464 260840 322516
rect 260892 322504 260898 322516
rect 306374 322504 306380 322516
rect 260892 322476 306380 322504
rect 260892 322464 260898 322476
rect 306374 322464 306380 322476
rect 306432 322464 306438 322516
rect 264514 322396 264520 322448
rect 264572 322436 264578 322448
rect 335354 322436 335360 322448
rect 264572 322408 335360 322436
rect 264572 322396 264578 322408
rect 335354 322396 335360 322408
rect 335412 322396 335418 322448
rect 146202 322328 146208 322380
rect 146260 322368 146266 322380
rect 244642 322368 244648 322380
rect 146260 322340 244648 322368
rect 146260 322328 146266 322340
rect 244642 322328 244648 322340
rect 244700 322328 244706 322380
rect 269666 322328 269672 322380
rect 269724 322368 269730 322380
rect 385034 322368 385040 322380
rect 269724 322340 385040 322368
rect 269724 322328 269730 322340
rect 385034 322328 385040 322340
rect 385092 322328 385098 322380
rect 103422 322260 103428 322312
rect 103480 322300 103486 322312
rect 241422 322300 241428 322312
rect 103480 322272 241428 322300
rect 103480 322260 103486 322272
rect 241422 322260 241428 322272
rect 241480 322260 241486 322312
rect 277302 322260 277308 322312
rect 277360 322300 277366 322312
rect 458174 322300 458180 322312
rect 277360 322272 458180 322300
rect 277360 322260 277366 322272
rect 458174 322260 458180 322272
rect 458232 322260 458238 322312
rect 56410 322192 56416 322244
rect 56468 322232 56474 322244
rect 235626 322232 235632 322244
rect 56468 322204 235632 322232
rect 56468 322192 56474 322204
rect 235626 322192 235632 322204
rect 235684 322192 235690 322244
rect 287146 322192 287152 322244
rect 287204 322232 287210 322244
rect 554866 322232 554872 322244
rect 287204 322204 554872 322232
rect 287204 322192 287210 322204
rect 554866 322192 554872 322204
rect 554924 322192 554930 322244
rect 289630 321716 289636 321768
rect 289688 321756 289694 321768
rect 298002 321756 298008 321768
rect 289688 321728 298008 321756
rect 289688 321716 289694 321728
rect 298002 321716 298008 321728
rect 298060 321716 298066 321768
rect 379422 321716 379428 321768
rect 379480 321756 379486 321768
rect 386322 321756 386328 321768
rect 379480 321728 386328 321756
rect 379480 321716 379486 321728
rect 386322 321716 386328 321728
rect 386380 321716 386386 321768
rect 287514 321580 287520 321632
rect 287572 321620 287578 321632
rect 287698 321620 287704 321632
rect 287572 321592 287704 321620
rect 287572 321580 287578 321592
rect 287698 321580 287704 321592
rect 287756 321580 287762 321632
rect 210970 321036 210976 321088
rect 211028 321076 211034 321088
rect 252278 321076 252284 321088
rect 211028 321048 252284 321076
rect 211028 321036 211034 321048
rect 252278 321036 252284 321048
rect 252336 321036 252342 321088
rect 272150 321036 272156 321088
rect 272208 321076 272214 321088
rect 418154 321076 418160 321088
rect 272208 321048 418160 321076
rect 272208 321036 272214 321048
rect 418154 321036 418160 321048
rect 418212 321036 418218 321088
rect 136542 320968 136548 321020
rect 136600 321008 136606 321020
rect 243906 321008 243912 321020
rect 136600 320980 243912 321008
rect 136600 320968 136606 320980
rect 243906 320968 243912 320980
rect 243964 320968 243970 321020
rect 278222 320968 278228 321020
rect 278280 321008 278286 321020
rect 466454 321008 466460 321020
rect 278280 320980 466460 321008
rect 278280 320968 278286 320980
rect 466454 320968 466460 320980
rect 466512 320968 466518 321020
rect 125410 320900 125416 320952
rect 125468 320940 125474 320952
rect 242526 320940 242532 320952
rect 125468 320912 242532 320940
rect 125468 320900 125474 320912
rect 242526 320900 242532 320912
rect 242584 320900 242590 320952
rect 279234 320900 279240 320952
rect 279292 320940 279298 320952
rect 476114 320940 476120 320952
rect 279292 320912 476120 320940
rect 279292 320900 279298 320912
rect 476114 320900 476120 320912
rect 476172 320900 476178 320952
rect 74442 320832 74448 320884
rect 74500 320872 74506 320884
rect 233878 320872 233884 320884
rect 74500 320844 233884 320872
rect 74500 320832 74506 320844
rect 233878 320832 233884 320844
rect 233936 320832 233942 320884
rect 286318 320832 286324 320884
rect 286376 320872 286382 320884
rect 540974 320872 540980 320884
rect 286376 320844 540980 320872
rect 286376 320832 286382 320844
rect 540974 320832 540980 320844
rect 541032 320832 541038 320884
rect 262582 319676 262588 319728
rect 262640 319716 262646 319728
rect 317414 319716 317420 319728
rect 262640 319688 317420 319716
rect 262640 319676 262646 319688
rect 317414 319676 317420 319688
rect 317472 319676 317478 319728
rect 215202 319608 215208 319660
rect 215260 319648 215266 319660
rect 251634 319648 251640 319660
rect 215260 319620 251640 319648
rect 215260 319608 215266 319620
rect 251634 319608 251640 319620
rect 251692 319608 251698 319660
rect 268194 319608 268200 319660
rect 268252 319648 268258 319660
rect 371234 319648 371240 319660
rect 268252 319620 371240 319648
rect 268252 319608 268258 319620
rect 371234 319608 371240 319620
rect 371292 319608 371298 319660
rect 154482 319540 154488 319592
rect 154540 319580 154546 319592
rect 246390 319580 246396 319592
rect 154540 319552 246396 319580
rect 154540 319540 154546 319552
rect 246390 319540 246396 319552
rect 246448 319540 246454 319592
rect 283466 319540 283472 319592
rect 283524 319580 283530 319592
rect 447134 319580 447140 319592
rect 283524 319552 447140 319580
rect 283524 319540 283530 319552
rect 447134 319540 447140 319552
rect 447192 319540 447198 319592
rect 67542 319472 67548 319524
rect 67600 319512 67606 319524
rect 229738 319512 229744 319524
rect 67600 319484 229744 319512
rect 67600 319472 67606 319484
rect 229738 319472 229744 319484
rect 229796 319472 229802 319524
rect 238938 319512 238944 319524
rect 238899 319484 238944 319512
rect 238938 319472 238944 319484
rect 238996 319472 239002 319524
rect 280706 319472 280712 319524
rect 280764 319512 280770 319524
rect 487154 319512 487160 319524
rect 280764 319484 487160 319512
rect 280764 319472 280770 319484
rect 487154 319472 487160 319484
rect 487212 319472 487218 319524
rect 50338 319404 50344 319456
rect 50396 319444 50402 319456
rect 234982 319444 234988 319456
rect 50396 319416 234988 319444
rect 50396 319404 50402 319416
rect 234982 319404 234988 319416
rect 235040 319404 235046 319456
rect 261570 319404 261576 319456
rect 261628 319444 261634 319456
rect 278774 319444 278780 319456
rect 261628 319416 278780 319444
rect 261628 319404 261634 319416
rect 278774 319404 278780 319416
rect 278832 319404 278838 319456
rect 287974 319404 287980 319456
rect 288032 319444 288038 319456
rect 556798 319444 556804 319456
rect 288032 319416 556804 319444
rect 288032 319404 288038 319416
rect 556798 319404 556804 319416
rect 556856 319404 556862 319456
rect 231486 318832 231492 318844
rect 231447 318804 231492 318832
rect 231486 318792 231492 318804
rect 231544 318792 231550 318844
rect 243354 318792 243360 318844
rect 243412 318832 243418 318844
rect 243538 318832 243544 318844
rect 243412 318804 243544 318832
rect 243412 318792 243418 318804
rect 243538 318792 243544 318804
rect 243596 318792 243602 318844
rect 254026 318792 254032 318844
rect 254084 318832 254090 318844
rect 254118 318832 254124 318844
rect 254084 318804 254124 318832
rect 254084 318792 254090 318804
rect 254118 318792 254124 318804
rect 254176 318792 254182 318844
rect 265342 318792 265348 318844
rect 265400 318832 265406 318844
rect 265526 318832 265532 318844
rect 265400 318804 265532 318832
rect 265400 318792 265406 318804
rect 265526 318792 265532 318804
rect 265584 318792 265590 318844
rect 283006 318792 283012 318844
rect 283064 318832 283070 318844
rect 283374 318832 283380 318844
rect 283064 318804 283380 318832
rect 283064 318792 283070 318804
rect 283374 318792 283380 318804
rect 283432 318792 283438 318844
rect 284570 318832 284576 318844
rect 284531 318804 284576 318832
rect 284570 318792 284576 318804
rect 284628 318792 284634 318844
rect 229465 318767 229523 318773
rect 229465 318733 229477 318767
rect 229511 318764 229523 318767
rect 229554 318764 229560 318776
rect 229511 318736 229560 318764
rect 229511 318733 229523 318736
rect 229465 318727 229523 318733
rect 229554 318724 229560 318736
rect 229612 318724 229618 318776
rect 249150 318764 249156 318776
rect 249111 318736 249156 318764
rect 249150 318724 249156 318736
rect 249208 318724 249214 318776
rect 269022 318656 269028 318708
rect 269080 318696 269086 318708
rect 269206 318696 269212 318708
rect 269080 318668 269212 318696
rect 269080 318656 269086 318668
rect 269206 318656 269212 318668
rect 269264 318656 269270 318708
rect 262398 318248 262404 318300
rect 262456 318288 262462 318300
rect 321554 318288 321560 318300
rect 262456 318260 321560 318288
rect 262456 318248 262462 318260
rect 321554 318248 321560 318260
rect 321612 318248 321618 318300
rect 276750 318180 276756 318232
rect 276808 318220 276814 318232
rect 454034 318220 454040 318232
rect 276808 318192 454040 318220
rect 276808 318180 276814 318192
rect 454034 318180 454040 318192
rect 454092 318180 454098 318232
rect 140682 318112 140688 318164
rect 140740 318152 140746 318164
rect 244550 318152 244556 318164
rect 140740 318124 244556 318152
rect 140740 318112 140746 318124
rect 244550 318112 244556 318124
rect 244608 318112 244614 318164
rect 281718 318112 281724 318164
rect 281776 318152 281782 318164
rect 505094 318152 505100 318164
rect 281776 318124 505100 318152
rect 281776 318112 281782 318124
rect 505094 318112 505100 318124
rect 505152 318112 505158 318164
rect 85482 318044 85488 318096
rect 85540 318084 85546 318096
rect 238662 318084 238668 318096
rect 85540 318056 238668 318084
rect 85540 318044 85546 318056
rect 238662 318044 238668 318056
rect 238720 318044 238726 318096
rect 258994 318044 259000 318096
rect 259052 318084 259058 318096
rect 281534 318084 281540 318096
rect 259052 318056 281540 318084
rect 259052 318044 259058 318056
rect 281534 318044 281540 318056
rect 281592 318044 281598 318096
rect 289262 318044 289268 318096
rect 289320 318084 289326 318096
rect 567838 318084 567844 318096
rect 289320 318056 567844 318084
rect 289320 318044 289326 318056
rect 567838 318044 567844 318056
rect 567896 318044 567902 318096
rect 233510 317472 233516 317484
rect 233471 317444 233516 317472
rect 233510 317432 233516 317444
rect 233568 317432 233574 317484
rect 237558 317472 237564 317484
rect 237519 317444 237564 317472
rect 237558 317432 237564 317444
rect 237616 317432 237622 317484
rect 238938 317472 238944 317484
rect 238899 317444 238944 317472
rect 238938 317432 238944 317444
rect 238996 317432 239002 317484
rect 272426 317432 272432 317484
rect 272484 317472 272490 317484
rect 272610 317472 272616 317484
rect 272484 317444 272616 317472
rect 272484 317432 272490 317444
rect 272610 317432 272616 317444
rect 272668 317432 272674 317484
rect 277854 317432 277860 317484
rect 277912 317472 277918 317484
rect 277946 317472 277952 317484
rect 277912 317444 277952 317472
rect 277912 317432 277918 317444
rect 277946 317432 277952 317444
rect 278004 317432 278010 317484
rect 283742 317404 283748 317416
rect 283703 317376 283748 317404
rect 283742 317364 283748 317376
rect 283800 317364 283806 317416
rect 288158 317404 288164 317416
rect 288119 317376 288164 317404
rect 288158 317364 288164 317376
rect 288216 317364 288222 317416
rect 267182 316888 267188 316940
rect 267240 316928 267246 316940
rect 364334 316928 364340 316940
rect 267240 316900 364340 316928
rect 267240 316888 267246 316900
rect 364334 316888 364340 316900
rect 364392 316888 364398 316940
rect 271690 316820 271696 316872
rect 271748 316860 271754 316872
rect 405734 316860 405740 316872
rect 271748 316832 405740 316860
rect 271748 316820 271754 316832
rect 405734 316820 405740 316832
rect 405792 316820 405798 316872
rect 143442 316752 143448 316804
rect 143500 316792 143506 316804
rect 245102 316792 245108 316804
rect 143500 316764 245108 316792
rect 143500 316752 143506 316764
rect 245102 316752 245108 316764
rect 245160 316752 245166 316804
rect 280614 316752 280620 316804
rect 280672 316792 280678 316804
rect 460934 316792 460940 316804
rect 280672 316764 460940 316792
rect 280672 316752 280678 316764
rect 460934 316752 460940 316764
rect 460992 316752 460998 316804
rect 107470 316684 107476 316736
rect 107528 316724 107534 316736
rect 240686 316724 240692 316736
rect 107528 316696 240692 316724
rect 107528 316684 107534 316696
rect 240686 316684 240692 316696
rect 240744 316684 240750 316736
rect 257154 316684 257160 316736
rect 257212 316724 257218 316736
rect 270494 316724 270500 316736
rect 257212 316696 270500 316724
rect 257212 316684 257218 316696
rect 270494 316684 270500 316696
rect 270552 316684 270558 316736
rect 283834 316684 283840 316736
rect 283892 316724 283898 316736
rect 516134 316724 516140 316736
rect 283892 316696 516140 316724
rect 283892 316684 283898 316696
rect 516134 316684 516140 316696
rect 516192 316684 516198 316736
rect 256418 316004 256424 316056
rect 256476 316044 256482 316056
rect 256602 316044 256608 316056
rect 256476 316016 256608 316044
rect 256476 316004 256482 316016
rect 256602 316004 256608 316016
rect 256660 316004 256666 316056
rect 268286 315460 268292 315512
rect 268344 315500 268350 315512
rect 373994 315500 374000 315512
rect 268344 315472 374000 315500
rect 268344 315460 268350 315472
rect 373994 315460 374000 315472
rect 374052 315460 374058 315512
rect 272058 315392 272064 315444
rect 272116 315432 272122 315444
rect 408586 315432 408592 315444
rect 272116 315404 408592 315432
rect 272116 315392 272122 315404
rect 408586 315392 408592 315404
rect 408644 315392 408650 315444
rect 147582 315324 147588 315376
rect 147640 315364 147646 315376
rect 245562 315364 245568 315376
rect 147640 315336 245568 315364
rect 147640 315324 147646 315336
rect 245562 315324 245568 315336
rect 245620 315324 245626 315376
rect 279786 315324 279792 315376
rect 279844 315364 279850 315376
rect 478874 315364 478880 315376
rect 279844 315336 478880 315364
rect 279844 315324 279850 315336
rect 478874 315324 478880 315336
rect 478932 315324 478938 315376
rect 19978 315256 19984 315308
rect 20036 315296 20042 315308
rect 231578 315296 231584 315308
rect 20036 315268 231584 315296
rect 20036 315256 20042 315268
rect 231578 315256 231584 315268
rect 231636 315256 231642 315308
rect 284294 315256 284300 315308
rect 284352 315296 284358 315308
rect 529934 315296 529940 315308
rect 284352 315268 529940 315296
rect 284352 315256 284358 315268
rect 529934 315256 529940 315268
rect 529992 315256 529998 315308
rect 269850 314100 269856 314152
rect 269908 314140 269914 314152
rect 389174 314140 389180 314152
rect 269908 314112 389180 314140
rect 269908 314100 269914 314112
rect 389174 314100 389180 314112
rect 389232 314100 389238 314152
rect 273530 314032 273536 314084
rect 273588 314072 273594 314084
rect 423674 314072 423680 314084
rect 273588 314044 423680 314072
rect 273588 314032 273594 314044
rect 423674 314032 423680 314044
rect 423732 314032 423738 314084
rect 158622 313964 158628 314016
rect 158680 314004 158686 314016
rect 246114 314004 246120 314016
rect 158680 313976 246120 314004
rect 158680 313964 158686 313976
rect 246114 313964 246120 313976
rect 246172 313964 246178 314016
rect 279510 313964 279516 314016
rect 279568 314004 279574 314016
rect 484394 314004 484400 314016
rect 279568 313976 484400 314004
rect 279568 313964 279574 313976
rect 484394 313964 484400 313976
rect 484452 313964 484458 314016
rect 24118 313896 24124 313948
rect 24176 313936 24182 313948
rect 232406 313936 232412 313948
rect 24176 313908 232412 313936
rect 24176 313896 24182 313908
rect 232406 313896 232412 313908
rect 232464 313896 232470 313948
rect 286686 313896 286692 313948
rect 286744 313936 286750 313948
rect 545114 313936 545120 313948
rect 286744 313908 545120 313936
rect 286744 313896 286750 313908
rect 545114 313896 545120 313908
rect 545172 313896 545178 313948
rect 275370 312672 275376 312724
rect 275428 312712 275434 312724
rect 437474 312712 437480 312724
rect 275428 312684 437480 312712
rect 275428 312672 275434 312684
rect 437474 312672 437480 312684
rect 437532 312672 437538 312724
rect 161382 312604 161388 312656
rect 161440 312644 161446 312656
rect 246298 312644 246304 312656
rect 161440 312616 246304 312644
rect 161440 312604 161446 312616
rect 246298 312604 246304 312616
rect 246356 312604 246362 312656
rect 280890 312604 280896 312656
rect 280948 312644 280954 312656
rect 491294 312644 491300 312656
rect 280948 312616 491300 312644
rect 280948 312604 280954 312616
rect 491294 312604 491300 312616
rect 491352 312604 491358 312656
rect 31662 312536 31668 312588
rect 31720 312576 31726 312588
rect 233142 312576 233148 312588
rect 31720 312548 233148 312576
rect 31720 312536 31726 312548
rect 233142 312536 233148 312548
rect 233200 312536 233206 312588
rect 286594 312536 286600 312588
rect 286652 312576 286658 312588
rect 552014 312576 552020 312588
rect 286652 312548 552020 312576
rect 286652 312536 286658 312548
rect 552014 312536 552020 312548
rect 552072 312536 552078 312588
rect 288986 311788 288992 311840
rect 289044 311828 289050 311840
rect 289262 311828 289268 311840
rect 289044 311800 289268 311828
rect 289044 311788 289050 311800
rect 289262 311788 289268 311800
rect 289320 311788 289326 311840
rect 271414 311176 271420 311228
rect 271472 311216 271478 311228
rect 401594 311216 401600 311228
rect 271472 311188 401600 311216
rect 271472 311176 271478 311188
rect 401594 311176 401600 311188
rect 401652 311176 401658 311228
rect 110322 311108 110328 311160
rect 110380 311148 110386 311160
rect 241146 311148 241152 311160
rect 110380 311120 241152 311148
rect 110380 311108 110386 311120
rect 241146 311108 241152 311120
rect 241204 311108 241210 311160
rect 274910 311108 274916 311160
rect 274968 311148 274974 311160
rect 441614 311148 441620 311160
rect 274968 311120 441620 311148
rect 274968 311108 274974 311120
rect 441614 311108 441620 311120
rect 441672 311108 441678 311160
rect 299566 310768 299572 310820
rect 299624 310808 299630 310820
rect 304350 310808 304356 310820
rect 299624 310780 304356 310808
rect 299624 310768 299630 310780
rect 304350 310768 304356 310780
rect 304408 310768 304414 310820
rect 320726 310768 320732 310820
rect 320784 310808 320790 310820
rect 328362 310808 328368 310820
rect 320784 310780 328368 310808
rect 320784 310768 320790 310780
rect 328362 310768 328368 310780
rect 328420 310768 328426 310820
rect 359642 310768 359648 310820
rect 359700 310808 359706 310820
rect 367002 310808 367008 310820
rect 359700 310780 367008 310808
rect 359700 310768 359706 310780
rect 367002 310768 367008 310780
rect 367060 310768 367066 310820
rect 475562 310768 475568 310820
rect 475620 310808 475626 310820
rect 482922 310808 482928 310820
rect 475620 310780 482928 310808
rect 475620 310768 475626 310780
rect 482922 310768 482928 310780
rect 482980 310768 482986 310820
rect 541066 310768 541072 310820
rect 541124 310808 541130 310820
rect 543826 310808 543832 310820
rect 541124 310780 543832 310808
rect 541124 310768 541130 310780
rect 543826 310768 543832 310780
rect 543884 310768 543890 310820
rect 288342 310700 288348 310752
rect 288400 310740 288406 310752
rect 296622 310740 296628 310752
rect 288400 310712 296628 310740
rect 288400 310700 288406 310712
rect 296622 310700 296628 310712
rect 296680 310700 296686 310752
rect 340782 310700 340788 310752
rect 340840 310740 340846 310752
rect 347682 310740 347688 310752
rect 340840 310712 347688 310740
rect 340840 310700 340846 310712
rect 347682 310700 347688 310712
rect 347740 310700 347746 310752
rect 379422 310700 379428 310752
rect 379480 310740 379486 310752
rect 386322 310740 386328 310752
rect 379480 310712 386328 310740
rect 379480 310700 379486 310712
rect 386322 310700 386328 310712
rect 386380 310700 386386 310752
rect 398742 310700 398748 310752
rect 398800 310740 398806 310752
rect 405642 310740 405648 310752
rect 398800 310712 405648 310740
rect 398800 310700 398806 310712
rect 405642 310700 405648 310712
rect 405700 310700 405706 310752
rect 418062 310700 418068 310752
rect 418120 310740 418126 310752
rect 424962 310740 424968 310752
rect 418120 310712 424968 310740
rect 418120 310700 418126 310712
rect 424962 310700 424968 310712
rect 425020 310700 425026 310752
rect 437382 310700 437388 310752
rect 437440 310740 437446 310752
rect 444282 310740 444288 310752
rect 437440 310712 444288 310740
rect 437440 310700 437446 310712
rect 444282 310700 444288 310712
rect 444340 310700 444346 310752
rect 456702 310700 456708 310752
rect 456760 310740 456766 310752
rect 463602 310740 463608 310752
rect 456760 310712 463608 310740
rect 456760 310700 456766 310712
rect 463602 310700 463608 310712
rect 463660 310700 463666 310752
rect 495342 310700 495348 310752
rect 495400 310740 495406 310752
rect 502242 310740 502248 310752
rect 495400 310712 502248 310740
rect 495400 310700 495406 310712
rect 502242 310700 502248 310712
rect 502300 310700 502306 310752
rect 514662 310700 514668 310752
rect 514720 310740 514726 310752
rect 521562 310740 521568 310752
rect 514720 310712 521568 310740
rect 514720 310700 514726 310712
rect 521562 310700 521568 310712
rect 521620 310700 521626 310752
rect 533982 310700 533988 310752
rect 534040 310740 534046 310752
rect 540882 310740 540888 310752
rect 534040 310712 540888 310740
rect 534040 310700 534046 310712
rect 540882 310700 540888 310712
rect 540940 310700 540946 310752
rect 261018 309952 261024 310004
rect 261076 309992 261082 310004
rect 310514 309992 310520 310004
rect 261076 309964 310520 309992
rect 261076 309952 261082 309964
rect 310514 309952 310520 309964
rect 310572 309952 310578 310004
rect 268654 309884 268660 309936
rect 268712 309924 268718 309936
rect 378134 309924 378140 309936
rect 268712 309896 378140 309924
rect 268712 309884 268718 309896
rect 378134 309884 378140 309896
rect 378192 309884 378198 309936
rect 280982 309816 280988 309868
rect 281040 309856 281046 309868
rect 494054 309856 494060 309868
rect 281040 309828 494060 309856
rect 281040 309816 281046 309828
rect 494054 309816 494060 309828
rect 494112 309816 494118 309868
rect 31018 309748 31024 309800
rect 31076 309788 31082 309800
rect 232314 309788 232320 309800
rect 31076 309760 232320 309788
rect 31076 309748 31082 309760
rect 232314 309748 232320 309760
rect 232372 309748 232378 309800
rect 287882 309748 287888 309800
rect 287940 309788 287946 309800
rect 563054 309788 563060 309800
rect 287940 309760 563060 309788
rect 287940 309748 287946 309760
rect 563054 309748 563060 309760
rect 563112 309748 563118 309800
rect 229462 309244 229468 309256
rect 229423 309216 229468 309244
rect 229462 309204 229468 309216
rect 229520 309204 229526 309256
rect 243354 309136 243360 309188
rect 243412 309176 243418 309188
rect 243538 309176 243544 309188
rect 243412 309148 243544 309176
rect 243412 309136 243418 309148
rect 243538 309136 243544 309148
rect 243596 309136 243602 309188
rect 249150 309176 249156 309188
rect 249111 309148 249156 309176
rect 249150 309136 249156 309148
rect 249208 309136 249214 309188
rect 3326 309068 3332 309120
rect 3384 309108 3390 309120
rect 213178 309108 213184 309120
rect 3384 309080 213184 309108
rect 3384 309068 3390 309080
rect 213178 309068 213184 309080
rect 213236 309068 213242 309120
rect 229462 309108 229468 309120
rect 229423 309080 229468 309108
rect 229462 309068 229468 309080
rect 229520 309068 229526 309120
rect 233510 309108 233516 309120
rect 233471 309080 233516 309108
rect 233510 309068 233516 309080
rect 233568 309068 233574 309120
rect 237558 309068 237564 309120
rect 237616 309068 237622 309120
rect 238938 309108 238944 309120
rect 238899 309080 238944 309108
rect 238938 309068 238944 309080
rect 238996 309068 239002 309120
rect 284662 309108 284668 309120
rect 284623 309080 284668 309108
rect 284662 309068 284668 309080
rect 284720 309068 284726 309120
rect 289170 309068 289176 309120
rect 289228 309108 289234 309120
rect 289262 309108 289268 309120
rect 289228 309080 289268 309108
rect 289228 309068 289234 309080
rect 289262 309068 289268 309080
rect 289320 309068 289326 309120
rect 237576 309040 237604 309068
rect 237650 309040 237656 309052
rect 237576 309012 237656 309040
rect 237650 309000 237656 309012
rect 237708 309000 237714 309052
rect 283006 309040 283012 309052
rect 282967 309012 283012 309040
rect 283006 309000 283012 309012
rect 283064 309000 283070 309052
rect 263962 308524 263968 308576
rect 264020 308564 264026 308576
rect 339494 308564 339500 308576
rect 264020 308536 339500 308564
rect 264020 308524 264026 308536
rect 339494 308524 339500 308536
rect 339552 308524 339558 308576
rect 281074 308456 281080 308508
rect 281132 308496 281138 308508
rect 498194 308496 498200 308508
rect 281132 308468 498200 308496
rect 281132 308456 281138 308468
rect 498194 308456 498200 308468
rect 498252 308456 498258 308508
rect 289354 308388 289360 308440
rect 289412 308428 289418 308440
rect 574830 308428 574836 308440
rect 289412 308400 574836 308428
rect 289412 308388 289418 308400
rect 574830 308388 574836 308400
rect 574888 308388 574894 308440
rect 278038 307776 278044 307828
rect 278096 307816 278102 307828
rect 278130 307816 278136 307828
rect 278096 307788 278136 307816
rect 278096 307776 278102 307788
rect 278130 307776 278136 307788
rect 278188 307776 278194 307828
rect 288158 307816 288164 307828
rect 288119 307788 288164 307816
rect 288158 307776 288164 307788
rect 288216 307776 288222 307828
rect 251729 307751 251787 307757
rect 251729 307717 251741 307751
rect 251775 307748 251787 307751
rect 251818 307748 251824 307760
rect 251775 307720 251824 307748
rect 251775 307717 251787 307720
rect 251729 307711 251787 307717
rect 251818 307708 251824 307720
rect 251876 307708 251882 307760
rect 260190 307748 260196 307760
rect 260151 307720 260196 307748
rect 260190 307708 260196 307720
rect 260248 307708 260254 307760
rect 260374 307708 260380 307760
rect 260432 307748 260438 307760
rect 260558 307748 260564 307760
rect 260432 307720 260564 307748
rect 260432 307708 260438 307720
rect 260558 307708 260564 307720
rect 260616 307708 260622 307760
rect 272702 307164 272708 307216
rect 272760 307204 272766 307216
rect 412634 307204 412640 307216
rect 272760 307176 412640 307204
rect 272760 307164 272766 307176
rect 412634 307164 412640 307176
rect 412692 307164 412698 307216
rect 277486 307096 277492 307148
rect 277544 307136 277550 307148
rect 473354 307136 473360 307148
rect 277544 307108 473360 307136
rect 277544 307096 277550 307108
rect 473354 307096 473360 307108
rect 473412 307096 473418 307148
rect 43438 307028 43444 307080
rect 43496 307068 43502 307080
rect 233694 307068 233700 307080
rect 43496 307040 233700 307068
rect 43496 307028 43502 307040
rect 233694 307028 233700 307040
rect 233752 307028 233758 307080
rect 282730 307028 282736 307080
rect 282788 307068 282794 307080
rect 511994 307068 512000 307080
rect 282788 307040 512000 307068
rect 282788 307028 282794 307040
rect 511994 307028 512000 307040
rect 512052 307028 512058 307080
rect 256418 306348 256424 306400
rect 256476 306388 256482 306400
rect 256694 306388 256700 306400
rect 256476 306360 256700 306388
rect 256476 306348 256482 306360
rect 256694 306348 256700 306360
rect 256752 306348 256758 306400
rect 272794 305668 272800 305720
rect 272852 305708 272858 305720
rect 416866 305708 416872 305720
rect 272852 305680 416872 305708
rect 272852 305668 272858 305680
rect 416866 305668 416872 305680
rect 416924 305668 416930 305720
rect 38470 305600 38476 305652
rect 38528 305640 38534 305652
rect 233513 305643 233571 305649
rect 233513 305640 233525 305643
rect 38528 305612 233525 305640
rect 38528 305600 38534 305612
rect 233513 305609 233525 305612
rect 233559 305609 233571 305643
rect 233513 305603 233571 305609
rect 282914 305600 282920 305652
rect 282972 305640 282978 305652
rect 520274 305640 520280 305652
rect 282972 305612 520280 305640
rect 282972 305600 282978 305612
rect 520274 305600 520280 305612
rect 520332 305600 520338 305652
rect 275186 304988 275192 305040
rect 275244 305028 275250 305040
rect 275278 305028 275284 305040
rect 275244 305000 275284 305028
rect 275244 304988 275250 305000
rect 275278 304988 275284 305000
rect 275336 304988 275342 305040
rect 277854 304920 277860 304972
rect 277912 304960 277918 304972
rect 278222 304960 278228 304972
rect 277912 304932 278228 304960
rect 277912 304920 277918 304932
rect 278222 304920 278228 304932
rect 278280 304920 278286 304972
rect 274082 304308 274088 304360
rect 274140 304348 274146 304360
rect 426434 304348 426440 304360
rect 274140 304320 426440 304348
rect 274140 304308 274146 304320
rect 426434 304308 426440 304320
rect 426492 304308 426498 304360
rect 42702 304240 42708 304292
rect 42760 304280 42766 304292
rect 234246 304280 234252 304292
rect 42760 304252 234252 304280
rect 42760 304240 42766 304252
rect 234246 304240 234252 304252
rect 234304 304240 234310 304292
rect 283926 304240 283932 304292
rect 283984 304280 283990 304292
rect 523034 304280 523040 304292
rect 283984 304252 523040 304280
rect 283984 304240 283990 304252
rect 523034 304240 523040 304252
rect 523092 304240 523098 304292
rect 275554 302948 275560 303000
rect 275612 302988 275618 303000
rect 444374 302988 444380 303000
rect 275612 302960 444380 302988
rect 275612 302948 275618 302960
rect 444374 302948 444380 302960
rect 444432 302948 444438 303000
rect 50982 302880 50988 302932
rect 51040 302920 51046 302932
rect 235074 302920 235080 302932
rect 51040 302892 235080 302920
rect 51040 302880 51046 302892
rect 235074 302880 235080 302892
rect 235132 302880 235138 302932
rect 283009 302923 283067 302929
rect 283009 302889 283021 302923
rect 283055 302920 283067 302923
rect 527174 302920 527180 302932
rect 283055 302892 527180 302920
rect 283055 302889 283067 302892
rect 283009 302883 283067 302889
rect 527174 302880 527180 302892
rect 527232 302880 527238 302932
rect 238110 302268 238116 302320
rect 238168 302268 238174 302320
rect 275278 302268 275284 302320
rect 275336 302268 275342 302320
rect 238128 302104 238156 302268
rect 238202 302104 238208 302116
rect 238128 302076 238208 302104
rect 238202 302064 238208 302076
rect 238260 302064 238266 302116
rect 256510 302064 256516 302116
rect 256568 302104 256574 302116
rect 256694 302104 256700 302116
rect 256568 302076 256700 302104
rect 256568 302064 256574 302076
rect 256694 302064 256700 302076
rect 256752 302064 256758 302116
rect 275296 302104 275324 302268
rect 284662 302172 284668 302184
rect 284623 302144 284668 302172
rect 284662 302132 284668 302144
rect 284720 302132 284726 302184
rect 275370 302104 275376 302116
rect 275296 302076 275376 302104
rect 275370 302064 275376 302076
rect 275428 302064 275434 302116
rect 277026 301520 277032 301572
rect 277084 301560 277090 301572
rect 448514 301560 448520 301572
rect 277084 301532 448520 301560
rect 277084 301520 277090 301532
rect 448514 301520 448520 301532
rect 448572 301520 448578 301572
rect 284386 301452 284392 301504
rect 284444 301492 284450 301504
rect 534074 301492 534080 301504
rect 284444 301464 534080 301492
rect 284444 301452 284450 301464
rect 534074 301452 534080 301464
rect 534132 301452 534138 301504
rect 276842 300160 276848 300212
rect 276900 300200 276906 300212
rect 455414 300200 455420 300212
rect 276900 300172 455420 300200
rect 276900 300160 276906 300172
rect 455414 300160 455420 300172
rect 455472 300160 455478 300212
rect 285306 300092 285312 300144
rect 285364 300132 285370 300144
rect 536926 300132 536932 300144
rect 285364 300104 536932 300132
rect 285364 300092 285370 300104
rect 536926 300092 536932 300104
rect 536984 300092 536990 300144
rect 283742 299588 283748 299600
rect 283703 299560 283748 299588
rect 283742 299548 283748 299560
rect 283800 299548 283806 299600
rect 229465 299523 229523 299529
rect 229465 299489 229477 299523
rect 229511 299520 229523 299523
rect 229554 299520 229560 299532
rect 229511 299492 229560 299520
rect 229511 299489 229523 299492
rect 229465 299483 229523 299489
rect 229554 299480 229560 299492
rect 229612 299480 229618 299532
rect 238938 299520 238944 299532
rect 238899 299492 238944 299520
rect 238938 299480 238944 299492
rect 238996 299480 239002 299532
rect 302970 299412 302976 299464
rect 303028 299452 303034 299464
rect 579798 299452 579804 299464
rect 303028 299424 579804 299452
rect 303028 299412 303034 299424
rect 579798 299412 579804 299424
rect 579856 299412 579862 299464
rect 260193 299387 260251 299393
rect 260193 299353 260205 299387
rect 260239 299384 260251 299387
rect 260282 299384 260288 299396
rect 260239 299356 260288 299384
rect 260239 299353 260251 299356
rect 260193 299347 260251 299353
rect 260282 299344 260288 299356
rect 260340 299344 260346 299396
rect 277578 298732 277584 298784
rect 277636 298772 277642 298784
rect 469214 298772 469220 298784
rect 277636 298744 469220 298772
rect 277636 298732 277642 298744
rect 469214 298732 469220 298744
rect 469272 298732 469278 298784
rect 254026 298256 254032 298308
rect 254084 298256 254090 298308
rect 254044 298172 254072 298256
rect 251726 298160 251732 298172
rect 251687 298132 251732 298160
rect 251726 298120 251732 298132
rect 251784 298120 251790 298172
rect 254026 298120 254032 298172
rect 254084 298120 254090 298172
rect 237561 298095 237619 298101
rect 237561 298061 237573 298095
rect 237607 298092 237619 298095
rect 237650 298092 237656 298104
rect 237607 298064 237656 298092
rect 237607 298061 237619 298064
rect 237561 298055 237619 298061
rect 237650 298052 237656 298064
rect 237708 298052 237714 298104
rect 283742 298092 283748 298104
rect 283703 298064 283748 298092
rect 283742 298052 283748 298064
rect 283800 298052 283806 298104
rect 288158 298092 288164 298104
rect 288119 298064 288164 298092
rect 288158 298052 288164 298064
rect 288216 298052 288222 298104
rect 282546 297440 282552 297492
rect 282604 297480 282610 297492
rect 502426 297480 502432 297492
rect 282604 297452 502432 297480
rect 282604 297440 282610 297452
rect 502426 297440 502432 297452
rect 502484 297440 502490 297492
rect 285950 297372 285956 297424
rect 286008 297412 286014 297424
rect 547874 297412 547880 297424
rect 286008 297384 547880 297412
rect 286008 297372 286014 297384
rect 547874 297372 547880 297384
rect 547932 297372 547938 297424
rect 278130 296692 278136 296744
rect 278188 296732 278194 296744
rect 278314 296732 278320 296744
rect 278188 296704 278320 296732
rect 278188 296692 278194 296704
rect 278314 296692 278320 296704
rect 278372 296692 278378 296744
rect 289446 296012 289452 296064
rect 289504 296052 289510 296064
rect 482278 296052 482284 296064
rect 289504 296024 482284 296052
rect 289504 296012 289510 296024
rect 482278 296012 482284 296024
rect 482336 296012 482342 296064
rect 288066 295944 288072 295996
rect 288124 295984 288130 295996
rect 565078 295984 565084 295996
rect 288124 295956 565084 295984
rect 288124 295944 288130 295956
rect 565078 295944 565084 295956
rect 565136 295944 565142 295996
rect 3510 295264 3516 295316
rect 3568 295304 3574 295316
rect 227162 295304 227168 295316
rect 3568 295276 227168 295304
rect 3568 295264 3574 295276
rect 227162 295264 227168 295276
rect 227220 295264 227226 295316
rect 289538 294652 289544 294704
rect 289596 294692 289602 294704
rect 475378 294692 475384 294704
rect 289596 294664 475384 294692
rect 289596 294652 289602 294664
rect 475378 294652 475384 294664
rect 475436 294652 475442 294704
rect 290550 294584 290556 294636
rect 290608 294624 290614 294636
rect 569954 294624 569960 294636
rect 290608 294596 569960 294624
rect 290608 294584 290614 294596
rect 569954 294584 569960 294596
rect 570012 294584 570018 294636
rect 263318 293292 263324 293344
rect 263376 293332 263382 293344
rect 324314 293332 324320 293344
rect 263376 293304 324320 293332
rect 263376 293292 263382 293304
rect 324314 293292 324320 293304
rect 324372 293292 324378 293344
rect 289354 293224 289360 293276
rect 289412 293264 289418 293276
rect 573450 293264 573456 293276
rect 289412 293236 573456 293264
rect 289412 293224 289418 293236
rect 573450 293224 573456 293236
rect 573508 293224 573514 293276
rect 275370 292652 275376 292664
rect 275296 292624 275376 292652
rect 275296 292528 275324 292624
rect 275370 292612 275376 292624
rect 275428 292612 275434 292664
rect 251637 292519 251695 292525
rect 251637 292485 251649 292519
rect 251683 292516 251695 292519
rect 251726 292516 251732 292528
rect 251683 292488 251732 292516
rect 251683 292485 251695 292488
rect 251637 292479 251695 292485
rect 251726 292476 251732 292488
rect 251784 292476 251790 292528
rect 275278 292476 275284 292528
rect 275336 292476 275342 292528
rect 272886 291864 272892 291916
rect 272944 291904 272950 291916
rect 419534 291904 419540 291916
rect 272944 291876 419540 291904
rect 272944 291864 272950 291876
rect 419534 291864 419540 291876
rect 419592 291864 419598 291916
rect 282638 291796 282644 291848
rect 282696 291836 282702 291848
rect 506474 291836 506480 291848
rect 282696 291808 506480 291836
rect 282696 291796 282702 291808
rect 506474 291796 506480 291808
rect 506532 291796 506538 291848
rect 274174 290504 274180 290556
rect 274232 290544 274238 290556
rect 430574 290544 430580 290556
rect 274232 290516 430580 290544
rect 274232 290504 274238 290516
rect 430574 290504 430580 290516
rect 430632 290504 430638 290556
rect 284938 290436 284944 290488
rect 284996 290476 285002 290488
rect 524414 290476 524420 290488
rect 284996 290448 524420 290476
rect 284996 290436 285002 290448
rect 524414 290436 524420 290448
rect 524472 290436 524478 290488
rect 256510 289824 256516 289876
rect 256568 289824 256574 289876
rect 238110 289756 238116 289808
rect 238168 289796 238174 289808
rect 238202 289796 238208 289808
rect 238168 289768 238208 289796
rect 238168 289756 238174 289768
rect 238202 289756 238208 289768
rect 238260 289756 238266 289808
rect 241054 289756 241060 289808
rect 241112 289796 241118 289808
rect 241146 289796 241152 289808
rect 241112 289768 241152 289796
rect 241112 289756 241118 289768
rect 241146 289756 241152 289768
rect 241204 289756 241210 289808
rect 243446 289796 243452 289808
rect 243407 289768 243452 289796
rect 243446 289756 243452 289768
rect 243504 289756 243510 289808
rect 256528 289728 256556 289824
rect 284386 289756 284392 289808
rect 284444 289796 284450 289808
rect 284662 289796 284668 289808
rect 284444 289768 284668 289796
rect 284444 289756 284450 289768
rect 284662 289756 284668 289768
rect 284720 289756 284726 289808
rect 256602 289728 256608 289740
rect 256528 289700 256608 289728
rect 256602 289688 256608 289700
rect 256660 289688 256666 289740
rect 277857 289595 277915 289601
rect 277857 289561 277869 289595
rect 277903 289592 277915 289595
rect 277946 289592 277952 289604
rect 277903 289564 277952 289592
rect 277903 289561 277915 289564
rect 277857 289555 277915 289561
rect 277946 289552 277952 289564
rect 278004 289552 278010 289604
rect 276014 289144 276020 289196
rect 276072 289184 276078 289196
rect 451366 289184 451372 289196
rect 276072 289156 451372 289184
rect 276072 289144 276078 289156
rect 451366 289144 451372 289156
rect 451424 289144 451430 289196
rect 286042 289076 286048 289128
rect 286100 289116 286106 289128
rect 549254 289116 549260 289128
rect 286100 289088 549260 289116
rect 286100 289076 286106 289088
rect 549254 289076 549260 289088
rect 549312 289076 549318 289128
rect 237558 288436 237564 288448
rect 237519 288408 237564 288436
rect 237558 288396 237564 288408
rect 237616 288396 237622 288448
rect 283745 288439 283803 288445
rect 283745 288405 283757 288439
rect 283791 288436 283803 288439
rect 283834 288436 283840 288448
rect 283791 288408 283840 288436
rect 283791 288405 283803 288408
rect 283745 288399 283803 288405
rect 283834 288396 283840 288408
rect 283892 288396 283898 288448
rect 288158 288436 288164 288448
rect 288119 288408 288164 288436
rect 288158 288396 288164 288408
rect 288216 288396 288222 288448
rect 276290 287716 276296 287768
rect 276348 287756 276354 287768
rect 459646 287756 459652 287768
rect 276348 287728 459652 287756
rect 276348 287716 276354 287728
rect 459646 287716 459652 287728
rect 459704 287716 459710 287768
rect 289354 287648 289360 287700
rect 289412 287688 289418 287700
rect 571426 287688 571432 287700
rect 289412 287660 571432 287688
rect 289412 287648 289418 287660
rect 571426 287648 571432 287660
rect 571484 287648 571490 287700
rect 251634 287076 251640 287088
rect 251595 287048 251640 287076
rect 251634 287036 251640 287048
rect 251692 287036 251698 287088
rect 253842 287036 253848 287088
rect 253900 287076 253906 287088
rect 254026 287076 254032 287088
rect 253900 287048 254032 287076
rect 253900 287036 253906 287048
rect 254026 287036 254032 287048
rect 254084 287036 254090 287088
rect 279602 286288 279608 286340
rect 279660 286328 279666 286340
rect 477494 286328 477500 286340
rect 279660 286300 477500 286328
rect 279660 286288 279666 286300
rect 477494 286288 477500 286300
rect 477552 286288 477558 286340
rect 279694 284928 279700 284980
rect 279752 284968 279758 284980
rect 480254 284968 480260 284980
rect 279752 284940 480260 284968
rect 279752 284928 279758 284940
rect 480254 284928 480260 284940
rect 480312 284928 480318 284980
rect 278866 283568 278872 283620
rect 278924 283608 278930 283620
rect 485774 283608 485780 283620
rect 278924 283580 485780 283608
rect 278924 283568 278930 283580
rect 485774 283568 485780 283580
rect 485832 283568 485838 283620
rect 275370 282928 275376 282940
rect 275296 282900 275376 282928
rect 275296 282872 275324 282900
rect 275370 282888 275376 282900
rect 275428 282888 275434 282940
rect 275278 282820 275284 282872
rect 275336 282820 275342 282872
rect 280246 282140 280252 282192
rect 280304 282180 280310 282192
rect 488534 282180 488540 282192
rect 280304 282152 488540 282180
rect 280304 282140 280310 282152
rect 488534 282140 488540 282152
rect 488592 282140 488598 282192
rect 260098 281936 260104 281988
rect 260156 281976 260162 281988
rect 260282 281976 260288 281988
rect 260156 281948 260288 281976
rect 260156 281936 260162 281948
rect 260282 281936 260288 281948
rect 260340 281936 260346 281988
rect 281258 280780 281264 280832
rect 281316 280820 281322 280832
rect 492674 280820 492680 280832
rect 281316 280792 492680 280820
rect 281316 280780 281322 280792
rect 492674 280780 492680 280792
rect 492732 280780 492738 280832
rect 243449 280211 243507 280217
rect 243449 280177 243461 280211
rect 243495 280208 243507 280211
rect 243538 280208 243544 280220
rect 243495 280180 243544 280208
rect 243495 280177 243507 280180
rect 243449 280171 243507 280177
rect 243538 280168 243544 280180
rect 243596 280168 243602 280220
rect 260282 280168 260288 280220
rect 260340 280208 260346 280220
rect 260558 280208 260564 280220
rect 260340 280180 260564 280208
rect 260340 280168 260346 280180
rect 260558 280168 260564 280180
rect 260616 280168 260622 280220
rect 229554 280140 229560 280152
rect 229515 280112 229560 280140
rect 229554 280100 229560 280112
rect 229612 280100 229618 280152
rect 259914 280100 259920 280152
rect 259972 280140 259978 280152
rect 260098 280140 260104 280152
rect 259972 280112 260104 280140
rect 259972 280100 259978 280112
rect 260098 280100 260104 280112
rect 260156 280100 260162 280152
rect 281350 279420 281356 279472
rect 281408 279460 281414 279472
rect 499574 279460 499580 279472
rect 281408 279432 499580 279460
rect 281408 279420 281414 279432
rect 499574 279420 499580 279432
rect 499632 279420 499638 279472
rect 284386 279148 284392 279200
rect 284444 279188 284450 279200
rect 284938 279188 284944 279200
rect 284444 279160 284944 279188
rect 284444 279148 284450 279160
rect 284938 279148 284944 279160
rect 284996 279148 285002 279200
rect 243449 278715 243507 278721
rect 243449 278681 243461 278715
rect 243495 278712 243507 278715
rect 243538 278712 243544 278724
rect 243495 278684 243544 278712
rect 243495 278681 243507 278684
rect 243449 278675 243507 278681
rect 243538 278672 243544 278684
rect 243596 278672 243602 278724
rect 259914 278712 259920 278724
rect 259875 278684 259920 278712
rect 259914 278672 259920 278684
rect 259972 278672 259978 278724
rect 281902 277992 281908 278044
rect 281960 278032 281966 278044
rect 510614 278032 510620 278044
rect 281960 278004 510620 278032
rect 281960 277992 281966 278004
rect 510614 277992 510620 278004
rect 510672 277992 510678 278044
rect 277854 277420 277860 277432
rect 277815 277392 277860 277420
rect 277854 277380 277860 277392
rect 277912 277380 277918 277432
rect 282086 276632 282092 276684
rect 282144 276672 282150 276684
rect 513374 276672 513380 276684
rect 282144 276644 513380 276672
rect 282144 276632 282150 276644
rect 513374 276632 513380 276644
rect 513432 276632 513438 276684
rect 393958 275952 393964 276004
rect 394016 275992 394022 276004
rect 580166 275992 580172 276004
rect 394016 275964 580172 275992
rect 394016 275952 394022 275964
rect 580166 275952 580172 275964
rect 580224 275952 580230 276004
rect 260282 275272 260288 275324
rect 260340 275312 260346 275324
rect 260558 275312 260564 275324
rect 260340 275284 260564 275312
rect 260340 275272 260346 275284
rect 260558 275272 260564 275284
rect 260616 275272 260622 275324
rect 284110 273912 284116 273964
rect 284168 273952 284174 273964
rect 517514 273952 517520 273964
rect 284168 273924 517520 273952
rect 284168 273912 284174 273924
rect 517514 273912 517520 273924
rect 517572 273912 517578 273964
rect 272426 273340 272432 273352
rect 272352 273312 272432 273340
rect 272352 273216 272380 273312
rect 272426 273300 272432 273312
rect 272484 273300 272490 273352
rect 272334 273164 272340 273216
rect 272392 273164 272398 273216
rect 283742 272484 283748 272536
rect 283800 272524 283806 272536
rect 520366 272524 520372 272536
rect 283800 272496 520372 272524
rect 283800 272484 283806 272496
rect 520366 272484 520372 272496
rect 520424 272484 520430 272536
rect 284478 271124 284484 271176
rect 284536 271164 284542 271176
rect 528646 271164 528652 271176
rect 284536 271136 528652 271164
rect 284536 271124 284542 271136
rect 528646 271124 528652 271136
rect 528704 271124 528710 271176
rect 229557 270555 229615 270561
rect 229557 270521 229569 270555
rect 229603 270552 229615 270555
rect 229646 270552 229652 270564
rect 229603 270524 229652 270552
rect 229603 270521 229615 270524
rect 229557 270515 229615 270521
rect 229646 270512 229652 270524
rect 229704 270512 229710 270564
rect 241146 270484 241152 270496
rect 241107 270456 241152 270484
rect 241146 270444 241152 270456
rect 241204 270444 241210 270496
rect 284938 269764 284944 269816
rect 284996 269804 285002 269816
rect 531314 269804 531320 269816
rect 284996 269776 531320 269804
rect 284996 269764 285002 269776
rect 531314 269764 531320 269776
rect 531372 269764 531378 269816
rect 270862 269084 270868 269136
rect 270920 269124 270926 269136
rect 270954 269124 270960 269136
rect 270920 269096 270960 269124
rect 270920 269084 270926 269096
rect 270954 269084 270960 269096
rect 271012 269084 271018 269136
rect 288066 269084 288072 269136
rect 288124 269124 288130 269136
rect 288158 269124 288164 269136
rect 288124 269096 288164 269124
rect 288124 269084 288130 269096
rect 288158 269084 288164 269096
rect 288216 269084 288222 269136
rect 284754 268336 284760 268388
rect 284812 268376 284818 268388
rect 535454 268376 535460 268388
rect 284812 268348 535460 268376
rect 284812 268336 284818 268348
rect 535454 268336 535460 268348
rect 535512 268336 535518 268388
rect 259917 267767 259975 267773
rect 259917 267733 259929 267767
rect 259963 267764 259975 267767
rect 260098 267764 260104 267776
rect 259963 267736 260104 267764
rect 259963 267733 259975 267736
rect 259917 267727 259975 267733
rect 260098 267724 260104 267736
rect 260156 267724 260162 267776
rect 284846 266976 284852 267028
rect 284904 267016 284910 267028
rect 538214 267016 538220 267028
rect 284904 266988 538220 267016
rect 284904 266976 284910 266988
rect 538214 266976 538220 266988
rect 538272 266976 538278 267028
rect 3510 266296 3516 266348
rect 3568 266336 3574 266348
rect 211798 266336 211804 266348
rect 3568 266308 211804 266336
rect 3568 266296 3574 266308
rect 211798 266296 211804 266308
rect 211856 266296 211862 266348
rect 286778 265616 286784 265668
rect 286836 265656 286842 265668
rect 542354 265656 542360 265668
rect 286836 265628 542360 265656
rect 286836 265616 286842 265628
rect 542354 265616 542360 265628
rect 542412 265616 542418 265668
rect 315298 264868 315304 264920
rect 315356 264908 315362 264920
rect 580166 264908 580172 264920
rect 315356 264880 580172 264908
rect 315356 264868 315362 264880
rect 580166 264868 580172 264880
rect 580224 264868 580230 264920
rect 286134 262828 286140 262880
rect 286192 262868 286198 262880
rect 546586 262868 546592 262880
rect 286192 262840 546592 262868
rect 286192 262828 286198 262840
rect 546586 262828 546592 262840
rect 546644 262828 546650 262880
rect 286226 261468 286232 261520
rect 286284 261508 286290 261520
rect 553394 261508 553400 261520
rect 286284 261480 553400 261508
rect 286284 261468 286290 261480
rect 553394 261468 553400 261480
rect 553452 261468 553458 261520
rect 275370 260964 275376 260976
rect 275296 260936 275376 260964
rect 241146 260896 241152 260908
rect 241107 260868 241152 260896
rect 241146 260856 241152 260868
rect 241204 260856 241210 260908
rect 253937 260899 253995 260905
rect 253937 260865 253949 260899
rect 253983 260896 253995 260899
rect 254026 260896 254032 260908
rect 253983 260868 254032 260896
rect 253983 260865 253995 260868
rect 253937 260859 253995 260865
rect 254026 260856 254032 260868
rect 254084 260856 254090 260908
rect 229554 260828 229560 260840
rect 229515 260800 229560 260828
rect 229554 260788 229560 260800
rect 229612 260788 229618 260840
rect 251358 260788 251364 260840
rect 251416 260828 251422 260840
rect 251634 260828 251640 260840
rect 251416 260800 251640 260828
rect 251416 260788 251422 260800
rect 251634 260788 251640 260800
rect 251692 260788 251698 260840
rect 275296 260772 275324 260936
rect 275370 260924 275376 260936
rect 275428 260924 275434 260976
rect 275278 260720 275284 260772
rect 275336 260720 275342 260772
rect 287238 260108 287244 260160
rect 287296 260148 287302 260160
rect 556154 260148 556160 260160
rect 287296 260120 556160 260148
rect 287296 260108 287302 260120
rect 556154 260108 556160 260120
rect 556212 260108 556218 260160
rect 237650 259564 237656 259616
rect 237708 259564 237714 259616
rect 237668 259480 237696 259564
rect 237650 259428 237656 259480
rect 237708 259428 237714 259480
rect 260374 259428 260380 259480
rect 260432 259468 260438 259480
rect 260558 259468 260564 259480
rect 260432 259440 260564 259468
rect 260432 259428 260438 259440
rect 260558 259428 260564 259440
rect 260616 259428 260622 259480
rect 270770 259428 270776 259480
rect 270828 259468 270834 259480
rect 270954 259468 270960 259480
rect 270828 259440 270960 259468
rect 270828 259428 270834 259440
rect 270954 259428 270960 259440
rect 271012 259428 271018 259480
rect 288158 258680 288164 258732
rect 288216 258720 288222 258732
rect 560294 258720 560300 258732
rect 288216 258692 560300 258720
rect 288216 258680 288222 258692
rect 560294 258680 560300 258692
rect 560352 258680 560358 258732
rect 253934 258108 253940 258120
rect 253895 258080 253940 258108
rect 253934 258068 253940 258080
rect 253992 258068 253998 258120
rect 260098 258040 260104 258052
rect 260059 258012 260104 258040
rect 260098 258000 260104 258012
rect 260156 258000 260162 258052
rect 260193 258043 260251 258049
rect 260193 258009 260205 258043
rect 260239 258040 260251 258043
rect 260374 258040 260380 258052
rect 260239 258012 260380 258040
rect 260239 258009 260251 258012
rect 260193 258003 260251 258009
rect 260374 258000 260380 258012
rect 260432 258000 260438 258052
rect 287514 257320 287520 257372
rect 287572 257360 287578 257372
rect 563146 257360 563152 257372
rect 287572 257332 563152 257360
rect 287572 257320 287578 257332
rect 563146 257320 563152 257332
rect 563204 257320 563210 257372
rect 243449 256751 243507 256757
rect 243449 256717 243461 256751
rect 243495 256748 243507 256751
rect 243538 256748 243544 256760
rect 243495 256720 243544 256748
rect 243495 256717 243507 256720
rect 243449 256711 243507 256717
rect 243538 256708 243544 256720
rect 243596 256708 243602 256760
rect 291102 255960 291108 256012
rect 291160 256000 291166 256012
rect 471238 256000 471244 256012
rect 291160 255972 471244 256000
rect 291160 255960 291166 255972
rect 471238 255960 471244 255972
rect 471296 255960 471302 256012
rect 243449 255255 243507 255261
rect 243449 255221 243461 255255
rect 243495 255252 243507 255255
rect 243538 255252 243544 255264
rect 243495 255224 243544 255252
rect 243495 255221 243507 255224
rect 243449 255215 243507 255221
rect 243538 255212 243544 255224
rect 243596 255212 243602 255264
rect 277854 254532 277860 254584
rect 277912 254572 277918 254584
rect 278038 254572 278044 254584
rect 277912 254544 278044 254572
rect 277912 254532 277918 254544
rect 278038 254532 278044 254544
rect 278096 254532 278102 254584
rect 237650 254028 237656 254040
rect 237576 254000 237656 254028
rect 237576 253904 237604 254000
rect 237650 253988 237656 254000
rect 237708 253988 237714 254040
rect 237558 253852 237564 253904
rect 237616 253852 237622 253904
rect 251358 253172 251364 253224
rect 251416 253212 251422 253224
rect 251542 253212 251548 253224
rect 251416 253184 251548 253212
rect 251416 253172 251422 253184
rect 251542 253172 251548 253184
rect 251600 253172 251606 253224
rect 3142 252492 3148 252544
rect 3200 252532 3206 252544
rect 225782 252532 225788 252544
rect 3200 252504 225788 252532
rect 3200 252492 3206 252504
rect 225782 252492 225788 252504
rect 225840 252492 225846 252544
rect 301590 252492 301596 252544
rect 301648 252532 301654 252544
rect 579798 252532 579804 252544
rect 301648 252504 579804 252532
rect 301648 252492 301654 252504
rect 579798 252492 579804 252504
rect 579856 252492 579862 252544
rect 229557 251243 229615 251249
rect 229557 251209 229569 251243
rect 229603 251240 229615 251243
rect 229646 251240 229652 251252
rect 229603 251212 229652 251240
rect 229603 251209 229615 251212
rect 229557 251203 229615 251209
rect 229646 251200 229652 251212
rect 229704 251200 229710 251252
rect 275278 249812 275284 249824
rect 275239 249784 275284 249812
rect 275278 249772 275284 249784
rect 275336 249772 275342 249824
rect 260098 249744 260104 249756
rect 260059 249716 260104 249744
rect 260098 249704 260104 249716
rect 260156 249704 260162 249756
rect 260190 248452 260196 248464
rect 260151 248424 260196 248452
rect 260190 248412 260196 248424
rect 260248 248412 260254 248464
rect 275278 248452 275284 248464
rect 275239 248424 275284 248452
rect 275278 248412 275284 248424
rect 275336 248412 275342 248464
rect 237558 248384 237564 248396
rect 237519 248356 237564 248384
rect 237558 248344 237564 248356
rect 237616 248344 237622 248396
rect 277854 248344 277860 248396
rect 277912 248384 277918 248396
rect 278038 248384 278044 248396
rect 277912 248356 278044 248384
rect 277912 248344 277918 248356
rect 278038 248344 278044 248356
rect 278096 248344 278102 248396
rect 240870 246984 240876 247036
rect 240928 247024 240934 247036
rect 241146 247024 241152 247036
rect 240928 246996 241152 247024
rect 240928 246984 240934 246996
rect 241146 246984 241152 246996
rect 241204 246984 241210 247036
rect 251542 244944 251548 244996
rect 251600 244984 251606 244996
rect 251726 244984 251732 244996
rect 251600 244956 251732 244984
rect 251600 244944 251606 244956
rect 251726 244944 251732 244956
rect 251784 244944 251790 244996
rect 259914 244944 259920 244996
rect 259972 244984 259978 244996
rect 260098 244984 260104 244996
rect 259972 244956 260104 244984
rect 259972 244944 259978 244956
rect 260098 244944 260104 244956
rect 260156 244944 260162 244996
rect 258537 244443 258595 244449
rect 258537 244409 258549 244443
rect 258583 244440 258595 244443
rect 258626 244440 258632 244452
rect 258583 244412 258632 244440
rect 258583 244409 258595 244412
rect 258537 244403 258595 244409
rect 258626 244400 258632 244412
rect 258684 244400 258690 244452
rect 259362 244304 259368 244316
rect 259288 244276 259368 244304
rect 259288 244248 259316 244276
rect 259362 244264 259368 244276
rect 259420 244264 259426 244316
rect 259270 244196 259276 244248
rect 259328 244196 259334 244248
rect 237561 244171 237619 244177
rect 237561 244137 237573 244171
rect 237607 244168 237619 244171
rect 237650 244168 237656 244180
rect 237607 244140 237656 244168
rect 237607 244137 237619 244140
rect 237561 244131 237619 244137
rect 237650 244128 237656 244140
rect 237708 244128 237714 244180
rect 272334 241476 272340 241528
rect 272392 241516 272398 241528
rect 272426 241516 272432 241528
rect 272392 241488 272432 241516
rect 272392 241476 272398 241488
rect 272426 241476 272432 241488
rect 272484 241476 272490 241528
rect 278222 241476 278228 241528
rect 278280 241516 278286 241528
rect 278314 241516 278320 241528
rect 278280 241488 278320 241516
rect 278280 241476 278286 241488
rect 278314 241476 278320 241488
rect 278372 241476 278378 241528
rect 243449 240227 243507 240233
rect 243449 240193 243461 240227
rect 243495 240224 243507 240227
rect 243538 240224 243544 240236
rect 243495 240196 243544 240224
rect 243495 240193 243507 240196
rect 243449 240187 243507 240193
rect 243538 240184 243544 240196
rect 243596 240184 243602 240236
rect 258534 240156 258540 240168
rect 258495 240128 258540 240156
rect 258534 240116 258540 240128
rect 258592 240116 258598 240168
rect 270770 240116 270776 240168
rect 270828 240156 270834 240168
rect 270954 240156 270960 240168
rect 270828 240128 270960 240156
rect 270828 240116 270834 240128
rect 270954 240116 270960 240128
rect 271012 240116 271018 240168
rect 275278 240116 275284 240168
rect 275336 240156 275342 240168
rect 275370 240156 275376 240168
rect 275336 240128 275376 240156
rect 275336 240116 275342 240128
rect 275370 240116 275376 240128
rect 275428 240116 275434 240168
rect 259178 240048 259184 240100
rect 259236 240088 259242 240100
rect 259270 240088 259276 240100
rect 259236 240060 259276 240088
rect 259236 240048 259242 240060
rect 259270 240048 259276 240060
rect 259328 240048 259334 240100
rect 260190 240048 260196 240100
rect 260248 240088 260254 240100
rect 260285 240091 260343 240097
rect 260285 240088 260297 240091
rect 260248 240060 260297 240088
rect 260248 240048 260254 240060
rect 260285 240057 260297 240060
rect 260331 240057 260343 240091
rect 260285 240051 260343 240057
rect 254026 238728 254032 238740
rect 253987 238700 254032 238728
rect 254026 238688 254032 238700
rect 254084 238688 254090 238740
rect 275370 238688 275376 238740
rect 275428 238728 275434 238740
rect 275554 238728 275560 238740
rect 275428 238700 275560 238728
rect 275428 238688 275434 238700
rect 275554 238688 275560 238700
rect 275612 238688 275618 238740
rect 277762 238688 277768 238740
rect 277820 238728 277826 238740
rect 278038 238728 278044 238740
rect 277820 238700 278044 238728
rect 277820 238688 277826 238700
rect 278038 238688 278044 238700
rect 278096 238688 278102 238740
rect 238110 237328 238116 237380
rect 238168 237368 238174 237380
rect 238294 237368 238300 237380
rect 238168 237340 238300 237368
rect 238168 237328 238174 237340
rect 238294 237328 238300 237340
rect 238352 237328 238358 237380
rect 243449 237371 243507 237377
rect 243449 237337 243461 237371
rect 243495 237368 243507 237371
rect 243538 237368 243544 237380
rect 243495 237340 243544 237368
rect 243495 237337 243507 237340
rect 243449 237331 243507 237337
rect 243538 237328 243544 237340
rect 243596 237328 243602 237380
rect 259914 235288 259920 235340
rect 259972 235328 259978 235340
rect 260190 235328 260196 235340
rect 259972 235300 260196 235328
rect 259972 235288 259978 235300
rect 260190 235288 260196 235300
rect 260248 235288 260254 235340
rect 237469 231999 237527 232005
rect 237469 231965 237481 231999
rect 237515 231996 237527 231999
rect 237650 231996 237656 232008
rect 237515 231968 237656 231996
rect 237515 231965 237527 231968
rect 237469 231959 237527 231965
rect 237650 231956 237656 231968
rect 237708 231956 237714 232008
rect 229646 231820 229652 231872
rect 229704 231860 229710 231872
rect 229830 231860 229836 231872
rect 229704 231832 229836 231860
rect 229704 231820 229710 231832
rect 229830 231820 229836 231832
rect 229888 231820 229894 231872
rect 258534 230460 258540 230512
rect 258592 230500 258598 230512
rect 258626 230500 258632 230512
rect 258592 230472 258632 230500
rect 258592 230460 258598 230472
rect 258626 230460 258632 230472
rect 258684 230460 258690 230512
rect 260282 230500 260288 230512
rect 260243 230472 260288 230500
rect 260282 230460 260288 230472
rect 260340 230460 260346 230512
rect 254026 230296 254032 230308
rect 253987 230268 254032 230296
rect 254026 230256 254032 230268
rect 254084 230256 254090 230308
rect 238938 229032 238944 229084
rect 238996 229072 239002 229084
rect 239122 229072 239128 229084
rect 238996 229044 239128 229072
rect 238996 229032 239002 229044
rect 239122 229032 239128 229044
rect 239180 229032 239186 229084
rect 240870 229032 240876 229084
rect 240928 229072 240934 229084
rect 241146 229072 241152 229084
rect 240928 229044 241152 229072
rect 240928 229032 240934 229044
rect 241146 229032 241152 229044
rect 241204 229032 241210 229084
rect 259454 227944 259460 227996
rect 259512 227984 259518 227996
rect 270402 227984 270408 227996
rect 259512 227956 270408 227984
rect 259512 227944 259518 227956
rect 270402 227944 270408 227956
rect 270460 227944 270466 227996
rect 321462 227876 321468 227928
rect 321520 227916 321526 227928
rect 323026 227916 323032 227928
rect 321520 227888 323032 227916
rect 321520 227876 321526 227888
rect 323026 227876 323032 227888
rect 323084 227876 323090 227928
rect 302142 227808 302148 227860
rect 302200 227848 302206 227860
rect 309042 227848 309048 227860
rect 302200 227820 309048 227848
rect 302200 227808 302206 227820
rect 309042 227808 309048 227820
rect 309100 227808 309106 227860
rect 437382 227808 437388 227860
rect 437440 227848 437446 227860
rect 444282 227848 444288 227860
rect 437440 227820 444288 227848
rect 437440 227808 437446 227820
rect 444282 227808 444288 227820
rect 444340 227808 444346 227860
rect 476022 227808 476028 227860
rect 476080 227848 476086 227860
rect 482922 227848 482928 227860
rect 476080 227820 482928 227848
rect 476080 227808 476086 227820
rect 482922 227808 482928 227820
rect 482980 227808 482986 227860
rect 533982 227808 533988 227860
rect 534040 227848 534046 227860
rect 540882 227848 540888 227860
rect 534040 227820 540888 227848
rect 534040 227808 534046 227820
rect 540882 227808 540888 227820
rect 540940 227808 540946 227860
rect 553302 227808 553308 227860
rect 553360 227848 553366 227860
rect 560202 227848 560208 227860
rect 553360 227820 560208 227848
rect 553360 227808 553366 227820
rect 560202 227808 560208 227820
rect 560260 227808 560266 227860
rect 572622 227808 572628 227860
rect 572680 227848 572686 227860
rect 579522 227848 579528 227860
rect 572680 227820 579528 227848
rect 572680 227808 572686 227820
rect 579522 227808 579528 227820
rect 579580 227808 579586 227860
rect 237466 227780 237472 227792
rect 237427 227752 237472 227780
rect 237466 227740 237472 227752
rect 237524 227740 237530 227792
rect 277946 225196 277952 225208
rect 277907 225168 277952 225196
rect 277946 225156 277952 225168
rect 278004 225156 278010 225208
rect 251818 224992 251824 225004
rect 251779 224964 251824 224992
rect 251818 224952 251824 224964
rect 251876 224952 251882 225004
rect 3142 223524 3148 223576
rect 3200 223564 3206 223576
rect 209038 223564 209044 223576
rect 3200 223536 209044 223564
rect 3200 223524 3206 223536
rect 209038 223524 209044 223536
rect 209096 223524 209102 223576
rect 260282 222300 260288 222352
rect 260340 222300 260346 222352
rect 260300 222216 260328 222300
rect 251818 222204 251824 222216
rect 251779 222176 251824 222204
rect 251818 222164 251824 222176
rect 251876 222164 251882 222216
rect 256510 222164 256516 222216
rect 256568 222204 256574 222216
rect 256602 222204 256608 222216
rect 256568 222176 256608 222204
rect 256568 222164 256574 222176
rect 256602 222164 256608 222176
rect 256660 222164 256666 222216
rect 260098 222164 260104 222216
rect 260156 222204 260162 222216
rect 260190 222204 260196 222216
rect 260156 222176 260196 222204
rect 260156 222164 260162 222176
rect 260190 222164 260196 222176
rect 260248 222164 260254 222216
rect 260282 222164 260288 222216
rect 260340 222164 260346 222216
rect 259546 220804 259552 220856
rect 259604 220844 259610 220856
rect 259638 220844 259644 220856
rect 259604 220816 259644 220844
rect 259604 220804 259610 220816
rect 259638 220804 259644 220816
rect 259696 220804 259702 220856
rect 277946 220844 277952 220856
rect 277907 220816 277952 220844
rect 277946 220804 277952 220816
rect 278004 220804 278010 220856
rect 270954 220776 270960 220788
rect 270915 220748 270960 220776
rect 270954 220736 270960 220748
rect 271012 220736 271018 220788
rect 243446 219484 243452 219496
rect 243407 219456 243452 219484
rect 243446 219444 243452 219456
rect 243504 219444 243510 219496
rect 277857 219419 277915 219425
rect 277857 219385 277869 219419
rect 277903 219416 277915 219419
rect 277946 219416 277952 219428
rect 277903 219388 277952 219416
rect 277903 219385 277915 219388
rect 277857 219379 277915 219385
rect 277946 219376 277952 219388
rect 278004 219376 278010 219428
rect 237650 219348 237656 219360
rect 237611 219320 237656 219348
rect 237650 219308 237656 219320
rect 237708 219308 237714 219360
rect 243446 219348 243452 219360
rect 243407 219320 243452 219348
rect 243446 219308 243452 219320
rect 243504 219308 243510 219360
rect 238846 218832 238852 218884
rect 238904 218872 238910 218884
rect 238941 218875 238999 218881
rect 238941 218872 238953 218875
rect 238904 218844 238953 218872
rect 238904 218832 238910 218844
rect 238941 218841 238953 218844
rect 238987 218841 238999 218875
rect 238941 218835 238999 218841
rect 312538 217948 312544 218000
rect 312596 217988 312602 218000
rect 580166 217988 580172 218000
rect 312596 217960 580172 217988
rect 312596 217948 312602 217960
rect 580166 217948 580172 217960
rect 580224 217948 580230 218000
rect 272426 215404 272432 215416
rect 272352 215376 272432 215404
rect 272352 215280 272380 215376
rect 272426 215364 272432 215376
rect 272484 215364 272490 215416
rect 272334 215228 272340 215280
rect 272392 215228 272398 215280
rect 237650 214588 237656 214600
rect 237611 214560 237656 214588
rect 237650 214548 237656 214560
rect 237708 214548 237714 214600
rect 260006 212576 260012 212628
rect 260064 212576 260070 212628
rect 229646 212508 229652 212560
rect 229704 212548 229710 212560
rect 229830 212548 229836 212560
rect 229704 212520 229836 212548
rect 229704 212508 229710 212520
rect 229830 212508 229836 212520
rect 229888 212508 229894 212560
rect 259362 212508 259368 212560
rect 259420 212548 259426 212560
rect 259638 212548 259644 212560
rect 259420 212520 259644 212548
rect 259420 212508 259426 212520
rect 259638 212508 259644 212520
rect 259696 212508 259702 212560
rect 260024 212492 260052 212576
rect 260006 212440 260012 212492
rect 260064 212440 260070 212492
rect 270954 211188 270960 211200
rect 270915 211160 270960 211188
rect 270954 211148 270960 211160
rect 271012 211148 271018 211200
rect 277854 209828 277860 209840
rect 277815 209800 277860 209828
rect 277854 209788 277860 209800
rect 277912 209788 277918 209840
rect 275278 209760 275284 209772
rect 275239 209732 275284 209760
rect 275278 209720 275284 209732
rect 275336 209720 275342 209772
rect 3510 208292 3516 208344
rect 3568 208332 3574 208344
rect 180058 208332 180064 208344
rect 3568 208304 180064 208332
rect 3568 208292 3574 208304
rect 180058 208292 180064 208304
rect 180116 208292 180122 208344
rect 230842 205640 230848 205692
rect 230900 205680 230906 205692
rect 231026 205680 231032 205692
rect 230900 205652 231032 205680
rect 230900 205640 230906 205652
rect 231026 205640 231032 205652
rect 231084 205640 231090 205692
rect 251542 205640 251548 205692
rect 251600 205640 251606 205692
rect 251560 205556 251588 205640
rect 275278 205612 275284 205624
rect 275239 205584 275284 205612
rect 275278 205572 275284 205584
rect 275336 205572 275342 205624
rect 298830 205572 298836 205624
rect 298888 205612 298894 205624
rect 579798 205612 579804 205624
rect 298888 205584 579804 205612
rect 298888 205572 298894 205584
rect 579798 205572 579804 205584
rect 579856 205572 579862 205624
rect 251542 205504 251548 205556
rect 251600 205504 251606 205556
rect 238938 205340 238944 205352
rect 238899 205312 238944 205340
rect 238938 205300 238944 205312
rect 238996 205300 239002 205352
rect 243449 202895 243507 202901
rect 243449 202861 243461 202895
rect 243495 202892 243507 202895
rect 243538 202892 243544 202904
rect 243495 202864 243544 202892
rect 243495 202861 243507 202864
rect 243449 202855 243507 202861
rect 243538 202852 243544 202864
rect 243596 202852 243602 202904
rect 258626 202852 258632 202904
rect 258684 202892 258690 202904
rect 258718 202892 258724 202904
rect 258684 202864 258724 202892
rect 258684 202852 258690 202864
rect 258718 202852 258724 202864
rect 258776 202852 258782 202904
rect 259914 202852 259920 202904
rect 259972 202892 259978 202904
rect 260098 202892 260104 202904
rect 259972 202864 260104 202892
rect 259972 202852 259978 202864
rect 260098 202852 260104 202864
rect 260156 202852 260162 202904
rect 260190 202852 260196 202904
rect 260248 202892 260254 202904
rect 260282 202892 260288 202904
rect 260248 202864 260288 202892
rect 260248 202852 260254 202864
rect 260282 202852 260288 202864
rect 260340 202852 260346 202904
rect 237558 201424 237564 201476
rect 237616 201464 237622 201476
rect 237650 201464 237656 201476
rect 237616 201436 237656 201464
rect 237616 201424 237622 201436
rect 237650 201424 237656 201436
rect 237708 201424 237714 201476
rect 241146 201424 241152 201476
rect 241204 201464 241210 201476
rect 241330 201464 241336 201476
rect 241204 201436 241336 201464
rect 241204 201424 241210 201436
rect 241330 201424 241336 201436
rect 241388 201424 241394 201476
rect 259730 201424 259736 201476
rect 259788 201464 259794 201476
rect 260098 201464 260104 201476
rect 259788 201436 260104 201464
rect 259788 201424 259794 201436
rect 260098 201424 260104 201436
rect 260156 201424 260162 201476
rect 260193 201467 260251 201473
rect 260193 201433 260205 201467
rect 260239 201464 260251 201467
rect 260282 201464 260288 201476
rect 260239 201436 260288 201464
rect 260239 201433 260251 201436
rect 260193 201427 260251 201433
rect 260282 201424 260288 201436
rect 260340 201424 260346 201476
rect 251634 197888 251640 197940
rect 251692 197928 251698 197940
rect 251726 197928 251732 197940
rect 251692 197900 251732 197928
rect 251692 197888 251698 197900
rect 251726 197888 251732 197900
rect 251784 197888 251790 197940
rect 230842 195916 230848 195968
rect 230900 195956 230906 195968
rect 231026 195956 231032 195968
rect 230900 195928 231032 195956
rect 230900 195916 230906 195928
rect 231026 195916 231032 195928
rect 231084 195916 231090 195968
rect 229646 193196 229652 193248
rect 229704 193236 229710 193248
rect 229830 193236 229836 193248
rect 229704 193208 229836 193236
rect 229704 193196 229710 193208
rect 229830 193196 229836 193208
rect 229888 193196 229894 193248
rect 260190 191876 260196 191888
rect 260151 191848 260196 191876
rect 260190 191836 260196 191848
rect 260248 191836 260254 191888
rect 277946 191836 277952 191888
rect 278004 191836 278010 191888
rect 243354 191808 243360 191820
rect 243315 191780 243360 191808
rect 243354 191768 243360 191780
rect 243412 191768 243418 191820
rect 270954 191808 270960 191820
rect 270915 191780 270960 191808
rect 270954 191768 270960 191780
rect 271012 191768 271018 191820
rect 277964 191740 277992 191836
rect 278038 191740 278044 191752
rect 277964 191712 278044 191740
rect 278038 191700 278044 191712
rect 278096 191700 278102 191752
rect 275281 190655 275339 190661
rect 275281 190621 275293 190655
rect 275327 190652 275339 190655
rect 275370 190652 275376 190664
rect 275327 190624 275376 190652
rect 275327 190621 275339 190624
rect 275281 190615 275339 190621
rect 275370 190612 275376 190624
rect 275428 190612 275434 190664
rect 275278 190516 275284 190528
rect 275239 190488 275284 190516
rect 275278 190476 275284 190488
rect 275336 190476 275342 190528
rect 277762 190408 277768 190460
rect 277820 190448 277826 190460
rect 278038 190448 278044 190460
rect 277820 190420 278044 190448
rect 277820 190408 277826 190420
rect 278038 190408 278044 190420
rect 278096 190408 278102 190460
rect 230842 186328 230848 186380
rect 230900 186368 230906 186380
rect 231026 186368 231032 186380
rect 230900 186340 231032 186368
rect 230900 186328 230906 186340
rect 231026 186328 231032 186340
rect 231084 186328 231090 186380
rect 237558 186328 237564 186380
rect 237616 186328 237622 186380
rect 275278 186328 275284 186380
rect 275336 186328 275342 186380
rect 237576 186232 237604 186328
rect 243357 186303 243415 186309
rect 243357 186269 243369 186303
rect 243403 186300 243415 186303
rect 243446 186300 243452 186312
rect 243403 186272 243452 186300
rect 243403 186269 243415 186272
rect 243357 186263 243415 186269
rect 243446 186260 243452 186272
rect 243504 186260 243510 186312
rect 259914 186260 259920 186312
rect 259972 186300 259978 186312
rect 260098 186300 260104 186312
rect 259972 186272 260104 186300
rect 259972 186260 259978 186272
rect 260098 186260 260104 186272
rect 260156 186260 260162 186312
rect 237650 186232 237656 186244
rect 237576 186204 237656 186232
rect 237650 186192 237656 186204
rect 237708 186192 237714 186244
rect 275296 186232 275324 186328
rect 278222 186260 278228 186312
rect 278280 186300 278286 186312
rect 278406 186300 278412 186312
rect 278280 186272 278412 186300
rect 278280 186260 278286 186272
rect 278406 186260 278412 186272
rect 278464 186260 278470 186312
rect 275370 186232 275376 186244
rect 275296 186204 275376 186232
rect 275370 186192 275376 186204
rect 275428 186192 275434 186244
rect 260282 183512 260288 183524
rect 260243 183484 260288 183512
rect 260282 183472 260288 183484
rect 260340 183472 260346 183524
rect 270954 182220 270960 182232
rect 270915 182192 270960 182220
rect 270954 182180 270960 182192
rect 271012 182180 271018 182232
rect 241146 182112 241152 182164
rect 241204 182152 241210 182164
rect 241330 182152 241336 182164
rect 241204 182124 241336 182152
rect 241204 182112 241210 182124
rect 241330 182112 241336 182124
rect 241388 182112 241394 182164
rect 308398 182112 308404 182164
rect 308456 182152 308462 182164
rect 580166 182152 580172 182164
rect 308456 182124 580172 182152
rect 308456 182112 308462 182124
rect 580166 182112 580172 182124
rect 580224 182112 580230 182164
rect 243449 182087 243507 182093
rect 243449 182053 243461 182087
rect 243495 182084 243507 182087
rect 243538 182084 243544 182096
rect 243495 182056 243544 182084
rect 243495 182053 243507 182056
rect 243449 182047 243507 182053
rect 243538 182044 243544 182056
rect 243596 182044 243602 182096
rect 3234 180752 3240 180804
rect 3292 180792 3298 180804
rect 207658 180792 207664 180804
rect 3292 180764 207664 180792
rect 3292 180752 3298 180764
rect 207658 180752 207664 180764
rect 207716 180752 207722 180804
rect 258626 180792 258632 180804
rect 258587 180764 258632 180792
rect 258626 180752 258632 180764
rect 258684 180752 258690 180804
rect 259270 180752 259276 180804
rect 259328 180792 259334 180804
rect 259362 180792 259368 180804
rect 259328 180764 259368 180792
rect 259328 180752 259334 180764
rect 259362 180752 259368 180764
rect 259420 180752 259426 180804
rect 270773 180795 270831 180801
rect 270773 180761 270785 180795
rect 270819 180792 270831 180795
rect 270954 180792 270960 180804
rect 270819 180764 270960 180792
rect 270819 180761 270831 180764
rect 270773 180755 270831 180761
rect 270954 180752 270960 180764
rect 271012 180752 271018 180804
rect 275189 180795 275247 180801
rect 275189 180761 275201 180795
rect 275235 180792 275247 180795
rect 275370 180792 275376 180804
rect 275235 180764 275376 180792
rect 275235 180761 275247 180764
rect 275189 180755 275247 180761
rect 275370 180752 275376 180764
rect 275428 180752 275434 180804
rect 259914 178712 259920 178764
rect 259972 178752 259978 178764
rect 260098 178752 260104 178764
rect 259972 178724 260104 178752
rect 259972 178712 259978 178724
rect 260098 178712 260104 178724
rect 260156 178712 260162 178764
rect 260282 178752 260288 178764
rect 260243 178724 260288 178752
rect 260282 178712 260288 178724
rect 260340 178712 260346 178764
rect 230842 176604 230848 176656
rect 230900 176644 230906 176656
rect 231026 176644 231032 176656
rect 230900 176616 231032 176644
rect 230900 176604 230906 176616
rect 231026 176604 231032 176616
rect 231084 176604 231090 176656
rect 243446 174400 243452 174412
rect 243407 174372 243452 174400
rect 243446 174360 243452 174372
rect 243504 174360 243510 174412
rect 237558 173952 237564 174004
rect 237616 173992 237622 174004
rect 237650 173992 237656 174004
rect 237616 173964 237656 173992
rect 237616 173952 237622 173964
rect 237650 173952 237656 173964
rect 237708 173952 237714 174004
rect 256513 173995 256571 174001
rect 256513 173961 256525 173995
rect 256559 173992 256571 173995
rect 256602 173992 256608 174004
rect 256559 173964 256608 173992
rect 256559 173961 256571 173964
rect 256513 173955 256571 173961
rect 256602 173952 256608 173964
rect 256660 173952 256666 174004
rect 229646 173884 229652 173936
rect 229704 173924 229710 173936
rect 229830 173924 229836 173936
rect 229704 173896 229836 173924
rect 229704 173884 229710 173896
rect 229830 173884 229836 173896
rect 229888 173884 229894 173936
rect 253934 173884 253940 173936
rect 253992 173884 253998 173936
rect 253952 173856 253980 173884
rect 254118 173856 254124 173868
rect 253952 173828 254124 173856
rect 254118 173816 254124 173828
rect 254176 173816 254182 173868
rect 237558 172496 237564 172508
rect 237519 172468 237564 172496
rect 237558 172456 237564 172468
rect 237616 172456 237622 172508
rect 238202 172496 238208 172508
rect 238163 172468 238208 172496
rect 238202 172456 238208 172468
rect 238260 172456 238266 172508
rect 258626 171204 258632 171216
rect 258587 171176 258632 171204
rect 258626 171164 258632 171176
rect 258684 171164 258690 171216
rect 270770 171136 270776 171148
rect 270731 171108 270776 171136
rect 270770 171096 270776 171108
rect 270828 171096 270834 171148
rect 275186 171136 275192 171148
rect 275147 171108 275192 171136
rect 275186 171096 275192 171108
rect 275244 171096 275250 171148
rect 277854 171096 277860 171148
rect 277912 171136 277918 171148
rect 277946 171136 277952 171148
rect 277912 171108 277952 171136
rect 277912 171096 277918 171108
rect 277946 171096 277952 171108
rect 278004 171096 278010 171148
rect 251634 171028 251640 171080
rect 251692 171068 251698 171080
rect 251818 171068 251824 171080
rect 251692 171040 251824 171068
rect 251692 171028 251698 171040
rect 251818 171028 251824 171040
rect 251876 171028 251882 171080
rect 258626 171068 258632 171080
rect 258587 171040 258632 171068
rect 258626 171028 258632 171040
rect 258684 171028 258690 171080
rect 259362 171068 259368 171080
rect 259323 171040 259368 171068
rect 259362 171028 259368 171040
rect 259420 171028 259426 171080
rect 485038 171028 485044 171080
rect 485096 171068 485102 171080
rect 580166 171068 580172 171080
rect 485096 171040 580172 171068
rect 485096 171028 485102 171040
rect 580166 171028 580172 171040
rect 580224 171028 580230 171080
rect 275186 171000 275192 171012
rect 275147 170972 275192 171000
rect 275186 170960 275192 170972
rect 275244 170960 275250 171012
rect 256510 169776 256516 169788
rect 256471 169748 256516 169776
rect 256510 169736 256516 169748
rect 256568 169736 256574 169788
rect 230842 167016 230848 167068
rect 230900 167056 230906 167068
rect 231026 167056 231032 167068
rect 230900 167028 231032 167056
rect 230900 167016 230906 167028
rect 231026 167016 231032 167028
rect 231084 167016 231090 167068
rect 243446 167016 243452 167068
rect 243504 167016 243510 167068
rect 237558 166988 237564 167000
rect 237519 166960 237564 166988
rect 237558 166948 237564 166960
rect 237616 166948 237622 167000
rect 243464 166920 243492 167016
rect 243538 166920 243544 166932
rect 243464 166892 243544 166920
rect 243538 166880 243544 166892
rect 243596 166880 243602 166932
rect 3510 165520 3516 165572
rect 3568 165560 3574 165572
rect 222838 165560 222844 165572
rect 3568 165532 222844 165560
rect 3568 165520 3574 165532
rect 222838 165520 222844 165532
rect 222896 165520 222902 165572
rect 229554 164160 229560 164212
rect 229612 164200 229618 164212
rect 229830 164200 229836 164212
rect 229612 164172 229836 164200
rect 229612 164160 229618 164172
rect 229830 164160 229836 164172
rect 229888 164160 229894 164212
rect 260098 164160 260104 164212
rect 260156 164200 260162 164212
rect 260190 164200 260196 164212
rect 260156 164172 260196 164200
rect 260156 164160 260162 164172
rect 260190 164160 260196 164172
rect 260248 164160 260254 164212
rect 260282 164160 260288 164212
rect 260340 164200 260346 164212
rect 260374 164200 260380 164212
rect 260340 164172 260380 164200
rect 260340 164160 260346 164172
rect 260374 164160 260380 164172
rect 260432 164160 260438 164212
rect 238202 162908 238208 162920
rect 238163 162880 238208 162908
rect 238202 162868 238208 162880
rect 238260 162868 238266 162920
rect 237558 162800 237564 162852
rect 237616 162840 237622 162852
rect 237650 162840 237656 162852
rect 237616 162812 237656 162840
rect 237616 162800 237622 162812
rect 237650 162800 237656 162812
rect 237708 162800 237714 162852
rect 238938 162800 238944 162852
rect 238996 162840 239002 162852
rect 239122 162840 239128 162852
rect 238996 162812 239128 162840
rect 238996 162800 239002 162812
rect 239122 162800 239128 162812
rect 239180 162800 239186 162852
rect 241146 162840 241152 162852
rect 241107 162812 241152 162840
rect 241146 162800 241152 162812
rect 241204 162800 241210 162852
rect 260190 162840 260196 162852
rect 260151 162812 260196 162840
rect 260190 162800 260196 162812
rect 260248 162800 260254 162852
rect 259362 161548 259368 161560
rect 259323 161520 259368 161548
rect 259362 161508 259368 161520
rect 259420 161508 259426 161560
rect 258626 161480 258632 161492
rect 258587 161452 258632 161480
rect 258626 161440 258632 161452
rect 258684 161440 258690 161492
rect 275189 161483 275247 161489
rect 275189 161449 275201 161483
rect 275235 161480 275247 161483
rect 275370 161480 275376 161492
rect 275235 161452 275376 161480
rect 275235 161449 275247 161452
rect 275189 161443 275247 161449
rect 275370 161440 275376 161452
rect 275428 161440 275434 161492
rect 277854 161440 277860 161492
rect 277912 161480 277918 161492
rect 278130 161480 278136 161492
rect 277912 161452 278136 161480
rect 277912 161440 277918 161452
rect 278130 161440 278136 161452
rect 278188 161440 278194 161492
rect 259273 160055 259331 160061
rect 259273 160021 259285 160055
rect 259319 160052 259331 160055
rect 259362 160052 259368 160064
rect 259319 160024 259368 160052
rect 259319 160021 259331 160024
rect 259273 160015 259331 160021
rect 259362 160012 259368 160024
rect 259420 160012 259426 160064
rect 297450 158652 297456 158704
rect 297508 158692 297514 158704
rect 579798 158692 579804 158704
rect 297508 158664 579804 158692
rect 297508 158652 297514 158664
rect 579798 158652 579804 158664
rect 579856 158652 579862 158704
rect 243449 157403 243507 157409
rect 243449 157369 243461 157403
rect 243495 157400 243507 157403
rect 243538 157400 243544 157412
rect 243495 157372 243544 157400
rect 243495 157369 243507 157372
rect 243449 157363 243507 157369
rect 243538 157360 243544 157372
rect 243596 157360 243602 157412
rect 230842 157292 230848 157344
rect 230900 157332 230906 157344
rect 231026 157332 231032 157344
rect 230900 157304 231032 157332
rect 230900 157292 230906 157304
rect 231026 157292 231032 157304
rect 231084 157292 231090 157344
rect 260374 154680 260380 154692
rect 260300 154652 260380 154680
rect 260300 154556 260328 154652
rect 260374 154640 260380 154652
rect 260432 154640 260438 154692
rect 260282 154504 260288 154556
rect 260340 154504 260346 154556
rect 243446 153320 243452 153332
rect 243407 153292 243452 153320
rect 243446 153280 243452 153292
rect 243504 153280 243510 153332
rect 260190 153320 260196 153332
rect 260151 153292 260196 153320
rect 260190 153280 260196 153292
rect 260248 153280 260254 153332
rect 241146 153252 241152 153264
rect 241107 153224 241152 153252
rect 241146 153212 241152 153224
rect 241204 153212 241210 153264
rect 237558 153184 237564 153196
rect 237519 153156 237564 153184
rect 237558 153144 237564 153156
rect 237616 153144 237622 153196
rect 238202 153184 238208 153196
rect 238163 153156 238208 153184
rect 238202 153144 238208 153156
rect 238260 153144 238266 153196
rect 238938 153184 238944 153196
rect 238899 153156 238944 153184
rect 238938 153144 238944 153156
rect 238996 153144 239002 153196
rect 251726 151784 251732 151836
rect 251784 151824 251790 151836
rect 251818 151824 251824 151836
rect 251784 151796 251824 151824
rect 251784 151784 251790 151796
rect 251818 151784 251824 151796
rect 251876 151784 251882 151836
rect 253934 151784 253940 151836
rect 253992 151824 253998 151836
rect 254118 151824 254124 151836
rect 253992 151796 254124 151824
rect 253992 151784 253998 151796
rect 254118 151784 254124 151796
rect 254176 151784 254182 151836
rect 256602 151784 256608 151836
rect 256660 151824 256666 151836
rect 256878 151824 256884 151836
rect 256660 151796 256884 151824
rect 256660 151784 256666 151796
rect 256878 151784 256884 151796
rect 256936 151784 256942 151836
rect 258626 151756 258632 151768
rect 258587 151728 258632 151756
rect 258626 151716 258632 151728
rect 258684 151716 258690 151768
rect 256421 149039 256479 149045
rect 256421 149005 256433 149039
rect 256467 149036 256479 149039
rect 256786 149036 256792 149048
rect 256467 149008 256792 149036
rect 256467 149005 256479 149008
rect 256421 148999 256479 149005
rect 256786 148996 256792 149008
rect 256844 148996 256850 149048
rect 243446 147704 243452 147756
rect 243504 147704 243510 147756
rect 243464 147620 243492 147704
rect 278130 147636 278136 147688
rect 278188 147676 278194 147688
rect 278314 147676 278320 147688
rect 278188 147648 278320 147676
rect 278188 147636 278194 147648
rect 278314 147636 278320 147648
rect 278372 147636 278378 147688
rect 237558 147608 237564 147620
rect 237519 147580 237564 147608
rect 237558 147568 237564 147580
rect 237616 147568 237622 147620
rect 243446 147568 243452 147620
rect 243504 147568 243510 147620
rect 238938 147200 238944 147212
rect 238899 147172 238944 147200
rect 238938 147160 238944 147172
rect 238996 147160 239002 147212
rect 260098 144848 260104 144900
rect 260156 144888 260162 144900
rect 260190 144888 260196 144900
rect 260156 144860 260196 144888
rect 260156 144848 260162 144860
rect 260190 144848 260196 144860
rect 260248 144848 260254 144900
rect 260282 144848 260288 144900
rect 260340 144888 260346 144900
rect 260374 144888 260380 144900
rect 260340 144860 260380 144888
rect 260340 144848 260346 144860
rect 260374 144848 260380 144860
rect 260432 144848 260438 144900
rect 276474 144888 276480 144900
rect 276435 144860 276480 144888
rect 276474 144848 276480 144860
rect 276532 144848 276538 144900
rect 238202 143596 238208 143608
rect 238163 143568 238208 143596
rect 238202 143556 238208 143568
rect 238260 143556 238266 143608
rect 237561 143463 237619 143469
rect 237561 143429 237573 143463
rect 237607 143460 237619 143463
rect 237650 143460 237656 143472
rect 237607 143432 237656 143460
rect 237607 143429 237619 143432
rect 237561 143423 237619 143429
rect 237650 143420 237656 143432
rect 237708 143420 237714 143472
rect 258626 142168 258632 142180
rect 258587 142140 258632 142168
rect 258626 142128 258632 142140
rect 258684 142128 258690 142180
rect 259270 142168 259276 142180
rect 259231 142140 259276 142168
rect 259270 142128 259276 142140
rect 259328 142128 259334 142180
rect 275370 142128 275376 142180
rect 275428 142168 275434 142180
rect 275462 142168 275468 142180
rect 275428 142140 275468 142168
rect 275428 142128 275434 142140
rect 275462 142128 275468 142140
rect 275520 142128 275526 142180
rect 243449 142103 243507 142109
rect 243449 142069 243461 142103
rect 243495 142100 243507 142103
rect 243538 142100 243544 142112
rect 243495 142072 243544 142100
rect 243495 142069 243507 142072
rect 243449 142063 243507 142069
rect 243538 142060 243544 142072
rect 243596 142060 243602 142112
rect 254029 142103 254087 142109
rect 254029 142069 254041 142103
rect 254075 142100 254087 142103
rect 254118 142100 254124 142112
rect 254075 142072 254124 142100
rect 254075 142069 254087 142072
rect 254029 142063 254087 142069
rect 254118 142060 254124 142072
rect 254176 142060 254182 142112
rect 256418 139448 256424 139460
rect 256379 139420 256424 139448
rect 256418 139408 256424 139420
rect 256476 139408 256482 139460
rect 260098 138660 260104 138712
rect 260156 138700 260162 138712
rect 260374 138700 260380 138712
rect 260156 138672 260380 138700
rect 260156 138660 260162 138672
rect 260374 138660 260380 138672
rect 260432 138660 260438 138712
rect 229554 137980 229560 138032
rect 229612 137980 229618 138032
rect 229462 137912 229468 137964
rect 229520 137952 229526 137964
rect 229572 137952 229600 137980
rect 229520 137924 229600 137952
rect 229520 137912 229526 137924
rect 251637 137139 251695 137145
rect 251637 137105 251649 137139
rect 251683 137136 251695 137139
rect 251726 137136 251732 137148
rect 251683 137108 251732 137136
rect 251683 137105 251695 137108
rect 251637 137099 251695 137105
rect 251726 137096 251732 137108
rect 251784 137096 251790 137148
rect 3510 136552 3516 136604
rect 3568 136592 3574 136604
rect 227070 136592 227076 136604
rect 3568 136564 227076 136592
rect 3568 136552 3574 136564
rect 227070 136552 227076 136564
rect 227128 136552 227134 136604
rect 275462 135300 275468 135312
rect 275388 135272 275468 135300
rect 275388 135244 275416 135272
rect 275462 135260 275468 135272
rect 275520 135260 275526 135312
rect 276474 135260 276480 135312
rect 276532 135300 276538 135312
rect 276532 135272 276577 135300
rect 276532 135260 276538 135272
rect 275370 135192 275376 135244
rect 275428 135192 275434 135244
rect 278130 135232 278136 135244
rect 278091 135204 278136 135232
rect 278130 135192 278136 135204
rect 278188 135192 278194 135244
rect 496078 135192 496084 135244
rect 496136 135232 496142 135244
rect 580166 135232 580172 135244
rect 496136 135204 580172 135232
rect 496136 135192 496142 135204
rect 580166 135192 580172 135204
rect 580224 135192 580230 135244
rect 281442 134512 281448 134564
rect 281500 134552 281506 134564
rect 495434 134552 495440 134564
rect 281500 134524 495440 134552
rect 281500 134512 281506 134524
rect 495434 134512 495440 134524
rect 495492 134512 495498 134564
rect 237558 134008 237564 134020
rect 237519 133980 237564 134008
rect 237558 133968 237564 133980
rect 237616 133968 237622 134020
rect 238110 133872 238116 133884
rect 238071 133844 238116 133872
rect 238110 133832 238116 133844
rect 238168 133832 238174 133884
rect 238662 133832 238668 133884
rect 238720 133872 238726 133884
rect 238938 133872 238944 133884
rect 238720 133844 238944 133872
rect 238720 133832 238726 133844
rect 238938 133832 238944 133844
rect 238996 133832 239002 133884
rect 260282 133872 260288 133884
rect 260243 133844 260288 133872
rect 260282 133832 260288 133844
rect 260340 133832 260346 133884
rect 275370 133872 275376 133884
rect 275331 133844 275376 133872
rect 275370 133832 275376 133844
rect 275428 133832 275434 133884
rect 251634 132512 251640 132524
rect 251595 132484 251640 132512
rect 251634 132472 251640 132484
rect 251692 132472 251698 132524
rect 254026 132512 254032 132524
rect 253987 132484 254032 132512
rect 254026 132472 254032 132484
rect 254084 132472 254090 132524
rect 258534 131084 258540 131096
rect 258495 131056 258540 131084
rect 258534 131044 258540 131056
rect 258592 131044 258598 131096
rect 278133 128299 278191 128305
rect 278133 128265 278145 128299
rect 278179 128296 278191 128299
rect 278222 128296 278228 128308
rect 278179 128268 278228 128296
rect 278179 128265 278191 128268
rect 278133 128259 278191 128265
rect 278222 128256 278228 128268
rect 278280 128256 278286 128308
rect 260098 125604 260104 125656
rect 260156 125644 260162 125656
rect 260190 125644 260196 125656
rect 260156 125616 260196 125644
rect 260156 125604 260162 125616
rect 260190 125604 260196 125616
rect 260248 125604 260254 125656
rect 272334 125536 272340 125588
rect 272392 125576 272398 125588
rect 272426 125576 272432 125588
rect 272392 125548 272432 125576
rect 272392 125536 272398 125548
rect 272426 125536 272432 125548
rect 272484 125536 272490 125588
rect 251634 124244 251640 124296
rect 251692 124244 251698 124296
rect 260282 124284 260288 124296
rect 260243 124256 260288 124284
rect 260282 124244 260288 124256
rect 260340 124244 260346 124296
rect 243446 124216 243452 124228
rect 243407 124188 243452 124216
rect 243446 124176 243452 124188
rect 243504 124176 243510 124228
rect 241054 124148 241060 124160
rect 241015 124120 241060 124148
rect 241054 124108 241060 124120
rect 241112 124108 241118 124160
rect 251652 124080 251680 124244
rect 253934 124176 253940 124228
rect 253992 124216 253998 124228
rect 254026 124216 254032 124228
rect 253992 124188 254032 124216
rect 253992 124176 253998 124188
rect 254026 124176 254032 124188
rect 254084 124176 254090 124228
rect 275370 124216 275376 124228
rect 275331 124188 275376 124216
rect 275370 124176 275376 124188
rect 275428 124176 275434 124228
rect 260098 124148 260104 124160
rect 260059 124120 260104 124148
rect 260098 124108 260104 124120
rect 260156 124108 260162 124160
rect 260282 124148 260288 124160
rect 260243 124120 260288 124148
rect 260282 124108 260288 124120
rect 260340 124108 260346 124160
rect 272426 124108 272432 124160
rect 272484 124148 272490 124160
rect 272610 124148 272616 124160
rect 272484 124120 272616 124148
rect 272484 124108 272490 124120
rect 272610 124108 272616 124120
rect 272668 124108 272674 124160
rect 309778 124108 309784 124160
rect 309836 124148 309842 124160
rect 580166 124148 580172 124160
rect 309836 124120 580172 124148
rect 309836 124108 309842 124120
rect 580166 124108 580172 124120
rect 580224 124108 580230 124160
rect 251726 124080 251732 124092
rect 251652 124052 251732 124080
rect 251726 124040 251732 124052
rect 251784 124040 251790 124092
rect 238110 122856 238116 122868
rect 238071 122828 238116 122856
rect 238110 122816 238116 122828
rect 238168 122816 238174 122868
rect 2958 122748 2964 122800
rect 3016 122788 3022 122800
rect 218698 122788 218704 122800
rect 3016 122760 218704 122788
rect 3016 122748 3022 122760
rect 218698 122748 218704 122760
rect 218756 122748 218762 122800
rect 253934 122788 253940 122800
rect 253895 122760 253940 122788
rect 253934 122748 253940 122760
rect 253992 122748 253998 122800
rect 256510 122788 256516 122800
rect 256471 122760 256516 122788
rect 256510 122748 256516 122760
rect 256568 122748 256574 122800
rect 259270 122748 259276 122800
rect 259328 122748 259334 122800
rect 259288 122720 259316 122748
rect 259362 122720 259368 122732
rect 259288 122692 259368 122720
rect 259362 122680 259368 122692
rect 259420 122680 259426 122732
rect 219250 122068 219256 122120
rect 219308 122108 219314 122120
rect 252186 122108 252192 122120
rect 219308 122080 252192 122108
rect 219308 122068 219314 122080
rect 252186 122068 252192 122080
rect 252244 122068 252250 122120
rect 258537 121499 258595 121505
rect 258537 121465 258549 121499
rect 258583 121496 258595 121499
rect 258626 121496 258632 121508
rect 258583 121468 258632 121496
rect 258583 121465 258595 121468
rect 258537 121459 258595 121465
rect 258626 121456 258632 121468
rect 258684 121456 258690 121508
rect 238021 121431 238079 121437
rect 238021 121397 238033 121431
rect 238067 121428 238079 121431
rect 238110 121428 238116 121440
rect 238067 121400 238116 121428
rect 238067 121397 238079 121400
rect 238021 121391 238079 121397
rect 238110 121388 238116 121400
rect 238168 121388 238174 121440
rect 238757 121431 238815 121437
rect 238757 121397 238769 121431
rect 238803 121428 238815 121431
rect 238846 121428 238852 121440
rect 238803 121400 238852 121428
rect 238803 121397 238815 121400
rect 238757 121391 238815 121397
rect 238846 121388 238852 121400
rect 238904 121388 238910 121440
rect 272429 121431 272487 121437
rect 272429 121397 272441 121431
rect 272475 121428 272487 121431
rect 272610 121428 272616 121440
rect 272475 121400 272616 121428
rect 272475 121397 272487 121400
rect 272429 121391 272487 121397
rect 272610 121388 272616 121400
rect 272668 121388 272674 121440
rect 276477 119391 276535 119397
rect 276477 119357 276489 119391
rect 276523 119388 276535 119391
rect 276566 119388 276572 119400
rect 276523 119360 276572 119388
rect 276523 119357 276535 119360
rect 276477 119351 276535 119357
rect 276566 119348 276572 119360
rect 276624 119348 276630 119400
rect 243446 118872 243452 118924
rect 243504 118912 243510 118924
rect 243541 118915 243599 118921
rect 243541 118912 243553 118915
rect 243504 118884 243553 118912
rect 243504 118872 243510 118884
rect 243541 118881 243553 118884
rect 243587 118881 243599 118915
rect 243541 118875 243599 118881
rect 229554 118668 229560 118720
rect 229612 118668 229618 118720
rect 270954 118668 270960 118720
rect 271012 118668 271018 118720
rect 229462 118600 229468 118652
rect 229520 118640 229526 118652
rect 229572 118640 229600 118668
rect 229520 118612 229600 118640
rect 229520 118600 229526 118612
rect 270972 118584 271000 118668
rect 270954 118532 270960 118584
rect 271012 118532 271018 118584
rect 238757 115379 238815 115385
rect 238757 115345 238769 115379
rect 238803 115376 238815 115379
rect 238846 115376 238852 115388
rect 238803 115348 238852 115376
rect 238803 115345 238815 115348
rect 238757 115339 238815 115345
rect 238846 115336 238852 115348
rect 238904 115336 238910 115388
rect 241057 114563 241115 114569
rect 241057 114529 241069 114563
rect 241103 114560 241115 114563
rect 241146 114560 241152 114572
rect 241103 114532 241152 114560
rect 241103 114529 241115 114532
rect 241057 114523 241115 114529
rect 241146 114520 241152 114532
rect 241204 114520 241210 114572
rect 260101 114563 260159 114569
rect 260101 114529 260113 114563
rect 260147 114560 260159 114563
rect 260190 114560 260196 114572
rect 260147 114532 260196 114560
rect 260147 114529 260159 114532
rect 260101 114523 260159 114529
rect 260190 114520 260196 114532
rect 260248 114520 260254 114572
rect 260285 114563 260343 114569
rect 260285 114529 260297 114563
rect 260331 114560 260343 114563
rect 260374 114560 260380 114572
rect 260331 114532 260380 114560
rect 260331 114529 260343 114532
rect 260285 114523 260343 114529
rect 260374 114520 260380 114532
rect 260432 114520 260438 114572
rect 278222 114520 278228 114572
rect 278280 114560 278286 114572
rect 278280 114532 278452 114560
rect 278280 114520 278286 114532
rect 278317 114495 278375 114501
rect 278317 114461 278329 114495
rect 278363 114492 278375 114495
rect 278424 114492 278452 114532
rect 278363 114464 278452 114492
rect 278363 114461 278375 114464
rect 278317 114455 278375 114461
rect 237558 113160 237564 113212
rect 237616 113200 237622 113212
rect 237650 113200 237656 113212
rect 237616 113172 237656 113200
rect 237616 113160 237622 113172
rect 237650 113160 237656 113172
rect 237708 113160 237714 113212
rect 256513 113203 256571 113209
rect 256513 113169 256525 113203
rect 256559 113200 256571 113203
rect 256602 113200 256608 113212
rect 256559 113172 256608 113200
rect 256559 113169 256571 113172
rect 256513 113163 256571 113169
rect 256602 113160 256608 113172
rect 256660 113160 256666 113212
rect 238021 113135 238079 113141
rect 238021 113101 238033 113135
rect 238067 113132 238079 113135
rect 238110 113132 238116 113144
rect 238067 113104 238116 113132
rect 238067 113101 238079 113104
rect 238021 113095 238079 113101
rect 238110 113092 238116 113104
rect 238168 113092 238174 113144
rect 253937 111843 253995 111849
rect 253937 111809 253949 111843
rect 253983 111840 253995 111843
rect 254118 111840 254124 111852
rect 253983 111812 254124 111840
rect 253983 111809 253995 111812
rect 253937 111803 253995 111809
rect 254118 111800 254124 111812
rect 254176 111800 254182 111852
rect 272426 111840 272432 111852
rect 272387 111812 272432 111840
rect 272426 111800 272432 111812
rect 272484 111800 272490 111852
rect 258626 111772 258632 111784
rect 258587 111744 258632 111772
rect 258626 111732 258632 111744
rect 258684 111732 258690 111784
rect 291930 111732 291936 111784
rect 291988 111772 291994 111784
rect 579798 111772 579804 111784
rect 291988 111744 579804 111772
rect 291988 111732 291994 111744
rect 579798 111732 579804 111744
rect 579856 111732 579862 111784
rect 272337 111707 272395 111713
rect 272337 111673 272349 111707
rect 272383 111704 272395 111707
rect 272426 111704 272432 111716
rect 272383 111676 272432 111704
rect 272383 111673 272395 111676
rect 272337 111667 272395 111673
rect 272426 111664 272432 111676
rect 272484 111664 272490 111716
rect 251729 110415 251787 110421
rect 251729 110381 251741 110415
rect 251775 110412 251787 110415
rect 251818 110412 251824 110424
rect 251775 110384 251824 110412
rect 251775 110381 251787 110384
rect 251729 110375 251787 110381
rect 251818 110372 251824 110384
rect 251876 110372 251882 110424
rect 243538 108984 243544 108996
rect 243499 108956 243544 108984
rect 243538 108944 243544 108956
rect 243596 108944 243602 108996
rect 276474 107624 276480 107636
rect 276435 107596 276480 107624
rect 276474 107584 276480 107596
rect 276532 107584 276538 107636
rect 238846 106292 238852 106344
rect 238904 106292 238910 106344
rect 238864 106208 238892 106292
rect 249058 106224 249064 106276
rect 249116 106224 249122 106276
rect 238846 106156 238852 106208
rect 238904 106156 238910 106208
rect 248966 106196 248972 106208
rect 248927 106168 248972 106196
rect 248966 106156 248972 106168
rect 249024 106156 249030 106208
rect 249076 106140 249104 106224
rect 249150 106156 249156 106208
rect 249208 106156 249214 106208
rect 249058 106088 249064 106140
rect 249116 106088 249122 106140
rect 249168 106072 249196 106156
rect 249150 106020 249156 106072
rect 249208 106020 249214 106072
rect 278314 104904 278320 104916
rect 278275 104876 278320 104904
rect 278314 104864 278320 104876
rect 278372 104864 278378 104916
rect 253934 103572 253940 103624
rect 253992 103612 253998 103624
rect 254118 103612 254124 103624
rect 253992 103584 254124 103612
rect 253992 103572 253998 103584
rect 254118 103572 254124 103584
rect 254176 103572 254182 103624
rect 238110 103504 238116 103556
rect 238168 103544 238174 103556
rect 238202 103544 238208 103556
rect 238168 103516 238208 103544
rect 238168 103504 238174 103516
rect 238202 103504 238208 103516
rect 238260 103504 238266 103556
rect 258626 102184 258632 102196
rect 258587 102156 258632 102184
rect 258626 102144 258632 102156
rect 258684 102144 258690 102196
rect 272334 102184 272340 102196
rect 272295 102156 272340 102184
rect 272334 102144 272340 102156
rect 272392 102144 272398 102196
rect 238113 102119 238171 102125
rect 238113 102085 238125 102119
rect 238159 102116 238171 102119
rect 238202 102116 238208 102128
rect 238159 102088 238208 102116
rect 238159 102085 238171 102088
rect 238113 102079 238171 102085
rect 238202 102076 238208 102088
rect 238260 102076 238266 102128
rect 260098 102116 260104 102128
rect 260059 102088 260104 102116
rect 260098 102076 260104 102088
rect 260156 102076 260162 102128
rect 243538 101396 243544 101448
rect 243596 101396 243602 101448
rect 243556 101312 243584 101396
rect 243538 101260 243544 101312
rect 243596 101260 243602 101312
rect 251726 100756 251732 100768
rect 251687 100728 251732 100756
rect 251726 100716 251732 100728
rect 251784 100716 251790 100768
rect 229554 99356 229560 99408
rect 229612 99356 229618 99408
rect 237650 99396 237656 99408
rect 237576 99368 237656 99396
rect 229462 99288 229468 99340
rect 229520 99328 229526 99340
rect 229572 99328 229600 99356
rect 237576 99340 237604 99368
rect 237650 99356 237656 99368
rect 237708 99356 237714 99408
rect 260282 99356 260288 99408
rect 260340 99356 260346 99408
rect 229520 99300 229600 99328
rect 229520 99288 229526 99300
rect 237558 99288 237564 99340
rect 237616 99288 237622 99340
rect 260300 99328 260328 99356
rect 260374 99328 260380 99340
rect 260300 99300 260380 99328
rect 260374 99288 260380 99300
rect 260432 99288 260438 99340
rect 248966 97832 248972 97844
rect 248927 97804 248972 97832
rect 248966 97792 248972 97804
rect 249024 97792 249030 97844
rect 258537 97291 258595 97297
rect 258537 97257 258549 97291
rect 258583 97288 258595 97291
rect 258626 97288 258632 97300
rect 258583 97260 258632 97288
rect 258583 97257 258595 97260
rect 258537 97251 258595 97257
rect 258626 97248 258632 97260
rect 258684 97248 258690 97300
rect 272337 97291 272395 97297
rect 272337 97257 272349 97291
rect 272383 97288 272395 97291
rect 272426 97288 272432 97300
rect 272383 97260 272432 97288
rect 272383 97257 272395 97260
rect 272337 97251 272395 97257
rect 272426 97248 272432 97260
rect 272484 97248 272490 97300
rect 253842 95248 253848 95260
rect 253803 95220 253848 95248
rect 253842 95208 253848 95220
rect 253900 95208 253906 95260
rect 237558 95180 237564 95192
rect 237519 95152 237564 95180
rect 237558 95140 237564 95152
rect 237616 95140 237622 95192
rect 238846 95140 238852 95192
rect 238904 95140 238910 95192
rect 238864 95112 238892 95140
rect 238938 95112 238944 95124
rect 238864 95084 238944 95112
rect 238938 95072 238944 95084
rect 238996 95072 239002 95124
rect 3510 93780 3516 93832
rect 3568 93820 3574 93832
rect 204898 93820 204904 93832
rect 3568 93792 204904 93820
rect 3568 93780 3574 93792
rect 204898 93780 204904 93792
rect 204956 93780 204962 93832
rect 275278 93820 275284 93832
rect 275239 93792 275284 93820
rect 275278 93780 275284 93792
rect 275336 93780 275342 93832
rect 238110 92528 238116 92540
rect 238071 92500 238116 92528
rect 238110 92488 238116 92500
rect 238168 92488 238174 92540
rect 260101 92531 260159 92537
rect 260101 92497 260113 92531
rect 260147 92528 260159 92531
rect 260190 92528 260196 92540
rect 260147 92500 260196 92528
rect 260147 92497 260159 92500
rect 260101 92491 260159 92497
rect 260190 92488 260196 92500
rect 260248 92488 260254 92540
rect 253842 91100 253848 91112
rect 253803 91072 253848 91100
rect 253842 91060 253848 91072
rect 253900 91060 253906 91112
rect 305638 88272 305644 88324
rect 305696 88312 305702 88324
rect 580166 88312 580172 88324
rect 305696 88284 580172 88312
rect 305696 88272 305702 88284
rect 580166 88272 580172 88284
rect 580224 88272 580230 88324
rect 243538 86952 243544 86964
rect 243499 86924 243544 86952
rect 243538 86912 243544 86924
rect 243596 86912 243602 86964
rect 248785 86955 248843 86961
rect 248785 86921 248797 86955
rect 248831 86952 248843 86955
rect 248874 86952 248880 86964
rect 248831 86924 248880 86952
rect 248831 86921 248843 86924
rect 248785 86915 248843 86921
rect 248874 86912 248880 86924
rect 248932 86912 248938 86964
rect 249150 86952 249156 86964
rect 249111 86924 249156 86952
rect 249150 86912 249156 86924
rect 249208 86912 249214 86964
rect 248966 86884 248972 86896
rect 248927 86856 248972 86884
rect 248966 86844 248972 86856
rect 249024 86844 249030 86896
rect 249058 86844 249064 86896
rect 249116 86844 249122 86896
rect 249076 86760 249104 86844
rect 249058 86708 249064 86760
rect 249116 86708 249122 86760
rect 260285 86547 260343 86553
rect 260285 86513 260297 86547
rect 260331 86544 260343 86547
rect 260374 86544 260380 86556
rect 260331 86516 260380 86544
rect 260331 86513 260343 86516
rect 260285 86507 260343 86513
rect 260374 86504 260380 86516
rect 260432 86504 260438 86556
rect 259362 85796 259368 85808
rect 259288 85768 259368 85796
rect 259288 85740 259316 85768
rect 259362 85756 259368 85768
rect 259420 85756 259426 85808
rect 259270 85688 259276 85740
rect 259328 85688 259334 85740
rect 237561 85595 237619 85601
rect 237561 85561 237573 85595
rect 237607 85592 237619 85595
rect 237650 85592 237656 85604
rect 237607 85564 237656 85592
rect 237607 85561 237619 85564
rect 237561 85555 237619 85561
rect 237650 85552 237656 85564
rect 237708 85552 237714 85604
rect 238110 85552 238116 85604
rect 238168 85592 238174 85604
rect 238202 85592 238208 85604
rect 238168 85564 238208 85592
rect 238168 85552 238174 85564
rect 238202 85552 238208 85564
rect 238260 85552 238266 85604
rect 253842 85552 253848 85604
rect 253900 85592 253906 85604
rect 253934 85592 253940 85604
rect 253900 85564 253940 85592
rect 253900 85552 253906 85564
rect 253934 85552 253940 85564
rect 253992 85552 253998 85604
rect 256510 85552 256516 85604
rect 256568 85592 256574 85604
rect 256694 85592 256700 85604
rect 256568 85564 256700 85592
rect 256568 85552 256574 85564
rect 256694 85552 256700 85564
rect 256752 85552 256758 85604
rect 258534 84232 258540 84244
rect 258495 84204 258540 84232
rect 258534 84192 258540 84204
rect 258592 84192 258598 84244
rect 275278 84232 275284 84244
rect 275239 84204 275284 84232
rect 275278 84192 275284 84204
rect 275336 84192 275342 84244
rect 251726 84164 251732 84176
rect 251687 84136 251732 84164
rect 251726 84124 251732 84136
rect 251784 84124 251790 84176
rect 259270 84164 259276 84176
rect 259231 84136 259276 84164
rect 259270 84124 259276 84136
rect 259328 84124 259334 84176
rect 237561 82807 237619 82813
rect 237561 82773 237573 82807
rect 237607 82804 237619 82807
rect 237650 82804 237656 82816
rect 237607 82776 237656 82804
rect 237607 82773 237619 82776
rect 237561 82767 237619 82773
rect 237650 82764 237656 82776
rect 237708 82764 237714 82816
rect 248785 82127 248843 82133
rect 248785 82093 248797 82127
rect 248831 82124 248843 82127
rect 248874 82124 248880 82136
rect 248831 82096 248880 82124
rect 248831 82093 248843 82096
rect 248785 82087 248843 82093
rect 248874 82084 248880 82096
rect 248932 82084 248938 82136
rect 229554 80152 229560 80164
rect 229515 80124 229560 80152
rect 229554 80112 229560 80124
rect 229612 80112 229618 80164
rect 253934 80152 253940 80164
rect 253895 80124 253940 80152
rect 253934 80112 253940 80124
rect 253992 80112 253998 80164
rect 256510 80044 256516 80096
rect 256568 80044 256574 80096
rect 3234 79976 3240 80028
rect 3292 80016 3298 80028
rect 215938 80016 215944 80028
rect 3292 79988 215944 80016
rect 3292 79976 3298 79988
rect 215938 79976 215944 79988
rect 215996 79976 216002 80028
rect 256528 79948 256556 80044
rect 256602 79948 256608 79960
rect 256528 79920 256608 79948
rect 256602 79908 256608 79920
rect 256660 79908 256666 79960
rect 248966 78452 248972 78464
rect 248927 78424 248972 78452
rect 248966 78412 248972 78424
rect 249024 78412 249030 78464
rect 229462 77324 229468 77376
rect 229520 77364 229526 77376
rect 229557 77367 229615 77373
rect 229557 77364 229569 77367
rect 229520 77336 229569 77364
rect 229520 77324 229526 77336
rect 229557 77333 229569 77336
rect 229603 77333 229615 77367
rect 229557 77327 229615 77333
rect 243538 77296 243544 77308
rect 243499 77268 243544 77296
rect 243538 77256 243544 77268
rect 243596 77256 243602 77308
rect 249150 77296 249156 77308
rect 249111 77268 249156 77296
rect 249150 77256 249156 77268
rect 249208 77256 249214 77308
rect 229554 77228 229560 77240
rect 229515 77200 229560 77228
rect 229554 77188 229560 77200
rect 229612 77188 229618 77240
rect 321462 76100 321468 76152
rect 321520 76140 321526 76152
rect 323026 76140 323032 76152
rect 321520 76112 323032 76140
rect 321520 76100 321526 76112
rect 323026 76100 323032 76112
rect 323084 76100 323090 76152
rect 280246 76032 280252 76084
rect 280304 76072 280310 76084
rect 289722 76072 289728 76084
rect 280304 76044 289728 76072
rect 280304 76032 280310 76044
rect 289722 76032 289728 76044
rect 289780 76032 289786 76084
rect 302142 76032 302148 76084
rect 302200 76072 302206 76084
rect 309042 76072 309048 76084
rect 302200 76044 309048 76072
rect 302200 76032 302206 76044
rect 309042 76032 309048 76044
rect 309100 76032 309106 76084
rect 437382 76032 437388 76084
rect 437440 76072 437446 76084
rect 444282 76072 444288 76084
rect 437440 76044 444288 76072
rect 437440 76032 437446 76044
rect 444282 76032 444288 76044
rect 444340 76032 444346 76084
rect 502242 76032 502248 76084
rect 502300 76072 502306 76084
rect 510522 76072 510528 76084
rect 502300 76044 510528 76072
rect 502300 76032 502306 76044
rect 510522 76032 510528 76044
rect 510580 76032 510586 76084
rect 533982 76032 533988 76084
rect 534040 76072 534046 76084
rect 540882 76072 540888 76084
rect 534040 76044 540888 76072
rect 534040 76032 534046 76044
rect 540882 76032 540888 76044
rect 540940 76032 540946 76084
rect 553302 76032 553308 76084
rect 553360 76072 553366 76084
rect 560202 76072 560208 76084
rect 553360 76044 560208 76072
rect 553360 76032 553366 76044
rect 560202 76032 560208 76044
rect 560260 76032 560266 76084
rect 572622 76032 572628 76084
rect 572680 76072 572686 76084
rect 579522 76072 579528 76084
rect 572680 76044 579528 76072
rect 572680 76032 572686 76044
rect 579522 76032 579528 76044
rect 579580 76032 579586 76084
rect 260285 75939 260343 75945
rect 260285 75905 260297 75939
rect 260331 75936 260343 75939
rect 260374 75936 260380 75948
rect 260331 75908 260380 75936
rect 260331 75905 260343 75908
rect 260285 75899 260343 75905
rect 260374 75896 260380 75908
rect 260432 75896 260438 75948
rect 253934 75868 253940 75880
rect 253895 75840 253940 75868
rect 253934 75828 253940 75840
rect 253992 75828 253998 75880
rect 251729 74579 251787 74585
rect 251729 74545 251741 74579
rect 251775 74576 251787 74579
rect 251818 74576 251824 74588
rect 251775 74548 251824 74576
rect 251775 74545 251787 74548
rect 251729 74539 251787 74545
rect 251818 74536 251824 74548
rect 251876 74536 251882 74588
rect 259273 74579 259331 74585
rect 259273 74545 259285 74579
rect 259319 74576 259331 74579
rect 259362 74576 259368 74588
rect 259319 74548 259368 74576
rect 259319 74545 259331 74548
rect 259273 74539 259331 74545
rect 259362 74536 259368 74548
rect 259420 74536 259426 74588
rect 272334 74576 272340 74588
rect 272295 74548 272340 74576
rect 272334 74536 272340 74548
rect 272392 74536 272398 74588
rect 238938 74508 238944 74520
rect 238899 74480 238944 74508
rect 238938 74468 238944 74480
rect 238996 74468 239002 74520
rect 258537 74511 258595 74517
rect 258537 74477 258549 74511
rect 258583 74508 258595 74511
rect 258626 74508 258632 74520
rect 258583 74480 258632 74508
rect 258583 74477 258595 74480
rect 258537 74471 258595 74477
rect 258626 74468 258632 74480
rect 258684 74468 258690 74520
rect 237558 73216 237564 73228
rect 237519 73188 237564 73216
rect 237558 73176 237564 73188
rect 237616 73176 237622 73228
rect 229557 67643 229615 67649
rect 229557 67609 229569 67643
rect 229603 67640 229615 67643
rect 229646 67640 229652 67652
rect 229603 67612 229652 67640
rect 229603 67609 229615 67612
rect 229557 67603 229615 67609
rect 229646 67600 229652 67612
rect 229704 67600 229710 67652
rect 278038 67600 278044 67652
rect 278096 67640 278102 67652
rect 278130 67640 278136 67652
rect 278096 67612 278136 67640
rect 278096 67600 278102 67612
rect 278130 67600 278136 67612
rect 278188 67600 278194 67652
rect 240502 67572 240508 67584
rect 240463 67544 240508 67572
rect 240502 67532 240508 67544
rect 240560 67532 240566 67584
rect 260098 67532 260104 67584
rect 260156 67532 260162 67584
rect 260116 67436 260144 67532
rect 260190 67436 260196 67448
rect 260116 67408 260196 67436
rect 260190 67396 260196 67408
rect 260248 67396 260254 67448
rect 237558 66348 237564 66360
rect 237484 66320 237564 66348
rect 237484 66224 237512 66320
rect 237558 66308 237564 66320
rect 237616 66308 237622 66360
rect 251634 66240 251640 66292
rect 251692 66280 251698 66292
rect 251818 66280 251824 66292
rect 251692 66252 251824 66280
rect 251692 66240 251698 66252
rect 251818 66240 251824 66252
rect 251876 66240 251882 66292
rect 256510 66240 256516 66292
rect 256568 66280 256574 66292
rect 256602 66280 256608 66292
rect 256568 66252 256608 66280
rect 256568 66240 256574 66252
rect 256602 66240 256608 66252
rect 256660 66240 256666 66292
rect 259270 66240 259276 66292
rect 259328 66280 259334 66292
rect 259362 66280 259368 66292
rect 259328 66252 259368 66280
rect 259328 66240 259334 66252
rect 259362 66240 259368 66252
rect 259420 66240 259426 66292
rect 237466 66172 237472 66224
rect 237524 66172 237530 66224
rect 258534 64988 258540 65000
rect 258495 64960 258540 64988
rect 258534 64948 258540 64960
rect 258592 64948 258598 65000
rect 238938 64880 238944 64932
rect 238996 64920 239002 64932
rect 238996 64892 239041 64920
rect 238996 64880 239002 64892
rect 238202 64852 238208 64864
rect 238163 64824 238208 64852
rect 238202 64812 238208 64824
rect 238260 64812 238266 64864
rect 241146 64852 241152 64864
rect 241107 64824 241152 64852
rect 241146 64812 241152 64824
rect 241204 64812 241210 64864
rect 258534 64812 258540 64864
rect 258592 64852 258598 64864
rect 258626 64852 258632 64864
rect 258592 64824 258632 64852
rect 258592 64812 258598 64824
rect 258626 64812 258632 64824
rect 258684 64812 258690 64864
rect 272426 64852 272432 64864
rect 272352 64824 272432 64852
rect 272352 64796 272380 64824
rect 272426 64812 272432 64824
rect 272484 64812 272490 64864
rect 294598 64812 294604 64864
rect 294656 64852 294662 64864
rect 579798 64852 579804 64864
rect 294656 64824 579804 64852
rect 294656 64812 294662 64824
rect 579798 64812 579804 64824
rect 579856 64812 579862 64864
rect 272334 64744 272340 64796
rect 272392 64744 272398 64796
rect 258626 63492 258632 63504
rect 258587 63464 258632 63492
rect 258626 63452 258632 63464
rect 258684 63452 258690 63504
rect 240502 57984 240508 57996
rect 240463 57956 240508 57984
rect 240502 57944 240508 57956
rect 240560 57944 240566 57996
rect 260282 57944 260288 57996
rect 260340 57984 260346 57996
rect 260374 57984 260380 57996
rect 260340 57956 260380 57984
rect 260340 57944 260346 57956
rect 260374 57944 260380 57956
rect 260432 57944 260438 57996
rect 229557 57919 229615 57925
rect 229557 57885 229569 57919
rect 229603 57916 229615 57919
rect 229646 57916 229652 57928
rect 229603 57888 229652 57916
rect 229603 57885 229615 57888
rect 229557 57879 229615 57885
rect 229646 57876 229652 57888
rect 229704 57876 229710 57928
rect 256510 56584 256516 56636
rect 256568 56624 256574 56636
rect 256602 56624 256608 56636
rect 256568 56596 256608 56624
rect 256568 56584 256574 56596
rect 256602 56584 256608 56596
rect 256660 56584 256666 56636
rect 275278 56556 275284 56568
rect 275239 56528 275284 56556
rect 275278 56516 275284 56528
rect 275336 56516 275342 56568
rect 238202 55264 238208 55276
rect 238163 55236 238208 55264
rect 238202 55224 238208 55236
rect 238260 55224 238266 55276
rect 241146 55264 241152 55276
rect 241107 55236 241152 55264
rect 241146 55224 241152 55236
rect 241204 55224 241210 55276
rect 238938 55196 238944 55208
rect 238899 55168 238944 55196
rect 238938 55156 238944 55168
rect 238996 55156 239002 55208
rect 243446 51144 243452 51196
rect 243504 51144 243510 51196
rect 230842 51076 230848 51128
rect 230900 51116 230906 51128
rect 231026 51116 231032 51128
rect 230900 51088 231032 51116
rect 230900 51076 230906 51088
rect 231026 51076 231032 51088
rect 231084 51076 231090 51128
rect 238202 51116 238208 51128
rect 238163 51088 238208 51116
rect 238202 51076 238208 51088
rect 238260 51076 238266 51128
rect 241146 51076 241152 51128
rect 241204 51076 241210 51128
rect 3050 51008 3056 51060
rect 3108 51048 3114 51060
rect 225598 51048 225604 51060
rect 3108 51020 225604 51048
rect 3108 51008 3114 51020
rect 225598 51008 225604 51020
rect 225656 51008 225662 51060
rect 241164 50980 241192 51076
rect 243464 51060 243492 51144
rect 243446 51008 243452 51060
rect 243504 51008 243510 51060
rect 275278 51048 275284 51060
rect 275239 51020 275284 51048
rect 275278 51008 275284 51020
rect 275336 51008 275342 51060
rect 278038 51008 278044 51060
rect 278096 51048 278102 51060
rect 278222 51048 278228 51060
rect 278096 51020 278228 51048
rect 278096 51008 278102 51020
rect 278222 51008 278228 51020
rect 278280 51008 278286 51060
rect 241238 50980 241244 50992
rect 241164 50952 241244 50980
rect 241238 50940 241244 50952
rect 241296 50940 241302 50992
rect 260101 48399 260159 48405
rect 260101 48365 260113 48399
rect 260147 48396 260159 48399
rect 260190 48396 260196 48408
rect 260147 48368 260196 48396
rect 260147 48365 260159 48368
rect 260101 48359 260159 48365
rect 260190 48356 260196 48368
rect 260248 48356 260254 48408
rect 260285 48399 260343 48405
rect 260285 48365 260297 48399
rect 260331 48396 260343 48399
rect 260374 48396 260380 48408
rect 260331 48368 260380 48396
rect 260331 48365 260343 48368
rect 260285 48359 260343 48365
rect 260374 48356 260380 48368
rect 260432 48356 260438 48408
rect 229554 48328 229560 48340
rect 229515 48300 229560 48328
rect 229554 48288 229560 48300
rect 229612 48288 229618 48340
rect 251542 48288 251548 48340
rect 251600 48328 251606 48340
rect 251634 48328 251640 48340
rect 251600 48300 251640 48328
rect 251600 48288 251606 48300
rect 251634 48288 251640 48300
rect 251692 48288 251698 48340
rect 243449 48263 243507 48269
rect 243449 48229 243461 48263
rect 243495 48260 243507 48263
rect 243538 48260 243544 48272
rect 243495 48232 243544 48260
rect 243495 48229 243507 48232
rect 243449 48223 243507 48229
rect 243538 48220 243544 48232
rect 243596 48220 243602 48272
rect 237466 46928 237472 46980
rect 237524 46968 237530 46980
rect 237558 46968 237564 46980
rect 237524 46940 237564 46968
rect 237524 46928 237530 46940
rect 237558 46928 237564 46940
rect 237616 46928 237622 46980
rect 238202 46968 238208 46980
rect 238163 46940 238208 46968
rect 238202 46928 238208 46940
rect 238260 46928 238266 46980
rect 260098 46968 260104 46980
rect 260059 46940 260104 46968
rect 260098 46928 260104 46940
rect 260156 46928 260162 46980
rect 260282 46968 260288 46980
rect 260243 46940 260288 46968
rect 260282 46928 260288 46940
rect 260340 46928 260346 46980
rect 278041 46903 278099 46909
rect 278041 46869 278053 46903
rect 278087 46900 278099 46903
rect 278222 46900 278228 46912
rect 278087 46872 278228 46900
rect 278087 46869 278099 46872
rect 278041 46863 278099 46869
rect 278222 46860 278228 46872
rect 278280 46860 278286 46912
rect 238938 45568 238944 45620
rect 238996 45608 239002 45620
rect 258626 45608 258632 45620
rect 238996 45580 239041 45608
rect 258587 45580 258632 45608
rect 238996 45568 239002 45580
rect 258626 45568 258632 45580
rect 258684 45568 258690 45620
rect 237558 45540 237564 45552
rect 237519 45512 237564 45540
rect 237558 45500 237564 45512
rect 237616 45500 237622 45552
rect 238202 45500 238208 45552
rect 238260 45540 238266 45552
rect 238297 45543 238355 45549
rect 238297 45540 238309 45543
rect 238260 45512 238309 45540
rect 238260 45500 238266 45512
rect 238297 45509 238309 45512
rect 238343 45509 238355 45543
rect 241238 45540 241244 45552
rect 241199 45512 241244 45540
rect 238297 45503 238355 45509
rect 241238 45500 241244 45512
rect 241296 45500 241302 45552
rect 251542 44956 251548 45008
rect 251600 44996 251606 45008
rect 251726 44996 251732 45008
rect 251600 44968 251732 44996
rect 251600 44956 251606 44968
rect 251726 44956 251732 44968
rect 251784 44956 251790 45008
rect 253934 43460 253940 43512
rect 253992 43500 253998 43512
rect 254118 43500 254124 43512
rect 253992 43472 254124 43500
rect 253992 43460 253998 43472
rect 254118 43460 254124 43472
rect 254176 43460 254182 43512
rect 259270 43460 259276 43512
rect 259328 43500 259334 43512
rect 259454 43500 259460 43512
rect 259328 43472 259460 43500
rect 259328 43460 259334 43472
rect 259454 43460 259460 43472
rect 259512 43460 259518 43512
rect 229462 41352 229468 41404
rect 229520 41392 229526 41404
rect 229646 41392 229652 41404
rect 229520 41364 229652 41392
rect 229520 41352 229526 41364
rect 229646 41352 229652 41364
rect 229704 41352 229710 41404
rect 230842 41352 230848 41404
rect 230900 41392 230906 41404
rect 231026 41392 231032 41404
rect 230900 41364 231032 41392
rect 230900 41352 230906 41364
rect 231026 41352 231032 41364
rect 231084 41352 231090 41404
rect 304258 41352 304264 41404
rect 304316 41392 304322 41404
rect 580166 41392 580172 41404
rect 304316 41364 580172 41392
rect 304316 41352 304322 41364
rect 580166 41352 580172 41364
rect 580224 41352 580230 41404
rect 238938 38672 238944 38684
rect 238864 38644 238944 38672
rect 238864 38616 238892 38644
rect 238938 38632 238944 38644
rect 238996 38632 239002 38684
rect 249150 38632 249156 38684
rect 249208 38672 249214 38684
rect 249242 38672 249248 38684
rect 249208 38644 249248 38672
rect 249208 38632 249214 38644
rect 249242 38632 249248 38644
rect 249300 38632 249306 38684
rect 229557 38607 229615 38613
rect 229557 38573 229569 38607
rect 229603 38604 229615 38607
rect 229646 38604 229652 38616
rect 229603 38576 229652 38604
rect 229603 38573 229615 38576
rect 229557 38567 229615 38573
rect 229646 38564 229652 38576
rect 229704 38564 229710 38616
rect 238846 38564 238852 38616
rect 238904 38564 238910 38616
rect 278038 37312 278044 37324
rect 277999 37284 278044 37312
rect 278038 37272 278044 37284
rect 278096 37272 278102 37324
rect 256602 37204 256608 37256
rect 256660 37244 256666 37256
rect 256694 37244 256700 37256
rect 256660 37216 256700 37244
rect 256660 37204 256666 37216
rect 256694 37204 256700 37216
rect 256752 37204 256758 37256
rect 238202 35980 238208 36032
rect 238260 36020 238266 36032
rect 238297 36023 238355 36029
rect 238297 36020 238309 36023
rect 238260 35992 238309 36020
rect 238260 35980 238266 35992
rect 238297 35989 238309 35992
rect 238343 35989 238355 36023
rect 238297 35983 238355 35989
rect 237561 35955 237619 35961
rect 237561 35921 237573 35955
rect 237607 35952 237619 35955
rect 237650 35952 237656 35964
rect 237607 35924 237656 35952
rect 237607 35921 237619 35924
rect 237561 35915 237619 35921
rect 237650 35912 237656 35924
rect 237708 35912 237714 35964
rect 241238 35952 241244 35964
rect 241199 35924 241244 35952
rect 241238 35912 241244 35924
rect 241296 35912 241302 35964
rect 3510 35844 3516 35896
rect 3568 35884 3574 35896
rect 214558 35884 214564 35896
rect 3568 35856 214564 35884
rect 3568 35844 3574 35856
rect 214558 35844 214564 35856
rect 214616 35844 214622 35896
rect 238113 35887 238171 35893
rect 238113 35853 238125 35887
rect 238159 35884 238171 35887
rect 238202 35884 238208 35896
rect 238159 35856 238208 35884
rect 238159 35853 238171 35856
rect 238113 35847 238171 35853
rect 238202 35844 238208 35856
rect 238260 35844 238266 35896
rect 256605 35887 256663 35893
rect 256605 35853 256617 35887
rect 256651 35884 256663 35887
rect 256694 35884 256700 35896
rect 256651 35856 256700 35884
rect 256651 35853 256663 35856
rect 256605 35847 256663 35853
rect 256694 35844 256700 35856
rect 256752 35844 256758 35896
rect 259273 35887 259331 35893
rect 259273 35853 259285 35887
rect 259319 35884 259331 35887
rect 259454 35884 259460 35896
rect 259319 35856 259460 35884
rect 259319 35853 259331 35856
rect 259273 35847 259331 35853
rect 259454 35844 259460 35856
rect 259512 35844 259518 35896
rect 230842 31764 230848 31816
rect 230900 31804 230906 31816
rect 231026 31804 231032 31816
rect 230900 31776 231032 31804
rect 230900 31764 230906 31776
rect 231026 31764 231032 31776
rect 231084 31764 231090 31816
rect 321462 29180 321468 29232
rect 321520 29220 321526 29232
rect 321646 29220 321652 29232
rect 321520 29192 321652 29220
rect 321520 29180 321526 29192
rect 321646 29180 321652 29192
rect 321704 29180 321710 29232
rect 302142 29112 302148 29164
rect 302200 29152 302206 29164
rect 308950 29152 308956 29164
rect 302200 29124 308956 29152
rect 302200 29112 302206 29124
rect 308950 29112 308956 29124
rect 309008 29112 309014 29164
rect 437382 29112 437388 29164
rect 437440 29152 437446 29164
rect 444190 29152 444196 29164
rect 437440 29124 444196 29152
rect 437440 29112 437446 29124
rect 444190 29112 444196 29124
rect 444248 29112 444254 29164
rect 514662 29112 514668 29164
rect 514720 29152 514726 29164
rect 521470 29152 521476 29164
rect 514720 29124 521476 29152
rect 514720 29112 514726 29124
rect 521470 29112 521476 29124
rect 521528 29112 521534 29164
rect 533982 29112 533988 29164
rect 534040 29152 534046 29164
rect 540790 29152 540796 29164
rect 534040 29124 540796 29152
rect 534040 29112 534046 29124
rect 540790 29112 540796 29124
rect 540848 29112 540854 29164
rect 553302 29112 553308 29164
rect 553360 29152 553366 29164
rect 560110 29152 560116 29164
rect 553360 29124 560116 29152
rect 553360 29112 553366 29124
rect 560110 29112 560116 29124
rect 560168 29112 560174 29164
rect 572622 29112 572628 29164
rect 572680 29152 572686 29164
rect 579430 29152 579436 29164
rect 572680 29124 579436 29152
rect 572680 29112 572686 29124
rect 579430 29112 579436 29124
rect 579488 29112 579494 29164
rect 254118 29084 254124 29096
rect 253952 29056 254124 29084
rect 229554 29016 229560 29028
rect 229515 28988 229560 29016
rect 229554 28976 229560 28988
rect 229612 28976 229618 29028
rect 238846 28976 238852 29028
rect 238904 29016 238910 29028
rect 238938 29016 238944 29028
rect 238904 28988 238944 29016
rect 238904 28976 238910 28988
rect 238938 28976 238944 28988
rect 238996 28976 239002 29028
rect 253952 28960 253980 29056
rect 254118 29044 254124 29056
rect 254176 29044 254182 29096
rect 253934 28908 253940 28960
rect 253992 28908 253998 28960
rect 243449 27659 243507 27665
rect 243449 27625 243461 27659
rect 243495 27656 243507 27659
rect 243538 27656 243544 27668
rect 243495 27628 243544 27656
rect 243495 27625 243507 27628
rect 243449 27619 243507 27625
rect 243538 27616 243544 27628
rect 243596 27616 243602 27668
rect 274910 27548 274916 27600
rect 274968 27588 274974 27600
rect 275370 27588 275376 27600
rect 274968 27560 275376 27588
rect 274968 27548 274974 27560
rect 275370 27548 275376 27560
rect 275428 27548 275434 27600
rect 243449 27523 243507 27529
rect 243449 27489 243461 27523
rect 243495 27520 243507 27523
rect 243538 27520 243544 27532
rect 243495 27492 243544 27520
rect 243495 27489 243507 27492
rect 243449 27483 243507 27489
rect 243538 27480 243544 27492
rect 243596 27480 243602 27532
rect 278038 27480 278044 27532
rect 278096 27520 278102 27532
rect 278225 27523 278283 27529
rect 278225 27520 278237 27523
rect 278096 27492 278237 27520
rect 278096 27480 278102 27492
rect 278225 27489 278237 27492
rect 278271 27489 278283 27523
rect 278225 27483 278283 27489
rect 238110 26296 238116 26308
rect 238071 26268 238116 26296
rect 238110 26256 238116 26268
rect 238168 26256 238174 26308
rect 256602 26296 256608 26308
rect 256563 26268 256608 26296
rect 256602 26256 256608 26268
rect 256660 26256 256666 26308
rect 259270 26296 259276 26308
rect 259231 26268 259276 26296
rect 259270 26256 259276 26268
rect 259328 26256 259334 26308
rect 274910 26228 274916 26240
rect 274871 26200 274916 26228
rect 274910 26188 274916 26200
rect 274968 26188 274974 26240
rect 287606 22720 287612 22772
rect 287664 22760 287670 22772
rect 567194 22760 567200 22772
rect 287664 22732 567200 22760
rect 287664 22720 287670 22732
rect 567194 22720 567200 22732
rect 567252 22720 567258 22772
rect 229554 22108 229560 22160
rect 229612 22108 229618 22160
rect 229572 22024 229600 22108
rect 230842 22040 230848 22092
rect 230900 22080 230906 22092
rect 231026 22080 231032 22092
rect 230900 22052 231032 22080
rect 230900 22040 230906 22052
rect 231026 22040 231032 22052
rect 231084 22040 231090 22092
rect 243446 22080 243452 22092
rect 243407 22052 243452 22080
rect 243446 22040 243452 22052
rect 243504 22040 243510 22092
rect 229554 21972 229560 22024
rect 229612 21972 229618 22024
rect 238849 21471 238907 21477
rect 238849 21437 238861 21471
rect 238895 21468 238907 21471
rect 238938 21468 238944 21480
rect 238895 21440 238944 21468
rect 238895 21437 238907 21440
rect 238849 21431 238907 21437
rect 238938 21428 238944 21440
rect 238996 21428 239002 21480
rect 320818 21360 320824 21412
rect 320876 21400 320882 21412
rect 543734 21400 543740 21412
rect 320876 21372 543740 21400
rect 320876 21360 320882 21372
rect 543734 21360 543740 21372
rect 543792 21360 543798 21412
rect 294690 19932 294696 19984
rect 294748 19972 294754 19984
rect 532694 19972 532700 19984
rect 294748 19944 532700 19972
rect 294748 19932 294754 19944
rect 532694 19932 532700 19944
rect 532752 19932 532758 19984
rect 259917 19499 259975 19505
rect 259917 19465 259929 19499
rect 259963 19496 259975 19499
rect 260098 19496 260104 19508
rect 259963 19468 260104 19496
rect 259963 19465 259975 19468
rect 259917 19459 259975 19465
rect 260098 19456 260104 19468
rect 260156 19456 260162 19508
rect 260006 19388 260012 19440
rect 260064 19388 260070 19440
rect 237558 19320 237564 19372
rect 237616 19360 237622 19372
rect 237650 19360 237656 19372
rect 237616 19332 237656 19360
rect 237616 19320 237622 19332
rect 237650 19320 237656 19332
rect 237708 19320 237714 19372
rect 260024 19304 260052 19388
rect 260098 19320 260104 19372
rect 260156 19360 260162 19372
rect 260282 19360 260288 19372
rect 260156 19332 260288 19360
rect 260156 19320 260162 19332
rect 260282 19320 260288 19332
rect 260340 19320 260346 19372
rect 260006 19252 260012 19304
rect 260064 19252 260070 19304
rect 276474 19292 276480 19304
rect 276435 19264 276480 19292
rect 276474 19252 276480 19264
rect 276532 19252 276538 19304
rect 297358 18572 297364 18624
rect 297416 18612 297422 18624
rect 525794 18612 525800 18624
rect 297416 18584 525800 18612
rect 297416 18572 297422 18584
rect 525794 18572 525800 18584
rect 525852 18572 525858 18624
rect 253934 18068 253940 18080
rect 253895 18040 253940 18068
rect 253934 18028 253940 18040
rect 253992 18028 253998 18080
rect 240870 17960 240876 18012
rect 240928 18000 240934 18012
rect 241054 18000 241060 18012
rect 240928 17972 241060 18000
rect 240928 17960 240934 17972
rect 241054 17960 241060 17972
rect 241112 17960 241118 18012
rect 251634 17960 251640 18012
rect 251692 18000 251698 18012
rect 251726 18000 251732 18012
rect 251692 17972 251732 18000
rect 251692 17960 251698 17972
rect 251726 17960 251732 17972
rect 251784 17960 251790 18012
rect 258534 17960 258540 18012
rect 258592 18000 258598 18012
rect 258626 18000 258632 18012
rect 258592 17972 258632 18000
rect 258592 17960 258598 17972
rect 258626 17960 258632 17972
rect 258684 17960 258690 18012
rect 259914 18000 259920 18012
rect 259875 17972 259920 18000
rect 259914 17960 259920 17972
rect 259972 17960 259978 18012
rect 229094 17892 229100 17944
rect 229152 17932 229158 17944
rect 579798 17932 579804 17944
rect 229152 17904 579804 17932
rect 229152 17892 229158 17904
rect 579798 17892 579804 17904
rect 579856 17892 579862 17944
rect 259914 17824 259920 17876
rect 259972 17864 259978 17876
rect 260098 17864 260104 17876
rect 259972 17836 260104 17864
rect 259972 17824 259978 17836
rect 260098 17824 260104 17836
rect 260156 17824 260162 17876
rect 260193 17867 260251 17873
rect 260193 17833 260205 17867
rect 260239 17864 260251 17867
rect 260374 17864 260380 17876
rect 260239 17836 260380 17864
rect 260239 17833 260251 17836
rect 260193 17827 260251 17833
rect 260374 17824 260380 17836
rect 260432 17824 260438 17876
rect 256510 16668 256516 16720
rect 256568 16708 256574 16720
rect 256568 16680 256648 16708
rect 256568 16668 256574 16680
rect 256620 16652 256648 16680
rect 238846 16640 238852 16652
rect 238807 16612 238852 16640
rect 238846 16600 238852 16612
rect 238904 16600 238910 16652
rect 253934 16640 253940 16652
rect 253895 16612 253940 16640
rect 253934 16600 253940 16612
rect 253992 16600 253998 16652
rect 256602 16600 256608 16652
rect 256660 16600 256666 16652
rect 274910 16640 274916 16652
rect 274871 16612 274916 16640
rect 274910 16600 274916 16612
rect 274968 16600 274974 16652
rect 237558 16572 237564 16584
rect 237519 16544 237564 16572
rect 237558 16532 237564 16544
rect 237616 16532 237622 16584
rect 151630 15852 151636 15904
rect 151688 15892 151694 15904
rect 245194 15892 245200 15904
rect 151688 15864 245200 15892
rect 151688 15852 151694 15864
rect 245194 15852 245200 15864
rect 245252 15852 245258 15904
rect 290458 15852 290464 15904
rect 290516 15892 290522 15904
rect 514754 15892 514760 15904
rect 290516 15864 514760 15892
rect 290516 15852 290522 15864
rect 514754 15852 514760 15864
rect 514812 15852 514818 15904
rect 164142 14424 164148 14476
rect 164200 14464 164206 14476
rect 228358 14464 228364 14476
rect 164200 14436 228364 14464
rect 164200 14424 164206 14436
rect 228358 14424 228364 14436
rect 228416 14424 228422 14476
rect 298738 14424 298744 14476
rect 298796 14464 298802 14476
rect 512086 14464 512092 14476
rect 298796 14436 512092 14464
rect 298796 14424 298802 14436
rect 512086 14424 512092 14436
rect 512144 14424 512150 14476
rect 148962 13064 148968 13116
rect 149020 13104 149026 13116
rect 225690 13104 225696 13116
rect 149020 13076 225696 13104
rect 149020 13064 149026 13076
rect 225690 13064 225696 13076
rect 225748 13064 225754 13116
rect 291838 13064 291844 13116
rect 291896 13104 291902 13116
rect 507854 13104 507860 13116
rect 291896 13076 507860 13104
rect 291896 13064 291902 13076
rect 507854 13064 507860 13076
rect 507912 13064 507918 13116
rect 230842 12452 230848 12504
rect 230900 12492 230906 12504
rect 231026 12492 231032 12504
rect 230900 12464 231032 12492
rect 230900 12452 230906 12464
rect 231026 12452 231032 12464
rect 231084 12452 231090 12504
rect 243446 12492 243452 12504
rect 243372 12464 243452 12492
rect 243372 12436 243400 12464
rect 243446 12452 243452 12464
rect 243504 12452 243510 12504
rect 243354 12384 243360 12436
rect 243412 12384 243418 12436
rect 166902 11704 166908 11756
rect 166960 11744 166966 11756
rect 226978 11744 226984 11756
rect 166960 11716 226984 11744
rect 166960 11704 166966 11716
rect 226978 11704 226984 11716
rect 227036 11704 227042 11756
rect 228910 11704 228916 11756
rect 228968 11744 228974 11756
rect 252002 11744 252008 11756
rect 228968 11716 252008 11744
rect 228968 11704 228974 11716
rect 252002 11704 252008 11716
rect 252060 11704 252066 11756
rect 301498 11704 301504 11756
rect 301556 11744 301562 11756
rect 503714 11744 503720 11756
rect 301556 11716 503720 11744
rect 301556 11704 301562 11716
rect 503714 11704 503720 11716
rect 503772 11704 503778 11756
rect 266538 10956 266544 11008
rect 266596 10996 266602 11008
rect 356146 10996 356152 11008
rect 266596 10968 356152 10996
rect 266596 10956 266602 10968
rect 356146 10956 356152 10968
rect 356204 10956 356210 11008
rect 267366 10888 267372 10940
rect 267424 10928 267430 10940
rect 358814 10928 358820 10940
rect 267424 10900 358820 10928
rect 267424 10888 267430 10900
rect 358814 10888 358820 10900
rect 358872 10888 358878 10940
rect 267274 10820 267280 10872
rect 267332 10860 267338 10872
rect 362954 10860 362960 10872
rect 267332 10832 362960 10860
rect 267332 10820 267338 10832
rect 362954 10820 362960 10832
rect 363012 10820 363018 10872
rect 266354 10752 266360 10804
rect 266412 10792 266418 10804
rect 365714 10792 365720 10804
rect 266412 10764 365720 10792
rect 266412 10752 266418 10764
rect 365714 10752 365720 10764
rect 365772 10752 365778 10804
rect 64782 10684 64788 10736
rect 64840 10724 64846 10736
rect 236730 10724 236736 10736
rect 64840 10696 236736 10724
rect 64840 10684 64846 10696
rect 236730 10684 236736 10696
rect 236788 10684 236794 10736
rect 268470 10684 268476 10736
rect 268528 10724 268534 10736
rect 369854 10724 369860 10736
rect 268528 10696 369860 10724
rect 268528 10684 268534 10696
rect 369854 10684 369860 10696
rect 369912 10684 369918 10736
rect 60642 10616 60648 10668
rect 60700 10656 60706 10668
rect 236822 10656 236828 10668
rect 60700 10628 236828 10656
rect 60700 10616 60706 10628
rect 236822 10616 236828 10628
rect 236880 10616 236886 10668
rect 268562 10616 268568 10668
rect 268620 10656 268626 10668
rect 374086 10656 374092 10668
rect 268620 10628 374092 10656
rect 268620 10616 268626 10628
rect 374086 10616 374092 10628
rect 374144 10616 374150 10668
rect 30282 10548 30288 10600
rect 30340 10588 30346 10600
rect 232222 10588 232228 10600
rect 30340 10560 232228 10588
rect 30340 10548 30346 10560
rect 232222 10548 232228 10560
rect 232280 10548 232286 10600
rect 268746 10548 268752 10600
rect 268804 10588 268810 10600
rect 376754 10588 376760 10600
rect 268804 10560 376760 10588
rect 268804 10548 268810 10560
rect 376754 10548 376760 10560
rect 376812 10548 376818 10600
rect 27522 10480 27528 10532
rect 27580 10520 27586 10532
rect 232130 10520 232136 10532
rect 27580 10492 232136 10520
rect 27580 10480 27586 10492
rect 232130 10480 232136 10492
rect 232188 10480 232194 10532
rect 269114 10480 269120 10532
rect 269172 10520 269178 10532
rect 380894 10520 380900 10532
rect 269172 10492 380900 10520
rect 269172 10480 269178 10492
rect 380894 10480 380900 10492
rect 380952 10480 380958 10532
rect 22002 10412 22008 10464
rect 22060 10452 22066 10464
rect 232038 10452 232044 10464
rect 22060 10424 232044 10452
rect 22060 10412 22066 10424
rect 232038 10412 232044 10424
rect 232096 10412 232102 10464
rect 235994 10412 236000 10464
rect 236052 10452 236058 10464
rect 253198 10452 253204 10464
rect 236052 10424 253204 10452
rect 236052 10412 236058 10424
rect 253198 10412 253204 10424
rect 253256 10412 253262 10464
rect 269942 10412 269948 10464
rect 270000 10452 270006 10464
rect 383654 10452 383660 10464
rect 270000 10424 383660 10452
rect 270000 10412 270006 10424
rect 383654 10412 383660 10424
rect 383712 10412 383718 10464
rect 9582 10344 9588 10396
rect 9640 10384 9646 10396
rect 230934 10384 230940 10396
rect 9640 10356 230940 10384
rect 9640 10344 9646 10356
rect 230934 10344 230940 10356
rect 230992 10344 230998 10396
rect 233142 10344 233148 10396
rect 233200 10384 233206 10396
rect 252922 10384 252928 10396
rect 233200 10356 252928 10384
rect 233200 10344 233206 10356
rect 252922 10344 252928 10356
rect 252980 10344 252986 10396
rect 269298 10344 269304 10396
rect 269356 10384 269362 10396
rect 387794 10384 387800 10396
rect 269356 10356 387800 10384
rect 269356 10344 269362 10356
rect 387794 10344 387800 10356
rect 387852 10344 387858 10396
rect 3970 10276 3976 10328
rect 4028 10316 4034 10328
rect 229554 10316 229560 10328
rect 4028 10288 229560 10316
rect 4028 10276 4034 10288
rect 229554 10276 229560 10288
rect 229612 10276 229618 10328
rect 231762 10276 231768 10328
rect 231820 10316 231826 10328
rect 251910 10316 251916 10328
rect 231820 10288 251916 10316
rect 231820 10276 231826 10288
rect 251910 10276 251916 10288
rect 251968 10276 251974 10328
rect 270034 10276 270040 10328
rect 270092 10316 270098 10328
rect 390554 10316 390560 10328
rect 270092 10288 390560 10316
rect 270092 10276 270098 10288
rect 390554 10276 390560 10288
rect 390612 10276 390618 10328
rect 265618 10208 265624 10260
rect 265676 10248 265682 10260
rect 351914 10248 351920 10260
rect 265676 10220 351920 10248
rect 265676 10208 265682 10220
rect 351914 10208 351920 10220
rect 351972 10208 351978 10260
rect 265710 10140 265716 10192
rect 265768 10180 265774 10192
rect 347774 10180 347780 10192
rect 265768 10152 347780 10180
rect 265768 10140 265774 10152
rect 347774 10140 347780 10152
rect 347832 10140 347838 10192
rect 265894 10072 265900 10124
rect 265952 10112 265958 10124
rect 345014 10112 345020 10124
rect 265952 10084 345020 10112
rect 265952 10072 265958 10084
rect 345014 10072 345020 10084
rect 345072 10072 345078 10124
rect 265066 10004 265072 10056
rect 265124 10044 265130 10056
rect 340874 10044 340880 10056
rect 265124 10016 340880 10044
rect 265124 10004 265130 10016
rect 340874 10004 340880 10016
rect 340932 10004 340938 10056
rect 276474 9704 276480 9716
rect 276435 9676 276480 9704
rect 276474 9664 276480 9676
rect 276532 9664 276538 9716
rect 278222 9704 278228 9716
rect 278183 9676 278228 9704
rect 278222 9664 278228 9676
rect 278280 9664 278286 9716
rect 90910 9596 90916 9648
rect 90968 9636 90974 9648
rect 239306 9636 239312 9648
rect 90968 9608 239312 9636
rect 90968 9596 90974 9608
rect 239306 9596 239312 9608
rect 239364 9596 239370 9648
rect 87322 9528 87328 9580
rect 87380 9568 87386 9580
rect 239030 9568 239036 9580
rect 87380 9540 239036 9568
rect 87380 9528 87386 9540
rect 239030 9528 239036 9540
rect 239088 9528 239094 9580
rect 274910 9528 274916 9580
rect 274968 9568 274974 9580
rect 275370 9568 275376 9580
rect 274968 9540 275376 9568
rect 274968 9528 274974 9540
rect 275370 9528 275376 9540
rect 275428 9528 275434 9580
rect 83826 9460 83832 9512
rect 83884 9500 83890 9512
rect 238570 9500 238576 9512
rect 83884 9472 238576 9500
rect 83884 9460 83890 9472
rect 238570 9460 238576 9472
rect 238628 9460 238634 9512
rect 80238 9392 80244 9444
rect 80296 9432 80302 9444
rect 237742 9432 237748 9444
rect 80296 9404 237748 9432
rect 80296 9392 80302 9404
rect 237742 9392 237748 9404
rect 237800 9392 237806 9444
rect 76650 9324 76656 9376
rect 76708 9364 76714 9376
rect 237834 9364 237840 9376
rect 76708 9336 237840 9364
rect 76708 9324 76714 9336
rect 237834 9324 237840 9336
rect 237892 9324 237898 9376
rect 73062 9256 73068 9308
rect 73120 9296 73126 9308
rect 237561 9299 237619 9305
rect 237561 9296 237573 9299
rect 73120 9268 237573 9296
rect 73120 9256 73126 9268
rect 237561 9265 237573 9268
rect 237607 9265 237619 9299
rect 237561 9259 237619 9265
rect 260466 9256 260472 9308
rect 260524 9296 260530 9308
rect 291930 9296 291936 9308
rect 260524 9268 291936 9296
rect 260524 9256 260530 9268
rect 291930 9256 291936 9268
rect 291988 9256 291994 9308
rect 69474 9188 69480 9240
rect 69532 9228 69538 9240
rect 237098 9228 237104 9240
rect 69532 9200 237104 9228
rect 69532 9188 69538 9200
rect 237098 9188 237104 9200
rect 237156 9188 237162 9240
rect 260006 9188 260012 9240
rect 260064 9228 260070 9240
rect 295518 9228 295524 9240
rect 260064 9200 295524 9228
rect 260064 9188 260070 9200
rect 295518 9188 295524 9200
rect 295576 9188 295582 9240
rect 65978 9120 65984 9172
rect 66036 9160 66042 9172
rect 236362 9160 236368 9172
rect 66036 9132 236368 9160
rect 66036 9120 66042 9132
rect 236362 9120 236368 9132
rect 236420 9120 236426 9172
rect 259822 9120 259828 9172
rect 259880 9160 259886 9172
rect 299106 9160 299112 9172
rect 259880 9132 299112 9160
rect 259880 9120 259886 9132
rect 299106 9120 299112 9132
rect 299164 9120 299170 9172
rect 62390 9052 62396 9104
rect 62448 9092 62454 9104
rect 236638 9092 236644 9104
rect 62448 9064 236644 9092
rect 62448 9052 62454 9064
rect 236638 9052 236644 9064
rect 236696 9052 236702 9104
rect 261386 9052 261392 9104
rect 261444 9092 261450 9104
rect 306190 9092 306196 9104
rect 261444 9064 306196 9092
rect 261444 9052 261450 9064
rect 306190 9052 306196 9064
rect 306248 9052 306254 9104
rect 58802 8984 58808 9036
rect 58860 9024 58866 9036
rect 236454 9024 236460 9036
rect 58860 8996 236460 9024
rect 58860 8984 58866 8996
rect 236454 8984 236460 8996
rect 236512 8984 236518 9036
rect 261294 8984 261300 9036
rect 261352 9024 261358 9036
rect 309778 9024 309784 9036
rect 261352 8996 309784 9024
rect 261352 8984 261358 8996
rect 309778 8984 309784 8996
rect 309836 8984 309842 9036
rect 17310 8916 17316 8968
rect 17368 8956 17374 8968
rect 231670 8956 231676 8968
rect 17368 8928 231676 8956
rect 17368 8916 17374 8928
rect 231670 8916 231676 8928
rect 231728 8916 231734 8968
rect 241974 8916 241980 8968
rect 242032 8956 242038 8968
rect 251634 8956 251640 8968
rect 242032 8928 251640 8956
rect 242032 8916 242038 8928
rect 251634 8916 251640 8928
rect 251692 8916 251698 8968
rect 261202 8916 261208 8968
rect 261260 8956 261266 8968
rect 302602 8956 302608 8968
rect 261260 8928 302608 8956
rect 261260 8916 261266 8928
rect 302602 8916 302608 8928
rect 302660 8916 302666 8968
rect 302878 8916 302884 8968
rect 302936 8956 302942 8968
rect 494146 8956 494152 8968
rect 302936 8928 494152 8956
rect 302936 8916 302942 8928
rect 494146 8916 494152 8928
rect 494204 8916 494210 8968
rect 94498 8848 94504 8900
rect 94556 8888 94562 8900
rect 239214 8888 239220 8900
rect 94556 8860 239220 8888
rect 94556 8848 94562 8860
rect 239214 8848 239220 8860
rect 239272 8848 239278 8900
rect 98086 8780 98092 8832
rect 98144 8820 98150 8832
rect 240042 8820 240048 8832
rect 98144 8792 240048 8820
rect 98144 8780 98150 8792
rect 240042 8780 240048 8792
rect 240100 8780 240106 8832
rect 101582 8712 101588 8764
rect 101640 8752 101646 8764
rect 240502 8752 240508 8764
rect 101640 8724 240508 8752
rect 101640 8712 101646 8724
rect 240502 8712 240508 8724
rect 240560 8712 240566 8764
rect 105170 8644 105176 8696
rect 105228 8684 105234 8696
rect 240410 8684 240416 8696
rect 105228 8656 240416 8684
rect 105228 8644 105234 8656
rect 240410 8644 240416 8656
rect 240468 8644 240474 8696
rect 108758 8576 108764 8628
rect 108816 8616 108822 8628
rect 240318 8616 240324 8628
rect 108816 8588 240324 8616
rect 108816 8576 108822 8588
rect 240318 8576 240324 8588
rect 240376 8576 240382 8628
rect 112346 8508 112352 8560
rect 112404 8548 112410 8560
rect 241882 8548 241888 8560
rect 112404 8520 241888 8548
rect 112404 8508 112410 8520
rect 241882 8508 241888 8520
rect 241940 8508 241946 8560
rect 115934 8440 115940 8492
rect 115992 8480 115998 8492
rect 241790 8480 241796 8492
rect 115992 8452 241796 8480
rect 115992 8440 115998 8452
rect 241790 8440 241796 8452
rect 241848 8440 241854 8492
rect 119430 8372 119436 8424
rect 119488 8412 119494 8424
rect 242250 8412 242256 8424
rect 119488 8384 242256 8412
rect 119488 8372 119494 8384
rect 242250 8372 242256 8384
rect 242308 8372 242314 8424
rect 123018 8304 123024 8356
rect 123076 8344 123082 8356
rect 242618 8344 242624 8356
rect 123076 8316 242624 8344
rect 123076 8304 123082 8316
rect 242618 8304 242624 8316
rect 242676 8304 242682 8356
rect 260190 8344 260196 8356
rect 260151 8316 260196 8344
rect 260190 8304 260196 8316
rect 260248 8304 260254 8356
rect 3418 8236 3424 8288
rect 3476 8276 3482 8288
rect 13078 8276 13084 8288
rect 3476 8248 13084 8276
rect 3476 8236 3482 8248
rect 13078 8236 13084 8248
rect 13136 8236 13142 8288
rect 200390 8236 200396 8288
rect 200448 8276 200454 8288
rect 250530 8276 250536 8288
rect 200448 8248 250536 8276
rect 200448 8236 200454 8248
rect 250530 8236 250536 8248
rect 250588 8236 250594 8288
rect 256510 8236 256516 8288
rect 256568 8276 256574 8288
rect 257430 8276 257436 8288
rect 256568 8248 257436 8276
rect 256568 8236 256574 8248
rect 257430 8236 257436 8248
rect 257488 8236 257494 8288
rect 261478 8236 261484 8288
rect 261536 8276 261542 8288
rect 266998 8276 267004 8288
rect 261536 8248 267004 8276
rect 261536 8236 261542 8248
rect 266998 8236 267004 8248
rect 267056 8236 267062 8288
rect 275370 8276 275376 8288
rect 275331 8248 275376 8276
rect 275370 8236 275376 8248
rect 275428 8236 275434 8288
rect 196802 8168 196808 8220
rect 196860 8208 196866 8220
rect 250714 8208 250720 8220
rect 196860 8180 250720 8208
rect 196860 8168 196866 8180
rect 250714 8168 250720 8180
rect 250772 8168 250778 8220
rect 193214 8100 193220 8152
rect 193272 8140 193278 8152
rect 250070 8140 250076 8152
rect 193272 8112 250076 8140
rect 193272 8100 193278 8112
rect 250070 8100 250076 8112
rect 250128 8100 250134 8152
rect 189626 8032 189632 8084
rect 189684 8072 189690 8084
rect 249058 8072 249064 8084
rect 189684 8044 249064 8072
rect 189684 8032 189690 8044
rect 249058 8032 249064 8044
rect 249116 8032 249122 8084
rect 279786 8032 279792 8084
rect 279844 8072 279850 8084
rect 279970 8072 279976 8084
rect 279844 8044 279976 8072
rect 279844 8032 279850 8044
rect 279970 8032 279976 8044
rect 280028 8032 280034 8084
rect 186038 7964 186044 8016
rect 186096 8004 186102 8016
rect 248966 8004 248972 8016
rect 186096 7976 248972 8004
rect 186096 7964 186102 7976
rect 248966 7964 248972 7976
rect 249024 7964 249030 8016
rect 182542 7896 182548 7948
rect 182600 7936 182606 7948
rect 249150 7936 249156 7948
rect 182600 7908 249156 7936
rect 182600 7896 182606 7908
rect 249150 7896 249156 7908
rect 249208 7896 249214 7948
rect 178954 7828 178960 7880
rect 179012 7868 179018 7880
rect 248322 7868 248328 7880
rect 179012 7840 248328 7868
rect 179012 7828 179018 7840
rect 248322 7828 248328 7840
rect 248380 7828 248386 7880
rect 175366 7760 175372 7812
rect 175424 7800 175430 7812
rect 247954 7800 247960 7812
rect 175424 7772 247960 7800
rect 175424 7760 175430 7772
rect 247954 7760 247960 7772
rect 248012 7760 248018 7812
rect 171778 7692 171784 7744
rect 171836 7732 171842 7744
rect 247402 7732 247408 7744
rect 171836 7704 247408 7732
rect 171836 7692 171842 7704
rect 247402 7692 247408 7704
rect 247460 7692 247466 7744
rect 168190 7624 168196 7676
rect 168248 7664 168254 7676
rect 247310 7664 247316 7676
rect 168248 7636 247316 7664
rect 168248 7624 168254 7636
rect 247310 7624 247316 7636
rect 247368 7624 247374 7676
rect 132586 7556 132592 7608
rect 132644 7596 132650 7608
rect 243354 7596 243360 7608
rect 132644 7568 243360 7596
rect 132644 7556 132650 7568
rect 243354 7556 243360 7568
rect 243412 7556 243418 7608
rect 270494 7556 270500 7608
rect 270552 7596 270558 7608
rect 271690 7596 271696 7608
rect 270552 7568 271696 7596
rect 270552 7556 270558 7568
rect 271690 7556 271696 7568
rect 271748 7556 271754 7608
rect 280798 7556 280804 7608
rect 280856 7596 280862 7608
rect 314562 7596 314568 7608
rect 280856 7568 314568 7596
rect 280856 7556 280862 7568
rect 314562 7556 314568 7568
rect 314620 7556 314626 7608
rect 319438 7556 319444 7608
rect 319496 7596 319502 7608
rect 490558 7596 490564 7608
rect 319496 7568 490564 7596
rect 319496 7556 319502 7568
rect 490558 7556 490564 7568
rect 490616 7556 490622 7608
rect 203886 7488 203892 7540
rect 203944 7528 203950 7540
rect 250898 7528 250904 7540
rect 203944 7500 250904 7528
rect 203944 7488 203950 7500
rect 250898 7488 250904 7500
rect 250956 7488 250962 7540
rect 262950 6876 262956 6928
rect 263008 6916 263014 6928
rect 268102 6916 268108 6928
rect 263008 6888 268108 6916
rect 263008 6876 263014 6888
rect 268102 6876 268108 6888
rect 268160 6876 268166 6928
rect 283558 6876 283564 6928
rect 283616 6916 283622 6928
rect 288342 6916 288348 6928
rect 283616 6888 288348 6916
rect 283616 6876 283622 6888
rect 288342 6876 288348 6888
rect 288400 6876 288406 6928
rect 199194 6808 199200 6860
rect 199252 6848 199258 6860
rect 249794 6848 249800 6860
rect 199252 6820 249800 6848
rect 199252 6808 199258 6820
rect 249794 6808 249800 6820
rect 249852 6808 249858 6860
rect 266446 6808 266452 6860
rect 266504 6848 266510 6860
rect 354950 6848 354956 6860
rect 266504 6820 354956 6848
rect 266504 6808 266510 6820
rect 354950 6808 354956 6820
rect 355008 6808 355014 6860
rect 195606 6740 195612 6792
rect 195664 6780 195670 6792
rect 250346 6780 250352 6792
rect 195664 6752 250352 6780
rect 195664 6740 195670 6752
rect 250346 6740 250352 6752
rect 250404 6740 250410 6792
rect 266814 6740 266820 6792
rect 266872 6780 266878 6792
rect 358538 6780 358544 6792
rect 266872 6752 358544 6780
rect 266872 6740 266878 6752
rect 358538 6740 358544 6752
rect 358596 6740 358602 6792
rect 192018 6672 192024 6724
rect 192076 6712 192082 6724
rect 248874 6712 248880 6724
rect 192076 6684 248880 6712
rect 192076 6672 192082 6684
rect 248874 6672 248880 6684
rect 248932 6672 248938 6724
rect 266722 6672 266728 6724
rect 266780 6712 266786 6724
rect 362126 6712 362132 6724
rect 266780 6684 362132 6712
rect 266780 6672 266786 6684
rect 362126 6672 362132 6684
rect 362184 6672 362190 6724
rect 188430 6604 188436 6656
rect 188488 6644 188494 6656
rect 248782 6644 248788 6656
rect 188488 6616 248788 6644
rect 188488 6604 188494 6616
rect 248782 6604 248788 6616
rect 248840 6604 248846 6656
rect 267458 6604 267464 6656
rect 267516 6644 267522 6656
rect 365806 6644 365812 6656
rect 267516 6616 365812 6644
rect 267516 6604 267522 6616
rect 365806 6604 365812 6616
rect 365864 6604 365870 6656
rect 184842 6536 184848 6588
rect 184900 6576 184906 6588
rect 248690 6576 248696 6588
rect 184900 6548 248696 6576
rect 184900 6536 184906 6548
rect 248690 6536 248696 6548
rect 248748 6536 248754 6588
rect 269022 6536 269028 6588
rect 269080 6576 269086 6588
rect 369210 6576 369216 6588
rect 269080 6548 369216 6576
rect 269080 6536 269086 6548
rect 369210 6536 369216 6548
rect 369268 6536 369274 6588
rect 181346 6468 181352 6520
rect 181404 6508 181410 6520
rect 248598 6508 248604 6520
rect 181404 6480 248604 6508
rect 181404 6468 181410 6480
rect 248598 6468 248604 6480
rect 248656 6468 248662 6520
rect 268838 6468 268844 6520
rect 268896 6508 268902 6520
rect 372798 6508 372804 6520
rect 268896 6480 372804 6508
rect 268896 6468 268902 6480
rect 372798 6468 372804 6480
rect 372856 6468 372862 6520
rect 177758 6400 177764 6452
rect 177816 6440 177822 6452
rect 248138 6440 248144 6452
rect 177816 6412 248144 6440
rect 177816 6400 177822 6412
rect 248138 6400 248144 6412
rect 248196 6400 248202 6452
rect 267918 6400 267924 6452
rect 267976 6440 267982 6452
rect 376386 6440 376392 6452
rect 267976 6412 376392 6440
rect 267976 6400 267982 6412
rect 376386 6400 376392 6412
rect 376444 6400 376450 6452
rect 174170 6332 174176 6384
rect 174228 6372 174234 6384
rect 247862 6372 247868 6384
rect 174228 6344 247868 6372
rect 174228 6332 174234 6344
rect 247862 6332 247868 6344
rect 247920 6332 247926 6384
rect 268194 6332 268200 6384
rect 268252 6372 268258 6384
rect 379974 6372 379980 6384
rect 268252 6344 379980 6372
rect 268252 6332 268258 6344
rect 379974 6332 379980 6344
rect 380032 6332 380038 6384
rect 134886 6264 134892 6316
rect 134944 6304 134950 6316
rect 243262 6304 243268 6316
rect 134944 6276 243268 6304
rect 134944 6264 134950 6276
rect 243262 6264 243268 6276
rect 243320 6264 243326 6316
rect 270126 6264 270132 6316
rect 270184 6304 270190 6316
rect 383562 6304 383568 6316
rect 270184 6276 383568 6304
rect 270184 6264 270190 6276
rect 383562 6264 383568 6276
rect 383620 6264 383626 6316
rect 131390 6196 131396 6248
rect 131448 6236 131454 6248
rect 243170 6236 243176 6248
rect 131448 6208 243176 6236
rect 131448 6196 131454 6208
rect 243170 6196 243176 6208
rect 243228 6196 243234 6248
rect 269482 6196 269488 6248
rect 269540 6236 269546 6248
rect 387058 6236 387064 6248
rect 269540 6208 387064 6236
rect 269540 6196 269546 6208
rect 387058 6196 387064 6208
rect 387116 6196 387122 6248
rect 12434 6128 12440 6180
rect 12492 6168 12498 6180
rect 230842 6168 230848 6180
rect 12492 6140 230848 6168
rect 12492 6128 12498 6140
rect 230842 6128 230848 6140
rect 230900 6128 230906 6180
rect 234798 6128 234804 6180
rect 234856 6168 234862 6180
rect 254486 6168 254492 6180
rect 234856 6140 254492 6168
rect 234856 6128 234862 6140
rect 254486 6128 254492 6140
rect 254544 6128 254550 6180
rect 270218 6128 270224 6180
rect 270276 6168 270282 6180
rect 390646 6168 390652 6180
rect 270276 6140 390652 6168
rect 270276 6128 270282 6140
rect 390646 6128 390652 6140
rect 390704 6128 390710 6180
rect 202690 6060 202696 6112
rect 202748 6100 202754 6112
rect 250806 6100 250812 6112
rect 202748 6072 250812 6100
rect 202748 6060 202754 6072
rect 250806 6060 250812 6072
rect 250864 6060 250870 6112
rect 265342 6060 265348 6112
rect 265400 6100 265406 6112
rect 351362 6100 351368 6112
rect 265400 6072 351368 6100
rect 265400 6060 265406 6072
rect 351362 6060 351368 6072
rect 351420 6060 351426 6112
rect 238386 5992 238392 6044
rect 238444 6032 238450 6044
rect 254578 6032 254584 6044
rect 238444 6004 254584 6032
rect 238444 5992 238450 6004
rect 254578 5992 254584 6004
rect 254636 5992 254642 6044
rect 266078 5992 266084 6044
rect 266136 6032 266142 6044
rect 347866 6032 347872 6044
rect 266136 6004 347872 6032
rect 266136 5992 266142 6004
rect 347866 5992 347872 6004
rect 347924 5992 347930 6044
rect 265526 5924 265532 5976
rect 265584 5964 265590 5976
rect 344278 5964 344284 5976
rect 265584 5936 344284 5964
rect 265584 5924 265590 5936
rect 344278 5924 344284 5936
rect 344336 5924 344342 5976
rect 265986 5856 265992 5908
rect 266044 5896 266050 5908
rect 340690 5896 340696 5908
rect 266044 5868 340696 5896
rect 266044 5856 266050 5868
rect 340690 5856 340696 5868
rect 340748 5856 340754 5908
rect 264330 5788 264336 5840
rect 264388 5828 264394 5840
rect 337102 5828 337108 5840
rect 264388 5800 337108 5828
rect 264388 5788 264394 5800
rect 337102 5788 337108 5800
rect 337160 5788 337166 5840
rect 264238 5720 264244 5772
rect 264296 5760 264302 5772
rect 333606 5760 333612 5772
rect 264296 5732 333612 5760
rect 264296 5720 264302 5732
rect 333606 5720 333612 5732
rect 333664 5720 333670 5772
rect 264054 5652 264060 5704
rect 264112 5692 264118 5704
rect 330018 5692 330024 5704
rect 264112 5664 330024 5692
rect 264112 5652 264118 5664
rect 330018 5652 330024 5664
rect 330076 5652 330082 5704
rect 262766 5584 262772 5636
rect 262824 5624 262830 5636
rect 326430 5624 326436 5636
rect 262824 5596 326436 5624
rect 262824 5584 262830 5596
rect 326430 5584 326436 5596
rect 326488 5584 326494 5636
rect 262674 5516 262680 5568
rect 262732 5556 262738 5568
rect 322842 5556 322848 5568
rect 262732 5528 322848 5556
rect 262732 5516 262738 5528
rect 322842 5516 322848 5528
rect 322900 5516 322906 5568
rect 197998 5448 198004 5500
rect 198056 5488 198062 5500
rect 244277 5491 244335 5497
rect 244277 5488 244289 5491
rect 198056 5460 244289 5488
rect 198056 5448 198062 5460
rect 244277 5457 244289 5460
rect 244323 5457 244335 5491
rect 244277 5451 244335 5457
rect 244366 5448 244372 5500
rect 244424 5488 244430 5500
rect 247678 5488 247684 5500
rect 244424 5460 247684 5488
rect 244424 5448 244430 5460
rect 247678 5448 247684 5460
rect 247736 5448 247742 5500
rect 257706 5448 257712 5500
rect 257764 5488 257770 5500
rect 270494 5488 270500 5500
rect 257764 5460 270500 5488
rect 257764 5448 257770 5460
rect 270494 5448 270500 5460
rect 270552 5448 270558 5500
rect 194410 5380 194416 5432
rect 194468 5420 194474 5432
rect 249978 5420 249984 5432
rect 194468 5392 249984 5420
rect 194468 5380 194474 5392
rect 249978 5380 249984 5392
rect 250036 5380 250042 5432
rect 258166 5380 258172 5432
rect 258224 5420 258230 5432
rect 274082 5420 274088 5432
rect 258224 5392 274088 5420
rect 258224 5380 258230 5392
rect 274082 5380 274088 5392
rect 274140 5380 274146 5432
rect 190822 5312 190828 5364
rect 190880 5352 190886 5364
rect 248506 5352 248512 5364
rect 190880 5324 248512 5352
rect 190880 5312 190886 5324
rect 248506 5312 248512 5324
rect 248564 5312 248570 5364
rect 257522 5312 257528 5364
rect 257580 5352 257586 5364
rect 272886 5352 272892 5364
rect 257580 5324 272892 5352
rect 257580 5312 257586 5324
rect 272886 5312 272892 5324
rect 272944 5312 272950 5364
rect 137278 5244 137284 5296
rect 137336 5284 137342 5296
rect 137336 5256 143948 5284
rect 137336 5244 137342 5256
rect 140866 5176 140872 5228
rect 140924 5216 140930 5228
rect 142062 5216 142068 5228
rect 140924 5188 142068 5216
rect 140924 5176 140930 5188
rect 142062 5176 142068 5188
rect 142120 5176 142126 5228
rect 143920 5216 143948 5256
rect 187234 5244 187240 5296
rect 187292 5284 187298 5296
rect 249610 5284 249616 5296
rect 187292 5256 249616 5284
rect 187292 5244 187298 5256
rect 249610 5244 249616 5256
rect 249668 5244 249674 5296
rect 259270 5244 259276 5296
rect 259328 5284 259334 5296
rect 276474 5284 276480 5296
rect 259328 5256 276480 5284
rect 259328 5244 259334 5256
rect 276474 5244 276480 5256
rect 276532 5244 276538 5296
rect 243998 5216 244004 5228
rect 143920 5188 244004 5216
rect 243998 5176 244004 5188
rect 244056 5176 244062 5228
rect 244277 5219 244335 5225
rect 244277 5185 244289 5219
rect 244323 5216 244335 5219
rect 251082 5216 251088 5228
rect 244323 5188 251088 5216
rect 244323 5185 244335 5188
rect 244277 5179 244335 5185
rect 251082 5176 251088 5188
rect 251140 5176 251146 5228
rect 258902 5176 258908 5228
rect 258960 5216 258966 5228
rect 277670 5216 277676 5228
rect 258960 5188 277676 5216
rect 258960 5176 258966 5188
rect 277670 5176 277676 5188
rect 277728 5176 277734 5228
rect 133782 5108 133788 5160
rect 133840 5148 133846 5160
rect 243722 5148 243728 5160
rect 133840 5120 243728 5148
rect 133840 5108 133846 5120
rect 243722 5108 243728 5120
rect 243780 5108 243786 5160
rect 258534 5108 258540 5160
rect 258592 5148 258598 5160
rect 280062 5148 280068 5160
rect 258592 5120 280068 5148
rect 258592 5108 258598 5120
rect 280062 5108 280068 5120
rect 280120 5108 280126 5160
rect 130194 5040 130200 5092
rect 130252 5080 130258 5092
rect 243630 5080 243636 5092
rect 130252 5052 243636 5080
rect 130252 5040 130258 5052
rect 243630 5040 243636 5052
rect 243688 5040 243694 5092
rect 258810 5040 258816 5092
rect 258868 5080 258874 5092
rect 281258 5080 281264 5092
rect 258868 5052 281264 5080
rect 258868 5040 258874 5052
rect 281258 5040 281264 5052
rect 281316 5040 281322 5092
rect 7650 4972 7656 5024
rect 7708 5012 7714 5024
rect 224129 5015 224187 5021
rect 224129 5012 224141 5015
rect 7708 4984 224141 5012
rect 7708 4972 7714 4984
rect 224129 4981 224141 4984
rect 224175 4981 224187 5015
rect 224129 4975 224187 4981
rect 224221 5015 224279 5021
rect 224221 4981 224233 5015
rect 224267 5012 224279 5015
rect 229186 5012 229192 5024
rect 224267 4984 229192 5012
rect 224267 4981 224279 4984
rect 224221 4975 224279 4981
rect 229186 4972 229192 4984
rect 229244 4972 229250 5024
rect 258350 4972 258356 5024
rect 258408 5012 258414 5024
rect 283650 5012 283656 5024
rect 258408 4984 283656 5012
rect 258408 4972 258414 4984
rect 283650 4972 283656 4984
rect 283708 4972 283714 5024
rect 2866 4904 2872 4956
rect 2924 4944 2930 4956
rect 229370 4944 229376 4956
rect 2924 4916 229376 4944
rect 2924 4904 2930 4916
rect 229370 4904 229376 4916
rect 229428 4904 229434 4956
rect 240778 4904 240784 4956
rect 240836 4944 240842 4956
rect 254302 4944 254308 4956
rect 240836 4916 254308 4944
rect 240836 4904 240842 4916
rect 254302 4904 254308 4916
rect 254360 4904 254366 4956
rect 258258 4904 258264 4956
rect 258316 4944 258322 4956
rect 284754 4944 284760 4956
rect 258316 4916 284760 4944
rect 258316 4904 258322 4916
rect 284754 4904 284760 4916
rect 284812 4904 284818 4956
rect 1670 4836 1676 4888
rect 1728 4876 1734 4888
rect 1728 4848 224356 4876
rect 1728 4836 1734 4848
rect 566 4768 572 4820
rect 624 4808 630 4820
rect 224221 4811 224279 4817
rect 224221 4808 224233 4811
rect 624 4780 224233 4808
rect 624 4768 630 4780
rect 224221 4777 224233 4780
rect 224267 4777 224279 4811
rect 224328 4808 224356 4848
rect 237282 4836 237288 4888
rect 237340 4876 237346 4888
rect 254210 4876 254216 4888
rect 237340 4848 254216 4876
rect 237340 4836 237346 4848
rect 254210 4836 254216 4848
rect 254268 4836 254274 4888
rect 260190 4836 260196 4888
rect 260248 4876 260254 4888
rect 287146 4876 287152 4888
rect 260248 4848 287152 4876
rect 260248 4836 260254 4848
rect 287146 4836 287152 4848
rect 287204 4836 287210 4888
rect 229278 4808 229284 4820
rect 224328 4780 229284 4808
rect 224221 4771 224279 4777
rect 229278 4768 229284 4780
rect 229336 4768 229342 4820
rect 233694 4768 233700 4820
rect 233752 4808 233758 4820
rect 254394 4808 254400 4820
rect 233752 4780 254400 4808
rect 233752 4768 233758 4780
rect 254394 4768 254400 4780
rect 254452 4768 254458 4820
rect 260098 4768 260104 4820
rect 260156 4808 260162 4820
rect 290734 4808 290740 4820
rect 260156 4780 290740 4808
rect 260156 4768 260162 4780
rect 290734 4768 290740 4780
rect 290792 4768 290798 4820
rect 316678 4768 316684 4820
rect 316736 4808 316742 4820
rect 486970 4808 486976 4820
rect 316736 4780 486976 4808
rect 316736 4768 316742 4780
rect 486970 4768 486976 4780
rect 487028 4768 487034 4820
rect 489178 4768 489184 4820
rect 489236 4808 489242 4820
rect 497734 4808 497740 4820
rect 489236 4780 497740 4808
rect 489236 4768 489242 4780
rect 497734 4768 497740 4780
rect 497792 4768 497798 4820
rect 201494 4700 201500 4752
rect 201552 4740 201558 4752
rect 249886 4740 249892 4752
rect 201552 4712 249892 4740
rect 201552 4700 201558 4712
rect 249886 4700 249892 4712
rect 249944 4700 249950 4752
rect 257062 4700 257068 4752
rect 257120 4740 257126 4752
rect 269298 4740 269304 4752
rect 257120 4712 269304 4740
rect 257120 4700 257126 4712
rect 269298 4700 269304 4712
rect 269356 4700 269362 4752
rect 205082 4632 205088 4684
rect 205140 4672 205146 4684
rect 250990 4672 250996 4684
rect 205140 4644 250996 4672
rect 205140 4632 205146 4644
rect 250990 4632 250996 4644
rect 251048 4632 251054 4684
rect 224129 4607 224187 4613
rect 224129 4573 224141 4607
rect 224175 4604 224187 4607
rect 230750 4604 230756 4616
rect 224175 4576 230756 4604
rect 224175 4573 224187 4576
rect 224129 4567 224187 4573
rect 230750 4564 230756 4576
rect 230808 4564 230814 4616
rect 124214 4156 124220 4208
rect 124272 4196 124278 4208
rect 125410 4196 125416 4208
rect 124272 4168 125416 4196
rect 124272 4156 124278 4168
rect 125410 4156 125416 4168
rect 125468 4156 125474 4208
rect 150434 4156 150440 4208
rect 150492 4196 150498 4208
rect 151630 4196 151636 4208
rect 150492 4168 151636 4196
rect 150492 4156 150498 4168
rect 151630 4156 151636 4168
rect 151688 4156 151694 4208
rect 158714 4156 158720 4208
rect 158772 4196 158778 4208
rect 160002 4196 160008 4208
rect 158772 4168 160008 4196
rect 158772 4156 158778 4168
rect 160002 4156 160008 4168
rect 160060 4156 160066 4208
rect 167086 4156 167092 4208
rect 167144 4196 167150 4208
rect 168282 4196 168288 4208
rect 167144 4168 168288 4196
rect 167144 4156 167150 4168
rect 168282 4156 168288 4168
rect 168340 4156 168346 4208
rect 209866 4156 209872 4208
rect 209924 4196 209930 4208
rect 211062 4196 211068 4208
rect 209924 4168 211068 4196
rect 209924 4156 209930 4168
rect 211062 4156 211068 4168
rect 211120 4156 211126 4208
rect 227714 4156 227720 4208
rect 227772 4196 227778 4208
rect 229002 4196 229008 4208
rect 227772 4168 229008 4196
rect 227772 4156 227778 4168
rect 229002 4156 229008 4168
rect 229060 4156 229066 4208
rect 272518 4156 272524 4208
rect 272576 4196 272582 4208
rect 275278 4196 275284 4208
rect 272576 4168 275284 4196
rect 272576 4156 272582 4168
rect 275278 4156 275284 4168
rect 275336 4156 275342 4208
rect 296714 4156 296720 4208
rect 296772 4196 296778 4208
rect 297910 4196 297916 4208
rect 296772 4168 297916 4196
rect 296772 4156 296778 4168
rect 297910 4156 297916 4168
rect 297968 4156 297974 4208
rect 347774 4156 347780 4208
rect 347832 4196 347838 4208
rect 349062 4196 349068 4208
rect 347832 4168 349068 4196
rect 347832 4156 347838 4168
rect 349062 4156 349068 4168
rect 349120 4156 349126 4208
rect 356054 4156 356060 4208
rect 356112 4196 356118 4208
rect 357342 4196 357348 4208
rect 356112 4168 357348 4196
rect 356112 4156 356118 4168
rect 357342 4156 357348 4168
rect 357400 4156 357406 4208
rect 365714 4156 365720 4208
rect 365772 4196 365778 4208
rect 366910 4196 366916 4208
rect 365772 4168 366916 4196
rect 365772 4156 365778 4168
rect 366910 4156 366916 4168
rect 366968 4156 366974 4208
rect 373994 4156 374000 4208
rect 374052 4196 374058 4208
rect 375190 4196 375196 4208
rect 374052 4168 375196 4196
rect 374052 4156 374058 4168
rect 375190 4156 375196 4168
rect 375248 4156 375254 4208
rect 20714 4088 20720 4140
rect 20772 4128 20778 4140
rect 28258 4128 28264 4140
rect 20772 4100 28264 4128
rect 20772 4088 20778 4100
rect 28258 4088 28264 4100
rect 28316 4088 28322 4140
rect 79042 4088 79048 4140
rect 79100 4128 79106 4140
rect 238018 4128 238024 4140
rect 79100 4100 238024 4128
rect 79100 4088 79106 4100
rect 238018 4088 238024 4100
rect 238076 4088 238082 4140
rect 255498 4088 255504 4140
rect 255556 4128 255562 4140
rect 256234 4128 256240 4140
rect 255556 4100 256240 4128
rect 255556 4088 255562 4100
rect 256234 4088 256240 4100
rect 256292 4088 256298 4140
rect 258442 4088 258448 4140
rect 258500 4128 258506 4140
rect 259822 4128 259828 4140
rect 258500 4100 259828 4128
rect 258500 4088 258506 4100
rect 259822 4088 259828 4100
rect 259880 4088 259886 4140
rect 262858 4088 262864 4140
rect 262916 4128 262922 4140
rect 264606 4128 264612 4140
rect 262916 4100 264612 4128
rect 262916 4088 262922 4100
rect 264606 4088 264612 4100
rect 264664 4088 264670 4140
rect 273898 4088 273904 4140
rect 273956 4128 273962 4140
rect 425054 4128 425060 4140
rect 273956 4100 425060 4128
rect 273956 4088 273962 4100
rect 425054 4088 425060 4100
rect 425112 4088 425118 4140
rect 556798 4088 556804 4140
rect 556856 4128 556862 4140
rect 559558 4128 559564 4140
rect 556856 4100 559564 4128
rect 556856 4088 556862 4100
rect 559558 4088 559564 4100
rect 559616 4088 559622 4140
rect 13630 4020 13636 4072
rect 13688 4060 13694 4072
rect 17218 4060 17224 4072
rect 13688 4032 17224 4060
rect 13688 4020 13694 4032
rect 17218 4020 17224 4032
rect 17276 4020 17282 4072
rect 84102 4020 84108 4072
rect 84160 4060 84166 4072
rect 93949 4063 94007 4069
rect 93949 4060 93961 4063
rect 84160 4032 93961 4060
rect 84160 4020 84166 4032
rect 93949 4029 93961 4032
rect 93995 4029 94007 4063
rect 93949 4023 94007 4029
rect 103333 4063 103391 4069
rect 103333 4029 103345 4063
rect 103379 4060 103391 4063
rect 232317 4063 232375 4069
rect 232317 4060 232329 4063
rect 103379 4032 232329 4060
rect 103379 4029 103391 4032
rect 103333 4023 103391 4029
rect 232317 4029 232329 4032
rect 232363 4029 232375 4063
rect 232317 4023 232375 4029
rect 232409 4063 232467 4069
rect 232409 4029 232421 4063
rect 232455 4060 232467 4063
rect 235810 4060 235816 4072
rect 232455 4032 235816 4060
rect 232455 4029 232467 4032
rect 232409 4023 232467 4029
rect 235810 4020 235816 4032
rect 235868 4020 235874 4072
rect 255038 4020 255044 4072
rect 255096 4060 255102 4072
rect 255866 4060 255872 4072
rect 255096 4032 255872 4060
rect 255096 4020 255102 4032
rect 255866 4020 255872 4032
rect 255924 4020 255930 4072
rect 257338 4020 257344 4072
rect 257396 4060 257402 4072
rect 258626 4060 258632 4072
rect 257396 4032 258632 4060
rect 257396 4020 257402 4032
rect 258626 4020 258632 4032
rect 258684 4020 258690 4072
rect 273714 4020 273720 4072
rect 273772 4060 273778 4072
rect 428734 4060 428740 4072
rect 273772 4032 428740 4060
rect 273772 4020 273778 4032
rect 428734 4020 428740 4032
rect 428792 4020 428798 4072
rect 71866 3952 71872 4004
rect 71924 3992 71930 4004
rect 74537 3995 74595 4001
rect 74537 3992 74549 3995
rect 71924 3964 74549 3992
rect 71924 3952 71930 3964
rect 74537 3961 74549 3964
rect 74583 3961 74595 3995
rect 74537 3955 74595 3961
rect 84013 3995 84071 4001
rect 84013 3961 84025 3995
rect 84059 3992 84071 3995
rect 93857 3995 93915 4001
rect 93857 3992 93869 3995
rect 84059 3964 93869 3992
rect 84059 3961 84071 3964
rect 84013 3955 84071 3961
rect 93857 3961 93869 3964
rect 93903 3961 93915 3995
rect 93857 3955 93915 3961
rect 103425 3995 103483 4001
rect 103425 3961 103437 3995
rect 103471 3992 103483 3995
rect 237006 3992 237012 4004
rect 103471 3964 237012 3992
rect 103471 3961 103483 3964
rect 103425 3955 103483 3961
rect 237006 3952 237012 3964
rect 237064 3952 237070 4004
rect 257798 3952 257804 4004
rect 257856 3992 257862 4004
rect 261018 3992 261024 4004
rect 257856 3964 261024 3992
rect 257856 3952 257862 3964
rect 261018 3952 261024 3964
rect 261076 3952 261082 4004
rect 273438 3952 273444 4004
rect 273496 3992 273502 4004
rect 432322 3992 432328 4004
rect 273496 3964 432328 3992
rect 273496 3952 273502 3964
rect 432322 3952 432328 3964
rect 432380 3952 432386 4004
rect 433337 3995 433395 4001
rect 433337 3961 433349 3995
rect 433383 3992 433395 3995
rect 439406 3992 439412 4004
rect 433383 3964 439412 3992
rect 433383 3961 433395 3964
rect 433337 3955 433395 3961
rect 439406 3952 439412 3964
rect 439464 3952 439470 4004
rect 68278 3884 68284 3936
rect 68336 3924 68342 3936
rect 236270 3924 236276 3936
rect 68336 3896 236276 3924
rect 68336 3884 68342 3896
rect 236270 3884 236276 3896
rect 236328 3884 236334 3936
rect 248969 3927 249027 3933
rect 248969 3893 248981 3927
rect 249015 3924 249027 3927
rect 254946 3924 254952 3936
rect 249015 3896 254952 3924
rect 249015 3893 249027 3896
rect 248969 3887 249027 3893
rect 254946 3884 254952 3896
rect 255004 3884 255010 3936
rect 257982 3884 257988 3936
rect 258040 3924 258046 3936
rect 262214 3924 262220 3936
rect 258040 3896 262220 3924
rect 258040 3884 258046 3896
rect 262214 3884 262220 3896
rect 262272 3884 262278 3936
rect 275738 3884 275744 3936
rect 275796 3924 275802 3936
rect 435818 3924 435824 3936
rect 275796 3896 435824 3924
rect 275796 3884 275802 3896
rect 435818 3884 435824 3896
rect 435876 3884 435882 3936
rect 64690 3816 64696 3868
rect 64748 3856 64754 3868
rect 236178 3856 236184 3868
rect 64748 3828 236184 3856
rect 64748 3816 64754 3828
rect 236178 3816 236184 3828
rect 236236 3816 236242 3868
rect 246758 3816 246764 3868
rect 246816 3856 246822 3868
rect 255314 3856 255320 3868
rect 246816 3828 255320 3856
rect 246816 3816 246822 3828
rect 255314 3816 255320 3828
rect 255372 3816 255378 3868
rect 257890 3816 257896 3868
rect 257948 3856 257954 3868
rect 263410 3856 263416 3868
rect 257948 3828 263416 3856
rect 257948 3816 257954 3828
rect 263410 3816 263416 3828
rect 263468 3816 263474 3868
rect 275094 3816 275100 3868
rect 275152 3856 275158 3868
rect 433337 3859 433395 3865
rect 433337 3856 433349 3859
rect 275152 3828 433349 3856
rect 275152 3816 275158 3828
rect 433337 3825 433349 3828
rect 433383 3825 433395 3859
rect 433337 3819 433395 3825
rect 433426 3816 433432 3868
rect 433484 3856 433490 3868
rect 434622 3856 434628 3868
rect 433484 3828 434628 3856
rect 433484 3816 433490 3828
rect 434622 3816 434628 3828
rect 434680 3816 434686 3868
rect 61194 3748 61200 3800
rect 61252 3788 61258 3800
rect 236086 3788 236092 3800
rect 61252 3760 236092 3788
rect 61252 3748 61258 3760
rect 236086 3748 236092 3760
rect 236144 3748 236150 3800
rect 275002 3748 275008 3800
rect 275060 3788 275066 3800
rect 442994 3788 443000 3800
rect 275060 3760 443000 3788
rect 275060 3748 275066 3760
rect 442994 3748 443000 3760
rect 443052 3748 443058 3800
rect 567838 3748 567844 3800
rect 567896 3788 567902 3800
rect 573818 3788 573824 3800
rect 567896 3760 573824 3788
rect 567896 3748 567902 3760
rect 573818 3748 573824 3760
rect 573876 3748 573882 3800
rect 44542 3680 44548 3732
rect 44600 3720 44606 3732
rect 46198 3720 46204 3732
rect 44600 3692 46204 3720
rect 44600 3680 44606 3692
rect 46198 3680 46204 3692
rect 46256 3680 46262 3732
rect 57606 3680 57612 3732
rect 57664 3720 57670 3732
rect 232409 3723 232467 3729
rect 232409 3720 232421 3723
rect 57664 3692 232421 3720
rect 57664 3680 57670 3692
rect 232409 3689 232421 3692
rect 232455 3689 232467 3723
rect 232409 3683 232467 3689
rect 233053 3723 233111 3729
rect 233053 3689 233065 3723
rect 233099 3720 233111 3723
rect 241054 3720 241060 3732
rect 233099 3692 241060 3720
rect 233099 3689 233111 3692
rect 233053 3683 233111 3689
rect 241054 3680 241060 3692
rect 241112 3680 241118 3732
rect 247954 3680 247960 3732
rect 248012 3720 248018 3732
rect 254670 3720 254676 3732
rect 248012 3692 254676 3720
rect 248012 3680 248018 3692
rect 254670 3680 254676 3692
rect 254728 3680 254734 3732
rect 275373 3723 275431 3729
rect 275373 3689 275385 3723
rect 275419 3720 275431 3723
rect 446582 3720 446588 3732
rect 275419 3692 446588 3720
rect 275419 3689 275431 3692
rect 275373 3683 275431 3689
rect 446582 3680 446588 3692
rect 446640 3680 446646 3732
rect 573358 3680 573364 3732
rect 573416 3720 573422 3732
rect 579798 3720 579804 3732
rect 573416 3692 579804 3720
rect 573416 3680 573422 3692
rect 579798 3680 579804 3692
rect 579856 3680 579862 3732
rect 46934 3612 46940 3664
rect 46992 3652 46998 3664
rect 46992 3624 53880 3652
rect 46992 3612 46998 3624
rect 34974 3544 34980 3596
rect 35032 3584 35038 3596
rect 35032 3556 37320 3584
rect 35032 3544 35038 3556
rect 8846 3476 8852 3528
rect 8904 3516 8910 3528
rect 9582 3516 9588 3528
rect 8904 3488 9588 3516
rect 8904 3476 8910 3488
rect 9582 3476 9588 3488
rect 9640 3476 9646 3528
rect 10042 3476 10048 3528
rect 10100 3516 10106 3528
rect 14458 3516 14464 3528
rect 10100 3488 14464 3516
rect 10100 3476 10106 3488
rect 14458 3476 14464 3488
rect 14516 3476 14522 3528
rect 18322 3476 18328 3528
rect 18380 3516 18386 3528
rect 19978 3516 19984 3528
rect 18380 3488 19984 3516
rect 18380 3476 18386 3488
rect 19978 3476 19984 3488
rect 20036 3476 20042 3528
rect 23106 3476 23112 3528
rect 23164 3516 23170 3528
rect 24118 3516 24124 3528
rect 23164 3488 24124 3516
rect 23164 3476 23170 3488
rect 24118 3476 24124 3488
rect 24176 3476 24182 3528
rect 26694 3476 26700 3528
rect 26752 3516 26758 3528
rect 27522 3516 27528 3528
rect 26752 3488 27528 3516
rect 26752 3476 26758 3488
rect 27522 3476 27528 3488
rect 27580 3476 27586 3528
rect 32398 3516 32404 3528
rect 28736 3488 32404 3516
rect 5258 3408 5264 3460
rect 5316 3448 5322 3460
rect 10318 3448 10324 3460
rect 5316 3420 10324 3448
rect 5316 3408 5322 3420
rect 10318 3408 10324 3420
rect 10376 3408 10382 3460
rect 19518 3408 19524 3460
rect 19576 3448 19582 3460
rect 28736 3448 28764 3488
rect 32398 3476 32404 3488
rect 32456 3476 32462 3528
rect 33870 3476 33876 3528
rect 33928 3516 33934 3528
rect 34422 3516 34428 3528
rect 33928 3488 34428 3516
rect 33928 3476 33934 3488
rect 34422 3476 34428 3488
rect 34480 3476 34486 3528
rect 37292 3516 37320 3556
rect 37366 3544 37372 3596
rect 37424 3584 37430 3596
rect 38562 3584 38568 3596
rect 37424 3556 38568 3584
rect 37424 3544 37430 3556
rect 38562 3544 38568 3556
rect 38620 3544 38626 3596
rect 43438 3584 43444 3596
rect 38672 3556 43444 3584
rect 38672 3516 38700 3556
rect 43438 3544 43444 3556
rect 43496 3544 43502 3596
rect 50522 3544 50528 3596
rect 50580 3584 50586 3596
rect 50982 3584 50988 3596
rect 50580 3556 50988 3584
rect 50580 3544 50586 3556
rect 50982 3544 50988 3556
rect 51040 3544 51046 3596
rect 51626 3544 51632 3596
rect 51684 3584 51690 3596
rect 52362 3584 52368 3596
rect 51684 3556 52368 3584
rect 51684 3544 51690 3556
rect 52362 3544 52368 3556
rect 52420 3544 52426 3596
rect 52822 3544 52828 3596
rect 52880 3584 52886 3596
rect 53742 3584 53748 3596
rect 52880 3556 53748 3584
rect 52880 3544 52886 3556
rect 53742 3544 53748 3556
rect 53800 3544 53806 3596
rect 53852 3584 53880 3624
rect 54018 3612 54024 3664
rect 54076 3652 54082 3664
rect 235166 3652 235172 3664
rect 54076 3624 235172 3652
rect 54076 3612 54082 3624
rect 235166 3612 235172 3624
rect 235224 3612 235230 3664
rect 245562 3612 245568 3664
rect 245620 3652 245626 3664
rect 255130 3652 255136 3664
rect 245620 3624 255136 3652
rect 245620 3612 245626 3624
rect 255130 3612 255136 3624
rect 255188 3612 255194 3664
rect 277118 3612 277124 3664
rect 277176 3652 277182 3664
rect 450170 3652 450176 3664
rect 277176 3624 450176 3652
rect 277176 3612 277182 3624
rect 450170 3612 450176 3624
rect 450228 3612 450234 3664
rect 502426 3612 502432 3664
rect 502484 3652 502490 3664
rect 503622 3652 503628 3664
rect 502484 3624 503628 3652
rect 502484 3612 502490 3624
rect 503622 3612 503628 3624
rect 503680 3612 503686 3664
rect 536926 3612 536932 3664
rect 536984 3652 536990 3664
rect 538122 3652 538128 3664
rect 536984 3624 538128 3652
rect 536984 3612 536990 3624
rect 538122 3612 538128 3624
rect 538180 3612 538186 3664
rect 546494 3612 546500 3664
rect 546552 3652 546558 3664
rect 547690 3652 547696 3664
rect 546552 3624 547696 3652
rect 546552 3612 546558 3624
rect 547690 3612 547696 3624
rect 547748 3612 547754 3664
rect 563146 3612 563152 3664
rect 563204 3652 563210 3664
rect 564342 3652 564348 3664
rect 563204 3624 564348 3652
rect 563204 3612 563210 3624
rect 564342 3612 564348 3624
rect 564400 3612 564406 3664
rect 565078 3612 565084 3664
rect 565136 3652 565142 3664
rect 566734 3652 566740 3664
rect 565136 3624 566740 3652
rect 565136 3612 565142 3624
rect 566734 3612 566740 3624
rect 566792 3612 566798 3664
rect 573450 3612 573456 3664
rect 573508 3652 573514 3664
rect 580994 3652 581000 3664
rect 573508 3624 581000 3652
rect 573508 3612 573514 3624
rect 580994 3612 581000 3624
rect 581052 3612 581058 3664
rect 231121 3587 231179 3593
rect 231121 3584 231133 3587
rect 53852 3556 231133 3584
rect 231121 3553 231133 3556
rect 231167 3553 231179 3587
rect 234062 3584 234068 3596
rect 231121 3547 231179 3553
rect 231228 3556 234068 3584
rect 37292 3488 38700 3516
rect 40954 3476 40960 3528
rect 41012 3516 41018 3528
rect 42058 3516 42064 3528
rect 41012 3488 42064 3516
rect 41012 3476 41018 3488
rect 42058 3476 42064 3488
rect 42116 3476 42122 3528
rect 42150 3476 42156 3528
rect 42208 3516 42214 3528
rect 42702 3516 42708 3528
rect 42208 3488 42708 3516
rect 42208 3476 42214 3488
rect 42702 3476 42708 3488
rect 42760 3476 42766 3528
rect 43346 3476 43352 3528
rect 43404 3516 43410 3528
rect 231228 3516 231256 3556
rect 234062 3544 234068 3556
rect 234120 3544 234126 3596
rect 238110 3584 238116 3596
rect 234172 3556 238116 3584
rect 43404 3488 231256 3516
rect 43404 3476 43410 3488
rect 231302 3476 231308 3528
rect 231360 3516 231366 3528
rect 231762 3516 231768 3528
rect 231360 3488 231768 3516
rect 231360 3476 231366 3488
rect 231762 3476 231768 3488
rect 231820 3476 231826 3528
rect 232498 3476 232504 3528
rect 232556 3516 232562 3528
rect 233142 3516 233148 3528
rect 232556 3488 233148 3516
rect 232556 3476 232562 3488
rect 233142 3476 233148 3488
rect 233200 3476 233206 3528
rect 233234 3476 233240 3528
rect 233292 3516 233298 3528
rect 234172 3516 234200 3556
rect 238110 3544 238116 3556
rect 238168 3544 238174 3596
rect 252646 3544 252652 3596
rect 252704 3584 252710 3596
rect 255774 3584 255780 3596
rect 252704 3556 255780 3584
rect 252704 3544 252710 3556
rect 255774 3544 255780 3556
rect 255832 3544 255838 3596
rect 276566 3544 276572 3596
rect 276624 3584 276630 3596
rect 453666 3584 453672 3596
rect 276624 3556 453672 3584
rect 276624 3544 276630 3556
rect 453666 3544 453672 3556
rect 453724 3544 453730 3596
rect 482278 3544 482284 3596
rect 482336 3584 482342 3596
rect 571061 3587 571119 3593
rect 571061 3584 571073 3587
rect 482336 3556 571073 3584
rect 482336 3544 482342 3556
rect 571061 3553 571073 3556
rect 571107 3553 571119 3587
rect 571061 3547 571119 3553
rect 571334 3544 571340 3596
rect 571392 3584 571398 3596
rect 572622 3584 572628 3596
rect 571392 3556 572628 3584
rect 571392 3544 571398 3556
rect 572622 3544 572628 3556
rect 572680 3544 572686 3596
rect 233292 3488 234200 3516
rect 233292 3476 233298 3488
rect 243170 3476 243176 3528
rect 243228 3516 243234 3528
rect 248969 3519 249027 3525
rect 248969 3516 248981 3519
rect 243228 3488 248981 3516
rect 243228 3476 243234 3488
rect 248969 3485 248981 3488
rect 249015 3485 249027 3519
rect 253934 3516 253940 3528
rect 248969 3479 249027 3485
rect 251008 3488 253940 3516
rect 19576 3420 28764 3448
rect 19576 3408 19582 3420
rect 29086 3408 29092 3460
rect 29144 3448 29150 3460
rect 35158 3448 35164 3460
rect 29144 3420 35164 3448
rect 29144 3408 29150 3420
rect 35158 3408 35164 3420
rect 35216 3408 35222 3460
rect 39758 3408 39764 3460
rect 39816 3448 39822 3460
rect 232317 3451 232375 3457
rect 39816 3420 231072 3448
rect 39816 3408 39822 3420
rect 55214 3340 55220 3392
rect 55272 3380 55278 3392
rect 56502 3380 56508 3392
rect 55272 3352 56508 3380
rect 55272 3340 55278 3352
rect 56502 3340 56508 3352
rect 56560 3340 56566 3392
rect 59998 3340 60004 3392
rect 60056 3380 60062 3392
rect 60642 3380 60648 3392
rect 60056 3352 60648 3380
rect 60056 3340 60062 3352
rect 60642 3340 60648 3352
rect 60700 3340 60706 3392
rect 63586 3340 63592 3392
rect 63644 3380 63650 3392
rect 64782 3380 64788 3392
rect 63644 3352 64788 3380
rect 63644 3340 63650 3352
rect 64782 3340 64788 3352
rect 64840 3340 64846 3392
rect 70670 3340 70676 3392
rect 70728 3380 70734 3392
rect 71682 3380 71688 3392
rect 70728 3352 71688 3380
rect 70728 3340 70734 3352
rect 71682 3340 71688 3352
rect 71740 3340 71746 3392
rect 77846 3340 77852 3392
rect 77904 3380 77910 3392
rect 78582 3380 78588 3392
rect 77904 3352 78588 3380
rect 77904 3340 77910 3352
rect 78582 3340 78588 3352
rect 78640 3340 78646 3392
rect 81434 3340 81440 3392
rect 81492 3380 81498 3392
rect 82722 3380 82728 3392
rect 81492 3352 82728 3380
rect 81492 3340 81498 3352
rect 82722 3340 82728 3352
rect 82780 3340 82786 3392
rect 230934 3380 230940 3392
rect 82832 3352 230940 3380
rect 27890 3204 27896 3256
rect 27948 3244 27954 3256
rect 31018 3244 31024 3256
rect 27948 3216 31024 3244
rect 27948 3204 27954 3216
rect 31018 3204 31024 3216
rect 31076 3204 31082 3256
rect 36170 3204 36176 3256
rect 36228 3244 36234 3256
rect 39298 3244 39304 3256
rect 36228 3216 39304 3244
rect 36228 3204 36234 3216
rect 39298 3204 39304 3216
rect 39356 3204 39362 3256
rect 82630 3204 82636 3256
rect 82688 3244 82694 3256
rect 82832 3244 82860 3352
rect 230934 3340 230940 3352
rect 230992 3340 230998 3392
rect 84930 3272 84936 3324
rect 84988 3312 84994 3324
rect 85482 3312 85488 3324
rect 84988 3284 85488 3312
rect 84988 3272 84994 3284
rect 85482 3272 85488 3284
rect 85540 3272 85546 3324
rect 229094 3312 229100 3324
rect 89640 3284 229100 3312
rect 82688 3216 82860 3244
rect 82688 3204 82694 3216
rect 86126 3204 86132 3256
rect 86184 3244 86190 3256
rect 89640 3244 89668 3284
rect 229094 3272 229100 3284
rect 229152 3272 229158 3324
rect 231044 3312 231072 3420
rect 232317 3417 232329 3451
rect 232363 3448 232375 3451
rect 238478 3448 238484 3460
rect 232363 3420 238484 3448
rect 232363 3417 232375 3420
rect 232317 3411 232375 3417
rect 238478 3408 238484 3420
rect 238536 3408 238542 3460
rect 239582 3408 239588 3460
rect 239640 3448 239646 3460
rect 251008 3448 251036 3488
rect 253934 3476 253940 3488
rect 253992 3476 253998 3528
rect 276382 3476 276388 3528
rect 276440 3516 276446 3528
rect 457254 3516 457260 3528
rect 276440 3488 457260 3516
rect 276440 3476 276446 3488
rect 457254 3476 457260 3488
rect 457312 3476 457318 3528
rect 467834 3476 467840 3528
rect 467892 3516 467898 3528
rect 469122 3516 469128 3528
rect 467892 3488 469128 3516
rect 467892 3476 467898 3488
rect 469122 3476 469128 3488
rect 469180 3476 469186 3528
rect 475378 3476 475384 3528
rect 475436 3516 475442 3528
rect 571981 3519 572039 3525
rect 571981 3516 571993 3519
rect 475436 3488 571993 3516
rect 475436 3476 475442 3488
rect 571981 3485 571993 3488
rect 572027 3485 572039 3519
rect 571981 3479 572039 3485
rect 239640 3420 251036 3448
rect 239640 3408 239646 3420
rect 253842 3408 253848 3460
rect 253900 3448 253906 3460
rect 255682 3448 255688 3460
rect 253900 3420 255688 3448
rect 253900 3408 253906 3420
rect 255682 3408 255688 3420
rect 255740 3408 255746 3460
rect 276106 3408 276112 3460
rect 276164 3448 276170 3460
rect 460842 3448 460848 3460
rect 276164 3420 460848 3448
rect 276164 3408 276170 3420
rect 460842 3408 460848 3420
rect 460900 3408 460906 3460
rect 471238 3408 471244 3460
rect 471296 3448 471302 3460
rect 582190 3448 582196 3460
rect 471296 3420 582196 3448
rect 471296 3408 471302 3420
rect 582190 3408 582196 3420
rect 582248 3408 582254 3460
rect 231121 3383 231179 3389
rect 231121 3349 231133 3383
rect 231167 3380 231179 3383
rect 234706 3380 234712 3392
rect 231167 3352 234712 3380
rect 231167 3349 231179 3352
rect 231121 3343 231179 3349
rect 234706 3340 234712 3352
rect 234764 3340 234770 3392
rect 249150 3340 249156 3392
rect 249208 3380 249214 3392
rect 255590 3380 255596 3392
rect 249208 3352 255596 3380
rect 249208 3340 249214 3352
rect 255590 3340 255596 3352
rect 255648 3340 255654 3392
rect 273806 3340 273812 3392
rect 273864 3380 273870 3392
rect 421558 3380 421564 3392
rect 273864 3352 421564 3380
rect 273864 3340 273870 3352
rect 421558 3340 421564 3352
rect 421616 3340 421622 3392
rect 494054 3340 494060 3392
rect 494112 3380 494118 3392
rect 495342 3380 495348 3392
rect 494112 3352 495348 3380
rect 494112 3340 494118 3352
rect 495342 3340 495348 3352
rect 495400 3340 495406 3392
rect 511994 3340 512000 3392
rect 512052 3380 512058 3392
rect 513190 3380 513196 3392
rect 512052 3352 513196 3380
rect 512052 3340 512058 3352
rect 513190 3340 513196 3352
rect 513248 3340 513254 3392
rect 528554 3340 528560 3392
rect 528612 3380 528618 3392
rect 529842 3380 529848 3392
rect 528612 3352 529848 3380
rect 528612 3340 528618 3352
rect 529842 3340 529848 3352
rect 529900 3340 529906 3392
rect 560938 3340 560944 3392
rect 560996 3380 561002 3392
rect 561950 3380 561956 3392
rect 560996 3352 561956 3380
rect 560996 3340 561002 3352
rect 561950 3340 561956 3352
rect 562008 3340 562014 3392
rect 571981 3383 572039 3389
rect 571981 3349 571993 3383
rect 572027 3380 572039 3383
rect 578602 3380 578608 3392
rect 572027 3352 578608 3380
rect 572027 3349 572039 3352
rect 571981 3343 572039 3349
rect 578602 3340 578608 3352
rect 578660 3340 578666 3392
rect 234154 3312 234160 3324
rect 231044 3284 234160 3312
rect 234154 3272 234160 3284
rect 234212 3272 234218 3324
rect 251450 3272 251456 3324
rect 251508 3312 251514 3324
rect 254762 3312 254768 3324
rect 251508 3284 254768 3312
rect 251508 3272 251514 3284
rect 254762 3272 254768 3284
rect 254820 3272 254826 3324
rect 272978 3272 272984 3324
rect 273036 3312 273042 3324
rect 417970 3312 417976 3324
rect 273036 3284 417976 3312
rect 273036 3272 273042 3284
rect 417970 3272 417976 3284
rect 418028 3272 418034 3324
rect 574830 3272 574836 3324
rect 574888 3312 574894 3324
rect 577406 3312 577412 3324
rect 574888 3284 577412 3312
rect 574888 3272 574894 3284
rect 577406 3272 577412 3284
rect 577464 3272 577470 3324
rect 86184 3216 89668 3244
rect 86184 3204 86190 3216
rect 89714 3204 89720 3256
rect 89772 3244 89778 3256
rect 89772 3216 233740 3244
rect 89772 3204 89778 3216
rect 75454 3136 75460 3188
rect 75512 3176 75518 3188
rect 84102 3176 84108 3188
rect 75512 3148 84108 3176
rect 75512 3136 75518 3148
rect 84102 3136 84108 3148
rect 84160 3136 84166 3188
rect 88518 3136 88524 3188
rect 88576 3176 88582 3188
rect 89622 3176 89628 3188
rect 88576 3148 89628 3176
rect 88576 3136 88582 3148
rect 89622 3136 89628 3148
rect 89680 3136 89686 3188
rect 93302 3136 93308 3188
rect 93360 3176 93366 3188
rect 233712 3176 233740 3216
rect 233786 3204 233792 3256
rect 233844 3244 233850 3256
rect 238754 3244 238760 3256
rect 233844 3216 238760 3244
rect 233844 3204 233850 3216
rect 238754 3204 238760 3216
rect 238812 3204 238818 3256
rect 272334 3204 272340 3256
rect 272392 3244 272398 3256
rect 414474 3244 414480 3256
rect 272392 3216 414480 3244
rect 272392 3204 272398 3216
rect 414474 3204 414480 3216
rect 414532 3204 414538 3256
rect 571061 3247 571119 3253
rect 571061 3213 571073 3247
rect 571107 3244 571119 3247
rect 575014 3244 575020 3256
rect 571107 3216 575020 3244
rect 571107 3213 571119 3216
rect 571061 3207 571119 3213
rect 575014 3204 575020 3216
rect 575072 3204 575078 3256
rect 238846 3176 238852 3188
rect 93360 3148 233372 3176
rect 233712 3148 238852 3176
rect 93360 3136 93366 3148
rect 74537 3111 74595 3117
rect 74537 3077 74549 3111
rect 74583 3108 74595 3111
rect 84013 3111 84071 3117
rect 84013 3108 84025 3111
rect 74583 3080 84025 3108
rect 74583 3077 74595 3080
rect 74537 3071 74595 3077
rect 84013 3077 84025 3080
rect 84059 3077 84071 3111
rect 84013 3071 84071 3077
rect 95694 3068 95700 3120
rect 95752 3108 95758 3120
rect 96522 3108 96528 3120
rect 95752 3080 96528 3108
rect 95752 3068 95758 3080
rect 96522 3068 96528 3080
rect 96580 3068 96586 3120
rect 102778 3068 102784 3120
rect 102836 3108 102842 3120
rect 103422 3108 103428 3120
rect 102836 3080 103428 3108
rect 102836 3068 102842 3080
rect 103422 3068 103428 3080
rect 103480 3068 103486 3120
rect 106366 3068 106372 3120
rect 106424 3108 106430 3120
rect 107470 3108 107476 3120
rect 106424 3080 107476 3108
rect 106424 3068 106430 3080
rect 107470 3068 107476 3080
rect 107528 3068 107534 3120
rect 233344 3108 233372 3148
rect 238846 3136 238852 3148
rect 238904 3136 238910 3188
rect 271966 3136 271972 3188
rect 272024 3176 272030 3188
rect 410886 3176 410892 3188
rect 272024 3148 410892 3176
rect 272024 3136 272030 3148
rect 410886 3136 410892 3148
rect 410944 3136 410950 3188
rect 239490 3108 239496 3120
rect 108316 3080 233280 3108
rect 233344 3080 239496 3108
rect 11238 3000 11244 3052
rect 11296 3040 11302 3052
rect 15838 3040 15844 3052
rect 11296 3012 15844 3040
rect 11296 3000 11302 3012
rect 15838 3000 15844 3012
rect 15896 3000 15902 3052
rect 96890 3000 96896 3052
rect 96948 3040 96954 3052
rect 108316 3040 108344 3080
rect 233252 3040 233280 3080
rect 239490 3068 239496 3080
rect 239548 3068 239554 3120
rect 272242 3068 272248 3120
rect 272300 3108 272306 3120
rect 407298 3108 407304 3120
rect 272300 3080 407304 3108
rect 272300 3068 272306 3080
rect 407298 3068 407304 3080
rect 407356 3068 407362 3120
rect 239858 3040 239864 3052
rect 96948 3012 108344 3040
rect 108408 3012 233188 3040
rect 233252 3012 239864 3040
rect 96948 3000 96954 3012
rect 93857 2975 93915 2981
rect 93857 2941 93869 2975
rect 93903 2972 93915 2975
rect 103425 2975 103483 2981
rect 103425 2972 103437 2975
rect 93903 2944 103437 2972
rect 93903 2941 93915 2944
rect 93857 2935 93915 2941
rect 103425 2941 103437 2944
rect 103471 2941 103483 2975
rect 103425 2935 103483 2941
rect 45738 2864 45744 2916
rect 45796 2904 45802 2916
rect 50338 2904 50344 2916
rect 45796 2876 50344 2904
rect 45796 2864 45802 2876
rect 50338 2864 50344 2876
rect 50396 2864 50402 2916
rect 93949 2907 94007 2913
rect 93949 2873 93961 2907
rect 93995 2904 94007 2907
rect 103333 2907 103391 2913
rect 103333 2904 103345 2907
rect 93995 2876 103345 2904
rect 93995 2873 94007 2876
rect 93949 2867 94007 2873
rect 103333 2873 103345 2876
rect 103379 2873 103391 2907
rect 103333 2867 103391 2873
rect 103974 2864 103980 2916
rect 104032 2904 104038 2916
rect 108408 2904 108436 3012
rect 113542 2932 113548 2984
rect 113600 2972 113606 2984
rect 114462 2972 114468 2984
rect 113600 2944 114468 2972
rect 113600 2932 113606 2944
rect 114462 2932 114468 2944
rect 114520 2932 114526 2984
rect 233053 2975 233111 2981
rect 233053 2972 233065 2975
rect 114572 2944 233065 2972
rect 104032 2876 108436 2904
rect 104032 2864 104038 2876
rect 111150 2864 111156 2916
rect 111208 2904 111214 2916
rect 114572 2904 114600 2944
rect 233053 2941 233065 2944
rect 233099 2941 233111 2975
rect 233160 2972 233188 3012
rect 239858 3000 239864 3012
rect 239916 3000 239922 3052
rect 271046 3000 271052 3052
rect 271104 3040 271110 3052
rect 403710 3040 403716 3052
rect 271104 3012 403716 3040
rect 271104 3000 271110 3012
rect 403710 3000 403716 3012
rect 403768 3000 403774 3052
rect 574738 3000 574744 3052
rect 574796 3040 574802 3052
rect 576210 3040 576216 3052
rect 574796 3012 576216 3040
rect 574796 3000 574802 3012
rect 576210 3000 576216 3012
rect 576268 3000 576274 3052
rect 240962 2972 240968 2984
rect 233160 2944 240968 2972
rect 233053 2935 233111 2941
rect 240962 2932 240968 2944
rect 241020 2932 241026 2984
rect 270678 2932 270684 2984
rect 270736 2972 270742 2984
rect 400214 2972 400220 2984
rect 270736 2944 400220 2972
rect 270736 2932 270742 2944
rect 400214 2932 400220 2944
rect 400272 2932 400278 2984
rect 111208 2876 114600 2904
rect 111208 2864 111214 2876
rect 114738 2864 114744 2916
rect 114796 2904 114802 2916
rect 115842 2904 115848 2916
rect 114796 2876 115848 2904
rect 114796 2864 114802 2876
rect 115842 2864 115848 2876
rect 115900 2864 115906 2916
rect 120626 2864 120632 2916
rect 120684 2904 120690 2916
rect 121362 2904 121368 2916
rect 120684 2876 121368 2904
rect 120684 2864 120690 2876
rect 121362 2864 121368 2876
rect 121420 2864 121426 2916
rect 242066 2904 242072 2916
rect 121472 2876 242072 2904
rect 118234 2796 118240 2848
rect 118292 2836 118298 2848
rect 121472 2836 121500 2876
rect 242066 2864 242072 2876
rect 242124 2864 242130 2916
rect 250346 2864 250352 2916
rect 250404 2904 250410 2916
rect 256050 2904 256056 2916
rect 250404 2876 256056 2904
rect 250404 2864 250410 2876
rect 256050 2864 256056 2876
rect 256108 2864 256114 2916
rect 270954 2864 270960 2916
rect 271012 2904 271018 2916
rect 396626 2904 396632 2916
rect 271012 2876 396632 2904
rect 271012 2864 271018 2876
rect 396626 2864 396632 2876
rect 396684 2864 396690 2916
rect 425146 2864 425152 2916
rect 425204 2904 425210 2916
rect 426342 2904 426348 2916
rect 425204 2876 426348 2904
rect 425204 2864 425210 2876
rect 426342 2864 426348 2876
rect 426400 2864 426406 2916
rect 118292 2808 121500 2836
rect 118292 2796 118298 2808
rect 121822 2796 121828 2848
rect 121880 2836 121886 2848
rect 242158 2836 242164 2848
rect 121880 2808 242164 2836
rect 121880 2796 121886 2808
rect 242158 2796 242164 2808
rect 242216 2796 242222 2848
rect 269574 2796 269580 2848
rect 269632 2836 269638 2848
rect 269632 2808 390508 2836
rect 269632 2796 269638 2808
rect 390480 2768 390508 2808
rect 390554 2796 390560 2848
rect 390612 2836 390618 2848
rect 391842 2836 391848 2848
rect 390612 2808 391848 2836
rect 390612 2796 390618 2808
rect 391842 2796 391848 2808
rect 391900 2796 391906 2848
rect 393038 2836 393044 2848
rect 391952 2808 393044 2836
rect 391952 2768 391980 2808
rect 393038 2796 393044 2808
rect 393096 2796 393102 2848
rect 390480 2740 391980 2768
rect 74258 552 74264 604
rect 74316 592 74322 604
rect 74442 592 74448 604
rect 74316 564 74448 592
rect 74316 552 74322 564
rect 74442 552 74448 564
rect 74500 552 74506 604
rect 92106 552 92112 604
rect 92164 592 92170 604
rect 92382 592 92388 604
rect 92164 564 92388 592
rect 92164 552 92170 564
rect 92382 552 92388 564
rect 92440 552 92446 604
rect 109954 552 109960 604
rect 110012 592 110018 604
rect 110322 592 110328 604
rect 110012 564 110328 592
rect 110012 552 110018 564
rect 110322 552 110328 564
rect 110380 552 110386 604
rect 183738 552 183744 604
rect 183796 592 183802 604
rect 184750 592 184756 604
rect 183796 564 184756 592
rect 183796 552 183802 564
rect 184750 552 184756 564
rect 184808 552 184814 604
rect 206278 552 206284 604
rect 206336 592 206342 604
rect 206922 592 206928 604
rect 206336 564 206928 592
rect 206336 552 206342 564
rect 206922 552 206928 564
rect 206980 552 206986 604
rect 207474 552 207480 604
rect 207532 592 207538 604
rect 208302 592 208308 604
rect 207532 564 208308 592
rect 207532 552 207538 564
rect 208302 552 208308 564
rect 208360 552 208366 604
rect 208670 552 208676 604
rect 208728 592 208734 604
rect 209682 592 209688 604
rect 208728 564 209688 592
rect 208728 552 208734 564
rect 209682 552 209688 564
rect 209740 552 209746 604
rect 230106 552 230112 604
rect 230164 592 230170 604
rect 230382 592 230388 604
rect 230164 564 230388 592
rect 230164 552 230170 564
rect 230382 552 230388 564
rect 230440 552 230446 604
rect 281534 552 281540 604
rect 281592 592 281598 604
rect 282454 592 282460 604
rect 281592 564 282460 592
rect 281592 552 281598 564
rect 282454 552 282460 564
rect 282512 552 282518 604
rect 285674 552 285680 604
rect 285732 592 285738 604
rect 285950 592 285956 604
rect 285732 564 285956 592
rect 285732 552 285738 564
rect 285950 552 285956 564
rect 286008 552 286014 604
rect 288434 552 288440 604
rect 288492 592 288498 604
rect 289538 592 289544 604
rect 288492 564 289544 592
rect 288492 552 288498 564
rect 289538 552 289544 564
rect 289596 552 289602 604
rect 292574 552 292580 604
rect 292632 592 292638 604
rect 293126 592 293132 604
rect 292632 564 293132 592
rect 292632 552 292638 564
rect 293126 552 293132 564
rect 293184 552 293190 604
rect 299474 552 299480 604
rect 299532 592 299538 604
rect 300302 592 300308 604
rect 299532 564 300308 592
rect 299532 552 299538 564
rect 300302 552 300308 564
rect 300360 552 300366 604
rect 300854 552 300860 604
rect 300912 592 300918 604
rect 301406 592 301412 604
rect 300912 564 301412 592
rect 300912 552 300918 564
rect 301406 552 301412 564
rect 301464 552 301470 604
rect 303614 552 303620 604
rect 303672 592 303678 604
rect 303798 592 303804 604
rect 303672 564 303804 592
rect 303672 552 303678 564
rect 303798 552 303804 564
rect 303856 552 303862 604
rect 492674 552 492680 604
rect 492732 592 492738 604
rect 492950 592 492956 604
rect 492732 564 492956 592
rect 492732 552 492738 564
rect 492950 552 492956 564
rect 493008 552 493014 604
rect 495434 552 495440 604
rect 495492 592 495498 604
rect 496538 592 496544 604
rect 495492 564 496544 592
rect 495492 552 495498 564
rect 496538 552 496544 564
rect 496596 552 496602 604
rect 498194 552 498200 604
rect 498252 592 498258 604
rect 498930 592 498936 604
rect 498252 564 498936 592
rect 498252 552 498258 564
rect 498930 552 498936 564
rect 498988 552 498994 604
<< via1 >>
rect 257896 700952 257948 701004
rect 397460 700952 397512 701004
rect 259368 700884 259420 700936
rect 413652 700884 413704 700936
rect 257988 700816 258040 700868
rect 429844 700816 429896 700868
rect 72976 700748 73028 700800
rect 265072 700748 265124 700800
rect 256516 700680 256568 700732
rect 462320 700680 462372 700732
rect 256608 700612 256660 700664
rect 478512 700612 478564 700664
rect 256424 700544 256476 700596
rect 494796 700544 494848 700596
rect 8116 700476 8168 700528
rect 266544 700476 266596 700528
rect 255228 700408 255280 700460
rect 527180 700408 527232 700460
rect 40500 700340 40552 700392
rect 41328 700340 41380 700392
rect 255136 700340 255188 700392
rect 543464 700340 543516 700392
rect 253848 700272 253900 700324
rect 559656 700272 559708 700324
rect 137836 700204 137888 700256
rect 263784 700204 263836 700256
rect 259276 700136 259328 700188
rect 364984 700136 365036 700188
rect 260656 700068 260708 700120
rect 348792 700068 348844 700120
rect 259184 700000 259236 700052
rect 332508 700000 332560 700052
rect 202788 699932 202840 699984
rect 262220 699932 262272 699984
rect 262128 699864 262180 699916
rect 283840 699864 283892 699916
rect 24308 699660 24360 699712
rect 24768 699660 24820 699712
rect 89168 699660 89220 699712
rect 89628 699660 89680 699712
rect 105452 699660 105504 699712
rect 106188 699660 106240 699712
rect 170312 699660 170364 699712
rect 171048 699660 171100 699712
rect 235172 699660 235224 699712
rect 235908 699660 235960 699712
rect 260748 699660 260800 699712
rect 267648 699660 267700 699712
rect 253756 696940 253808 696992
rect 580172 696940 580224 696992
rect 154120 695512 154172 695564
rect 154212 695512 154264 695564
rect 219164 695444 219216 695496
rect 154212 688576 154264 688628
rect 154396 688576 154448 688628
rect 299664 688576 299716 688628
rect 300124 688576 300176 688628
rect 219072 685899 219124 685908
rect 219072 685865 219081 685899
rect 219081 685865 219115 685899
rect 219115 685865 219124 685899
rect 219072 685856 219124 685865
rect 253664 685856 253716 685908
rect 580172 685856 580224 685908
rect 154396 685788 154448 685840
rect 299572 684428 299624 684480
rect 154304 676243 154356 676252
rect 154304 676209 154313 676243
rect 154313 676209 154347 676243
rect 154347 676209 154356 676243
rect 154304 676200 154356 676209
rect 218980 676175 219032 676184
rect 218980 676141 218989 676175
rect 218989 676141 219023 676175
rect 219023 676141 219032 676175
rect 218980 676132 219032 676141
rect 154304 673480 154356 673532
rect 154488 673480 154540 673532
rect 252468 673480 252520 673532
rect 580172 673480 580224 673532
rect 219072 666544 219124 666596
rect 299940 666544 299992 666596
rect 219164 659608 219216 659660
rect 219348 659608 219400 659660
rect 219348 656820 219400 656872
rect 154304 654100 154356 654152
rect 154488 654100 154540 654152
rect 3332 652740 3384 652792
rect 267832 652740 267884 652792
rect 252376 650020 252428 650072
rect 580172 650020 580224 650072
rect 219256 647275 219308 647284
rect 219256 647241 219265 647275
rect 219265 647241 219299 647275
rect 219299 647241 219308 647275
rect 219256 647232 219308 647241
rect 299664 647232 299716 647284
rect 299756 647232 299808 647284
rect 219256 640364 219308 640416
rect 299664 640364 299716 640416
rect 299756 640364 299808 640416
rect 219072 640228 219124 640280
rect 252284 638936 252336 638988
rect 580172 638936 580224 638988
rect 219072 637508 219124 637560
rect 219164 637508 219216 637560
rect 154304 634788 154356 634840
rect 154488 634788 154540 634840
rect 299572 630640 299624 630692
rect 299756 630640 299808 630692
rect 251088 626560 251140 626612
rect 580172 626560 580224 626612
rect 219348 626535 219400 626544
rect 219348 626501 219357 626535
rect 219357 626501 219391 626535
rect 219391 626501 219400 626535
rect 219348 626492 219400 626501
rect 219348 616879 219400 616888
rect 219348 616845 219357 616879
rect 219357 616845 219391 616879
rect 219391 616845 219400 616879
rect 219348 616836 219400 616845
rect 154304 615476 154356 615528
rect 154488 615476 154540 615528
rect 219348 611396 219400 611448
rect 299572 611328 299624 611380
rect 299756 611328 299808 611380
rect 219072 608719 219124 608728
rect 219072 608685 219081 608719
rect 219081 608685 219115 608719
rect 219115 608685 219124 608719
rect 219072 608676 219124 608685
rect 219072 608540 219124 608592
rect 299664 608583 299716 608592
rect 299664 608549 299673 608583
rect 299673 608549 299707 608583
rect 299707 608549 299716 608583
rect 299664 608540 299716 608549
rect 249708 603100 249760 603152
rect 580172 603100 580224 603152
rect 299848 601672 299900 601724
rect 219256 601579 219308 601588
rect 219256 601545 219265 601579
rect 219265 601545 219299 601579
rect 219299 601545 219308 601579
rect 219256 601536 219308 601545
rect 219256 598884 219308 598936
rect 299848 598927 299900 598936
rect 299848 598893 299857 598927
rect 299857 598893 299891 598927
rect 299891 598893 299900 598927
rect 299848 598884 299900 598893
rect 154304 596164 154356 596216
rect 154488 596164 154540 596216
rect 3056 594804 3108 594856
rect 269304 594804 269356 594856
rect 250996 592016 251048 592068
rect 580172 592016 580224 592068
rect 219164 589339 219216 589348
rect 219164 589305 219173 589339
rect 219173 589305 219207 589339
rect 219207 589305 219216 589339
rect 219164 589296 219216 589305
rect 299940 589296 299992 589348
rect 154304 589271 154356 589280
rect 154304 589237 154313 589271
rect 154313 589237 154347 589271
rect 154347 589237 154356 589271
rect 154304 589228 154356 589237
rect 218980 582360 219032 582412
rect 219164 582360 219216 582412
rect 299940 582428 299992 582480
rect 299848 582292 299900 582344
rect 154304 579751 154356 579760
rect 154304 579717 154313 579751
rect 154313 579717 154347 579751
rect 154347 579717 154356 579751
rect 154304 579708 154356 579717
rect 249616 579640 249668 579692
rect 580172 579640 580224 579692
rect 154212 579572 154264 579624
rect 154396 579572 154448 579624
rect 218980 579572 219032 579624
rect 218888 569959 218940 569968
rect 218888 569925 218897 569959
rect 218897 569925 218931 569959
rect 218931 569925 218940 569959
rect 218888 569916 218940 569925
rect 299572 563116 299624 563168
rect 218888 563048 218940 563100
rect 154212 562912 154264 562964
rect 154396 562912 154448 562964
rect 299572 562980 299624 563032
rect 218980 562912 219032 562964
rect 248328 556180 248380 556232
rect 580172 556180 580224 556232
rect 218888 553435 218940 553444
rect 218888 553401 218897 553435
rect 218897 553401 218931 553435
rect 218931 553401 218940 553435
rect 218888 553392 218940 553401
rect 299572 553460 299624 553512
rect 299480 553324 299532 553376
rect 2964 552032 3016 552084
rect 262864 552032 262916 552084
rect 218888 550647 218940 550656
rect 218888 550613 218897 550647
rect 218897 550613 218931 550647
rect 218931 550613 218940 550647
rect 218888 550604 218940 550613
rect 249524 545096 249576 545148
rect 580172 545096 580224 545148
rect 218888 543736 218940 543788
rect 299296 543668 299348 543720
rect 299480 543668 299532 543720
rect 218980 543600 219032 543652
rect 3148 538228 3200 538280
rect 270776 538228 270828 538280
rect 248236 532720 248288 532772
rect 580172 532720 580224 532772
rect 299572 531292 299624 531344
rect 299756 531292 299808 531344
rect 154396 531267 154448 531276
rect 154396 531233 154405 531267
rect 154405 531233 154439 531267
rect 154439 531233 154448 531267
rect 154396 531224 154448 531233
rect 299756 524424 299808 524476
rect 299848 524356 299900 524408
rect 218980 524288 219032 524340
rect 219164 524288 219216 524340
rect 154488 521636 154540 521688
rect 218796 514632 218848 514684
rect 219072 514632 219124 514684
rect 299664 511980 299716 512032
rect 299940 511980 299992 512032
rect 154396 511955 154448 511964
rect 154396 511921 154405 511955
rect 154405 511921 154439 511955
rect 154439 511921 154448 511955
rect 154396 511912 154448 511921
rect 219072 510595 219124 510604
rect 219072 510561 219081 510595
rect 219081 510561 219115 510595
rect 219115 510561 219124 510595
rect 219072 510552 219124 510561
rect 246948 509260 247000 509312
rect 580172 509260 580224 509312
rect 219072 505087 219124 505096
rect 219072 505053 219081 505087
rect 219081 505053 219115 505087
rect 219115 505053 219124 505087
rect 219072 505044 219124 505053
rect 154488 502324 154540 502376
rect 299756 502324 299808 502376
rect 299940 502324 299992 502376
rect 248144 498176 248196 498228
rect 580172 498176 580224 498228
rect 3332 495456 3384 495508
rect 264244 495456 264296 495508
rect 219072 492668 219124 492720
rect 219164 492668 219216 492720
rect 154212 492600 154264 492652
rect 154396 492600 154448 492652
rect 299664 492643 299716 492652
rect 299664 492609 299673 492643
rect 299673 492609 299707 492643
rect 299707 492609 299716 492643
rect 299664 492600 299716 492609
rect 219164 485800 219216 485852
rect 246856 485800 246908 485852
rect 580172 485800 580224 485852
rect 299664 485775 299716 485784
rect 299664 485741 299673 485775
rect 299673 485741 299707 485775
rect 299707 485741 299716 485775
rect 299664 485732 299716 485741
rect 219256 485664 219308 485716
rect 3148 480224 3200 480276
rect 272524 480224 272576 480276
rect 299572 476076 299624 476128
rect 299756 476076 299808 476128
rect 299664 473331 299716 473340
rect 299664 473297 299673 473331
rect 299673 473297 299707 473331
rect 299707 473297 299716 473331
rect 299664 473288 299716 473297
rect 154304 466420 154356 466472
rect 154488 466420 154540 466472
rect 218980 466420 219032 466472
rect 299664 466395 299716 466404
rect 299664 466361 299673 466395
rect 299673 466361 299707 466395
rect 299707 466361 299716 466395
rect 299664 466352 299716 466361
rect 219348 466284 219400 466336
rect 245568 462340 245620 462392
rect 580172 462340 580224 462392
rect 299388 460844 299440 460896
rect 299756 460844 299808 460896
rect 154304 453976 154356 454028
rect 219072 453976 219124 454028
rect 245476 451256 245528 451308
rect 580172 451256 580224 451308
rect 299480 449871 299532 449880
rect 299480 449837 299489 449871
rect 299489 449837 299523 449871
rect 299523 449837 299532 449871
rect 299480 449828 299532 449837
rect 154212 444431 154264 444440
rect 154212 444397 154221 444431
rect 154221 444397 154255 444431
rect 154255 444397 154264 444431
rect 154212 444388 154264 444397
rect 218980 444431 219032 444440
rect 218980 444397 218989 444431
rect 218989 444397 219023 444431
rect 219023 444397 219032 444431
rect 218980 444388 219032 444397
rect 299572 440240 299624 440292
rect 245384 438880 245436 438932
rect 580172 438880 580224 438932
rect 2964 437452 3016 437504
rect 265624 437452 265676 437504
rect 299572 436815 299624 436824
rect 299572 436781 299581 436815
rect 299581 436781 299615 436815
rect 299615 436781 299624 436815
rect 299572 436772 299624 436781
rect 218980 434664 219032 434716
rect 219072 434664 219124 434716
rect 154304 427796 154356 427848
rect 154396 427728 154448 427780
rect 299572 427771 299624 427780
rect 299572 427737 299581 427771
rect 299581 427737 299615 427771
rect 299615 427737 299624 427771
rect 299572 427728 299624 427737
rect 154120 425008 154172 425060
rect 154396 425008 154448 425060
rect 3332 423648 3384 423700
rect 273904 423648 273956 423700
rect 244188 415420 244240 415472
rect 580172 415420 580224 415472
rect 299756 415352 299808 415404
rect 154488 408484 154540 408536
rect 154488 408348 154540 408400
rect 299664 405739 299716 405748
rect 299664 405705 299673 405739
rect 299673 405705 299707 405739
rect 299707 405705 299716 405739
rect 299664 405696 299716 405705
rect 243820 404336 243872 404388
rect 580172 404336 580224 404388
rect 106188 403112 106240 403164
rect 264888 402976 264940 403028
rect 264244 402908 264296 402960
rect 273812 402908 273864 402960
rect 273904 402908 273956 402960
rect 274916 402908 274968 402960
rect 89628 402840 89680 402892
rect 41328 402772 41380 402824
rect 255412 402840 255464 402892
rect 256424 402840 256476 402892
rect 256976 402840 257028 402892
rect 257988 402840 258040 402892
rect 258540 402840 258592 402892
rect 259276 402840 259328 402892
rect 259644 402840 259696 402892
rect 260656 402840 260708 402892
rect 261208 402840 261260 402892
rect 262128 402840 262180 402892
rect 265624 402840 265676 402892
rect 275376 402840 275428 402892
rect 265900 402772 265952 402824
rect 24768 402704 24820 402756
rect 254400 402704 254452 402756
rect 255228 402704 255280 402756
rect 262772 402704 262824 402756
rect 3424 402636 3476 402688
rect 268016 402636 268068 402688
rect 3608 402568 3660 402620
rect 266452 402568 266504 402620
rect 3516 402500 3568 402552
rect 269120 402500 269172 402552
rect 3884 402432 3936 402484
rect 271236 402432 271288 402484
rect 3700 402364 3752 402416
rect 270684 402364 270736 402416
rect 4068 402296 4120 402348
rect 272800 402296 272852 402348
rect 3240 402228 3292 402280
rect 274364 402228 274416 402280
rect 154488 402160 154540 402212
rect 258080 402160 258132 402212
rect 259368 402160 259420 402212
rect 171048 402092 171100 402144
rect 269580 402160 269632 402212
rect 219348 402024 219400 402076
rect 242256 401956 242308 402008
rect 244924 401956 244976 402008
rect 245568 401956 245620 402008
rect 247040 401956 247092 402008
rect 248144 401956 248196 402008
rect 248604 401956 248656 402008
rect 249524 401956 249576 402008
rect 250168 401956 250220 402008
rect 250996 401956 251048 402008
rect 251180 401956 251232 402008
rect 252376 401956 252428 402008
rect 252744 401956 252796 402008
rect 253756 401956 253808 402008
rect 261760 402092 261812 402144
rect 262864 402092 262916 402144
rect 272248 402092 272300 402144
rect 267556 402024 267608 402076
rect 277032 402024 277084 402076
rect 235908 401888 235960 401940
rect 260196 401956 260248 402008
rect 299664 401956 299716 402008
rect 264336 401888 264388 401940
rect 264980 401888 265032 401940
rect 272524 401888 272576 401940
rect 273260 401888 273312 401940
rect 243268 401820 243320 401872
rect 244188 401820 244240 401872
rect 244372 401820 244424 401872
rect 245384 401820 245436 401872
rect 245936 401820 245988 401872
rect 246856 401820 246908 401872
rect 247500 401820 247552 401872
rect 248236 401820 248288 401872
rect 489184 401820 489236 401872
rect 3332 401752 3384 401804
rect 278596 401752 278648 401804
rect 3976 401684 4028 401736
rect 280160 401684 280212 401736
rect 3792 401616 3844 401668
rect 281724 401616 281776 401668
rect 262956 401548 263008 401600
rect 10968 401412 11020 401464
rect 275928 401412 275980 401464
rect 14556 401344 14608 401396
rect 277492 401344 277544 401396
rect 227168 401276 227220 401328
rect 279056 401276 279108 401328
rect 225788 401208 225840 401260
rect 280712 401208 280764 401260
rect 227076 401140 227128 401192
rect 284392 401140 284444 401192
rect 233332 401072 233384 401124
rect 291936 401072 291988 401124
rect 222844 401004 222896 401056
rect 283840 401004 283892 401056
rect 225604 400936 225656 400988
rect 287520 400936 287572 400988
rect 234896 400868 234948 400920
rect 297456 400868 297508 400920
rect 231768 400800 231820 400852
rect 294604 400800 294656 400852
rect 238024 400732 238076 400784
rect 301596 400732 301648 400784
rect 211804 400664 211856 400716
rect 279608 400664 279660 400716
rect 215944 400596 215996 400648
rect 286968 400596 287020 400648
rect 209044 400528 209096 400580
rect 281172 400528 281224 400580
rect 235448 400460 235500 400512
rect 308404 400460 308456 400512
rect 230664 400392 230716 400444
rect 304264 400392 304316 400444
rect 233884 400324 233936 400376
rect 496084 400324 496136 400376
rect 241704 400256 241756 400308
rect 290556 400256 290608 400308
rect 241244 400188 241296 400240
rect 290464 400188 290516 400240
rect 238576 400120 238628 400172
rect 226984 400052 227036 400104
rect 276480 400052 276532 400104
rect 242624 399984 242676 400036
rect 290648 399984 290700 400036
rect 236736 399916 236788 399968
rect 298836 399916 298888 399968
rect 239864 399848 239916 399900
rect 302976 399848 303028 399900
rect 213184 399780 213236 399832
rect 277676 399780 277728 399832
rect 218704 399712 218756 399764
rect 285036 399712 285088 399764
rect 232504 399644 232556 399696
rect 305644 399644 305696 399696
rect 214564 399576 214616 399628
rect 288348 399576 288400 399628
rect 207664 399508 207716 399560
rect 282460 399508 282512 399560
rect 285588 399508 285640 399560
rect 3424 399440 3476 399492
rect 264980 399440 265032 399492
rect 204904 399372 204956 399424
rect 180064 399304 180116 399356
rect 281908 399304 281960 399356
rect 288716 399304 288768 399356
rect 13084 399168 13136 399220
rect 393964 398148 394016 398200
rect 3148 395972 3200 396024
rect 10968 395972 11020 396024
rect 290648 393252 290700 393304
rect 579804 393252 579856 393304
rect 290556 369792 290608 369844
rect 580172 369792 580224 369844
rect 2964 367004 3016 367056
rect 226984 367004 227036 367056
rect 489184 358708 489236 358760
rect 580080 358708 580132 358760
rect 290464 346332 290516 346384
rect 579804 346332 579856 346384
rect 277860 338104 277912 338156
rect 278136 338104 278188 338156
rect 3424 338036 3476 338088
rect 14556 338036 14608 338088
rect 125508 338036 125560 338088
rect 240232 338036 240284 338088
rect 240876 338036 240928 338088
rect 243084 338079 243136 338088
rect 243084 338045 243093 338079
rect 243093 338045 243127 338079
rect 243127 338045 243136 338079
rect 243084 338036 243136 338045
rect 267556 338036 267608 338088
rect 274916 338036 274968 338088
rect 278780 338036 278832 338088
rect 279700 338036 279752 338088
rect 290004 338036 290056 338088
rect 107568 337968 107620 338020
rect 115848 337900 115900 337952
rect 241704 337968 241756 338020
rect 277492 337968 277544 338020
rect 278504 337968 278556 338020
rect 284852 337968 284904 338020
rect 294696 337968 294748 338020
rect 253204 337900 253256 337952
rect 254216 337900 254268 337952
rect 263600 337900 263652 337952
rect 267740 337900 267792 337952
rect 271972 337900 272024 337952
rect 100668 337832 100720 337884
rect 245108 337832 245160 337884
rect 257160 337832 257212 337884
rect 263416 337832 263468 337884
rect 39304 337764 39356 337816
rect 233608 337764 233660 337816
rect 242808 337764 242860 337816
rect 262404 337764 262456 337816
rect 265532 337764 265584 337816
rect 266360 337764 266412 337816
rect 267004 337764 267056 337816
rect 267924 337807 267976 337816
rect 267924 337773 267933 337807
rect 267933 337773 267967 337807
rect 267967 337773 267976 337807
rect 267924 337764 267976 337773
rect 273904 337764 273956 337816
rect 274548 337764 274600 337816
rect 32404 337696 32456 337748
rect 231952 337696 232004 337748
rect 240968 337696 241020 337748
rect 246948 337696 247000 337748
rect 257528 337696 257580 337748
rect 262220 337696 262272 337748
rect 262312 337696 262364 337748
rect 279240 337900 279292 337952
rect 283564 337900 283616 337952
rect 285956 337900 286008 337952
rect 297364 337900 297416 337952
rect 282644 337832 282696 337884
rect 298744 337832 298796 337884
rect 276020 337764 276072 337816
rect 283012 337764 283064 337816
rect 301504 337764 301556 337816
rect 279608 337696 279660 337748
rect 35164 337628 35216 337680
rect 232872 337628 232924 337680
rect 246580 337628 246632 337680
rect 257252 337628 257304 337680
rect 275192 337628 275244 337680
rect 302884 337696 302936 337748
rect 283564 337628 283616 337680
rect 286324 337628 286376 337680
rect 286600 337628 286652 337680
rect 287428 337628 287480 337680
rect 290832 337628 290884 337680
rect 320824 337628 320876 337680
rect 28264 337560 28316 337612
rect 232044 337560 232096 337612
rect 258264 337560 258316 337612
rect 277492 337560 277544 337612
rect 278688 337560 278740 337612
rect 281172 337560 281224 337612
rect 15844 337492 15896 337544
rect 231032 337492 231084 337544
rect 241152 337492 241204 337544
rect 242992 337492 243044 337544
rect 260932 337492 260984 337544
rect 271144 337492 271196 337544
rect 280712 337492 280764 337544
rect 316684 337560 316736 337612
rect 319444 337492 319496 337544
rect 14464 337424 14516 337476
rect 230940 337424 230992 337476
rect 242900 337424 242952 337476
rect 253296 337424 253348 337476
rect 259644 337424 259696 337476
rect 265624 337424 265676 337476
rect 346400 337424 346452 337476
rect 10324 337356 10376 337408
rect 230480 337356 230532 337408
rect 245568 337356 245620 337408
rect 251272 337356 251324 337408
rect 260196 337356 260248 337408
rect 260564 337288 260616 337340
rect 225696 337220 225748 337272
rect 257436 337220 257488 337272
rect 261484 337220 261536 337272
rect 261668 337220 261720 337272
rect 228364 337152 228416 337204
rect 231952 337084 232004 337136
rect 234896 337084 234948 337136
rect 251272 337152 251324 337204
rect 254860 337152 254912 337204
rect 260472 337152 260524 337204
rect 262128 337152 262180 337204
rect 246764 337084 246816 337136
rect 256700 337084 256752 337136
rect 258448 337084 258500 337136
rect 258632 337084 258684 337136
rect 260932 337084 260984 337136
rect 261300 337084 261352 337136
rect 261668 337084 261720 337136
rect 247684 337016 247736 337068
rect 255044 337016 255096 337068
rect 256884 337016 256936 337068
rect 258080 337016 258132 337068
rect 260104 337016 260156 337068
rect 260564 337016 260616 337068
rect 260840 337016 260892 337068
rect 261852 337016 261904 337068
rect 230388 336948 230440 337000
rect 236828 336948 236880 337000
rect 248512 336948 248564 337000
rect 251364 336948 251416 337000
rect 253572 336948 253624 337000
rect 257068 336948 257120 337000
rect 257804 336948 257856 337000
rect 258356 336948 258408 337000
rect 259184 336948 259236 337000
rect 261024 336948 261076 337000
rect 261944 336948 261996 337000
rect 233240 336880 233292 336932
rect 234436 336880 234488 336932
rect 249616 336880 249668 336932
rect 252836 336880 252888 336932
rect 257160 336880 257212 336932
rect 257896 336880 257948 336932
rect 258264 336880 258316 336932
rect 259276 336880 259328 336932
rect 259828 336880 259880 336932
rect 260656 336880 260708 336932
rect 261208 336880 261260 336932
rect 262036 336880 262088 336932
rect 252284 336812 252336 336864
rect 253756 336812 253808 336864
rect 254860 336812 254912 336864
rect 255780 336812 255832 336864
rect 257068 336812 257120 336864
rect 257620 336812 257672 336864
rect 258356 336812 258408 336864
rect 259092 336812 259144 336864
rect 260840 336812 260892 336864
rect 261576 336812 261628 336864
rect 261944 336812 261996 336864
rect 262772 337016 262824 337068
rect 262956 337016 263008 337068
rect 262404 336948 262456 337000
rect 263048 336948 263100 337000
rect 277768 337356 277820 337408
rect 278320 337356 278372 337408
rect 281908 337356 281960 337408
rect 489184 337356 489236 337408
rect 263968 337288 264020 337340
rect 271328 337288 271380 337340
rect 273444 337288 273496 337340
rect 274548 337288 274600 337340
rect 277860 337288 277912 337340
rect 278596 337288 278648 337340
rect 265256 337220 265308 337272
rect 271236 337220 271288 337272
rect 278780 337220 278832 337272
rect 280068 337220 280120 337272
rect 282276 337220 282328 337272
rect 289912 337288 289964 337340
rect 283012 337220 283064 337272
rect 284208 337220 284260 337272
rect 284300 337220 284352 337272
rect 262772 336880 262824 336932
rect 263508 336880 263560 336932
rect 272524 337152 272576 337204
rect 273076 337152 273128 337204
rect 282552 337152 282604 337204
rect 282828 337152 282880 337204
rect 282920 337152 282972 337204
rect 283472 337152 283524 337204
rect 286048 337152 286100 337204
rect 286968 337152 287020 337204
rect 287428 337152 287480 337204
rect 288348 337152 288400 337204
rect 264980 337084 265032 337136
rect 265900 337084 265952 337136
rect 270500 337084 270552 337136
rect 274824 337127 274876 337136
rect 274824 337093 274833 337127
rect 274833 337093 274867 337127
rect 274867 337093 274876 337127
rect 274824 337084 274876 337093
rect 279240 337084 279292 337136
rect 279884 337084 279936 337136
rect 280804 337084 280856 337136
rect 291844 337084 291896 337136
rect 265164 337016 265216 337068
rect 265992 337016 266044 337068
rect 266728 337016 266780 337068
rect 262680 336812 262732 336864
rect 263140 336812 263192 336864
rect 264980 336948 265032 337000
rect 265256 336948 265308 337000
rect 266084 336948 266136 337000
rect 266360 336948 266412 337000
rect 267648 336948 267700 337000
rect 265440 336880 265492 336932
rect 266268 336880 266320 336932
rect 266728 336880 266780 336932
rect 267188 336880 267240 336932
rect 272340 337016 272392 337068
rect 273076 337016 273128 337068
rect 273352 337016 273404 337068
rect 274364 337016 274416 337068
rect 274732 337016 274784 337068
rect 275652 337016 275704 337068
rect 278136 337016 278188 337068
rect 278228 337016 278280 337068
rect 278780 337016 278832 337068
rect 279148 337016 279200 337068
rect 280068 337016 280120 337068
rect 280436 337016 280488 337068
rect 283472 337016 283524 337068
rect 283748 337016 283800 337068
rect 284024 337016 284076 337068
rect 267924 336948 267976 337000
rect 268660 336948 268712 337000
rect 273444 336948 273496 337000
rect 274456 336948 274508 337000
rect 276112 336948 276164 337000
rect 277032 336948 277084 337000
rect 278596 336948 278648 337000
rect 279056 336948 279108 337000
rect 279700 336948 279752 337000
rect 280344 336948 280396 337000
rect 280896 336948 280948 337000
rect 281540 336948 281592 337000
rect 283196 336948 283248 337000
rect 284116 336948 284168 337000
rect 268292 336880 268344 336932
rect 268844 336880 268896 336932
rect 270592 336880 270644 336932
rect 271236 336880 271288 336932
rect 272340 336880 272392 336932
rect 272708 336880 272760 336932
rect 273260 336880 273312 336932
rect 274088 336880 274140 336932
rect 274824 336880 274876 336932
rect 275376 336880 275428 336932
rect 276940 336880 276992 336932
rect 279332 336880 279384 336932
rect 279884 336880 279936 336932
rect 280620 336880 280672 336932
rect 281172 336880 281224 336932
rect 263968 336812 264020 336864
rect 264888 336812 264940 336864
rect 265624 336812 265676 336864
rect 266176 336812 266228 336864
rect 266912 336812 266964 336864
rect 267372 336812 267424 336864
rect 267648 336812 267700 336864
rect 271880 336812 271932 336864
rect 272156 336812 272208 336864
rect 273352 336812 273404 336864
rect 273812 336812 273864 336864
rect 274916 336812 274968 336864
rect 275468 336812 275520 336864
rect 276020 336812 276072 336864
rect 276480 336812 276532 336864
rect 233240 336744 233292 336796
rect 235264 336744 235316 336796
rect 240232 336744 240284 336796
rect 241612 336744 241664 336796
rect 245292 336744 245344 336796
rect 245844 336744 245896 336796
rect 247040 336744 247092 336796
rect 248420 336744 248472 336796
rect 251916 336744 251968 336796
rect 253480 336744 253532 336796
rect 254768 336744 254820 336796
rect 255412 336744 255464 336796
rect 256516 336744 256568 336796
rect 257344 336744 257396 336796
rect 257528 336744 257580 336796
rect 257988 336744 258040 336796
rect 258540 336744 258592 336796
rect 258908 336744 258960 336796
rect 260012 336744 260064 336796
rect 260472 336744 260524 336796
rect 260656 336787 260708 336796
rect 260656 336753 260665 336787
rect 260665 336753 260699 336787
rect 260699 336753 260708 336787
rect 260656 336744 260708 336753
rect 260932 336744 260984 336796
rect 261300 336744 261352 336796
rect 261760 336744 261812 336796
rect 262220 336744 262272 336796
rect 261576 336676 261628 336728
rect 261208 336651 261260 336660
rect 261208 336617 261217 336651
rect 261217 336617 261251 336651
rect 261251 336617 261260 336651
rect 261208 336608 261260 336617
rect 262496 336744 262548 336796
rect 262864 336744 262916 336796
rect 263784 336744 263836 336796
rect 264152 336744 264204 336796
rect 264336 336744 264388 336796
rect 264612 336744 264664 336796
rect 265716 336744 265768 336796
rect 265900 336744 265952 336796
rect 266084 336787 266136 336796
rect 266084 336753 266093 336787
rect 266093 336753 266127 336787
rect 266127 336753 266136 336787
rect 266084 336744 266136 336753
rect 266636 336744 266688 336796
rect 267096 336744 267148 336796
rect 267188 336744 267240 336796
rect 267464 336744 267516 336796
rect 268292 336744 268344 336796
rect 268568 336744 268620 336796
rect 268660 336744 268712 336796
rect 268936 336744 268988 336796
rect 269488 336744 269540 336796
rect 269764 336744 269816 336796
rect 270040 336744 270092 336796
rect 270224 336744 270276 336796
rect 270684 336787 270736 336796
rect 270684 336753 270693 336787
rect 270693 336753 270727 336787
rect 270727 336753 270736 336787
rect 270684 336744 270736 336753
rect 271052 336744 271104 336796
rect 271512 336744 271564 336796
rect 271972 336744 272024 336796
rect 272248 336744 272300 336796
rect 272432 336744 272484 336796
rect 272708 336744 272760 336796
rect 272892 336744 272944 336796
rect 273168 336744 273220 336796
rect 273628 336744 273680 336796
rect 274180 336744 274232 336796
rect 275008 336744 275060 336796
rect 275376 336744 275428 336796
rect 276388 336744 276440 336796
rect 276664 336744 276716 336796
rect 276112 336676 276164 336728
rect 277308 336812 277360 336864
rect 276940 336744 276992 336796
rect 277216 336744 277268 336796
rect 277584 336744 277636 336796
rect 277768 336744 277820 336796
rect 277952 336744 278004 336796
rect 278228 336744 278280 336796
rect 278504 336744 278556 336796
rect 262864 336608 262916 336660
rect 279516 336744 279568 336796
rect 279976 336744 280028 336796
rect 280160 336744 280212 336796
rect 280436 336744 280488 336796
rect 280528 336744 280580 336796
rect 280804 336787 280856 336796
rect 280804 336753 280813 336787
rect 280813 336753 280847 336787
rect 280847 336753 280856 336787
rect 280804 336744 280856 336753
rect 280988 336744 281040 336796
rect 281448 336744 281500 336796
rect 281632 336744 281684 336796
rect 280896 336676 280948 336728
rect 282092 336744 282144 336796
rect 282644 336744 282696 336796
rect 290464 337016 290516 337068
rect 284484 336948 284536 337000
rect 285496 336948 285548 337000
rect 286232 336948 286284 337000
rect 286876 336948 286928 337000
rect 288532 336948 288584 337000
rect 290740 336948 290792 337000
rect 285680 336880 285732 336932
rect 286324 336880 286376 336932
rect 288624 336880 288676 336932
rect 290556 336880 290608 336932
rect 285956 336812 286008 336864
rect 286416 336812 286468 336864
rect 287520 336812 287572 336864
rect 288072 336812 288124 336864
rect 288900 336812 288952 336864
rect 290648 336812 290700 336864
rect 284300 336744 284352 336796
rect 284576 336744 284628 336796
rect 286048 336744 286100 336796
rect 286508 336744 286560 336796
rect 286692 336744 286744 336796
rect 286876 336744 286928 336796
rect 287704 336744 287756 336796
rect 287980 336744 288032 336796
rect 289084 336744 289136 336796
rect 289452 336744 289504 336796
rect 289820 336744 289872 336796
rect 291108 336744 291160 336796
rect 282828 336676 282880 336728
rect 283288 336676 283340 336728
rect 280160 336608 280212 336660
rect 280712 336608 280764 336660
rect 293960 336608 294012 336660
rect 239036 336540 239088 336592
rect 279608 336540 279660 336592
rect 296720 336540 296772 336592
rect 227628 336472 227680 336524
rect 242900 336472 242952 336524
rect 261668 336472 261720 336524
rect 305000 336472 305052 336524
rect 220728 336404 220780 336456
rect 252652 336404 252704 336456
rect 265532 336404 265584 336456
rect 314660 336404 314712 336456
rect 216588 336336 216640 336388
rect 252100 336336 252152 336388
rect 267740 336336 267792 336388
rect 327080 336336 327132 336388
rect 209688 336268 209740 336320
rect 248512 336268 248564 336320
rect 265348 336268 265400 336320
rect 265532 336268 265584 336320
rect 267004 336268 267056 336320
rect 353300 336268 353352 336320
rect 162768 336200 162820 336252
rect 275284 336200 275336 336252
rect 440240 336200 440292 336252
rect 176568 336132 176620 336184
rect 248052 336132 248104 336184
rect 290004 336132 290056 336184
rect 483020 336132 483072 336184
rect 153200 336064 153252 336116
rect 153292 336064 153344 336116
rect 211252 336064 211304 336116
rect 211344 336064 211396 336116
rect 236276 336064 236328 336116
rect 236552 336064 236604 336116
rect 248696 336107 248748 336116
rect 248696 336073 248705 336107
rect 248705 336073 248739 336107
rect 248739 336073 248748 336107
rect 248696 336064 248748 336073
rect 284024 336064 284076 336116
rect 521660 336064 521712 336116
rect 52368 335996 52420 336048
rect 89628 335996 89680 336048
rect 153108 335996 153160 336048
rect 232044 335996 232096 336048
rect 232688 335996 232740 336048
rect 287060 335996 287112 336048
rect 554780 335996 554832 336048
rect 153108 335860 153160 335912
rect 232228 335928 232280 335980
rect 232780 335928 232832 335980
rect 233240 335860 233292 335912
rect 244648 335860 244700 335912
rect 245108 335860 245160 335912
rect 251364 335860 251416 335912
rect 251732 335860 251784 335912
rect 233516 335792 233568 335844
rect 233700 335792 233752 335844
rect 240508 335792 240560 335844
rect 241428 335792 241480 335844
rect 244280 335792 244332 335844
rect 244740 335792 244792 335844
rect 246212 335835 246264 335844
rect 246212 335801 246221 335835
rect 246221 335801 246255 335835
rect 246255 335801 246264 335835
rect 246212 335792 246264 335801
rect 248512 335792 248564 335844
rect 249524 335792 249576 335844
rect 236460 335724 236512 335776
rect 236736 335724 236788 335776
rect 237748 335724 237800 335776
rect 238484 335724 238536 335776
rect 245568 335767 245620 335776
rect 245568 335733 245577 335767
rect 245577 335733 245611 335767
rect 245611 335733 245620 335767
rect 245568 335724 245620 335733
rect 250352 335724 250404 335776
rect 251088 335724 251140 335776
rect 251456 335724 251508 335776
rect 252192 335724 252244 335776
rect 284944 335724 284996 335776
rect 230204 335656 230256 335708
rect 236368 335656 236420 335708
rect 236644 335656 236696 335708
rect 240324 335656 240376 335708
rect 241060 335656 241112 335708
rect 244464 335656 244516 335708
rect 245752 335656 245804 335708
rect 246028 335656 246080 335708
rect 246672 335656 246724 335708
rect 248420 335656 248472 335708
rect 248788 335656 248840 335708
rect 248972 335656 249024 335708
rect 249340 335656 249392 335708
rect 250168 335656 250220 335708
rect 250720 335656 250772 335708
rect 251548 335699 251600 335708
rect 251548 335665 251557 335699
rect 251557 335665 251591 335699
rect 251591 335665 251600 335699
rect 251548 335656 251600 335665
rect 251640 335656 251692 335708
rect 252100 335656 252152 335708
rect 252284 335656 252336 335708
rect 254032 335656 254084 335708
rect 254400 335656 254452 335708
rect 269304 335656 269356 335708
rect 269856 335656 269908 335708
rect 287612 335699 287664 335708
rect 287612 335665 287621 335699
rect 287621 335665 287655 335699
rect 287655 335665 287664 335699
rect 287612 335656 287664 335665
rect 229376 335588 229428 335640
rect 230664 335588 230716 335640
rect 231400 335588 231452 335640
rect 236092 335588 236144 335640
rect 236828 335588 236880 335640
rect 237748 335588 237800 335640
rect 238116 335588 238168 335640
rect 238852 335588 238904 335640
rect 239772 335588 239824 335640
rect 240692 335588 240744 335640
rect 240968 335588 241020 335640
rect 241520 335588 241572 335640
rect 241888 335588 241940 335640
rect 242164 335588 242216 335640
rect 242440 335588 242492 335640
rect 242532 335588 242584 335640
rect 242716 335588 242768 335640
rect 240416 335520 240468 335572
rect 240784 335520 240836 335572
rect 233332 335452 233384 335504
rect 234160 335452 234212 335504
rect 236000 335452 236052 335504
rect 236460 335452 236512 335504
rect 244648 335588 244700 335640
rect 244924 335588 244976 335640
rect 245016 335588 245068 335640
rect 245568 335588 245620 335640
rect 247408 335588 247460 335640
rect 247592 335588 247644 335640
rect 249248 335588 249300 335640
rect 249616 335588 249668 335640
rect 245936 335452 245988 335504
rect 246212 335452 246264 335504
rect 246396 335452 246448 335504
rect 249800 335452 249852 335504
rect 250076 335452 250128 335504
rect 251916 335452 251968 335504
rect 252928 335588 252980 335640
rect 253848 335588 253900 335640
rect 255504 335588 255556 335640
rect 256240 335588 256292 335640
rect 254124 335520 254176 335572
rect 244280 335316 244332 335368
rect 244372 335316 244424 335368
rect 245200 335316 245252 335368
rect 248880 335316 248932 335368
rect 249708 335316 249760 335368
rect 249800 335316 249852 335368
rect 250444 335316 250496 335368
rect 251732 335359 251784 335368
rect 251732 335325 251741 335359
rect 251741 335325 251775 335359
rect 251775 335325 251784 335359
rect 251732 335316 251784 335325
rect 249892 335248 249944 335300
rect 250628 335248 250680 335300
rect 254308 335316 254360 335368
rect 254676 335316 254728 335368
rect 254492 335180 254544 335232
rect 256056 335520 256108 335572
rect 277676 335520 277728 335572
rect 256792 335452 256844 335504
rect 257804 335452 257856 335504
rect 269580 335452 269632 335504
rect 269948 335452 270000 335504
rect 272156 335452 272208 335504
rect 272524 335452 272576 335504
rect 269396 335384 269448 335436
rect 270132 335384 270184 335436
rect 279516 335452 279568 335504
rect 279792 335452 279844 335504
rect 255688 335316 255740 335368
rect 256056 335316 256108 335368
rect 269580 335316 269632 335368
rect 270316 335316 270368 335368
rect 277676 335316 277728 335368
rect 280160 335316 280212 335368
rect 280528 335316 280580 335368
rect 256424 335291 256476 335300
rect 256424 335257 256433 335291
rect 256433 335257 256467 335291
rect 256467 335257 256476 335291
rect 256424 335248 256476 335257
rect 280436 335291 280488 335300
rect 280436 335257 280445 335291
rect 280445 335257 280479 335291
rect 280479 335257 280488 335291
rect 280436 335248 280488 335257
rect 255688 335180 255740 335232
rect 278872 335180 278924 335232
rect 279332 335180 279384 335232
rect 280160 335223 280212 335232
rect 280160 335189 280169 335223
rect 280169 335189 280203 335223
rect 280203 335189 280212 335223
rect 280160 335180 280212 335189
rect 229008 335112 229060 335164
rect 253388 335112 253440 335164
rect 278964 335155 279016 335164
rect 278964 335121 278973 335155
rect 278973 335121 279007 335155
rect 279007 335121 279016 335155
rect 278964 335112 279016 335121
rect 223488 335044 223540 335096
rect 249524 335044 249576 335096
rect 281632 335044 281684 335096
rect 282552 335044 282604 335096
rect 300860 335044 300912 335096
rect 208308 334976 208360 335028
rect 262128 334976 262180 335028
rect 311900 334976 311952 335028
rect 212448 334908 212500 334960
rect 251364 334908 251416 334960
rect 262312 334908 262364 334960
rect 316040 334908 316092 334960
rect 169668 334840 169720 334892
rect 247316 334840 247368 334892
rect 264428 334840 264480 334892
rect 333980 334840 334032 334892
rect 160008 334772 160060 334824
rect 259920 334772 259972 334824
rect 260196 334772 260248 334824
rect 274548 334772 274600 334824
rect 422300 334772 422352 334824
rect 126888 334704 126940 334756
rect 241152 334704 241204 334756
rect 289912 334704 289964 334756
rect 500960 334704 501012 334756
rect 117228 334636 117280 334688
rect 241980 334636 242032 334688
rect 285496 334636 285548 334688
rect 528560 334636 528612 334688
rect 56508 334568 56560 334620
rect 235632 334568 235684 334620
rect 289268 334568 289320 334620
rect 574744 334568 574796 334620
rect 276204 334500 276256 334552
rect 277124 334500 277176 334552
rect 230296 334160 230348 334212
rect 231676 333888 231728 333940
rect 232136 334024 232188 334076
rect 259460 334024 259512 334076
rect 260380 334024 260432 334076
rect 232044 333820 232096 333872
rect 231676 333752 231728 333804
rect 239220 333752 239272 333804
rect 239588 333752 239640 333804
rect 233608 333684 233660 333736
rect 233884 333684 233936 333736
rect 236276 333684 236328 333736
rect 236920 333684 236972 333736
rect 260564 333684 260616 333736
rect 292580 333684 292632 333736
rect 219348 333616 219400 333668
rect 252376 333616 252428 333668
rect 261484 333616 261536 333668
rect 307760 333616 307812 333668
rect 184848 333548 184900 333600
rect 248420 333548 248472 333600
rect 262956 333548 263008 333600
rect 318800 333548 318852 333600
rect 173808 333480 173860 333532
rect 247776 333480 247828 333532
rect 261208 333480 261260 333532
rect 261484 333480 261536 333532
rect 266084 333480 266136 333532
rect 342260 333480 342312 333532
rect 155868 333412 155920 333464
rect 245292 333412 245344 333464
rect 271604 333412 271656 333464
rect 404360 333412 404412 333464
rect 129648 333344 129700 333396
rect 243176 333344 243228 333396
rect 278596 333344 278648 333396
rect 465080 333344 465132 333396
rect 114468 333276 114520 333328
rect 240232 333276 240284 333328
rect 241060 333276 241112 333328
rect 241336 333276 241388 333328
rect 262864 333276 262916 333328
rect 263416 333276 263468 333328
rect 283380 333276 283432 333328
rect 518900 333276 518952 333328
rect 49608 333208 49660 333260
rect 234988 333208 235040 333260
rect 238944 333208 238996 333260
rect 239128 333208 239180 333260
rect 284024 333208 284076 333260
rect 284944 333208 284996 333260
rect 286600 333208 286652 333260
rect 546500 333208 546552 333260
rect 231584 333140 231636 333192
rect 231768 333140 231820 333192
rect 232228 333140 232280 333192
rect 233056 333140 233108 333192
rect 233884 333140 233936 333192
rect 237564 333140 237616 333192
rect 278044 333140 278096 333192
rect 287428 333140 287480 333192
rect 288164 333140 288216 333192
rect 234620 333072 234672 333124
rect 234988 333072 235040 333124
rect 277952 333072 278004 333124
rect 278044 333004 278096 333056
rect 278412 333004 278464 333056
rect 235172 332936 235224 332988
rect 235448 332936 235500 332988
rect 285864 332868 285916 332920
rect 286784 332868 286836 332920
rect 234068 332392 234120 332444
rect 234344 332392 234396 332444
rect 278780 332392 278832 332444
rect 260656 332324 260708 332376
rect 296812 332324 296864 332376
rect 230388 332256 230440 332308
rect 251732 332256 251784 332308
rect 261944 332256 261996 332308
rect 313280 332256 313332 332308
rect 224868 332188 224920 332240
rect 253020 332188 253072 332240
rect 271328 332188 271380 332240
rect 331220 332188 331272 332240
rect 180708 332120 180760 332172
rect 247040 332120 247092 332172
rect 267648 332120 267700 332172
rect 356060 332120 356112 332172
rect 142068 332052 142120 332104
rect 244280 332052 244332 332104
rect 397460 332052 397512 332104
rect 139308 331984 139360 332036
rect 48228 331916 48280 331968
rect 231952 331916 232004 331968
rect 243360 331984 243412 332036
rect 243636 331984 243688 332036
rect 273904 331984 273956 332036
rect 433340 331984 433392 332036
rect 244188 331916 244240 331968
rect 289176 331916 289228 331968
rect 289728 331916 289780 331968
rect 536840 331916 536892 331968
rect 17224 331848 17276 331900
rect 231308 331848 231360 331900
rect 244740 331848 244792 331900
rect 245476 331848 245528 331900
rect 287796 331848 287848 331900
rect 560944 331848 560996 331900
rect 285220 331780 285272 331832
rect 256608 331712 256660 331764
rect 243268 331304 243320 331356
rect 243820 331304 243872 331356
rect 237012 331236 237064 331288
rect 237288 331236 237340 331288
rect 239404 331236 239456 331288
rect 240508 331236 240560 331288
rect 268016 331236 268068 331288
rect 239588 331168 239640 331220
rect 268476 331168 268528 331220
rect 272524 331168 272576 331220
rect 240508 331100 240560 331152
rect 275744 331100 275796 331152
rect 283196 331100 283248 331152
rect 283840 331100 283892 331152
rect 262496 330896 262548 330948
rect 320180 330896 320232 330948
rect 211068 330828 211120 330880
rect 263692 330828 263744 330880
rect 328460 330828 328512 330880
rect 165528 330760 165580 330812
rect 246856 330760 246908 330812
rect 269212 330760 269264 330812
rect 382280 330760 382332 330812
rect 144828 330692 144880 330744
rect 244464 330692 244516 330744
rect 273076 330692 273128 330744
rect 411260 330692 411312 330744
rect 128268 330624 128320 330676
rect 276664 330624 276716 330676
rect 451280 330624 451332 330676
rect 121368 330556 121420 330608
rect 242348 330556 242400 330608
rect 71688 330488 71740 330540
rect 237196 330488 237248 330540
rect 259736 330420 259788 330472
rect 285588 330556 285640 330608
rect 539600 330556 539652 330608
rect 288440 330488 288492 330540
rect 289636 330488 289688 330540
rect 573364 330488 573416 330540
rect 279148 330012 279200 330064
rect 279884 330012 279936 330064
rect 238116 329740 238168 329792
rect 238392 329740 238444 329792
rect 226984 329468 227036 329520
rect 262036 329468 262088 329520
rect 303620 329468 303672 329520
rect 264888 329400 264940 329452
rect 338120 329400 338172 329452
rect 206928 329332 206980 329384
rect 251180 329332 251232 329384
rect 267832 329332 267884 329384
rect 367100 329332 367152 329384
rect 153108 329264 153160 329316
rect 246028 329264 246080 329316
rect 276388 329307 276440 329316
rect 276388 329273 276397 329307
rect 276397 329273 276431 329307
rect 276431 329273 276440 329307
rect 276388 329264 276440 329273
rect 280160 329264 280212 329316
rect 393320 329264 393372 329316
rect 151728 329196 151780 329248
rect 244740 329196 244792 329248
rect 272340 329196 272392 329248
rect 415400 329196 415452 329248
rect 78588 329128 78640 329180
rect 237932 329128 237984 329180
rect 268016 329128 268068 329180
rect 269028 329128 269080 329180
rect 279056 329128 279108 329180
rect 467840 329128 467892 329180
rect 34428 329060 34480 329112
rect 233240 329060 233292 329112
rect 286876 329060 286928 329112
rect 550640 329060 550692 329112
rect 249064 328992 249116 329044
rect 249432 328992 249484 329044
rect 284392 328899 284444 328908
rect 284392 328865 284401 328899
rect 284401 328865 284435 328899
rect 284435 328865 284444 328899
rect 284392 328856 284444 328865
rect 283656 328559 283708 328568
rect 283656 328525 283665 328559
rect 283665 328525 283699 328559
rect 283699 328525 283708 328559
rect 283656 328516 283708 328525
rect 229560 328491 229612 328500
rect 229560 328457 229569 328491
rect 229569 328457 229603 328491
rect 229603 328457 229612 328491
rect 229560 328448 229612 328457
rect 240692 328491 240744 328500
rect 240692 328457 240701 328491
rect 240701 328457 240735 328491
rect 240735 328457 240744 328491
rect 240692 328448 240744 328457
rect 249156 328448 249208 328500
rect 267464 328491 267516 328500
rect 267464 328457 267473 328491
rect 267473 328457 267507 328491
rect 267507 328457 267516 328491
rect 267464 328448 267516 328457
rect 231584 328380 231636 328432
rect 258540 328380 258592 328432
rect 258632 328380 258684 328432
rect 284576 328423 284628 328432
rect 284576 328389 284585 328423
rect 284585 328389 284619 328423
rect 284619 328389 284628 328423
rect 284576 328380 284628 328389
rect 261852 328040 261904 328092
rect 299480 328040 299532 328092
rect 222108 327972 222160 328024
rect 252744 327972 252796 328024
rect 283288 327972 283340 328024
rect 400312 327972 400364 328024
rect 168288 327904 168340 327956
rect 247132 327904 247184 327956
rect 273352 327904 273404 327956
rect 425152 327904 425204 327956
rect 150348 327836 150400 327888
rect 244372 327836 244424 327888
rect 277400 327836 277452 327888
rect 462320 327836 462372 327888
rect 82728 327768 82780 327820
rect 238300 327768 238352 327820
rect 282828 327768 282880 327820
rect 502340 327768 502392 327820
rect 38568 327700 38620 327752
rect 233516 327700 233568 327752
rect 290832 327700 290884 327752
rect 557540 327700 557592 327752
rect 288164 327088 288216 327140
rect 233608 327020 233660 327072
rect 237656 327020 237708 327072
rect 274640 326748 274692 326800
rect 263232 326680 263284 326732
rect 322940 326680 322992 326732
rect 226248 326612 226300 326664
rect 253112 326612 253164 326664
rect 266636 326612 266688 326664
rect 360200 326612 360252 326664
rect 171048 326544 171100 326596
rect 247592 326544 247644 326596
rect 274732 326544 274784 326596
rect 157248 326476 157300 326528
rect 246672 326476 246724 326528
rect 96528 326408 96580 326460
rect 238852 326408 238904 326460
rect 272524 326408 272576 326460
rect 279608 326408 279660 326460
rect 280436 326544 280488 326596
rect 408500 326544 408552 326596
rect 433432 326476 433484 326528
rect 53748 326340 53800 326392
rect 235356 326340 235408 326392
rect 251272 326340 251324 326392
rect 251732 326340 251784 326392
rect 252100 326340 252152 326392
rect 252284 326340 252336 326392
rect 265900 326340 265952 326392
rect 266084 326340 266136 326392
rect 273260 326340 273312 326392
rect 273720 326340 273772 326392
rect 273812 326340 273864 326392
rect 274364 326340 274416 326392
rect 276296 326340 276348 326392
rect 276940 326340 276992 326392
rect 443092 326408 443144 326460
rect 280344 326340 280396 326392
rect 280988 326340 281040 326392
rect 281080 326340 281132 326392
rect 281264 326340 281316 326392
rect 286692 326340 286744 326392
rect 286968 326340 287020 326392
rect 288900 326340 288952 326392
rect 289176 326340 289228 326392
rect 287428 326272 287480 326324
rect 564440 326340 564492 326392
rect 265900 326204 265952 326256
rect 266268 326204 266320 326256
rect 272524 326204 272576 326256
rect 279700 326204 279752 326256
rect 269028 325660 269080 325712
rect 269120 325660 269172 325712
rect 269212 325660 269264 325712
rect 263784 325184 263836 325236
rect 331312 325184 331364 325236
rect 213828 325116 213880 325168
rect 251548 325116 251600 325168
rect 271236 325116 271288 325168
rect 394700 325116 394752 325168
rect 141976 325048 142028 325100
rect 244832 325048 244884 325100
rect 273628 325048 273680 325100
rect 429200 325048 429252 325100
rect 92388 324980 92440 325032
rect 239588 324980 239640 325032
rect 277860 324980 277912 325032
rect 471980 324980 472032 325032
rect 42064 324912 42116 324964
rect 233332 324912 233384 324964
rect 290740 324912 290792 324964
rect 568580 324912 568632 324964
rect 284852 324232 284904 324284
rect 285404 324232 285456 324284
rect 265164 323824 265216 323876
rect 349160 323824 349212 323876
rect 217968 323756 218020 323808
rect 251456 323756 251508 323808
rect 270960 323756 271012 323808
rect 398840 323756 398892 323808
rect 159916 323688 159968 323740
rect 245936 323688 245988 323740
rect 278964 323688 279016 323740
rect 436100 323688 436152 323740
rect 99288 323620 99340 323672
rect 240232 323620 240284 323672
rect 281816 323620 281868 323672
rect 509240 323620 509292 323672
rect 46204 323552 46256 323604
rect 234528 323552 234580 323604
rect 259368 323552 259420 323604
rect 285680 323552 285732 323604
rect 290648 323552 290700 323604
rect 571340 323552 571392 323604
rect 259184 323416 259236 323468
rect 259368 323416 259420 323468
rect 260840 322464 260892 322516
rect 306380 322464 306432 322516
rect 264520 322396 264572 322448
rect 335360 322396 335412 322448
rect 146208 322328 146260 322380
rect 244648 322328 244700 322380
rect 269672 322328 269724 322380
rect 385040 322328 385092 322380
rect 103428 322260 103480 322312
rect 241428 322260 241480 322312
rect 277308 322260 277360 322312
rect 458180 322260 458232 322312
rect 56416 322192 56468 322244
rect 235632 322192 235684 322244
rect 287152 322192 287204 322244
rect 554872 322192 554924 322244
rect 289636 321716 289688 321768
rect 298008 321716 298060 321768
rect 379428 321716 379480 321768
rect 386328 321716 386380 321768
rect 287520 321580 287572 321632
rect 287704 321580 287756 321632
rect 210976 321036 211028 321088
rect 252284 321036 252336 321088
rect 272156 321036 272208 321088
rect 418160 321036 418212 321088
rect 136548 320968 136600 321020
rect 243912 320968 243964 321020
rect 278228 320968 278280 321020
rect 466460 320968 466512 321020
rect 125416 320900 125468 320952
rect 242532 320900 242584 320952
rect 279240 320900 279292 320952
rect 476120 320900 476172 320952
rect 74448 320832 74500 320884
rect 233884 320832 233936 320884
rect 286324 320832 286376 320884
rect 540980 320832 541032 320884
rect 262588 319676 262640 319728
rect 317420 319676 317472 319728
rect 215208 319608 215260 319660
rect 251640 319608 251692 319660
rect 268200 319608 268252 319660
rect 371240 319608 371292 319660
rect 154488 319540 154540 319592
rect 246396 319540 246448 319592
rect 283472 319540 283524 319592
rect 447140 319540 447192 319592
rect 67548 319472 67600 319524
rect 229744 319472 229796 319524
rect 238944 319515 238996 319524
rect 238944 319481 238953 319515
rect 238953 319481 238987 319515
rect 238987 319481 238996 319515
rect 238944 319472 238996 319481
rect 280712 319472 280764 319524
rect 487160 319472 487212 319524
rect 50344 319404 50396 319456
rect 234988 319404 235040 319456
rect 261576 319404 261628 319456
rect 278780 319404 278832 319456
rect 287980 319404 288032 319456
rect 556804 319404 556856 319456
rect 231492 318835 231544 318844
rect 231492 318801 231501 318835
rect 231501 318801 231535 318835
rect 231535 318801 231544 318835
rect 231492 318792 231544 318801
rect 243360 318792 243412 318844
rect 243544 318792 243596 318844
rect 254032 318792 254084 318844
rect 254124 318792 254176 318844
rect 265348 318792 265400 318844
rect 265532 318792 265584 318844
rect 283012 318792 283064 318844
rect 283380 318792 283432 318844
rect 284576 318835 284628 318844
rect 284576 318801 284585 318835
rect 284585 318801 284619 318835
rect 284619 318801 284628 318835
rect 284576 318792 284628 318801
rect 229560 318724 229612 318776
rect 249156 318767 249208 318776
rect 249156 318733 249165 318767
rect 249165 318733 249199 318767
rect 249199 318733 249208 318767
rect 249156 318724 249208 318733
rect 269028 318656 269080 318708
rect 269212 318656 269264 318708
rect 262404 318248 262456 318300
rect 321560 318248 321612 318300
rect 276756 318180 276808 318232
rect 454040 318180 454092 318232
rect 140688 318112 140740 318164
rect 244556 318112 244608 318164
rect 281724 318112 281776 318164
rect 505100 318112 505152 318164
rect 85488 318044 85540 318096
rect 238668 318044 238720 318096
rect 259000 318044 259052 318096
rect 281540 318044 281592 318096
rect 289268 318044 289320 318096
rect 567844 318044 567896 318096
rect 233516 317475 233568 317484
rect 233516 317441 233525 317475
rect 233525 317441 233559 317475
rect 233559 317441 233568 317475
rect 233516 317432 233568 317441
rect 237564 317475 237616 317484
rect 237564 317441 237573 317475
rect 237573 317441 237607 317475
rect 237607 317441 237616 317475
rect 237564 317432 237616 317441
rect 238944 317475 238996 317484
rect 238944 317441 238953 317475
rect 238953 317441 238987 317475
rect 238987 317441 238996 317475
rect 238944 317432 238996 317441
rect 272432 317432 272484 317484
rect 272616 317432 272668 317484
rect 277860 317432 277912 317484
rect 277952 317432 278004 317484
rect 283748 317407 283800 317416
rect 283748 317373 283757 317407
rect 283757 317373 283791 317407
rect 283791 317373 283800 317407
rect 283748 317364 283800 317373
rect 288164 317407 288216 317416
rect 288164 317373 288173 317407
rect 288173 317373 288207 317407
rect 288207 317373 288216 317407
rect 288164 317364 288216 317373
rect 267188 316888 267240 316940
rect 364340 316888 364392 316940
rect 271696 316820 271748 316872
rect 405740 316820 405792 316872
rect 143448 316752 143500 316804
rect 245108 316752 245160 316804
rect 280620 316752 280672 316804
rect 460940 316752 460992 316804
rect 107476 316684 107528 316736
rect 240692 316684 240744 316736
rect 257160 316684 257212 316736
rect 270500 316684 270552 316736
rect 283840 316684 283892 316736
rect 516140 316684 516192 316736
rect 256424 316004 256476 316056
rect 256608 316004 256660 316056
rect 268292 315460 268344 315512
rect 374000 315460 374052 315512
rect 272064 315392 272116 315444
rect 408592 315392 408644 315444
rect 147588 315324 147640 315376
rect 245568 315324 245620 315376
rect 279792 315324 279844 315376
rect 478880 315324 478932 315376
rect 19984 315256 20036 315308
rect 231584 315256 231636 315308
rect 284300 315256 284352 315308
rect 529940 315256 529992 315308
rect 269856 314100 269908 314152
rect 389180 314100 389232 314152
rect 273536 314032 273588 314084
rect 423680 314032 423732 314084
rect 158628 313964 158680 314016
rect 246120 313964 246172 314016
rect 279516 313964 279568 314016
rect 484400 313964 484452 314016
rect 24124 313896 24176 313948
rect 232412 313896 232464 313948
rect 286692 313896 286744 313948
rect 545120 313896 545172 313948
rect 275376 312672 275428 312724
rect 437480 312672 437532 312724
rect 161388 312604 161440 312656
rect 246304 312604 246356 312656
rect 280896 312604 280948 312656
rect 491300 312604 491352 312656
rect 31668 312536 31720 312588
rect 233148 312536 233200 312588
rect 286600 312536 286652 312588
rect 552020 312536 552072 312588
rect 288992 311788 289044 311840
rect 289268 311788 289320 311840
rect 271420 311176 271472 311228
rect 401600 311176 401652 311228
rect 110328 311108 110380 311160
rect 241152 311108 241204 311160
rect 274916 311108 274968 311160
rect 441620 311108 441672 311160
rect 299572 310768 299624 310820
rect 304356 310768 304408 310820
rect 320732 310768 320784 310820
rect 328368 310768 328420 310820
rect 359648 310768 359700 310820
rect 367008 310768 367060 310820
rect 475568 310768 475620 310820
rect 482928 310768 482980 310820
rect 541072 310768 541124 310820
rect 543832 310768 543884 310820
rect 288348 310700 288400 310752
rect 296628 310700 296680 310752
rect 340788 310700 340840 310752
rect 347688 310700 347740 310752
rect 379428 310700 379480 310752
rect 386328 310700 386380 310752
rect 398748 310700 398800 310752
rect 405648 310700 405700 310752
rect 418068 310700 418120 310752
rect 424968 310700 425020 310752
rect 437388 310700 437440 310752
rect 444288 310700 444340 310752
rect 456708 310700 456760 310752
rect 463608 310700 463660 310752
rect 495348 310700 495400 310752
rect 502248 310700 502300 310752
rect 514668 310700 514720 310752
rect 521568 310700 521620 310752
rect 533988 310700 534040 310752
rect 540888 310700 540940 310752
rect 261024 309952 261076 310004
rect 310520 309952 310572 310004
rect 268660 309884 268712 309936
rect 378140 309884 378192 309936
rect 280988 309816 281040 309868
rect 494060 309816 494112 309868
rect 31024 309748 31076 309800
rect 232320 309748 232372 309800
rect 287888 309748 287940 309800
rect 563060 309748 563112 309800
rect 229468 309247 229520 309256
rect 229468 309213 229477 309247
rect 229477 309213 229511 309247
rect 229511 309213 229520 309247
rect 229468 309204 229520 309213
rect 243360 309136 243412 309188
rect 243544 309136 243596 309188
rect 249156 309179 249208 309188
rect 249156 309145 249165 309179
rect 249165 309145 249199 309179
rect 249199 309145 249208 309179
rect 249156 309136 249208 309145
rect 3332 309068 3384 309120
rect 213184 309068 213236 309120
rect 229468 309111 229520 309120
rect 229468 309077 229477 309111
rect 229477 309077 229511 309111
rect 229511 309077 229520 309111
rect 229468 309068 229520 309077
rect 233516 309111 233568 309120
rect 233516 309077 233525 309111
rect 233525 309077 233559 309111
rect 233559 309077 233568 309111
rect 233516 309068 233568 309077
rect 237564 309068 237616 309120
rect 238944 309111 238996 309120
rect 238944 309077 238953 309111
rect 238953 309077 238987 309111
rect 238987 309077 238996 309111
rect 238944 309068 238996 309077
rect 284668 309111 284720 309120
rect 284668 309077 284677 309111
rect 284677 309077 284711 309111
rect 284711 309077 284720 309111
rect 284668 309068 284720 309077
rect 289176 309068 289228 309120
rect 289268 309068 289320 309120
rect 237656 309000 237708 309052
rect 283012 309043 283064 309052
rect 283012 309009 283021 309043
rect 283021 309009 283055 309043
rect 283055 309009 283064 309043
rect 283012 309000 283064 309009
rect 263968 308524 264020 308576
rect 339500 308524 339552 308576
rect 281080 308456 281132 308508
rect 498200 308456 498252 308508
rect 289360 308388 289412 308440
rect 574836 308388 574888 308440
rect 278044 307776 278096 307828
rect 278136 307776 278188 307828
rect 288164 307819 288216 307828
rect 288164 307785 288173 307819
rect 288173 307785 288207 307819
rect 288207 307785 288216 307819
rect 288164 307776 288216 307785
rect 251824 307708 251876 307760
rect 260196 307751 260248 307760
rect 260196 307717 260205 307751
rect 260205 307717 260239 307751
rect 260239 307717 260248 307751
rect 260196 307708 260248 307717
rect 260380 307708 260432 307760
rect 260564 307708 260616 307760
rect 272708 307164 272760 307216
rect 412640 307164 412692 307216
rect 277492 307096 277544 307148
rect 473360 307096 473412 307148
rect 43444 307028 43496 307080
rect 233700 307028 233752 307080
rect 282736 307028 282788 307080
rect 512000 307028 512052 307080
rect 256424 306348 256476 306400
rect 256700 306348 256752 306400
rect 272800 305668 272852 305720
rect 416872 305668 416924 305720
rect 38476 305600 38528 305652
rect 282920 305600 282972 305652
rect 520280 305600 520332 305652
rect 275192 304988 275244 305040
rect 275284 304988 275336 305040
rect 277860 304920 277912 304972
rect 278228 304920 278280 304972
rect 274088 304308 274140 304360
rect 426440 304308 426492 304360
rect 42708 304240 42760 304292
rect 234252 304240 234304 304292
rect 283932 304240 283984 304292
rect 523040 304240 523092 304292
rect 275560 302948 275612 303000
rect 444380 302948 444432 303000
rect 50988 302880 51040 302932
rect 235080 302880 235132 302932
rect 527180 302880 527232 302932
rect 238116 302268 238168 302320
rect 275284 302268 275336 302320
rect 238208 302064 238260 302116
rect 256516 302064 256568 302116
rect 256700 302064 256752 302116
rect 284668 302175 284720 302184
rect 284668 302141 284677 302175
rect 284677 302141 284711 302175
rect 284711 302141 284720 302175
rect 284668 302132 284720 302141
rect 275376 302064 275428 302116
rect 277032 301520 277084 301572
rect 448520 301520 448572 301572
rect 284392 301452 284444 301504
rect 534080 301452 534132 301504
rect 276848 300160 276900 300212
rect 455420 300160 455472 300212
rect 285312 300092 285364 300144
rect 536932 300092 536984 300144
rect 283748 299591 283800 299600
rect 283748 299557 283757 299591
rect 283757 299557 283791 299591
rect 283791 299557 283800 299591
rect 283748 299548 283800 299557
rect 229560 299480 229612 299532
rect 238944 299523 238996 299532
rect 238944 299489 238953 299523
rect 238953 299489 238987 299523
rect 238987 299489 238996 299523
rect 238944 299480 238996 299489
rect 302976 299412 303028 299464
rect 579804 299412 579856 299464
rect 260288 299344 260340 299396
rect 277584 298732 277636 298784
rect 469220 298732 469272 298784
rect 254032 298256 254084 298308
rect 251732 298163 251784 298172
rect 251732 298129 251741 298163
rect 251741 298129 251775 298163
rect 251775 298129 251784 298163
rect 251732 298120 251784 298129
rect 254032 298120 254084 298172
rect 237656 298052 237708 298104
rect 283748 298095 283800 298104
rect 283748 298061 283757 298095
rect 283757 298061 283791 298095
rect 283791 298061 283800 298095
rect 283748 298052 283800 298061
rect 288164 298095 288216 298104
rect 288164 298061 288173 298095
rect 288173 298061 288207 298095
rect 288207 298061 288216 298095
rect 288164 298052 288216 298061
rect 282552 297440 282604 297492
rect 502432 297440 502484 297492
rect 285956 297372 286008 297424
rect 547880 297372 547932 297424
rect 278136 296692 278188 296744
rect 278320 296692 278372 296744
rect 289452 296012 289504 296064
rect 482284 296012 482336 296064
rect 288072 295944 288124 295996
rect 565084 295944 565136 295996
rect 3516 295264 3568 295316
rect 227168 295264 227220 295316
rect 289544 294652 289596 294704
rect 475384 294652 475436 294704
rect 290556 294584 290608 294636
rect 569960 294584 570012 294636
rect 263324 293292 263376 293344
rect 324320 293292 324372 293344
rect 289360 293224 289412 293276
rect 573456 293224 573508 293276
rect 275376 292612 275428 292664
rect 251732 292476 251784 292528
rect 275284 292476 275336 292528
rect 272892 291864 272944 291916
rect 419540 291864 419592 291916
rect 282644 291796 282696 291848
rect 506480 291796 506532 291848
rect 274180 290504 274232 290556
rect 430580 290504 430632 290556
rect 284944 290436 284996 290488
rect 524420 290436 524472 290488
rect 256516 289824 256568 289876
rect 238116 289756 238168 289808
rect 238208 289756 238260 289808
rect 241060 289756 241112 289808
rect 241152 289756 241204 289808
rect 243452 289799 243504 289808
rect 243452 289765 243461 289799
rect 243461 289765 243495 289799
rect 243495 289765 243504 289799
rect 243452 289756 243504 289765
rect 284392 289756 284444 289808
rect 284668 289756 284720 289808
rect 256608 289688 256660 289740
rect 277952 289552 278004 289604
rect 276020 289144 276072 289196
rect 451372 289144 451424 289196
rect 286048 289076 286100 289128
rect 549260 289076 549312 289128
rect 237564 288439 237616 288448
rect 237564 288405 237573 288439
rect 237573 288405 237607 288439
rect 237607 288405 237616 288439
rect 237564 288396 237616 288405
rect 283840 288396 283892 288448
rect 288164 288439 288216 288448
rect 288164 288405 288173 288439
rect 288173 288405 288207 288439
rect 288207 288405 288216 288439
rect 288164 288396 288216 288405
rect 276296 287716 276348 287768
rect 459652 287716 459704 287768
rect 289360 287648 289412 287700
rect 571432 287648 571484 287700
rect 251640 287079 251692 287088
rect 251640 287045 251649 287079
rect 251649 287045 251683 287079
rect 251683 287045 251692 287079
rect 251640 287036 251692 287045
rect 253848 287036 253900 287088
rect 254032 287036 254084 287088
rect 279608 286288 279660 286340
rect 477500 286288 477552 286340
rect 279700 284928 279752 284980
rect 480260 284928 480312 284980
rect 278872 283568 278924 283620
rect 485780 283568 485832 283620
rect 275376 282888 275428 282940
rect 275284 282820 275336 282872
rect 280252 282140 280304 282192
rect 488540 282140 488592 282192
rect 260104 281936 260156 281988
rect 260288 281936 260340 281988
rect 281264 280780 281316 280832
rect 492680 280780 492732 280832
rect 243544 280168 243596 280220
rect 260288 280168 260340 280220
rect 260564 280168 260616 280220
rect 229560 280143 229612 280152
rect 229560 280109 229569 280143
rect 229569 280109 229603 280143
rect 229603 280109 229612 280143
rect 229560 280100 229612 280109
rect 259920 280100 259972 280152
rect 260104 280100 260156 280152
rect 281356 279420 281408 279472
rect 499580 279420 499632 279472
rect 284392 279148 284444 279200
rect 284944 279148 284996 279200
rect 243544 278672 243596 278724
rect 259920 278715 259972 278724
rect 259920 278681 259929 278715
rect 259929 278681 259963 278715
rect 259963 278681 259972 278715
rect 259920 278672 259972 278681
rect 281908 277992 281960 278044
rect 510620 277992 510672 278044
rect 277860 277423 277912 277432
rect 277860 277389 277869 277423
rect 277869 277389 277903 277423
rect 277903 277389 277912 277423
rect 277860 277380 277912 277389
rect 282092 276632 282144 276684
rect 513380 276632 513432 276684
rect 393964 275952 394016 276004
rect 580172 275952 580224 276004
rect 260288 275272 260340 275324
rect 260564 275272 260616 275324
rect 284116 273912 284168 273964
rect 517520 273912 517572 273964
rect 272432 273300 272484 273352
rect 272340 273164 272392 273216
rect 283748 272484 283800 272536
rect 520372 272484 520424 272536
rect 284484 271124 284536 271176
rect 528652 271124 528704 271176
rect 229652 270512 229704 270564
rect 241152 270487 241204 270496
rect 241152 270453 241161 270487
rect 241161 270453 241195 270487
rect 241195 270453 241204 270487
rect 241152 270444 241204 270453
rect 284944 269764 284996 269816
rect 531320 269764 531372 269816
rect 270868 269084 270920 269136
rect 270960 269084 271012 269136
rect 288072 269084 288124 269136
rect 288164 269084 288216 269136
rect 284760 268336 284812 268388
rect 535460 268336 535512 268388
rect 260104 267724 260156 267776
rect 284852 266976 284904 267028
rect 538220 266976 538272 267028
rect 3516 266296 3568 266348
rect 211804 266296 211856 266348
rect 286784 265616 286836 265668
rect 542360 265616 542412 265668
rect 315304 264868 315356 264920
rect 580172 264868 580224 264920
rect 286140 262828 286192 262880
rect 546592 262828 546644 262880
rect 286232 261468 286284 261520
rect 553400 261468 553452 261520
rect 241152 260899 241204 260908
rect 241152 260865 241161 260899
rect 241161 260865 241195 260899
rect 241195 260865 241204 260899
rect 241152 260856 241204 260865
rect 254032 260856 254084 260908
rect 229560 260831 229612 260840
rect 229560 260797 229569 260831
rect 229569 260797 229603 260831
rect 229603 260797 229612 260831
rect 229560 260788 229612 260797
rect 251364 260788 251416 260840
rect 251640 260788 251692 260840
rect 275376 260924 275428 260976
rect 275284 260720 275336 260772
rect 287244 260108 287296 260160
rect 556160 260108 556212 260160
rect 237656 259564 237708 259616
rect 237656 259428 237708 259480
rect 260380 259428 260432 259480
rect 260564 259428 260616 259480
rect 270776 259428 270828 259480
rect 270960 259428 271012 259480
rect 288164 258680 288216 258732
rect 560300 258680 560352 258732
rect 253940 258111 253992 258120
rect 253940 258077 253949 258111
rect 253949 258077 253983 258111
rect 253983 258077 253992 258111
rect 253940 258068 253992 258077
rect 260104 258043 260156 258052
rect 260104 258009 260113 258043
rect 260113 258009 260147 258043
rect 260147 258009 260156 258043
rect 260104 258000 260156 258009
rect 260380 258000 260432 258052
rect 287520 257320 287572 257372
rect 563152 257320 563204 257372
rect 243544 256708 243596 256760
rect 291108 255960 291160 256012
rect 471244 255960 471296 256012
rect 243544 255212 243596 255264
rect 277860 254532 277912 254584
rect 278044 254532 278096 254584
rect 237656 253988 237708 254040
rect 237564 253852 237616 253904
rect 251364 253172 251416 253224
rect 251548 253172 251600 253224
rect 3148 252492 3200 252544
rect 225788 252492 225840 252544
rect 301596 252492 301648 252544
rect 579804 252492 579856 252544
rect 229652 251200 229704 251252
rect 275284 249815 275336 249824
rect 275284 249781 275293 249815
rect 275293 249781 275327 249815
rect 275327 249781 275336 249815
rect 275284 249772 275336 249781
rect 260104 249747 260156 249756
rect 260104 249713 260113 249747
rect 260113 249713 260147 249747
rect 260147 249713 260156 249747
rect 260104 249704 260156 249713
rect 260196 248455 260248 248464
rect 260196 248421 260205 248455
rect 260205 248421 260239 248455
rect 260239 248421 260248 248455
rect 260196 248412 260248 248421
rect 275284 248455 275336 248464
rect 275284 248421 275293 248455
rect 275293 248421 275327 248455
rect 275327 248421 275336 248455
rect 275284 248412 275336 248421
rect 237564 248387 237616 248396
rect 237564 248353 237573 248387
rect 237573 248353 237607 248387
rect 237607 248353 237616 248387
rect 237564 248344 237616 248353
rect 277860 248344 277912 248396
rect 278044 248344 278096 248396
rect 240876 246984 240928 247036
rect 241152 246984 241204 247036
rect 251548 244944 251600 244996
rect 251732 244944 251784 244996
rect 259920 244944 259972 244996
rect 260104 244944 260156 244996
rect 258632 244400 258684 244452
rect 259368 244264 259420 244316
rect 259276 244196 259328 244248
rect 237656 244128 237708 244180
rect 272340 241476 272392 241528
rect 272432 241476 272484 241528
rect 278228 241476 278280 241528
rect 278320 241476 278372 241528
rect 243544 240184 243596 240236
rect 258540 240159 258592 240168
rect 258540 240125 258549 240159
rect 258549 240125 258583 240159
rect 258583 240125 258592 240159
rect 258540 240116 258592 240125
rect 270776 240116 270828 240168
rect 270960 240116 271012 240168
rect 275284 240116 275336 240168
rect 275376 240116 275428 240168
rect 259184 240048 259236 240100
rect 259276 240048 259328 240100
rect 260196 240048 260248 240100
rect 254032 238731 254084 238740
rect 254032 238697 254041 238731
rect 254041 238697 254075 238731
rect 254075 238697 254084 238731
rect 254032 238688 254084 238697
rect 275376 238688 275428 238740
rect 275560 238688 275612 238740
rect 277768 238688 277820 238740
rect 278044 238688 278096 238740
rect 238116 237328 238168 237380
rect 238300 237328 238352 237380
rect 243544 237328 243596 237380
rect 259920 235288 259972 235340
rect 260196 235288 260248 235340
rect 237656 231956 237708 232008
rect 229652 231820 229704 231872
rect 229836 231820 229888 231872
rect 258540 230460 258592 230512
rect 258632 230460 258684 230512
rect 260288 230503 260340 230512
rect 260288 230469 260297 230503
rect 260297 230469 260331 230503
rect 260331 230469 260340 230503
rect 260288 230460 260340 230469
rect 254032 230299 254084 230308
rect 254032 230265 254041 230299
rect 254041 230265 254075 230299
rect 254075 230265 254084 230299
rect 254032 230256 254084 230265
rect 238944 229032 238996 229084
rect 239128 229032 239180 229084
rect 240876 229032 240928 229084
rect 241152 229032 241204 229084
rect 259460 227944 259512 227996
rect 270408 227944 270460 227996
rect 321468 227876 321520 227928
rect 323032 227876 323084 227928
rect 302148 227808 302200 227860
rect 309048 227808 309100 227860
rect 437388 227808 437440 227860
rect 444288 227808 444340 227860
rect 476028 227808 476080 227860
rect 482928 227808 482980 227860
rect 533988 227808 534040 227860
rect 540888 227808 540940 227860
rect 553308 227808 553360 227860
rect 560208 227808 560260 227860
rect 572628 227808 572680 227860
rect 579528 227808 579580 227860
rect 237472 227783 237524 227792
rect 237472 227749 237481 227783
rect 237481 227749 237515 227783
rect 237515 227749 237524 227783
rect 237472 227740 237524 227749
rect 277952 225199 278004 225208
rect 277952 225165 277961 225199
rect 277961 225165 277995 225199
rect 277995 225165 278004 225199
rect 277952 225156 278004 225165
rect 251824 224995 251876 225004
rect 251824 224961 251833 224995
rect 251833 224961 251867 224995
rect 251867 224961 251876 224995
rect 251824 224952 251876 224961
rect 3148 223524 3200 223576
rect 209044 223524 209096 223576
rect 260288 222300 260340 222352
rect 251824 222207 251876 222216
rect 251824 222173 251833 222207
rect 251833 222173 251867 222207
rect 251867 222173 251876 222207
rect 251824 222164 251876 222173
rect 256516 222164 256568 222216
rect 256608 222164 256660 222216
rect 260104 222164 260156 222216
rect 260196 222164 260248 222216
rect 260288 222164 260340 222216
rect 259552 220804 259604 220856
rect 259644 220804 259696 220856
rect 277952 220847 278004 220856
rect 277952 220813 277961 220847
rect 277961 220813 277995 220847
rect 277995 220813 278004 220847
rect 277952 220804 278004 220813
rect 270960 220779 271012 220788
rect 270960 220745 270969 220779
rect 270969 220745 271003 220779
rect 271003 220745 271012 220779
rect 270960 220736 271012 220745
rect 243452 219487 243504 219496
rect 243452 219453 243461 219487
rect 243461 219453 243495 219487
rect 243495 219453 243504 219487
rect 243452 219444 243504 219453
rect 277952 219376 278004 219428
rect 237656 219351 237708 219360
rect 237656 219317 237665 219351
rect 237665 219317 237699 219351
rect 237699 219317 237708 219351
rect 237656 219308 237708 219317
rect 243452 219351 243504 219360
rect 243452 219317 243461 219351
rect 243461 219317 243495 219351
rect 243495 219317 243504 219351
rect 243452 219308 243504 219317
rect 238852 218832 238904 218884
rect 312544 217948 312596 218000
rect 580172 217948 580224 218000
rect 272432 215364 272484 215416
rect 272340 215228 272392 215280
rect 237656 214591 237708 214600
rect 237656 214557 237665 214591
rect 237665 214557 237699 214591
rect 237699 214557 237708 214591
rect 237656 214548 237708 214557
rect 260012 212576 260064 212628
rect 229652 212508 229704 212560
rect 229836 212508 229888 212560
rect 259368 212508 259420 212560
rect 259644 212508 259696 212560
rect 260012 212440 260064 212492
rect 270960 211191 271012 211200
rect 270960 211157 270969 211191
rect 270969 211157 271003 211191
rect 271003 211157 271012 211191
rect 270960 211148 271012 211157
rect 277860 209831 277912 209840
rect 277860 209797 277869 209831
rect 277869 209797 277903 209831
rect 277903 209797 277912 209831
rect 277860 209788 277912 209797
rect 275284 209763 275336 209772
rect 275284 209729 275293 209763
rect 275293 209729 275327 209763
rect 275327 209729 275336 209763
rect 275284 209720 275336 209729
rect 3516 208292 3568 208344
rect 180064 208292 180116 208344
rect 230848 205640 230900 205692
rect 231032 205640 231084 205692
rect 251548 205640 251600 205692
rect 275284 205615 275336 205624
rect 275284 205581 275293 205615
rect 275293 205581 275327 205615
rect 275327 205581 275336 205615
rect 275284 205572 275336 205581
rect 298836 205572 298888 205624
rect 579804 205572 579856 205624
rect 251548 205504 251600 205556
rect 238944 205343 238996 205352
rect 238944 205309 238953 205343
rect 238953 205309 238987 205343
rect 238987 205309 238996 205343
rect 238944 205300 238996 205309
rect 243544 202852 243596 202904
rect 258632 202852 258684 202904
rect 258724 202852 258776 202904
rect 259920 202852 259972 202904
rect 260104 202852 260156 202904
rect 260196 202852 260248 202904
rect 260288 202852 260340 202904
rect 237564 201424 237616 201476
rect 237656 201424 237708 201476
rect 241152 201424 241204 201476
rect 241336 201424 241388 201476
rect 259736 201424 259788 201476
rect 260104 201424 260156 201476
rect 260288 201424 260340 201476
rect 251640 197888 251692 197940
rect 251732 197888 251784 197940
rect 230848 195916 230900 195968
rect 231032 195916 231084 195968
rect 229652 193196 229704 193248
rect 229836 193196 229888 193248
rect 260196 191879 260248 191888
rect 260196 191845 260205 191879
rect 260205 191845 260239 191879
rect 260239 191845 260248 191879
rect 260196 191836 260248 191845
rect 277952 191836 278004 191888
rect 243360 191811 243412 191820
rect 243360 191777 243369 191811
rect 243369 191777 243403 191811
rect 243403 191777 243412 191811
rect 243360 191768 243412 191777
rect 270960 191811 271012 191820
rect 270960 191777 270969 191811
rect 270969 191777 271003 191811
rect 271003 191777 271012 191811
rect 270960 191768 271012 191777
rect 278044 191700 278096 191752
rect 275376 190612 275428 190664
rect 275284 190519 275336 190528
rect 275284 190485 275293 190519
rect 275293 190485 275327 190519
rect 275327 190485 275336 190519
rect 275284 190476 275336 190485
rect 277768 190408 277820 190460
rect 278044 190408 278096 190460
rect 230848 186328 230900 186380
rect 231032 186328 231084 186380
rect 237564 186328 237616 186380
rect 275284 186328 275336 186380
rect 243452 186260 243504 186312
rect 259920 186260 259972 186312
rect 260104 186260 260156 186312
rect 237656 186192 237708 186244
rect 278228 186260 278280 186312
rect 278412 186260 278464 186312
rect 275376 186192 275428 186244
rect 260288 183515 260340 183524
rect 260288 183481 260297 183515
rect 260297 183481 260331 183515
rect 260331 183481 260340 183515
rect 260288 183472 260340 183481
rect 270960 182223 271012 182232
rect 270960 182189 270969 182223
rect 270969 182189 271003 182223
rect 271003 182189 271012 182223
rect 270960 182180 271012 182189
rect 241152 182112 241204 182164
rect 241336 182112 241388 182164
rect 308404 182112 308456 182164
rect 580172 182112 580224 182164
rect 243544 182044 243596 182096
rect 3240 180752 3292 180804
rect 207664 180752 207716 180804
rect 258632 180795 258684 180804
rect 258632 180761 258641 180795
rect 258641 180761 258675 180795
rect 258675 180761 258684 180795
rect 258632 180752 258684 180761
rect 259276 180752 259328 180804
rect 259368 180752 259420 180804
rect 270960 180752 271012 180804
rect 275376 180752 275428 180804
rect 259920 178712 259972 178764
rect 260104 178712 260156 178764
rect 260288 178755 260340 178764
rect 260288 178721 260297 178755
rect 260297 178721 260331 178755
rect 260331 178721 260340 178755
rect 260288 178712 260340 178721
rect 230848 176604 230900 176656
rect 231032 176604 231084 176656
rect 243452 174403 243504 174412
rect 243452 174369 243461 174403
rect 243461 174369 243495 174403
rect 243495 174369 243504 174403
rect 243452 174360 243504 174369
rect 237564 173952 237616 174004
rect 237656 173952 237708 174004
rect 256608 173952 256660 174004
rect 229652 173884 229704 173936
rect 229836 173884 229888 173936
rect 253940 173884 253992 173936
rect 254124 173816 254176 173868
rect 237564 172499 237616 172508
rect 237564 172465 237573 172499
rect 237573 172465 237607 172499
rect 237607 172465 237616 172499
rect 237564 172456 237616 172465
rect 238208 172499 238260 172508
rect 238208 172465 238217 172499
rect 238217 172465 238251 172499
rect 238251 172465 238260 172499
rect 238208 172456 238260 172465
rect 258632 171207 258684 171216
rect 258632 171173 258641 171207
rect 258641 171173 258675 171207
rect 258675 171173 258684 171207
rect 258632 171164 258684 171173
rect 270776 171139 270828 171148
rect 270776 171105 270785 171139
rect 270785 171105 270819 171139
rect 270819 171105 270828 171139
rect 270776 171096 270828 171105
rect 275192 171139 275244 171148
rect 275192 171105 275201 171139
rect 275201 171105 275235 171139
rect 275235 171105 275244 171139
rect 275192 171096 275244 171105
rect 277860 171096 277912 171148
rect 277952 171096 278004 171148
rect 251640 171028 251692 171080
rect 251824 171028 251876 171080
rect 258632 171071 258684 171080
rect 258632 171037 258641 171071
rect 258641 171037 258675 171071
rect 258675 171037 258684 171071
rect 258632 171028 258684 171037
rect 259368 171071 259420 171080
rect 259368 171037 259377 171071
rect 259377 171037 259411 171071
rect 259411 171037 259420 171071
rect 259368 171028 259420 171037
rect 485044 171028 485096 171080
rect 580172 171028 580224 171080
rect 275192 171003 275244 171012
rect 275192 170969 275201 171003
rect 275201 170969 275235 171003
rect 275235 170969 275244 171003
rect 275192 170960 275244 170969
rect 256516 169779 256568 169788
rect 256516 169745 256525 169779
rect 256525 169745 256559 169779
rect 256559 169745 256568 169779
rect 256516 169736 256568 169745
rect 230848 167016 230900 167068
rect 231032 167016 231084 167068
rect 243452 167016 243504 167068
rect 237564 166991 237616 167000
rect 237564 166957 237573 166991
rect 237573 166957 237607 166991
rect 237607 166957 237616 166991
rect 237564 166948 237616 166957
rect 243544 166880 243596 166932
rect 3516 165520 3568 165572
rect 222844 165520 222896 165572
rect 229560 164160 229612 164212
rect 229836 164160 229888 164212
rect 260104 164160 260156 164212
rect 260196 164160 260248 164212
rect 260288 164160 260340 164212
rect 260380 164160 260432 164212
rect 238208 162911 238260 162920
rect 238208 162877 238217 162911
rect 238217 162877 238251 162911
rect 238251 162877 238260 162911
rect 238208 162868 238260 162877
rect 237564 162800 237616 162852
rect 237656 162800 237708 162852
rect 238944 162800 238996 162852
rect 239128 162800 239180 162852
rect 241152 162843 241204 162852
rect 241152 162809 241161 162843
rect 241161 162809 241195 162843
rect 241195 162809 241204 162843
rect 241152 162800 241204 162809
rect 260196 162843 260248 162852
rect 260196 162809 260205 162843
rect 260205 162809 260239 162843
rect 260239 162809 260248 162843
rect 260196 162800 260248 162809
rect 259368 161551 259420 161560
rect 259368 161517 259377 161551
rect 259377 161517 259411 161551
rect 259411 161517 259420 161551
rect 259368 161508 259420 161517
rect 258632 161483 258684 161492
rect 258632 161449 258641 161483
rect 258641 161449 258675 161483
rect 258675 161449 258684 161483
rect 258632 161440 258684 161449
rect 275376 161440 275428 161492
rect 277860 161440 277912 161492
rect 278136 161440 278188 161492
rect 259368 160012 259420 160064
rect 297456 158652 297508 158704
rect 579804 158652 579856 158704
rect 243544 157360 243596 157412
rect 230848 157292 230900 157344
rect 231032 157292 231084 157344
rect 260380 154640 260432 154692
rect 260288 154504 260340 154556
rect 243452 153323 243504 153332
rect 243452 153289 243461 153323
rect 243461 153289 243495 153323
rect 243495 153289 243504 153323
rect 243452 153280 243504 153289
rect 260196 153323 260248 153332
rect 260196 153289 260205 153323
rect 260205 153289 260239 153323
rect 260239 153289 260248 153323
rect 260196 153280 260248 153289
rect 241152 153255 241204 153264
rect 241152 153221 241161 153255
rect 241161 153221 241195 153255
rect 241195 153221 241204 153255
rect 241152 153212 241204 153221
rect 237564 153187 237616 153196
rect 237564 153153 237573 153187
rect 237573 153153 237607 153187
rect 237607 153153 237616 153187
rect 237564 153144 237616 153153
rect 238208 153187 238260 153196
rect 238208 153153 238217 153187
rect 238217 153153 238251 153187
rect 238251 153153 238260 153187
rect 238208 153144 238260 153153
rect 238944 153187 238996 153196
rect 238944 153153 238953 153187
rect 238953 153153 238987 153187
rect 238987 153153 238996 153187
rect 238944 153144 238996 153153
rect 251732 151784 251784 151836
rect 251824 151784 251876 151836
rect 253940 151784 253992 151836
rect 254124 151784 254176 151836
rect 256608 151784 256660 151836
rect 256884 151784 256936 151836
rect 258632 151759 258684 151768
rect 258632 151725 258641 151759
rect 258641 151725 258675 151759
rect 258675 151725 258684 151759
rect 258632 151716 258684 151725
rect 256792 148996 256844 149048
rect 243452 147704 243504 147756
rect 278136 147636 278188 147688
rect 278320 147636 278372 147688
rect 237564 147611 237616 147620
rect 237564 147577 237573 147611
rect 237573 147577 237607 147611
rect 237607 147577 237616 147611
rect 237564 147568 237616 147577
rect 243452 147568 243504 147620
rect 238944 147203 238996 147212
rect 238944 147169 238953 147203
rect 238953 147169 238987 147203
rect 238987 147169 238996 147203
rect 238944 147160 238996 147169
rect 260104 144848 260156 144900
rect 260196 144848 260248 144900
rect 260288 144848 260340 144900
rect 260380 144848 260432 144900
rect 276480 144891 276532 144900
rect 276480 144857 276489 144891
rect 276489 144857 276523 144891
rect 276523 144857 276532 144891
rect 276480 144848 276532 144857
rect 238208 143599 238260 143608
rect 238208 143565 238217 143599
rect 238217 143565 238251 143599
rect 238251 143565 238260 143599
rect 238208 143556 238260 143565
rect 237656 143420 237708 143472
rect 258632 142171 258684 142180
rect 258632 142137 258641 142171
rect 258641 142137 258675 142171
rect 258675 142137 258684 142171
rect 258632 142128 258684 142137
rect 259276 142171 259328 142180
rect 259276 142137 259285 142171
rect 259285 142137 259319 142171
rect 259319 142137 259328 142171
rect 259276 142128 259328 142137
rect 275376 142128 275428 142180
rect 275468 142128 275520 142180
rect 243544 142060 243596 142112
rect 254124 142060 254176 142112
rect 256424 139451 256476 139460
rect 256424 139417 256433 139451
rect 256433 139417 256467 139451
rect 256467 139417 256476 139451
rect 256424 139408 256476 139417
rect 260104 138660 260156 138712
rect 260380 138660 260432 138712
rect 229560 137980 229612 138032
rect 229468 137912 229520 137964
rect 251732 137096 251784 137148
rect 3516 136552 3568 136604
rect 227076 136552 227128 136604
rect 275468 135260 275520 135312
rect 276480 135303 276532 135312
rect 276480 135269 276489 135303
rect 276489 135269 276523 135303
rect 276523 135269 276532 135303
rect 276480 135260 276532 135269
rect 275376 135192 275428 135244
rect 278136 135235 278188 135244
rect 278136 135201 278145 135235
rect 278145 135201 278179 135235
rect 278179 135201 278188 135235
rect 278136 135192 278188 135201
rect 496084 135192 496136 135244
rect 580172 135192 580224 135244
rect 281448 134512 281500 134564
rect 495440 134512 495492 134564
rect 237564 134011 237616 134020
rect 237564 133977 237573 134011
rect 237573 133977 237607 134011
rect 237607 133977 237616 134011
rect 237564 133968 237616 133977
rect 238116 133875 238168 133884
rect 238116 133841 238125 133875
rect 238125 133841 238159 133875
rect 238159 133841 238168 133875
rect 238116 133832 238168 133841
rect 238668 133832 238720 133884
rect 238944 133832 238996 133884
rect 260288 133875 260340 133884
rect 260288 133841 260297 133875
rect 260297 133841 260331 133875
rect 260331 133841 260340 133875
rect 260288 133832 260340 133841
rect 275376 133875 275428 133884
rect 275376 133841 275385 133875
rect 275385 133841 275419 133875
rect 275419 133841 275428 133875
rect 275376 133832 275428 133841
rect 251640 132515 251692 132524
rect 251640 132481 251649 132515
rect 251649 132481 251683 132515
rect 251683 132481 251692 132515
rect 251640 132472 251692 132481
rect 254032 132515 254084 132524
rect 254032 132481 254041 132515
rect 254041 132481 254075 132515
rect 254075 132481 254084 132515
rect 254032 132472 254084 132481
rect 258540 131087 258592 131096
rect 258540 131053 258549 131087
rect 258549 131053 258583 131087
rect 258583 131053 258592 131087
rect 258540 131044 258592 131053
rect 278228 128256 278280 128308
rect 260104 125604 260156 125656
rect 260196 125604 260248 125656
rect 272340 125536 272392 125588
rect 272432 125536 272484 125588
rect 251640 124244 251692 124296
rect 260288 124287 260340 124296
rect 260288 124253 260297 124287
rect 260297 124253 260331 124287
rect 260331 124253 260340 124287
rect 260288 124244 260340 124253
rect 243452 124219 243504 124228
rect 243452 124185 243461 124219
rect 243461 124185 243495 124219
rect 243495 124185 243504 124219
rect 243452 124176 243504 124185
rect 241060 124151 241112 124160
rect 241060 124117 241069 124151
rect 241069 124117 241103 124151
rect 241103 124117 241112 124151
rect 241060 124108 241112 124117
rect 253940 124176 253992 124228
rect 254032 124176 254084 124228
rect 275376 124219 275428 124228
rect 275376 124185 275385 124219
rect 275385 124185 275419 124219
rect 275419 124185 275428 124219
rect 275376 124176 275428 124185
rect 260104 124151 260156 124160
rect 260104 124117 260113 124151
rect 260113 124117 260147 124151
rect 260147 124117 260156 124151
rect 260104 124108 260156 124117
rect 260288 124151 260340 124160
rect 260288 124117 260297 124151
rect 260297 124117 260331 124151
rect 260331 124117 260340 124151
rect 260288 124108 260340 124117
rect 272432 124108 272484 124160
rect 272616 124108 272668 124160
rect 309784 124108 309836 124160
rect 580172 124108 580224 124160
rect 251732 124040 251784 124092
rect 238116 122859 238168 122868
rect 238116 122825 238125 122859
rect 238125 122825 238159 122859
rect 238159 122825 238168 122859
rect 238116 122816 238168 122825
rect 2964 122748 3016 122800
rect 218704 122748 218756 122800
rect 253940 122791 253992 122800
rect 253940 122757 253949 122791
rect 253949 122757 253983 122791
rect 253983 122757 253992 122791
rect 253940 122748 253992 122757
rect 256516 122791 256568 122800
rect 256516 122757 256525 122791
rect 256525 122757 256559 122791
rect 256559 122757 256568 122791
rect 256516 122748 256568 122757
rect 259276 122748 259328 122800
rect 259368 122680 259420 122732
rect 219256 122068 219308 122120
rect 252192 122068 252244 122120
rect 258632 121456 258684 121508
rect 238116 121388 238168 121440
rect 238852 121388 238904 121440
rect 272616 121388 272668 121440
rect 276572 119348 276624 119400
rect 243452 118872 243504 118924
rect 229560 118668 229612 118720
rect 270960 118668 271012 118720
rect 229468 118600 229520 118652
rect 270960 118532 271012 118584
rect 238852 115336 238904 115388
rect 241152 114520 241204 114572
rect 260196 114520 260248 114572
rect 260380 114520 260432 114572
rect 278228 114520 278280 114572
rect 237564 113160 237616 113212
rect 237656 113160 237708 113212
rect 256608 113160 256660 113212
rect 238116 113092 238168 113144
rect 254124 111800 254176 111852
rect 272432 111843 272484 111852
rect 272432 111809 272441 111843
rect 272441 111809 272475 111843
rect 272475 111809 272484 111843
rect 272432 111800 272484 111809
rect 258632 111775 258684 111784
rect 258632 111741 258641 111775
rect 258641 111741 258675 111775
rect 258675 111741 258684 111775
rect 258632 111732 258684 111741
rect 291936 111732 291988 111784
rect 579804 111732 579856 111784
rect 272432 111664 272484 111716
rect 251824 110372 251876 110424
rect 243544 108987 243596 108996
rect 243544 108953 243553 108987
rect 243553 108953 243587 108987
rect 243587 108953 243596 108987
rect 243544 108944 243596 108953
rect 276480 107627 276532 107636
rect 276480 107593 276489 107627
rect 276489 107593 276523 107627
rect 276523 107593 276532 107627
rect 276480 107584 276532 107593
rect 238852 106292 238904 106344
rect 249064 106224 249116 106276
rect 238852 106156 238904 106208
rect 248972 106199 249024 106208
rect 248972 106165 248981 106199
rect 248981 106165 249015 106199
rect 249015 106165 249024 106199
rect 248972 106156 249024 106165
rect 249156 106156 249208 106208
rect 249064 106088 249116 106140
rect 249156 106020 249208 106072
rect 278320 104907 278372 104916
rect 278320 104873 278329 104907
rect 278329 104873 278363 104907
rect 278363 104873 278372 104907
rect 278320 104864 278372 104873
rect 253940 103572 253992 103624
rect 254124 103572 254176 103624
rect 238116 103504 238168 103556
rect 238208 103504 238260 103556
rect 258632 102187 258684 102196
rect 258632 102153 258641 102187
rect 258641 102153 258675 102187
rect 258675 102153 258684 102187
rect 258632 102144 258684 102153
rect 272340 102187 272392 102196
rect 272340 102153 272349 102187
rect 272349 102153 272383 102187
rect 272383 102153 272392 102187
rect 272340 102144 272392 102153
rect 238208 102076 238260 102128
rect 260104 102119 260156 102128
rect 260104 102085 260113 102119
rect 260113 102085 260147 102119
rect 260147 102085 260156 102119
rect 260104 102076 260156 102085
rect 243544 101396 243596 101448
rect 243544 101260 243596 101312
rect 251732 100759 251784 100768
rect 251732 100725 251741 100759
rect 251741 100725 251775 100759
rect 251775 100725 251784 100759
rect 251732 100716 251784 100725
rect 229560 99356 229612 99408
rect 229468 99288 229520 99340
rect 237656 99356 237708 99408
rect 260288 99356 260340 99408
rect 237564 99288 237616 99340
rect 260380 99288 260432 99340
rect 248972 97835 249024 97844
rect 248972 97801 248981 97835
rect 248981 97801 249015 97835
rect 249015 97801 249024 97835
rect 248972 97792 249024 97801
rect 258632 97248 258684 97300
rect 272432 97248 272484 97300
rect 253848 95251 253900 95260
rect 253848 95217 253857 95251
rect 253857 95217 253891 95251
rect 253891 95217 253900 95251
rect 253848 95208 253900 95217
rect 237564 95183 237616 95192
rect 237564 95149 237573 95183
rect 237573 95149 237607 95183
rect 237607 95149 237616 95183
rect 237564 95140 237616 95149
rect 238852 95140 238904 95192
rect 238944 95072 238996 95124
rect 3516 93780 3568 93832
rect 204904 93780 204956 93832
rect 275284 93823 275336 93832
rect 275284 93789 275293 93823
rect 275293 93789 275327 93823
rect 275327 93789 275336 93823
rect 275284 93780 275336 93789
rect 238116 92531 238168 92540
rect 238116 92497 238125 92531
rect 238125 92497 238159 92531
rect 238159 92497 238168 92531
rect 238116 92488 238168 92497
rect 260196 92488 260248 92540
rect 253848 91103 253900 91112
rect 253848 91069 253857 91103
rect 253857 91069 253891 91103
rect 253891 91069 253900 91103
rect 253848 91060 253900 91069
rect 305644 88272 305696 88324
rect 580172 88272 580224 88324
rect 243544 86955 243596 86964
rect 243544 86921 243553 86955
rect 243553 86921 243587 86955
rect 243587 86921 243596 86955
rect 243544 86912 243596 86921
rect 248880 86912 248932 86964
rect 249156 86955 249208 86964
rect 249156 86921 249165 86955
rect 249165 86921 249199 86955
rect 249199 86921 249208 86955
rect 249156 86912 249208 86921
rect 248972 86887 249024 86896
rect 248972 86853 248981 86887
rect 248981 86853 249015 86887
rect 249015 86853 249024 86887
rect 248972 86844 249024 86853
rect 249064 86844 249116 86896
rect 249064 86708 249116 86760
rect 260380 86504 260432 86556
rect 259368 85756 259420 85808
rect 259276 85688 259328 85740
rect 237656 85552 237708 85604
rect 238116 85552 238168 85604
rect 238208 85552 238260 85604
rect 253848 85552 253900 85604
rect 253940 85552 253992 85604
rect 256516 85552 256568 85604
rect 256700 85552 256752 85604
rect 258540 84235 258592 84244
rect 258540 84201 258549 84235
rect 258549 84201 258583 84235
rect 258583 84201 258592 84235
rect 258540 84192 258592 84201
rect 275284 84235 275336 84244
rect 275284 84201 275293 84235
rect 275293 84201 275327 84235
rect 275327 84201 275336 84235
rect 275284 84192 275336 84201
rect 251732 84167 251784 84176
rect 251732 84133 251741 84167
rect 251741 84133 251775 84167
rect 251775 84133 251784 84167
rect 251732 84124 251784 84133
rect 259276 84167 259328 84176
rect 259276 84133 259285 84167
rect 259285 84133 259319 84167
rect 259319 84133 259328 84167
rect 259276 84124 259328 84133
rect 237656 82764 237708 82816
rect 248880 82084 248932 82136
rect 229560 80155 229612 80164
rect 229560 80121 229569 80155
rect 229569 80121 229603 80155
rect 229603 80121 229612 80155
rect 229560 80112 229612 80121
rect 253940 80155 253992 80164
rect 253940 80121 253949 80155
rect 253949 80121 253983 80155
rect 253983 80121 253992 80155
rect 253940 80112 253992 80121
rect 256516 80044 256568 80096
rect 3240 79976 3292 80028
rect 215944 79976 215996 80028
rect 256608 79908 256660 79960
rect 248972 78455 249024 78464
rect 248972 78421 248981 78455
rect 248981 78421 249015 78455
rect 249015 78421 249024 78455
rect 248972 78412 249024 78421
rect 229468 77324 229520 77376
rect 243544 77299 243596 77308
rect 243544 77265 243553 77299
rect 243553 77265 243587 77299
rect 243587 77265 243596 77299
rect 243544 77256 243596 77265
rect 249156 77299 249208 77308
rect 249156 77265 249165 77299
rect 249165 77265 249199 77299
rect 249199 77265 249208 77299
rect 249156 77256 249208 77265
rect 229560 77231 229612 77240
rect 229560 77197 229569 77231
rect 229569 77197 229603 77231
rect 229603 77197 229612 77231
rect 229560 77188 229612 77197
rect 321468 76100 321520 76152
rect 323032 76100 323084 76152
rect 280252 76032 280304 76084
rect 289728 76032 289780 76084
rect 302148 76032 302200 76084
rect 309048 76032 309100 76084
rect 437388 76032 437440 76084
rect 444288 76032 444340 76084
rect 502248 76032 502300 76084
rect 510528 76032 510580 76084
rect 533988 76032 534040 76084
rect 540888 76032 540940 76084
rect 553308 76032 553360 76084
rect 560208 76032 560260 76084
rect 572628 76032 572680 76084
rect 579528 76032 579580 76084
rect 260380 75896 260432 75948
rect 253940 75871 253992 75880
rect 253940 75837 253949 75871
rect 253949 75837 253983 75871
rect 253983 75837 253992 75871
rect 253940 75828 253992 75837
rect 251824 74536 251876 74588
rect 259368 74536 259420 74588
rect 272340 74579 272392 74588
rect 272340 74545 272349 74579
rect 272349 74545 272383 74579
rect 272383 74545 272392 74579
rect 272340 74536 272392 74545
rect 238944 74511 238996 74520
rect 238944 74477 238953 74511
rect 238953 74477 238987 74511
rect 238987 74477 238996 74511
rect 238944 74468 238996 74477
rect 258632 74468 258684 74520
rect 237564 73219 237616 73228
rect 237564 73185 237573 73219
rect 237573 73185 237607 73219
rect 237607 73185 237616 73219
rect 237564 73176 237616 73185
rect 229652 67600 229704 67652
rect 278044 67600 278096 67652
rect 278136 67600 278188 67652
rect 240508 67575 240560 67584
rect 240508 67541 240517 67575
rect 240517 67541 240551 67575
rect 240551 67541 240560 67575
rect 240508 67532 240560 67541
rect 260104 67532 260156 67584
rect 260196 67396 260248 67448
rect 237564 66308 237616 66360
rect 251640 66240 251692 66292
rect 251824 66240 251876 66292
rect 256516 66240 256568 66292
rect 256608 66240 256660 66292
rect 259276 66240 259328 66292
rect 259368 66240 259420 66292
rect 237472 66172 237524 66224
rect 258540 64991 258592 65000
rect 258540 64957 258549 64991
rect 258549 64957 258583 64991
rect 258583 64957 258592 64991
rect 258540 64948 258592 64957
rect 238944 64923 238996 64932
rect 238944 64889 238953 64923
rect 238953 64889 238987 64923
rect 238987 64889 238996 64923
rect 238944 64880 238996 64889
rect 238208 64855 238260 64864
rect 238208 64821 238217 64855
rect 238217 64821 238251 64855
rect 238251 64821 238260 64855
rect 238208 64812 238260 64821
rect 241152 64855 241204 64864
rect 241152 64821 241161 64855
rect 241161 64821 241195 64855
rect 241195 64821 241204 64855
rect 241152 64812 241204 64821
rect 258540 64812 258592 64864
rect 258632 64812 258684 64864
rect 272432 64812 272484 64864
rect 294604 64812 294656 64864
rect 579804 64812 579856 64864
rect 272340 64744 272392 64796
rect 258632 63495 258684 63504
rect 258632 63461 258641 63495
rect 258641 63461 258675 63495
rect 258675 63461 258684 63495
rect 258632 63452 258684 63461
rect 240508 57987 240560 57996
rect 240508 57953 240517 57987
rect 240517 57953 240551 57987
rect 240551 57953 240560 57987
rect 240508 57944 240560 57953
rect 260288 57944 260340 57996
rect 260380 57944 260432 57996
rect 229652 57876 229704 57928
rect 256516 56584 256568 56636
rect 256608 56584 256660 56636
rect 275284 56559 275336 56568
rect 275284 56525 275293 56559
rect 275293 56525 275327 56559
rect 275327 56525 275336 56559
rect 275284 56516 275336 56525
rect 238208 55267 238260 55276
rect 238208 55233 238217 55267
rect 238217 55233 238251 55267
rect 238251 55233 238260 55267
rect 238208 55224 238260 55233
rect 241152 55267 241204 55276
rect 241152 55233 241161 55267
rect 241161 55233 241195 55267
rect 241195 55233 241204 55267
rect 241152 55224 241204 55233
rect 238944 55199 238996 55208
rect 238944 55165 238953 55199
rect 238953 55165 238987 55199
rect 238987 55165 238996 55199
rect 238944 55156 238996 55165
rect 243452 51144 243504 51196
rect 230848 51076 230900 51128
rect 231032 51076 231084 51128
rect 238208 51119 238260 51128
rect 238208 51085 238217 51119
rect 238217 51085 238251 51119
rect 238251 51085 238260 51119
rect 238208 51076 238260 51085
rect 241152 51076 241204 51128
rect 3056 51008 3108 51060
rect 225604 51008 225656 51060
rect 243452 51008 243504 51060
rect 275284 51051 275336 51060
rect 275284 51017 275293 51051
rect 275293 51017 275327 51051
rect 275327 51017 275336 51051
rect 275284 51008 275336 51017
rect 278044 51008 278096 51060
rect 278228 51008 278280 51060
rect 241244 50940 241296 50992
rect 260196 48356 260248 48408
rect 260380 48356 260432 48408
rect 229560 48331 229612 48340
rect 229560 48297 229569 48331
rect 229569 48297 229603 48331
rect 229603 48297 229612 48331
rect 229560 48288 229612 48297
rect 251548 48288 251600 48340
rect 251640 48288 251692 48340
rect 243544 48220 243596 48272
rect 237472 46928 237524 46980
rect 237564 46928 237616 46980
rect 238208 46971 238260 46980
rect 238208 46937 238217 46971
rect 238217 46937 238251 46971
rect 238251 46937 238260 46971
rect 238208 46928 238260 46937
rect 260104 46971 260156 46980
rect 260104 46937 260113 46971
rect 260113 46937 260147 46971
rect 260147 46937 260156 46971
rect 260104 46928 260156 46937
rect 260288 46971 260340 46980
rect 260288 46937 260297 46971
rect 260297 46937 260331 46971
rect 260331 46937 260340 46971
rect 260288 46928 260340 46937
rect 278228 46860 278280 46912
rect 238944 45611 238996 45620
rect 238944 45577 238953 45611
rect 238953 45577 238987 45611
rect 238987 45577 238996 45611
rect 258632 45611 258684 45620
rect 238944 45568 238996 45577
rect 258632 45577 258641 45611
rect 258641 45577 258675 45611
rect 258675 45577 258684 45611
rect 258632 45568 258684 45577
rect 237564 45543 237616 45552
rect 237564 45509 237573 45543
rect 237573 45509 237607 45543
rect 237607 45509 237616 45543
rect 237564 45500 237616 45509
rect 238208 45500 238260 45552
rect 241244 45543 241296 45552
rect 241244 45509 241253 45543
rect 241253 45509 241287 45543
rect 241287 45509 241296 45543
rect 241244 45500 241296 45509
rect 251548 44956 251600 45008
rect 251732 44956 251784 45008
rect 253940 43460 253992 43512
rect 254124 43460 254176 43512
rect 259276 43460 259328 43512
rect 259460 43460 259512 43512
rect 229468 41352 229520 41404
rect 229652 41352 229704 41404
rect 230848 41352 230900 41404
rect 231032 41352 231084 41404
rect 304264 41352 304316 41404
rect 580172 41352 580224 41404
rect 238944 38632 238996 38684
rect 249156 38632 249208 38684
rect 249248 38632 249300 38684
rect 229652 38564 229704 38616
rect 238852 38564 238904 38616
rect 278044 37315 278096 37324
rect 278044 37281 278053 37315
rect 278053 37281 278087 37315
rect 278087 37281 278096 37315
rect 278044 37272 278096 37281
rect 256608 37204 256660 37256
rect 256700 37204 256752 37256
rect 238208 35980 238260 36032
rect 237656 35912 237708 35964
rect 241244 35955 241296 35964
rect 241244 35921 241253 35955
rect 241253 35921 241287 35955
rect 241287 35921 241296 35955
rect 241244 35912 241296 35921
rect 3516 35844 3568 35896
rect 214564 35844 214616 35896
rect 238208 35844 238260 35896
rect 256700 35844 256752 35896
rect 259460 35844 259512 35896
rect 230848 31764 230900 31816
rect 231032 31764 231084 31816
rect 321468 29180 321520 29232
rect 321652 29180 321704 29232
rect 302148 29112 302200 29164
rect 308956 29112 309008 29164
rect 437388 29112 437440 29164
rect 444196 29112 444248 29164
rect 514668 29112 514720 29164
rect 521476 29112 521528 29164
rect 533988 29112 534040 29164
rect 540796 29112 540848 29164
rect 553308 29112 553360 29164
rect 560116 29112 560168 29164
rect 572628 29112 572680 29164
rect 579436 29112 579488 29164
rect 229560 29019 229612 29028
rect 229560 28985 229569 29019
rect 229569 28985 229603 29019
rect 229603 28985 229612 29019
rect 229560 28976 229612 28985
rect 238852 28976 238904 29028
rect 238944 28976 238996 29028
rect 254124 29044 254176 29096
rect 253940 28908 253992 28960
rect 243544 27616 243596 27668
rect 274916 27548 274968 27600
rect 275376 27548 275428 27600
rect 243544 27480 243596 27532
rect 278044 27480 278096 27532
rect 238116 26299 238168 26308
rect 238116 26265 238125 26299
rect 238125 26265 238159 26299
rect 238159 26265 238168 26299
rect 238116 26256 238168 26265
rect 256608 26299 256660 26308
rect 256608 26265 256617 26299
rect 256617 26265 256651 26299
rect 256651 26265 256660 26299
rect 256608 26256 256660 26265
rect 259276 26299 259328 26308
rect 259276 26265 259285 26299
rect 259285 26265 259319 26299
rect 259319 26265 259328 26299
rect 259276 26256 259328 26265
rect 274916 26231 274968 26240
rect 274916 26197 274925 26231
rect 274925 26197 274959 26231
rect 274959 26197 274968 26231
rect 274916 26188 274968 26197
rect 287612 22720 287664 22772
rect 567200 22720 567252 22772
rect 229560 22108 229612 22160
rect 230848 22040 230900 22092
rect 231032 22040 231084 22092
rect 243452 22083 243504 22092
rect 243452 22049 243461 22083
rect 243461 22049 243495 22083
rect 243495 22049 243504 22083
rect 243452 22040 243504 22049
rect 229560 21972 229612 22024
rect 238944 21428 238996 21480
rect 320824 21360 320876 21412
rect 543740 21360 543792 21412
rect 294696 19932 294748 19984
rect 532700 19932 532752 19984
rect 260104 19456 260156 19508
rect 260012 19388 260064 19440
rect 237564 19320 237616 19372
rect 237656 19320 237708 19372
rect 260104 19320 260156 19372
rect 260288 19320 260340 19372
rect 260012 19252 260064 19304
rect 276480 19295 276532 19304
rect 276480 19261 276489 19295
rect 276489 19261 276523 19295
rect 276523 19261 276532 19295
rect 276480 19252 276532 19261
rect 297364 18572 297416 18624
rect 525800 18572 525852 18624
rect 253940 18071 253992 18080
rect 253940 18037 253949 18071
rect 253949 18037 253983 18071
rect 253983 18037 253992 18071
rect 253940 18028 253992 18037
rect 240876 17960 240928 18012
rect 241060 17960 241112 18012
rect 251640 17960 251692 18012
rect 251732 17960 251784 18012
rect 258540 17960 258592 18012
rect 258632 17960 258684 18012
rect 259920 18003 259972 18012
rect 259920 17969 259929 18003
rect 259929 17969 259963 18003
rect 259963 17969 259972 18003
rect 259920 17960 259972 17969
rect 229100 17892 229152 17944
rect 579804 17892 579856 17944
rect 259920 17824 259972 17876
rect 260104 17824 260156 17876
rect 260380 17824 260432 17876
rect 256516 16668 256568 16720
rect 238852 16643 238904 16652
rect 238852 16609 238861 16643
rect 238861 16609 238895 16643
rect 238895 16609 238904 16643
rect 238852 16600 238904 16609
rect 253940 16643 253992 16652
rect 253940 16609 253949 16643
rect 253949 16609 253983 16643
rect 253983 16609 253992 16643
rect 253940 16600 253992 16609
rect 256608 16600 256660 16652
rect 274916 16643 274968 16652
rect 274916 16609 274925 16643
rect 274925 16609 274959 16643
rect 274959 16609 274968 16643
rect 274916 16600 274968 16609
rect 237564 16575 237616 16584
rect 237564 16541 237573 16575
rect 237573 16541 237607 16575
rect 237607 16541 237616 16575
rect 237564 16532 237616 16541
rect 151636 15852 151688 15904
rect 245200 15852 245252 15904
rect 290464 15852 290516 15904
rect 514760 15852 514812 15904
rect 164148 14424 164200 14476
rect 228364 14424 228416 14476
rect 298744 14424 298796 14476
rect 512092 14424 512144 14476
rect 148968 13064 149020 13116
rect 225696 13064 225748 13116
rect 291844 13064 291896 13116
rect 507860 13064 507912 13116
rect 230848 12452 230900 12504
rect 231032 12452 231084 12504
rect 243452 12452 243504 12504
rect 243360 12384 243412 12436
rect 166908 11704 166960 11756
rect 226984 11704 227036 11756
rect 228916 11704 228968 11756
rect 252008 11704 252060 11756
rect 301504 11704 301556 11756
rect 503720 11704 503772 11756
rect 266544 10956 266596 11008
rect 356152 10956 356204 11008
rect 267372 10888 267424 10940
rect 358820 10888 358872 10940
rect 267280 10820 267332 10872
rect 362960 10820 363012 10872
rect 266360 10752 266412 10804
rect 365720 10752 365772 10804
rect 64788 10684 64840 10736
rect 236736 10684 236788 10736
rect 268476 10684 268528 10736
rect 369860 10684 369912 10736
rect 60648 10616 60700 10668
rect 236828 10616 236880 10668
rect 268568 10616 268620 10668
rect 374092 10616 374144 10668
rect 30288 10548 30340 10600
rect 232228 10548 232280 10600
rect 268752 10548 268804 10600
rect 376760 10548 376812 10600
rect 27528 10480 27580 10532
rect 232136 10480 232188 10532
rect 269120 10480 269172 10532
rect 380900 10480 380952 10532
rect 22008 10412 22060 10464
rect 232044 10412 232096 10464
rect 236000 10412 236052 10464
rect 253204 10412 253256 10464
rect 269948 10412 270000 10464
rect 383660 10412 383712 10464
rect 9588 10344 9640 10396
rect 230940 10344 230992 10396
rect 233148 10344 233200 10396
rect 252928 10344 252980 10396
rect 269304 10344 269356 10396
rect 387800 10344 387852 10396
rect 3976 10276 4028 10328
rect 229560 10276 229612 10328
rect 231768 10276 231820 10328
rect 251916 10276 251968 10328
rect 270040 10276 270092 10328
rect 390560 10276 390612 10328
rect 265624 10208 265676 10260
rect 351920 10208 351972 10260
rect 265716 10140 265768 10192
rect 347780 10140 347832 10192
rect 265900 10072 265952 10124
rect 345020 10072 345072 10124
rect 265072 10004 265124 10056
rect 340880 10004 340932 10056
rect 276480 9707 276532 9716
rect 276480 9673 276489 9707
rect 276489 9673 276523 9707
rect 276523 9673 276532 9707
rect 276480 9664 276532 9673
rect 278228 9707 278280 9716
rect 278228 9673 278237 9707
rect 278237 9673 278271 9707
rect 278271 9673 278280 9707
rect 278228 9664 278280 9673
rect 90916 9596 90968 9648
rect 239312 9596 239364 9648
rect 87328 9528 87380 9580
rect 239036 9528 239088 9580
rect 274916 9528 274968 9580
rect 275376 9528 275428 9580
rect 83832 9460 83884 9512
rect 238576 9460 238628 9512
rect 80244 9392 80296 9444
rect 237748 9392 237800 9444
rect 76656 9324 76708 9376
rect 237840 9324 237892 9376
rect 73068 9256 73120 9308
rect 260472 9256 260524 9308
rect 291936 9256 291988 9308
rect 69480 9188 69532 9240
rect 237104 9188 237156 9240
rect 260012 9188 260064 9240
rect 295524 9188 295576 9240
rect 65984 9120 66036 9172
rect 236368 9120 236420 9172
rect 259828 9120 259880 9172
rect 299112 9120 299164 9172
rect 62396 9052 62448 9104
rect 236644 9052 236696 9104
rect 261392 9052 261444 9104
rect 306196 9052 306248 9104
rect 58808 8984 58860 9036
rect 236460 8984 236512 9036
rect 261300 8984 261352 9036
rect 309784 8984 309836 9036
rect 17316 8916 17368 8968
rect 231676 8916 231728 8968
rect 241980 8916 242032 8968
rect 251640 8916 251692 8968
rect 261208 8916 261260 8968
rect 302608 8916 302660 8968
rect 302884 8916 302936 8968
rect 494152 8916 494204 8968
rect 94504 8848 94556 8900
rect 239220 8848 239272 8900
rect 98092 8780 98144 8832
rect 240048 8780 240100 8832
rect 101588 8712 101640 8764
rect 240508 8712 240560 8764
rect 105176 8644 105228 8696
rect 240416 8644 240468 8696
rect 108764 8576 108816 8628
rect 240324 8576 240376 8628
rect 112352 8508 112404 8560
rect 241888 8508 241940 8560
rect 115940 8440 115992 8492
rect 241796 8440 241848 8492
rect 119436 8372 119488 8424
rect 242256 8372 242308 8424
rect 123024 8304 123076 8356
rect 242624 8304 242676 8356
rect 260196 8347 260248 8356
rect 260196 8313 260205 8347
rect 260205 8313 260239 8347
rect 260239 8313 260248 8347
rect 260196 8304 260248 8313
rect 3424 8236 3476 8288
rect 13084 8236 13136 8288
rect 200396 8236 200448 8288
rect 250536 8236 250588 8288
rect 256516 8236 256568 8288
rect 257436 8236 257488 8288
rect 261484 8236 261536 8288
rect 267004 8236 267056 8288
rect 275376 8279 275428 8288
rect 275376 8245 275385 8279
rect 275385 8245 275419 8279
rect 275419 8245 275428 8279
rect 275376 8236 275428 8245
rect 196808 8168 196860 8220
rect 250720 8168 250772 8220
rect 193220 8100 193272 8152
rect 250076 8100 250128 8152
rect 189632 8032 189684 8084
rect 249064 8032 249116 8084
rect 279792 8032 279844 8084
rect 279976 8032 280028 8084
rect 186044 7964 186096 8016
rect 248972 7964 249024 8016
rect 182548 7896 182600 7948
rect 249156 7896 249208 7948
rect 178960 7828 179012 7880
rect 248328 7828 248380 7880
rect 175372 7760 175424 7812
rect 247960 7760 248012 7812
rect 171784 7692 171836 7744
rect 247408 7692 247460 7744
rect 168196 7624 168248 7676
rect 247316 7624 247368 7676
rect 132592 7556 132644 7608
rect 243360 7556 243412 7608
rect 270500 7556 270552 7608
rect 271696 7556 271748 7608
rect 280804 7556 280856 7608
rect 314568 7556 314620 7608
rect 319444 7556 319496 7608
rect 490564 7556 490616 7608
rect 203892 7488 203944 7540
rect 250904 7488 250956 7540
rect 262956 6876 263008 6928
rect 268108 6876 268160 6928
rect 283564 6876 283616 6928
rect 288348 6876 288400 6928
rect 199200 6808 199252 6860
rect 249800 6808 249852 6860
rect 266452 6808 266504 6860
rect 354956 6808 355008 6860
rect 195612 6740 195664 6792
rect 250352 6740 250404 6792
rect 266820 6740 266872 6792
rect 358544 6740 358596 6792
rect 192024 6672 192076 6724
rect 248880 6672 248932 6724
rect 266728 6672 266780 6724
rect 362132 6672 362184 6724
rect 188436 6604 188488 6656
rect 248788 6604 248840 6656
rect 267464 6604 267516 6656
rect 365812 6604 365864 6656
rect 184848 6536 184900 6588
rect 248696 6536 248748 6588
rect 269028 6536 269080 6588
rect 369216 6536 369268 6588
rect 181352 6468 181404 6520
rect 248604 6468 248656 6520
rect 268844 6468 268896 6520
rect 372804 6468 372856 6520
rect 177764 6400 177816 6452
rect 248144 6400 248196 6452
rect 267924 6400 267976 6452
rect 376392 6400 376444 6452
rect 174176 6332 174228 6384
rect 247868 6332 247920 6384
rect 268200 6332 268252 6384
rect 379980 6332 380032 6384
rect 134892 6264 134944 6316
rect 243268 6264 243320 6316
rect 270132 6264 270184 6316
rect 383568 6264 383620 6316
rect 131396 6196 131448 6248
rect 243176 6196 243228 6248
rect 269488 6196 269540 6248
rect 387064 6196 387116 6248
rect 12440 6128 12492 6180
rect 230848 6128 230900 6180
rect 234804 6128 234856 6180
rect 254492 6128 254544 6180
rect 270224 6128 270276 6180
rect 390652 6128 390704 6180
rect 202696 6060 202748 6112
rect 250812 6060 250864 6112
rect 265348 6060 265400 6112
rect 351368 6060 351420 6112
rect 238392 5992 238444 6044
rect 254584 5992 254636 6044
rect 266084 5992 266136 6044
rect 347872 5992 347924 6044
rect 265532 5924 265584 5976
rect 344284 5924 344336 5976
rect 265992 5856 266044 5908
rect 340696 5856 340748 5908
rect 264336 5788 264388 5840
rect 337108 5788 337160 5840
rect 264244 5720 264296 5772
rect 333612 5720 333664 5772
rect 264060 5652 264112 5704
rect 330024 5652 330076 5704
rect 262772 5584 262824 5636
rect 326436 5584 326488 5636
rect 262680 5516 262732 5568
rect 322848 5516 322900 5568
rect 198004 5448 198056 5500
rect 244372 5448 244424 5500
rect 247684 5448 247736 5500
rect 257712 5448 257764 5500
rect 270500 5448 270552 5500
rect 194416 5380 194468 5432
rect 249984 5380 250036 5432
rect 258172 5380 258224 5432
rect 274088 5380 274140 5432
rect 190828 5312 190880 5364
rect 248512 5312 248564 5364
rect 257528 5312 257580 5364
rect 272892 5312 272944 5364
rect 137284 5244 137336 5296
rect 140872 5176 140924 5228
rect 142068 5176 142120 5228
rect 187240 5244 187292 5296
rect 249616 5244 249668 5296
rect 259276 5244 259328 5296
rect 276480 5244 276532 5296
rect 244004 5176 244056 5228
rect 251088 5176 251140 5228
rect 258908 5176 258960 5228
rect 277676 5176 277728 5228
rect 133788 5108 133840 5160
rect 243728 5108 243780 5160
rect 258540 5108 258592 5160
rect 280068 5108 280120 5160
rect 130200 5040 130252 5092
rect 243636 5040 243688 5092
rect 258816 5040 258868 5092
rect 281264 5040 281316 5092
rect 7656 4972 7708 5024
rect 229192 4972 229244 5024
rect 258356 4972 258408 5024
rect 283656 4972 283708 5024
rect 2872 4904 2924 4956
rect 229376 4904 229428 4956
rect 240784 4904 240836 4956
rect 254308 4904 254360 4956
rect 258264 4904 258316 4956
rect 284760 4904 284812 4956
rect 1676 4836 1728 4888
rect 572 4768 624 4820
rect 237288 4836 237340 4888
rect 254216 4836 254268 4888
rect 260196 4836 260248 4888
rect 287152 4836 287204 4888
rect 229284 4768 229336 4820
rect 233700 4768 233752 4820
rect 254400 4768 254452 4820
rect 260104 4768 260156 4820
rect 290740 4768 290792 4820
rect 316684 4768 316736 4820
rect 486976 4768 487028 4820
rect 489184 4768 489236 4820
rect 497740 4768 497792 4820
rect 201500 4700 201552 4752
rect 249892 4700 249944 4752
rect 257068 4700 257120 4752
rect 269304 4700 269356 4752
rect 205088 4632 205140 4684
rect 250996 4632 251048 4684
rect 230756 4564 230808 4616
rect 124220 4156 124272 4208
rect 125416 4156 125468 4208
rect 150440 4156 150492 4208
rect 151636 4156 151688 4208
rect 158720 4156 158772 4208
rect 160008 4156 160060 4208
rect 167092 4156 167144 4208
rect 168288 4156 168340 4208
rect 209872 4156 209924 4208
rect 211068 4156 211120 4208
rect 227720 4156 227772 4208
rect 229008 4156 229060 4208
rect 272524 4156 272576 4208
rect 275284 4156 275336 4208
rect 296720 4156 296772 4208
rect 297916 4156 297968 4208
rect 347780 4156 347832 4208
rect 349068 4156 349120 4208
rect 356060 4156 356112 4208
rect 357348 4156 357400 4208
rect 365720 4156 365772 4208
rect 366916 4156 366968 4208
rect 374000 4156 374052 4208
rect 375196 4156 375248 4208
rect 20720 4088 20772 4140
rect 28264 4088 28316 4140
rect 79048 4088 79100 4140
rect 238024 4088 238076 4140
rect 255504 4088 255556 4140
rect 256240 4088 256292 4140
rect 258448 4088 258500 4140
rect 259828 4088 259880 4140
rect 262864 4088 262916 4140
rect 264612 4088 264664 4140
rect 273904 4088 273956 4140
rect 425060 4088 425112 4140
rect 556804 4088 556856 4140
rect 559564 4088 559616 4140
rect 13636 4020 13688 4072
rect 17224 4020 17276 4072
rect 84108 4020 84160 4072
rect 235816 4020 235868 4072
rect 255044 4020 255096 4072
rect 255872 4020 255924 4072
rect 257344 4020 257396 4072
rect 258632 4020 258684 4072
rect 273720 4020 273772 4072
rect 428740 4020 428792 4072
rect 71872 3952 71924 4004
rect 237012 3952 237064 4004
rect 257804 3952 257856 4004
rect 261024 3952 261076 4004
rect 273444 3952 273496 4004
rect 432328 3952 432380 4004
rect 439412 3952 439464 4004
rect 68284 3884 68336 3936
rect 236276 3884 236328 3936
rect 254952 3884 255004 3936
rect 257988 3884 258040 3936
rect 262220 3884 262272 3936
rect 275744 3884 275796 3936
rect 435824 3884 435876 3936
rect 64696 3816 64748 3868
rect 236184 3816 236236 3868
rect 246764 3816 246816 3868
rect 255320 3816 255372 3868
rect 257896 3816 257948 3868
rect 263416 3816 263468 3868
rect 275100 3816 275152 3868
rect 433432 3816 433484 3868
rect 434628 3816 434680 3868
rect 61200 3748 61252 3800
rect 236092 3748 236144 3800
rect 275008 3748 275060 3800
rect 443000 3748 443052 3800
rect 567844 3748 567896 3800
rect 573824 3748 573876 3800
rect 44548 3680 44600 3732
rect 46204 3680 46256 3732
rect 57612 3680 57664 3732
rect 241060 3680 241112 3732
rect 247960 3680 248012 3732
rect 254676 3680 254728 3732
rect 446588 3680 446640 3732
rect 573364 3680 573416 3732
rect 579804 3680 579856 3732
rect 46940 3612 46992 3664
rect 34980 3544 35032 3596
rect 8852 3476 8904 3528
rect 9588 3476 9640 3528
rect 10048 3476 10100 3528
rect 14464 3476 14516 3528
rect 18328 3476 18380 3528
rect 19984 3476 20036 3528
rect 23112 3476 23164 3528
rect 24124 3476 24176 3528
rect 26700 3476 26752 3528
rect 27528 3476 27580 3528
rect 5264 3408 5316 3460
rect 10324 3408 10376 3460
rect 19524 3408 19576 3460
rect 32404 3476 32456 3528
rect 33876 3476 33928 3528
rect 34428 3476 34480 3528
rect 37372 3544 37424 3596
rect 38568 3544 38620 3596
rect 43444 3544 43496 3596
rect 50528 3544 50580 3596
rect 50988 3544 51040 3596
rect 51632 3544 51684 3596
rect 52368 3544 52420 3596
rect 52828 3544 52880 3596
rect 53748 3544 53800 3596
rect 54024 3612 54076 3664
rect 235172 3612 235224 3664
rect 245568 3612 245620 3664
rect 255136 3612 255188 3664
rect 277124 3612 277176 3664
rect 450176 3612 450228 3664
rect 502432 3612 502484 3664
rect 503628 3612 503680 3664
rect 536932 3612 536984 3664
rect 538128 3612 538180 3664
rect 546500 3612 546552 3664
rect 547696 3612 547748 3664
rect 563152 3612 563204 3664
rect 564348 3612 564400 3664
rect 565084 3612 565136 3664
rect 566740 3612 566792 3664
rect 573456 3612 573508 3664
rect 581000 3612 581052 3664
rect 40960 3476 41012 3528
rect 42064 3476 42116 3528
rect 42156 3476 42208 3528
rect 42708 3476 42760 3528
rect 43352 3476 43404 3528
rect 234068 3544 234120 3596
rect 231308 3476 231360 3528
rect 231768 3476 231820 3528
rect 232504 3476 232556 3528
rect 233148 3476 233200 3528
rect 233240 3476 233292 3528
rect 238116 3544 238168 3596
rect 252652 3544 252704 3596
rect 255780 3544 255832 3596
rect 276572 3544 276624 3596
rect 453672 3544 453724 3596
rect 482284 3544 482336 3596
rect 571340 3544 571392 3596
rect 572628 3544 572680 3596
rect 243176 3476 243228 3528
rect 29092 3408 29144 3460
rect 35164 3408 35216 3460
rect 39764 3408 39816 3460
rect 55220 3340 55272 3392
rect 56508 3340 56560 3392
rect 60004 3340 60056 3392
rect 60648 3340 60700 3392
rect 63592 3340 63644 3392
rect 64788 3340 64840 3392
rect 70676 3340 70728 3392
rect 71688 3340 71740 3392
rect 77852 3340 77904 3392
rect 78588 3340 78640 3392
rect 81440 3340 81492 3392
rect 82728 3340 82780 3392
rect 27896 3204 27948 3256
rect 31024 3204 31076 3256
rect 36176 3204 36228 3256
rect 39304 3204 39356 3256
rect 82636 3204 82688 3256
rect 230940 3340 230992 3392
rect 84936 3272 84988 3324
rect 85488 3272 85540 3324
rect 86132 3204 86184 3256
rect 229100 3272 229152 3324
rect 238484 3408 238536 3460
rect 239588 3408 239640 3460
rect 253940 3476 253992 3528
rect 276388 3476 276440 3528
rect 457260 3476 457312 3528
rect 467840 3476 467892 3528
rect 469128 3476 469180 3528
rect 475384 3476 475436 3528
rect 253848 3408 253900 3460
rect 255688 3408 255740 3460
rect 276112 3408 276164 3460
rect 460848 3408 460900 3460
rect 471244 3408 471296 3460
rect 582196 3408 582248 3460
rect 234712 3340 234764 3392
rect 249156 3340 249208 3392
rect 255596 3340 255648 3392
rect 273812 3340 273864 3392
rect 421564 3340 421616 3392
rect 494060 3340 494112 3392
rect 495348 3340 495400 3392
rect 512000 3340 512052 3392
rect 513196 3340 513248 3392
rect 528560 3340 528612 3392
rect 529848 3340 529900 3392
rect 560944 3340 560996 3392
rect 561956 3340 562008 3392
rect 578608 3340 578660 3392
rect 234160 3272 234212 3324
rect 251456 3272 251508 3324
rect 254768 3272 254820 3324
rect 272984 3272 273036 3324
rect 417976 3272 418028 3324
rect 574836 3272 574888 3324
rect 577412 3272 577464 3324
rect 89720 3204 89772 3256
rect 75460 3136 75512 3188
rect 84108 3136 84160 3188
rect 88524 3136 88576 3188
rect 89628 3136 89680 3188
rect 93308 3136 93360 3188
rect 233792 3204 233844 3256
rect 238760 3204 238812 3256
rect 272340 3204 272392 3256
rect 414480 3204 414532 3256
rect 575020 3204 575072 3256
rect 95700 3068 95752 3120
rect 96528 3068 96580 3120
rect 102784 3068 102836 3120
rect 103428 3068 103480 3120
rect 106372 3068 106424 3120
rect 107476 3068 107528 3120
rect 238852 3136 238904 3188
rect 271972 3136 272024 3188
rect 410892 3136 410944 3188
rect 11244 3000 11296 3052
rect 15844 3000 15896 3052
rect 96896 3000 96948 3052
rect 239496 3068 239548 3120
rect 272248 3068 272300 3120
rect 407304 3068 407356 3120
rect 45744 2864 45796 2916
rect 50344 2864 50396 2916
rect 103980 2864 104032 2916
rect 113548 2932 113600 2984
rect 114468 2932 114520 2984
rect 111156 2864 111208 2916
rect 239864 3000 239916 3052
rect 271052 3000 271104 3052
rect 403716 3000 403768 3052
rect 574744 3000 574796 3052
rect 576216 3000 576268 3052
rect 240968 2932 241020 2984
rect 270684 2932 270736 2984
rect 400220 2932 400272 2984
rect 114744 2864 114796 2916
rect 115848 2864 115900 2916
rect 120632 2864 120684 2916
rect 121368 2864 121420 2916
rect 118240 2796 118292 2848
rect 242072 2864 242124 2916
rect 250352 2864 250404 2916
rect 256056 2864 256108 2916
rect 270960 2864 271012 2916
rect 396632 2864 396684 2916
rect 425152 2864 425204 2916
rect 426348 2864 426400 2916
rect 121828 2796 121880 2848
rect 242164 2796 242216 2848
rect 269580 2796 269632 2848
rect 390560 2796 390612 2848
rect 391848 2796 391900 2848
rect 393044 2796 393096 2848
rect 74264 552 74316 604
rect 74448 552 74500 604
rect 92112 552 92164 604
rect 92388 552 92440 604
rect 109960 552 110012 604
rect 110328 552 110380 604
rect 183744 552 183796 604
rect 184756 552 184808 604
rect 206284 552 206336 604
rect 206928 552 206980 604
rect 207480 552 207532 604
rect 208308 552 208360 604
rect 208676 552 208728 604
rect 209688 552 209740 604
rect 230112 552 230164 604
rect 230388 552 230440 604
rect 281540 552 281592 604
rect 282460 552 282512 604
rect 285680 552 285732 604
rect 285956 552 286008 604
rect 288440 552 288492 604
rect 289544 552 289596 604
rect 292580 552 292632 604
rect 293132 552 293184 604
rect 299480 552 299532 604
rect 300308 552 300360 604
rect 300860 552 300912 604
rect 301412 552 301464 604
rect 303620 552 303672 604
rect 303804 552 303856 604
rect 492680 552 492732 604
rect 492956 552 493008 604
rect 495440 552 495492 604
rect 496544 552 496596 604
rect 498200 552 498252 604
rect 498936 552 498988 604
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 8128 700534 8156 703520
rect 8116 700528 8168 700534
rect 8116 700470 8168 700476
rect 24320 699718 24348 703520
rect 40512 700398 40540 703520
rect 72988 700806 73016 703520
rect 72976 700800 73028 700806
rect 72976 700742 73028 700748
rect 40500 700392 40552 700398
rect 40500 700334 40552 700340
rect 41328 700392 41380 700398
rect 41328 700334 41380 700340
rect 24308 699712 24360 699718
rect 24308 699654 24360 699660
rect 24768 699712 24820 699718
rect 24768 699654 24820 699660
rect 3422 682272 3478 682281
rect 3422 682207 3478 682216
rect 3330 653576 3386 653585
rect 3330 653511 3386 653520
rect 3344 652798 3372 653511
rect 3332 652792 3384 652798
rect 3332 652734 3384 652740
rect 3054 596048 3110 596057
rect 3054 595983 3110 595992
rect 3068 594862 3096 595983
rect 3056 594856 3108 594862
rect 3056 594798 3108 594804
rect 2962 553072 3018 553081
rect 2962 553007 3018 553016
rect 2976 552090 3004 553007
rect 2964 552084 3016 552090
rect 2964 552026 3016 552032
rect 3146 538656 3202 538665
rect 3146 538591 3202 538600
rect 3160 538286 3188 538591
rect 3148 538280 3200 538286
rect 3148 538222 3200 538228
rect 3330 495544 3386 495553
rect 3330 495479 3332 495488
rect 3384 495479 3386 495488
rect 3332 495450 3384 495456
rect 3146 481128 3202 481137
rect 3146 481063 3202 481072
rect 3160 480282 3188 481063
rect 3148 480276 3200 480282
rect 3148 480218 3200 480224
rect 3238 452432 3294 452441
rect 3238 452367 3294 452376
rect 2962 438016 3018 438025
rect 2962 437951 3018 437960
rect 2976 437510 3004 437951
rect 2964 437504 3016 437510
rect 2964 437446 3016 437452
rect 3252 402286 3280 452367
rect 3330 423736 3386 423745
rect 3330 423671 3332 423680
rect 3384 423671 3386 423680
rect 3332 423642 3384 423648
rect 3436 402694 3464 682207
rect 3514 667992 3570 668001
rect 3514 667927 3570 667936
rect 3424 402688 3476 402694
rect 3424 402630 3476 402636
rect 3528 402558 3556 667927
rect 3606 624880 3662 624889
rect 3606 624815 3662 624824
rect 3620 402626 3648 624815
rect 3698 610464 3754 610473
rect 3698 610399 3754 610408
rect 3608 402620 3660 402626
rect 3608 402562 3660 402568
rect 3516 402552 3568 402558
rect 3516 402494 3568 402500
rect 3712 402422 3740 610399
rect 3882 567352 3938 567361
rect 3882 567287 3938 567296
rect 3896 402490 3924 567287
rect 4066 509960 4122 509969
rect 4066 509895 4122 509904
rect 3884 402484 3936 402490
rect 3884 402426 3936 402432
rect 3700 402416 3752 402422
rect 3700 402358 3752 402364
rect 4080 402354 4108 509895
rect 24780 402762 24808 699654
rect 41340 402830 41368 700334
rect 89180 699718 89208 703520
rect 105464 699718 105492 703520
rect 137848 700262 137876 703520
rect 137836 700256 137888 700262
rect 137836 700198 137888 700204
rect 89168 699712 89220 699718
rect 89168 699654 89220 699660
rect 89628 699712 89680 699718
rect 89628 699654 89680 699660
rect 105452 699712 105504 699718
rect 105452 699654 105504 699660
rect 106188 699712 106240 699718
rect 106188 699654 106240 699660
rect 89640 402898 89668 699654
rect 106200 403170 106228 699654
rect 154132 695570 154160 703520
rect 170324 699718 170352 703520
rect 202800 699990 202828 703520
rect 218992 703474 219020 703520
rect 218900 703446 219020 703474
rect 202788 699984 202840 699990
rect 202788 699926 202840 699932
rect 170312 699712 170364 699718
rect 170312 699654 170364 699660
rect 171048 699712 171100 699718
rect 171048 699654 171100 699660
rect 154120 695564 154172 695570
rect 154120 695506 154172 695512
rect 154212 695564 154264 695570
rect 154212 695506 154264 695512
rect 154224 688634 154252 695506
rect 154212 688628 154264 688634
rect 154212 688570 154264 688576
rect 154396 688628 154448 688634
rect 154396 688570 154448 688576
rect 154408 685846 154436 688570
rect 154396 685840 154448 685846
rect 154396 685782 154448 685788
rect 154304 676252 154356 676258
rect 154304 676194 154356 676200
rect 154316 673538 154344 676194
rect 154304 673532 154356 673538
rect 154304 673474 154356 673480
rect 154488 673532 154540 673538
rect 154488 673474 154540 673480
rect 154500 663762 154528 673474
rect 154316 663734 154528 663762
rect 154316 654158 154344 663734
rect 154304 654152 154356 654158
rect 154304 654094 154356 654100
rect 154488 654152 154540 654158
rect 154488 654094 154540 654100
rect 154500 644450 154528 654094
rect 154316 644422 154528 644450
rect 154316 634846 154344 644422
rect 154304 634840 154356 634846
rect 154304 634782 154356 634788
rect 154488 634840 154540 634846
rect 154488 634782 154540 634788
rect 154500 625138 154528 634782
rect 154316 625110 154528 625138
rect 154316 615534 154344 625110
rect 154304 615528 154356 615534
rect 154304 615470 154356 615476
rect 154488 615528 154540 615534
rect 154488 615470 154540 615476
rect 154500 605826 154528 615470
rect 154316 605798 154528 605826
rect 154316 596222 154344 605798
rect 154304 596216 154356 596222
rect 154488 596216 154540 596222
rect 154304 596158 154356 596164
rect 154408 596164 154488 596170
rect 154408 596158 154540 596164
rect 154408 596142 154528 596158
rect 154408 591954 154436 596142
rect 154316 591926 154436 591954
rect 154316 589286 154344 591926
rect 154304 589280 154356 589286
rect 154304 589222 154356 589228
rect 154304 579760 154356 579766
rect 154224 579708 154304 579714
rect 154224 579702 154356 579708
rect 154224 579686 154344 579702
rect 154224 579630 154252 579686
rect 154212 579624 154264 579630
rect 154212 579566 154264 579572
rect 154396 579624 154448 579630
rect 154396 579566 154448 579572
rect 154408 562970 154436 579566
rect 154212 562964 154264 562970
rect 154212 562906 154264 562912
rect 154396 562964 154448 562970
rect 154396 562906 154448 562912
rect 154224 553330 154252 562906
rect 154224 553302 154344 553330
rect 154316 543810 154344 553302
rect 154316 543782 154528 543810
rect 154500 534018 154528 543782
rect 154408 533990 154528 534018
rect 154408 531282 154436 533990
rect 154396 531276 154448 531282
rect 154396 531218 154448 531224
rect 154488 521688 154540 521694
rect 154488 521630 154540 521636
rect 154500 514706 154528 521630
rect 154408 514678 154528 514706
rect 154408 511970 154436 514678
rect 154396 511964 154448 511970
rect 154396 511906 154448 511912
rect 154488 502376 154540 502382
rect 154488 502318 154540 502324
rect 154500 495394 154528 502318
rect 154408 495366 154528 495394
rect 154408 492658 154436 495366
rect 154212 492652 154264 492658
rect 154212 492594 154264 492600
rect 154396 492652 154448 492658
rect 154396 492594 154448 492600
rect 154224 483041 154252 492594
rect 154210 483032 154266 483041
rect 154210 482967 154266 482976
rect 154486 483032 154542 483041
rect 154486 482967 154542 482976
rect 154500 476082 154528 482967
rect 154316 476054 154528 476082
rect 154316 466478 154344 476054
rect 154304 466472 154356 466478
rect 154304 466414 154356 466420
rect 154488 466472 154540 466478
rect 154488 466414 154540 466420
rect 154500 456770 154528 466414
rect 154316 456742 154528 456770
rect 154316 454034 154344 456742
rect 154304 454028 154356 454034
rect 154304 453970 154356 453976
rect 154212 444440 154264 444446
rect 154212 444382 154264 444388
rect 154224 437458 154252 444382
rect 154224 437430 154344 437458
rect 154316 427854 154344 437430
rect 154304 427848 154356 427854
rect 154304 427790 154356 427796
rect 154396 427780 154448 427786
rect 154396 427722 154448 427728
rect 154408 425066 154436 427722
rect 154120 425060 154172 425066
rect 154120 425002 154172 425008
rect 154396 425060 154448 425066
rect 154396 425002 154448 425008
rect 154132 415449 154160 425002
rect 154118 415440 154174 415449
rect 154118 415375 154174 415384
rect 154302 415440 154358 415449
rect 154302 415375 154358 415384
rect 154316 415313 154344 415375
rect 154302 415304 154358 415313
rect 154302 415239 154358 415248
rect 154486 415304 154542 415313
rect 154486 415239 154542 415248
rect 154500 408542 154528 415239
rect 154488 408536 154540 408542
rect 154488 408478 154540 408484
rect 154488 408400 154540 408406
rect 154488 408342 154540 408348
rect 106188 403164 106240 403170
rect 106188 403106 106240 403112
rect 89628 402892 89680 402898
rect 89628 402834 89680 402840
rect 41328 402824 41380 402830
rect 41328 402766 41380 402772
rect 24768 402756 24820 402762
rect 24768 402698 24820 402704
rect 4068 402348 4120 402354
rect 4068 402290 4120 402296
rect 3240 402280 3292 402286
rect 3240 402222 3292 402228
rect 154500 402218 154528 408342
rect 154488 402212 154540 402218
rect 154488 402154 154540 402160
rect 171060 402150 171088 699654
rect 218900 695745 218928 703446
rect 235184 699718 235212 703520
rect 257896 701004 257948 701010
rect 257896 700946 257948 700952
rect 256516 700732 256568 700738
rect 256516 700674 256568 700680
rect 256424 700596 256476 700602
rect 256424 700538 256476 700544
rect 255228 700460 255280 700466
rect 255228 700402 255280 700408
rect 255136 700392 255188 700398
rect 255136 700334 255188 700340
rect 253848 700324 253900 700330
rect 253848 700266 253900 700272
rect 235172 699712 235224 699718
rect 235172 699654 235224 699660
rect 235908 699712 235960 699718
rect 235908 699654 235960 699660
rect 218886 695736 218942 695745
rect 218886 695671 218942 695680
rect 219254 695600 219310 695609
rect 219176 695558 219254 695586
rect 219176 695502 219204 695558
rect 219254 695535 219310 695544
rect 219164 695496 219216 695502
rect 219164 695438 219216 695444
rect 219072 685908 219124 685914
rect 219072 685850 219124 685856
rect 219084 678994 219112 685850
rect 218992 678966 219112 678994
rect 218992 676190 219020 678966
rect 218980 676184 219032 676190
rect 218980 676126 219032 676132
rect 219072 666596 219124 666602
rect 219072 666538 219124 666544
rect 219084 659682 219112 666538
rect 219084 659666 219204 659682
rect 219084 659660 219216 659666
rect 219084 659654 219164 659660
rect 219164 659602 219216 659608
rect 219348 659660 219400 659666
rect 219348 659602 219400 659608
rect 219360 656878 219388 659602
rect 219348 656872 219400 656878
rect 219348 656814 219400 656820
rect 219256 647284 219308 647290
rect 219256 647226 219308 647232
rect 219268 640422 219296 647226
rect 219256 640416 219308 640422
rect 219256 640358 219308 640364
rect 219072 640280 219124 640286
rect 219072 640222 219124 640228
rect 219084 637566 219112 640222
rect 219072 637560 219124 637566
rect 219072 637502 219124 637508
rect 219164 637560 219216 637566
rect 219164 637502 219216 637508
rect 219176 630578 219204 637502
rect 219176 630550 219388 630578
rect 219360 626550 219388 630550
rect 219348 626544 219400 626550
rect 219348 626486 219400 626492
rect 219348 616888 219400 616894
rect 219348 616830 219400 616836
rect 219360 611454 219388 616830
rect 219348 611448 219400 611454
rect 219348 611390 219400 611396
rect 219072 608728 219124 608734
rect 219072 608670 219124 608676
rect 219084 608598 219112 608670
rect 219072 608592 219124 608598
rect 219072 608534 219124 608540
rect 219256 601588 219308 601594
rect 219256 601530 219308 601536
rect 219268 598942 219296 601530
rect 219256 598936 219308 598942
rect 219256 598878 219308 598884
rect 219164 589348 219216 589354
rect 219164 589290 219216 589296
rect 219176 582418 219204 589290
rect 218980 582412 219032 582418
rect 218980 582354 219032 582360
rect 219164 582412 219216 582418
rect 219164 582354 219216 582360
rect 218992 579630 219020 582354
rect 218980 579624 219032 579630
rect 218980 579566 219032 579572
rect 218888 569968 218940 569974
rect 218888 569910 218940 569916
rect 218900 563106 218928 569910
rect 218888 563100 218940 563106
rect 218888 563042 218940 563048
rect 218980 562964 219032 562970
rect 218980 562906 219032 562912
rect 218992 560266 219020 562906
rect 218900 560238 219020 560266
rect 218900 553450 218928 560238
rect 218888 553444 218940 553450
rect 218888 553386 218940 553392
rect 218888 550656 218940 550662
rect 218888 550598 218940 550604
rect 218900 543794 218928 550598
rect 218888 543788 218940 543794
rect 218888 543730 218940 543736
rect 218980 543652 219032 543658
rect 218980 543594 219032 543600
rect 218992 540977 219020 543594
rect 218978 540968 219034 540977
rect 218978 540903 219034 540912
rect 219162 540968 219218 540977
rect 219162 540903 219218 540912
rect 219176 533882 219204 540903
rect 218992 533854 219204 533882
rect 218992 531321 219020 533854
rect 218978 531312 219034 531321
rect 218978 531247 219034 531256
rect 219162 531312 219218 531321
rect 219162 531247 219218 531256
rect 219176 524346 219204 531247
rect 218980 524340 219032 524346
rect 218980 524282 219032 524288
rect 219164 524340 219216 524346
rect 219164 524282 219216 524288
rect 218992 521665 219020 524282
rect 218794 521656 218850 521665
rect 218794 521591 218850 521600
rect 218978 521656 219034 521665
rect 218978 521591 219034 521600
rect 218808 514690 218836 521591
rect 218796 514684 218848 514690
rect 218796 514626 218848 514632
rect 219072 514684 219124 514690
rect 219072 514626 219124 514632
rect 219084 510610 219112 514626
rect 219072 510604 219124 510610
rect 219072 510546 219124 510552
rect 219072 505096 219124 505102
rect 219072 505038 219124 505044
rect 219084 492726 219112 505038
rect 219072 492720 219124 492726
rect 219072 492662 219124 492668
rect 219164 492720 219216 492726
rect 219164 492662 219216 492668
rect 219176 485858 219204 492662
rect 219164 485852 219216 485858
rect 219164 485794 219216 485800
rect 219256 485716 219308 485722
rect 219256 485658 219308 485664
rect 219268 473385 219296 485658
rect 218978 473376 219034 473385
rect 218978 473311 219034 473320
rect 219254 473376 219310 473385
rect 219254 473311 219310 473320
rect 218992 466478 219020 473311
rect 218980 466472 219032 466478
rect 218980 466414 219032 466420
rect 219348 466336 219400 466342
rect 219348 466278 219400 466284
rect 219360 456770 219388 466278
rect 219084 456742 219388 456770
rect 219084 454034 219112 456742
rect 219072 454028 219124 454034
rect 219072 453970 219124 453976
rect 218980 444440 219032 444446
rect 218980 444382 219032 444388
rect 218992 437458 219020 444382
rect 218992 437430 219112 437458
rect 219084 434722 219112 437430
rect 218980 434716 219032 434722
rect 218980 434658 219032 434664
rect 219072 434716 219124 434722
rect 219072 434658 219124 434664
rect 218992 425105 219020 434658
rect 218978 425096 219034 425105
rect 218978 425031 219034 425040
rect 219346 425096 219402 425105
rect 219346 425031 219402 425040
rect 171048 402144 171100 402150
rect 171048 402086 171100 402092
rect 219360 402082 219388 425031
rect 219348 402076 219400 402082
rect 219348 402018 219400 402024
rect 235814 401976 235870 401985
rect 235920 401946 235948 699654
rect 253756 696992 253808 696998
rect 253756 696934 253808 696940
rect 253664 685908 253716 685914
rect 253664 685850 253716 685856
rect 252468 673532 252520 673538
rect 252468 673474 252520 673480
rect 252376 650072 252428 650078
rect 252376 650014 252428 650020
rect 252284 638988 252336 638994
rect 252284 638930 252336 638936
rect 251088 626612 251140 626618
rect 251088 626554 251140 626560
rect 249708 603152 249760 603158
rect 249708 603094 249760 603100
rect 249616 579692 249668 579698
rect 249616 579634 249668 579640
rect 248328 556232 248380 556238
rect 248328 556174 248380 556180
rect 248236 532772 248288 532778
rect 248236 532714 248288 532720
rect 246948 509312 247000 509318
rect 246948 509254 247000 509260
rect 246856 485852 246908 485858
rect 246856 485794 246908 485800
rect 245568 462392 245620 462398
rect 245568 462334 245620 462340
rect 245476 451308 245528 451314
rect 245476 451250 245528 451256
rect 245384 438932 245436 438938
rect 245384 438874 245436 438880
rect 244188 415472 244240 415478
rect 244188 415414 244240 415420
rect 243820 404388 243872 404394
rect 243820 404330 243872 404336
rect 242256 402008 242308 402014
rect 242256 401950 242308 401956
rect 235814 401911 235870 401920
rect 235908 401940 235960 401946
rect 3332 401804 3384 401810
rect 3332 401746 3384 401752
rect 3148 396024 3200 396030
rect 3148 395966 3200 395972
rect 3160 395049 3188 395966
rect 3146 395040 3202 395049
rect 3146 394975 3202 394984
rect 2964 367056 3016 367062
rect 2964 366998 3016 367004
rect 2976 366217 3004 366998
rect 2962 366208 3018 366217
rect 2962 366143 3018 366152
rect 3344 323105 3372 401746
rect 3976 401736 4028 401742
rect 3976 401678 4028 401684
rect 3792 401668 3844 401674
rect 3792 401610 3844 401616
rect 3424 399492 3476 399498
rect 3424 399434 3476 399440
rect 3436 380633 3464 399434
rect 3422 380624 3478 380633
rect 3422 380559 3478 380568
rect 3424 338088 3476 338094
rect 3424 338030 3476 338036
rect 3436 337521 3464 338030
rect 3422 337512 3478 337521
rect 3422 337447 3478 337456
rect 3422 336016 3478 336025
rect 3422 335951 3478 335960
rect 3330 323096 3386 323105
rect 3330 323031 3386 323040
rect 3332 309120 3384 309126
rect 3332 309062 3384 309068
rect 3344 308825 3372 309062
rect 3330 308816 3386 308825
rect 3330 308751 3386 308760
rect 3148 252544 3200 252550
rect 3148 252486 3200 252492
rect 3160 251297 3188 252486
rect 3146 251288 3202 251297
rect 3146 251223 3202 251232
rect 3148 223576 3200 223582
rect 3148 223518 3200 223524
rect 3160 222601 3188 223518
rect 3146 222592 3202 222601
rect 3146 222527 3202 222536
rect 3240 180804 3292 180810
rect 3240 180746 3292 180752
rect 3252 179489 3280 180746
rect 3238 179480 3294 179489
rect 3238 179415 3294 179424
rect 2964 122800 3016 122806
rect 2964 122742 3016 122748
rect 2976 122097 3004 122742
rect 2962 122088 3018 122097
rect 2962 122023 3018 122032
rect 3240 80028 3292 80034
rect 3240 79970 3292 79976
rect 3252 78985 3280 79970
rect 3238 78976 3294 78985
rect 3238 78911 3294 78920
rect 3056 51060 3108 51066
rect 3056 51002 3108 51008
rect 3068 50153 3096 51002
rect 3054 50144 3110 50153
rect 3054 50079 3110 50088
rect 3436 21457 3464 335951
rect 3516 295316 3568 295322
rect 3516 295258 3568 295264
rect 3528 294409 3556 295258
rect 3514 294400 3570 294409
rect 3514 294335 3570 294344
rect 3516 266348 3568 266354
rect 3516 266290 3568 266296
rect 3528 265713 3556 266290
rect 3514 265704 3570 265713
rect 3514 265639 3570 265648
rect 3804 237017 3832 401610
rect 3988 280129 4016 401678
rect 10968 401464 11020 401470
rect 10968 401406 11020 401412
rect 10980 396030 11008 401406
rect 14556 401396 14608 401402
rect 14556 401338 14608 401344
rect 13084 399220 13136 399226
rect 13084 399162 13136 399168
rect 10968 396024 11020 396030
rect 10968 395966 11020 395972
rect 10324 337408 10376 337414
rect 10324 337350 10376 337356
rect 3974 280120 4030 280129
rect 3974 280055 4030 280064
rect 3790 237008 3846 237017
rect 3790 236943 3846 236952
rect 3516 208344 3568 208350
rect 3516 208286 3568 208292
rect 3528 208185 3556 208286
rect 3514 208176 3570 208185
rect 3514 208111 3570 208120
rect 3514 194576 3570 194585
rect 3514 194511 3570 194520
rect 3528 193905 3556 194511
rect 3514 193896 3570 193905
rect 3514 193831 3570 193840
rect 3516 165572 3568 165578
rect 3516 165514 3568 165520
rect 3528 165073 3556 165514
rect 3514 165064 3570 165073
rect 3514 164999 3570 165008
rect 3514 151736 3570 151745
rect 3514 151671 3570 151680
rect 3528 150793 3556 151671
rect 3514 150784 3570 150793
rect 3514 150719 3570 150728
rect 3516 136604 3568 136610
rect 3516 136546 3568 136552
rect 3528 136377 3556 136546
rect 3514 136368 3570 136377
rect 3514 136303 3570 136312
rect 3514 109032 3570 109041
rect 3514 108967 3570 108976
rect 3528 107681 3556 108967
rect 3514 107672 3570 107681
rect 3514 107607 3570 107616
rect 3516 93832 3568 93838
rect 3516 93774 3568 93780
rect 3528 93265 3556 93774
rect 3514 93256 3570 93265
rect 3514 93191 3570 93200
rect 3516 35896 3568 35902
rect 3514 35864 3516 35873
rect 3568 35864 3570 35873
rect 3514 35799 3570 35808
rect 3422 21448 3478 21457
rect 3422 21383 3478 21392
rect 9588 10396 9640 10402
rect 9588 10338 9640 10344
rect 3976 10328 4028 10334
rect 3976 10270 4028 10276
rect 3424 8288 3476 8294
rect 3424 8230 3476 8236
rect 3436 7177 3464 8230
rect 3422 7168 3478 7177
rect 3422 7103 3478 7112
rect 2872 4956 2924 4962
rect 2872 4898 2924 4904
rect 1676 4888 1728 4894
rect 1676 4830 1728 4836
rect 572 4820 624 4826
rect 572 4762 624 4768
rect 584 480 612 4762
rect 1688 480 1716 4830
rect 2884 480 2912 4898
rect 3988 626 4016 10270
rect 7656 5024 7708 5030
rect 7656 4966 7708 4972
rect 5264 3460 5316 3466
rect 5264 3402 5316 3408
rect 3988 598 4108 626
rect 4080 480 4108 598
rect 5276 480 5304 3402
rect 6458 3360 6514 3369
rect 6458 3295 6514 3304
rect 6472 480 6500 3295
rect 7668 480 7696 4966
rect 9600 3534 9628 10338
rect 8852 3528 8904 3534
rect 8852 3470 8904 3476
rect 9588 3528 9640 3534
rect 9588 3470 9640 3476
rect 10048 3528 10100 3534
rect 10048 3470 10100 3476
rect 8864 480 8892 3470
rect 10060 480 10088 3470
rect 10336 3466 10364 337350
rect 13096 8294 13124 399162
rect 14568 338094 14596 401338
rect 227168 401328 227220 401334
rect 227168 401270 227220 401276
rect 225788 401260 225840 401266
rect 225788 401202 225840 401208
rect 222844 401056 222896 401062
rect 222844 400998 222896 401004
rect 211804 400716 211856 400722
rect 211804 400658 211856 400664
rect 209044 400580 209096 400586
rect 209044 400522 209096 400528
rect 207664 399560 207716 399566
rect 207664 399502 207716 399508
rect 204904 399424 204956 399430
rect 204904 399366 204956 399372
rect 180064 399356 180116 399362
rect 180064 399298 180116 399304
rect 14556 338088 14608 338094
rect 14556 338030 14608 338036
rect 125508 338088 125560 338094
rect 125508 338030 125560 338036
rect 107568 338020 107620 338026
rect 107568 337962 107620 337968
rect 100668 337884 100720 337890
rect 100668 337826 100720 337832
rect 39304 337816 39356 337822
rect 39304 337758 39356 337764
rect 32404 337748 32456 337754
rect 32404 337690 32456 337696
rect 28264 337612 28316 337618
rect 28264 337554 28316 337560
rect 15844 337544 15896 337550
rect 15844 337486 15896 337492
rect 14464 337476 14516 337482
rect 14464 337418 14516 337424
rect 13084 8288 13136 8294
rect 13084 8230 13136 8236
rect 12440 6180 12492 6186
rect 12440 6122 12492 6128
rect 10324 3460 10376 3466
rect 10324 3402 10376 3408
rect 11244 3052 11296 3058
rect 11244 2994 11296 3000
rect 11256 480 11284 2994
rect 12452 480 12480 6122
rect 13636 4072 13688 4078
rect 13636 4014 13688 4020
rect 13648 480 13676 4014
rect 14476 3534 14504 337418
rect 14464 3528 14516 3534
rect 14464 3470 14516 3476
rect 14830 3496 14886 3505
rect 14830 3431 14886 3440
rect 14844 480 14872 3431
rect 15856 3058 15884 337486
rect 17224 331900 17276 331906
rect 17224 331842 17276 331848
rect 17236 4078 17264 331842
rect 19984 315308 20036 315314
rect 19984 315250 20036 315256
rect 17316 8968 17368 8974
rect 17316 8910 17368 8916
rect 17224 4072 17276 4078
rect 17224 4014 17276 4020
rect 16026 3632 16082 3641
rect 16026 3567 16082 3576
rect 15844 3052 15896 3058
rect 15844 2994 15896 3000
rect 16040 480 16068 3567
rect 17328 1442 17356 8910
rect 19996 3534 20024 315250
rect 24124 313948 24176 313954
rect 24124 313890 24176 313896
rect 22008 10464 22060 10470
rect 22008 10406 22060 10412
rect 20720 4140 20772 4146
rect 20720 4082 20772 4088
rect 18328 3528 18380 3534
rect 18328 3470 18380 3476
rect 19984 3528 20036 3534
rect 19984 3470 20036 3476
rect 17236 1414 17356 1442
rect 17236 480 17264 1414
rect 18340 480 18368 3470
rect 19524 3460 19576 3466
rect 19524 3402 19576 3408
rect 19536 480 19564 3402
rect 20732 480 20760 4082
rect 22020 3482 22048 10406
rect 24136 3534 24164 313890
rect 27528 10532 27580 10538
rect 27528 10474 27580 10480
rect 25502 3904 25558 3913
rect 25502 3839 25558 3848
rect 24306 3768 24362 3777
rect 24306 3703 24362 3712
rect 21928 3454 22048 3482
rect 23112 3528 23164 3534
rect 23112 3470 23164 3476
rect 24124 3528 24176 3534
rect 24124 3470 24176 3476
rect 21928 480 21956 3454
rect 23124 480 23152 3470
rect 24320 480 24348 3703
rect 25516 480 25544 3839
rect 27540 3534 27568 10474
rect 28276 4146 28304 337554
rect 31668 312588 31720 312594
rect 31668 312530 31720 312536
rect 31024 309800 31076 309806
rect 31024 309742 31076 309748
rect 30288 10600 30340 10606
rect 30288 10542 30340 10548
rect 28264 4140 28316 4146
rect 28264 4082 28316 4088
rect 26700 3528 26752 3534
rect 26700 3470 26752 3476
rect 27528 3528 27580 3534
rect 27528 3470 27580 3476
rect 26712 480 26740 3470
rect 29092 3460 29144 3466
rect 29092 3402 29144 3408
rect 27896 3256 27948 3262
rect 27896 3198 27948 3204
rect 27908 480 27936 3198
rect 29104 480 29132 3402
rect 30300 480 30328 10542
rect 31036 3262 31064 309742
rect 31680 3482 31708 312530
rect 32416 3534 32444 337690
rect 35164 337680 35216 337686
rect 35164 337622 35216 337628
rect 34428 329112 34480 329118
rect 34428 329054 34480 329060
rect 32678 4040 32734 4049
rect 32678 3975 32734 3984
rect 31496 3454 31708 3482
rect 32404 3528 32456 3534
rect 32404 3470 32456 3476
rect 31024 3256 31076 3262
rect 31024 3198 31076 3204
rect 31496 480 31524 3454
rect 32692 480 32720 3975
rect 34440 3534 34468 329054
rect 34980 3596 35032 3602
rect 34980 3538 35032 3544
rect 33876 3528 33928 3534
rect 33876 3470 33928 3476
rect 34428 3528 34480 3534
rect 34428 3470 34480 3476
rect 33888 480 33916 3470
rect 34992 480 35020 3538
rect 35176 3466 35204 337622
rect 38568 327752 38620 327758
rect 38568 327694 38620 327700
rect 38476 305652 38528 305658
rect 38476 305594 38528 305600
rect 37372 3596 37424 3602
rect 37372 3538 37424 3544
rect 35164 3460 35216 3466
rect 35164 3402 35216 3408
rect 36176 3256 36228 3262
rect 36176 3198 36228 3204
rect 36188 480 36216 3198
rect 37384 480 37412 3538
rect 38488 3482 38516 305594
rect 38580 3602 38608 327694
rect 38568 3596 38620 3602
rect 38568 3538 38620 3544
rect 38488 3454 38608 3482
rect 38580 480 38608 3454
rect 39316 3262 39344 337758
rect 52368 336048 52420 336054
rect 52368 335990 52420 335996
rect 89628 336048 89680 336054
rect 89628 335990 89680 335996
rect 49608 333260 49660 333266
rect 49608 333202 49660 333208
rect 48228 331968 48280 331974
rect 48228 331910 48280 331916
rect 42064 324964 42116 324970
rect 42064 324906 42116 324912
rect 42076 3534 42104 324906
rect 46204 323604 46256 323610
rect 46204 323546 46256 323552
rect 43444 307080 43496 307086
rect 43444 307022 43496 307028
rect 42708 304292 42760 304298
rect 42708 304234 42760 304240
rect 42720 3534 42748 304234
rect 43456 3602 43484 307022
rect 46216 3738 46244 323546
rect 44548 3732 44600 3738
rect 44548 3674 44600 3680
rect 46204 3732 46256 3738
rect 46204 3674 46256 3680
rect 43444 3596 43496 3602
rect 43444 3538 43496 3544
rect 40960 3528 41012 3534
rect 40960 3470 41012 3476
rect 42064 3528 42116 3534
rect 42064 3470 42116 3476
rect 42156 3528 42208 3534
rect 42156 3470 42208 3476
rect 42708 3528 42760 3534
rect 42708 3470 42760 3476
rect 43352 3528 43404 3534
rect 43352 3470 43404 3476
rect 39764 3460 39816 3466
rect 39764 3402 39816 3408
rect 39304 3256 39356 3262
rect 39304 3198 39356 3204
rect 39776 480 39804 3402
rect 40972 480 41000 3470
rect 42168 480 42196 3470
rect 43364 480 43392 3470
rect 44560 480 44588 3674
rect 46940 3664 46992 3670
rect 46940 3606 46992 3612
rect 45744 2916 45796 2922
rect 45744 2858 45796 2864
rect 45756 480 45784 2858
rect 46952 480 46980 3606
rect 48240 3482 48268 331910
rect 49620 3482 49648 333202
rect 50344 319456 50396 319462
rect 50344 319398 50396 319404
rect 48148 3454 48268 3482
rect 49344 3454 49648 3482
rect 48148 480 48176 3454
rect 49344 480 49372 3454
rect 50356 2922 50384 319398
rect 50988 302932 51040 302938
rect 50988 302874 51040 302880
rect 51000 3602 51028 302874
rect 52380 3602 52408 335990
rect 56508 334620 56560 334626
rect 56508 334562 56560 334568
rect 53748 326392 53800 326398
rect 53748 326334 53800 326340
rect 53760 3602 53788 326334
rect 56416 322244 56468 322250
rect 56416 322186 56468 322192
rect 54024 3664 54076 3670
rect 54024 3606 54076 3612
rect 50528 3596 50580 3602
rect 50528 3538 50580 3544
rect 50988 3596 51040 3602
rect 50988 3538 51040 3544
rect 51632 3596 51684 3602
rect 51632 3538 51684 3544
rect 52368 3596 52420 3602
rect 52368 3538 52420 3544
rect 52828 3596 52880 3602
rect 52828 3538 52880 3544
rect 53748 3596 53800 3602
rect 53748 3538 53800 3544
rect 50344 2916 50396 2922
rect 50344 2858 50396 2864
rect 50540 480 50568 3538
rect 51644 480 51672 3538
rect 52840 480 52868 3538
rect 54036 480 54064 3606
rect 55220 3392 55272 3398
rect 55220 3334 55272 3340
rect 55232 480 55260 3334
rect 56428 480 56456 322186
rect 56520 3398 56548 334562
rect 71688 330540 71740 330546
rect 71688 330482 71740 330488
rect 67548 319524 67600 319530
rect 67548 319466 67600 319472
rect 64788 10736 64840 10742
rect 64788 10678 64840 10684
rect 60648 10668 60700 10674
rect 60648 10610 60700 10616
rect 58808 9036 58860 9042
rect 58808 8978 58860 8984
rect 57612 3732 57664 3738
rect 57612 3674 57664 3680
rect 56508 3392 56560 3398
rect 56508 3334 56560 3340
rect 57624 480 57652 3674
rect 58820 480 58848 8978
rect 60660 3398 60688 10610
rect 62396 9104 62448 9110
rect 62396 9046 62448 9052
rect 61200 3800 61252 3806
rect 61200 3742 61252 3748
rect 60004 3392 60056 3398
rect 60004 3334 60056 3340
rect 60648 3392 60700 3398
rect 60648 3334 60700 3340
rect 60016 480 60044 3334
rect 61212 480 61240 3742
rect 62408 480 62436 9046
rect 64696 3868 64748 3874
rect 64696 3810 64748 3816
rect 63592 3392 63644 3398
rect 63592 3334 63644 3340
rect 63604 480 63632 3334
rect 64708 1986 64736 3810
rect 64800 3398 64828 10678
rect 65984 9172 66036 9178
rect 65984 9114 66036 9120
rect 64788 3392 64840 3398
rect 64788 3334 64840 3340
rect 64708 1958 64828 1986
rect 64800 480 64828 1958
rect 65996 480 66024 9114
rect 67560 626 67588 319466
rect 69480 9240 69532 9246
rect 69480 9182 69532 9188
rect 68284 3936 68336 3942
rect 68284 3878 68336 3884
rect 67192 598 67588 626
rect 67192 480 67220 598
rect 68296 480 68324 3878
rect 69492 480 69520 9182
rect 71700 3398 71728 330482
rect 78588 329180 78640 329186
rect 78588 329122 78640 329128
rect 74448 320884 74500 320890
rect 74448 320826 74500 320832
rect 73068 9308 73120 9314
rect 73068 9250 73120 9256
rect 71872 4004 71924 4010
rect 71872 3946 71924 3952
rect 70676 3392 70728 3398
rect 70676 3334 70728 3340
rect 71688 3392 71740 3398
rect 71688 3334 71740 3340
rect 70688 480 70716 3334
rect 71884 480 71912 3946
rect 73080 480 73108 9250
rect 74460 610 74488 320826
rect 76656 9376 76708 9382
rect 76656 9318 76708 9324
rect 75460 3188 75512 3194
rect 75460 3130 75512 3136
rect 74264 604 74316 610
rect 74264 546 74316 552
rect 74448 604 74500 610
rect 74448 546 74500 552
rect 74276 480 74304 546
rect 75472 480 75500 3130
rect 76668 480 76696 9318
rect 78600 3398 78628 329122
rect 82728 327820 82780 327826
rect 82728 327762 82780 327768
rect 80244 9444 80296 9450
rect 80244 9386 80296 9392
rect 79048 4140 79100 4146
rect 79048 4082 79100 4088
rect 77852 3392 77904 3398
rect 77852 3334 77904 3340
rect 78588 3392 78640 3398
rect 78588 3334 78640 3340
rect 77864 480 77892 3334
rect 79060 480 79088 4082
rect 80256 480 80284 9386
rect 82740 3398 82768 327762
rect 85488 318096 85540 318102
rect 85488 318038 85540 318044
rect 83832 9512 83884 9518
rect 83832 9454 83884 9460
rect 81440 3392 81492 3398
rect 81440 3334 81492 3340
rect 82728 3392 82780 3398
rect 82728 3334 82780 3340
rect 81452 480 81480 3334
rect 82636 3256 82688 3262
rect 82636 3198 82688 3204
rect 82648 480 82676 3198
rect 83844 480 83872 9454
rect 84108 4072 84160 4078
rect 84108 4014 84160 4020
rect 84120 3194 84148 4014
rect 85500 3330 85528 318038
rect 87328 9580 87380 9586
rect 87328 9522 87380 9528
rect 84936 3324 84988 3330
rect 84936 3266 84988 3272
rect 85488 3324 85540 3330
rect 85488 3266 85540 3272
rect 84108 3188 84160 3194
rect 84108 3130 84160 3136
rect 84948 480 84976 3266
rect 86132 3256 86184 3262
rect 86132 3198 86184 3204
rect 86144 480 86172 3198
rect 87340 480 87368 9522
rect 89640 3194 89668 335990
rect 96528 326460 96580 326466
rect 96528 326402 96580 326408
rect 92388 325032 92440 325038
rect 92388 324974 92440 324980
rect 90916 9648 90968 9654
rect 90916 9590 90968 9596
rect 89720 3256 89772 3262
rect 89720 3198 89772 3204
rect 88524 3188 88576 3194
rect 88524 3130 88576 3136
rect 89628 3188 89680 3194
rect 89628 3130 89680 3136
rect 88536 480 88564 3130
rect 89732 480 89760 3198
rect 90928 480 90956 9590
rect 92400 610 92428 324974
rect 94504 8900 94556 8906
rect 94504 8842 94556 8848
rect 93308 3188 93360 3194
rect 93308 3130 93360 3136
rect 92112 604 92164 610
rect 92112 546 92164 552
rect 92388 604 92440 610
rect 92388 546 92440 552
rect 92124 480 92152 546
rect 93320 480 93348 3130
rect 94516 480 94544 8842
rect 96540 3126 96568 326402
rect 99288 323672 99340 323678
rect 99288 323614 99340 323620
rect 98092 8832 98144 8838
rect 98092 8774 98144 8780
rect 95700 3120 95752 3126
rect 95700 3062 95752 3068
rect 96528 3120 96580 3126
rect 96528 3062 96580 3068
rect 95712 480 95740 3062
rect 96896 3052 96948 3058
rect 96896 2994 96948 3000
rect 96908 480 96936 2994
rect 98104 480 98132 8774
rect 99300 480 99328 323614
rect 100680 626 100708 337826
rect 103428 322312 103480 322318
rect 103428 322254 103480 322260
rect 101588 8764 101640 8770
rect 101588 8706 101640 8712
rect 100496 598 100708 626
rect 100496 480 100524 598
rect 101600 480 101628 8706
rect 103440 3126 103468 322254
rect 107476 316736 107528 316742
rect 107476 316678 107528 316684
rect 105176 8696 105228 8702
rect 105176 8638 105228 8644
rect 102784 3120 102836 3126
rect 102784 3062 102836 3068
rect 103428 3120 103480 3126
rect 103428 3062 103480 3068
rect 102796 480 102824 3062
rect 103980 2916 104032 2922
rect 103980 2858 104032 2864
rect 103992 480 104020 2858
rect 105188 480 105216 8638
rect 107488 3126 107516 316678
rect 106372 3120 106424 3126
rect 106372 3062 106424 3068
rect 107476 3120 107528 3126
rect 107476 3062 107528 3068
rect 106384 480 106412 3062
rect 107580 480 107608 337962
rect 115848 337952 115900 337958
rect 115848 337894 115900 337900
rect 114468 333328 114520 333334
rect 114468 333270 114520 333276
rect 110328 311160 110380 311166
rect 110328 311102 110380 311108
rect 108764 8628 108816 8634
rect 108764 8570 108816 8576
rect 108776 480 108804 8570
rect 110340 610 110368 311102
rect 112352 8560 112404 8566
rect 112352 8502 112404 8508
rect 111156 2916 111208 2922
rect 111156 2858 111208 2864
rect 109960 604 110012 610
rect 109960 546 110012 552
rect 110328 604 110380 610
rect 110328 546 110380 552
rect 109972 480 110000 546
rect 111168 480 111196 2858
rect 112364 480 112392 8502
rect 114480 2990 114508 333270
rect 113548 2984 113600 2990
rect 113548 2926 113600 2932
rect 114468 2984 114520 2990
rect 114468 2926 114520 2932
rect 113560 480 113588 2926
rect 115860 2922 115888 337894
rect 117228 334688 117280 334694
rect 117228 334630 117280 334636
rect 115940 8492 115992 8498
rect 115940 8434 115992 8440
rect 114744 2916 114796 2922
rect 114744 2858 114796 2864
rect 115848 2916 115900 2922
rect 115848 2858 115900 2864
rect 114756 480 114784 2858
rect 115952 480 115980 8434
rect 117240 4842 117268 334630
rect 121368 330608 121420 330614
rect 121368 330550 121420 330556
rect 119436 8424 119488 8430
rect 119436 8366 119488 8372
rect 117148 4814 117268 4842
rect 117148 480 117176 4814
rect 118240 2848 118292 2854
rect 118240 2790 118292 2796
rect 118252 480 118280 2790
rect 119448 480 119476 8366
rect 121380 2922 121408 330550
rect 125416 320952 125468 320958
rect 125416 320894 125468 320900
rect 123024 8356 123076 8362
rect 123024 8298 123076 8304
rect 120632 2916 120684 2922
rect 120632 2858 120684 2864
rect 121368 2916 121420 2922
rect 121368 2858 121420 2864
rect 120644 480 120672 2858
rect 121828 2848 121880 2854
rect 121828 2790 121880 2796
rect 121840 480 121868 2790
rect 123036 480 123064 8298
rect 125428 4214 125456 320894
rect 124220 4208 124272 4214
rect 124220 4150 124272 4156
rect 125416 4208 125468 4214
rect 125416 4150 125468 4156
rect 124232 480 124260 4150
rect 125520 3482 125548 338030
rect 162768 336252 162820 336258
rect 153212 336212 153332 336240
rect 153212 336122 153240 336212
rect 153304 336122 153332 336212
rect 162768 336194 162820 336200
rect 153200 336116 153252 336122
rect 153200 336058 153252 336064
rect 153292 336116 153344 336122
rect 153292 336058 153344 336064
rect 153108 336048 153160 336054
rect 153108 335990 153160 335996
rect 153120 335918 153148 335990
rect 153108 335912 153160 335918
rect 153108 335854 153160 335860
rect 160008 334824 160060 334830
rect 160008 334766 160060 334772
rect 126888 334756 126940 334762
rect 126888 334698 126940 334704
rect 126900 3482 126928 334698
rect 155868 333464 155920 333470
rect 155868 333406 155920 333412
rect 129648 333396 129700 333402
rect 129648 333338 129700 333344
rect 128268 330676 128320 330682
rect 128268 330618 128320 330624
rect 128280 3482 128308 330618
rect 129660 3482 129688 333338
rect 142068 332104 142120 332110
rect 142068 332046 142120 332052
rect 139308 332036 139360 332042
rect 139308 331978 139360 331984
rect 136548 321020 136600 321026
rect 136548 320962 136600 320968
rect 132592 7608 132644 7614
rect 132592 7550 132644 7556
rect 131396 6248 131448 6254
rect 131396 6190 131448 6196
rect 130200 5092 130252 5098
rect 130200 5034 130252 5040
rect 125428 3454 125548 3482
rect 126624 3454 126928 3482
rect 127820 3454 128308 3482
rect 129016 3454 129688 3482
rect 125428 480 125456 3454
rect 126624 480 126652 3454
rect 127820 480 127848 3454
rect 129016 480 129044 3454
rect 130212 480 130240 5034
rect 131408 480 131436 6190
rect 132604 480 132632 7550
rect 134892 6316 134944 6322
rect 134892 6258 134944 6264
rect 133788 5160 133840 5166
rect 133788 5102 133840 5108
rect 133800 480 133828 5102
rect 134904 480 134932 6258
rect 136560 4842 136588 320962
rect 137284 5296 137336 5302
rect 137284 5238 137336 5244
rect 136100 4814 136588 4842
rect 136100 480 136128 4814
rect 137296 480 137324 5238
rect 139320 4842 139348 331978
rect 141976 325100 142028 325106
rect 141976 325042 142028 325048
rect 140688 318164 140740 318170
rect 140688 318106 140740 318112
rect 140700 4842 140728 318106
rect 140872 5228 140924 5234
rect 140872 5170 140924 5176
rect 138492 4814 139348 4842
rect 139688 4814 140728 4842
rect 138492 480 138520 4814
rect 139688 480 139716 4814
rect 140884 480 140912 5170
rect 141988 4842 142016 325042
rect 142080 5234 142108 332046
rect 144828 330744 144880 330750
rect 144828 330686 144880 330692
rect 143448 316804 143500 316810
rect 143448 316746 143500 316752
rect 142068 5228 142120 5234
rect 142068 5170 142120 5176
rect 141988 4814 142108 4842
rect 142080 480 142108 4814
rect 143460 3346 143488 316746
rect 144840 3346 144868 330686
rect 153108 329316 153160 329322
rect 153108 329258 153160 329264
rect 151728 329248 151780 329254
rect 151728 329190 151780 329196
rect 150348 327888 150400 327894
rect 150348 327830 150400 327836
rect 146208 322380 146260 322386
rect 146208 322322 146260 322328
rect 146220 3346 146248 322322
rect 147588 315376 147640 315382
rect 147588 315318 147640 315324
rect 147600 3346 147628 315318
rect 148968 13116 149020 13122
rect 148968 13058 149020 13064
rect 148980 3346 149008 13058
rect 150360 3346 150388 327830
rect 151636 15904 151688 15910
rect 151636 15846 151688 15852
rect 151648 4214 151676 15846
rect 150440 4208 150492 4214
rect 150440 4150 150492 4156
rect 151636 4208 151688 4214
rect 151636 4150 151688 4156
rect 143276 3318 143488 3346
rect 144472 3318 144868 3346
rect 145668 3318 146248 3346
rect 146864 3318 147628 3346
rect 148060 3318 149008 3346
rect 149256 3318 150388 3346
rect 143276 480 143304 3318
rect 144472 480 144500 3318
rect 145668 480 145696 3318
rect 146864 480 146892 3318
rect 148060 480 148088 3318
rect 149256 480 149284 3318
rect 150452 480 150480 4150
rect 151740 3482 151768 329190
rect 153120 3618 153148 329258
rect 154488 319592 154540 319598
rect 154488 319534 154540 319540
rect 154500 3618 154528 319534
rect 155880 3618 155908 333406
rect 157248 326528 157300 326534
rect 157248 326470 157300 326476
rect 157260 3618 157288 326470
rect 159916 323740 159968 323746
rect 159916 323682 159968 323688
rect 158628 314016 158680 314022
rect 158628 313958 158680 313964
rect 158640 3618 158668 313958
rect 158720 4208 158772 4214
rect 158720 4150 158772 4156
rect 151556 3454 151768 3482
rect 152752 3590 153148 3618
rect 153948 3590 154528 3618
rect 155144 3590 155908 3618
rect 156340 3590 157288 3618
rect 157536 3590 158668 3618
rect 151556 480 151584 3454
rect 152752 480 152780 3590
rect 153948 480 153976 3590
rect 155144 480 155172 3590
rect 156340 480 156368 3590
rect 157536 480 157564 3590
rect 158732 480 158760 4150
rect 159928 480 159956 323682
rect 160020 4214 160048 334766
rect 161388 312656 161440 312662
rect 161388 312598 161440 312604
rect 160008 4208 160060 4214
rect 160008 4150 160060 4156
rect 161400 3618 161428 312598
rect 161124 3590 161428 3618
rect 161124 480 161152 3590
rect 162780 3482 162808 336194
rect 176568 336184 176620 336190
rect 176568 336126 176620 336132
rect 169668 334892 169720 334898
rect 169668 334834 169720 334840
rect 165528 330812 165580 330818
rect 165528 330754 165580 330760
rect 164148 14476 164200 14482
rect 164148 14418 164200 14424
rect 164160 3482 164188 14418
rect 165540 3482 165568 330754
rect 168288 327956 168340 327962
rect 168288 327898 168340 327904
rect 166908 11756 166960 11762
rect 166908 11698 166960 11704
rect 166920 3482 166948 11698
rect 168196 7676 168248 7682
rect 168196 7618 168248 7624
rect 167092 4208 167144 4214
rect 167092 4150 167144 4156
rect 162320 3454 162808 3482
rect 163516 3454 164188 3482
rect 164712 3454 165568 3482
rect 165908 3454 166948 3482
rect 162320 480 162348 3454
rect 163516 480 163544 3454
rect 164712 480 164740 3454
rect 165908 480 165936 3454
rect 167104 480 167132 4150
rect 168208 480 168236 7618
rect 168300 4214 168328 327898
rect 168288 4208 168340 4214
rect 168288 4150 168340 4156
rect 169680 3482 169708 334834
rect 173808 333532 173860 333538
rect 173808 333474 173860 333480
rect 171048 326596 171100 326602
rect 171048 326538 171100 326544
rect 171060 3482 171088 326538
rect 171784 7744 171836 7750
rect 171784 7686 171836 7692
rect 169404 3454 169708 3482
rect 170600 3454 171088 3482
rect 169404 480 169432 3454
rect 170600 480 170628 3454
rect 171796 480 171824 7686
rect 173820 4842 173848 333474
rect 175372 7812 175424 7818
rect 175372 7754 175424 7760
rect 174176 6384 174228 6390
rect 174176 6326 174228 6332
rect 172992 4814 173848 4842
rect 172992 480 173020 4814
rect 174188 480 174216 6326
rect 175384 480 175412 7754
rect 176580 480 176608 336126
rect 180076 208350 180104 399298
rect 184848 333600 184900 333606
rect 184848 333542 184900 333548
rect 180708 332172 180760 332178
rect 180708 332114 180760 332120
rect 180064 208344 180116 208350
rect 180064 208286 180116 208292
rect 178960 7880 179012 7886
rect 178960 7822 179012 7828
rect 177764 6452 177816 6458
rect 177764 6394 177816 6400
rect 177776 480 177804 6394
rect 178972 480 179000 7822
rect 180720 4842 180748 332114
rect 182548 7948 182600 7954
rect 182548 7890 182600 7896
rect 181352 6520 181404 6526
rect 181352 6462 181404 6468
rect 180168 4814 180748 4842
rect 180168 480 180196 4814
rect 181364 480 181392 6462
rect 182560 480 182588 7890
rect 184860 6746 184888 333542
rect 204916 93838 204944 399366
rect 206928 329384 206980 329390
rect 206928 329326 206980 329332
rect 204904 93832 204956 93838
rect 204904 93774 204956 93780
rect 200396 8288 200448 8294
rect 200396 8230 200448 8236
rect 196808 8220 196860 8226
rect 196808 8162 196860 8168
rect 193220 8152 193272 8158
rect 193220 8094 193272 8100
rect 189632 8084 189684 8090
rect 189632 8026 189684 8032
rect 186044 8016 186096 8022
rect 186044 7958 186096 7964
rect 184768 6718 184888 6746
rect 184768 610 184796 6718
rect 184848 6588 184900 6594
rect 184848 6530 184900 6536
rect 183744 604 183796 610
rect 183744 546 183796 552
rect 184756 604 184808 610
rect 184756 546 184808 552
rect 183756 480 183784 546
rect 184860 480 184888 6530
rect 186056 480 186084 7958
rect 188436 6656 188488 6662
rect 188436 6598 188488 6604
rect 187240 5296 187292 5302
rect 187240 5238 187292 5244
rect 187252 480 187280 5238
rect 188448 480 188476 6598
rect 189644 480 189672 8026
rect 192024 6724 192076 6730
rect 192024 6666 192076 6672
rect 190828 5364 190880 5370
rect 190828 5306 190880 5312
rect 190840 480 190868 5306
rect 192036 480 192064 6666
rect 193232 480 193260 8094
rect 195612 6792 195664 6798
rect 195612 6734 195664 6740
rect 194416 5432 194468 5438
rect 194416 5374 194468 5380
rect 194428 480 194456 5374
rect 195624 480 195652 6734
rect 196820 480 196848 8162
rect 199200 6860 199252 6866
rect 199200 6802 199252 6808
rect 198004 5500 198056 5506
rect 198004 5442 198056 5448
rect 198016 480 198044 5442
rect 199212 480 199240 6802
rect 200408 480 200436 8230
rect 203892 7540 203944 7546
rect 203892 7482 203944 7488
rect 202696 6112 202748 6118
rect 202696 6054 202748 6060
rect 201500 4752 201552 4758
rect 201500 4694 201552 4700
rect 201512 480 201540 4694
rect 202708 480 202736 6054
rect 203904 480 203932 7482
rect 205088 4684 205140 4690
rect 205088 4626 205140 4632
rect 205100 480 205128 4626
rect 206940 610 206968 329326
rect 207676 180810 207704 399502
rect 208308 335028 208360 335034
rect 208308 334970 208360 334976
rect 207664 180804 207716 180810
rect 207664 180746 207716 180752
rect 208320 610 208348 334970
rect 209056 223582 209084 400522
rect 209688 336320 209740 336326
rect 209688 336262 209740 336268
rect 209044 223576 209096 223582
rect 209044 223518 209096 223524
rect 209700 610 209728 336262
rect 211264 336122 211384 336138
rect 211252 336116 211396 336122
rect 211304 336110 211344 336116
rect 211252 336058 211304 336064
rect 211344 336058 211396 336064
rect 211068 330880 211120 330886
rect 211068 330822 211120 330828
rect 210976 321088 211028 321094
rect 210976 321030 211028 321036
rect 209872 4208 209924 4214
rect 209872 4150 209924 4156
rect 206284 604 206336 610
rect 206284 546 206336 552
rect 206928 604 206980 610
rect 206928 546 206980 552
rect 207480 604 207532 610
rect 207480 546 207532 552
rect 208308 604 208360 610
rect 208308 546 208360 552
rect 208676 604 208728 610
rect 208676 546 208728 552
rect 209688 604 209740 610
rect 209688 546 209740 552
rect 206296 480 206324 546
rect 207492 480 207520 546
rect 208688 480 208716 546
rect 209884 480 209912 4150
rect 210988 3482 211016 321030
rect 211080 4214 211108 330822
rect 211816 266354 211844 400658
rect 215944 400648 215996 400654
rect 215944 400590 215996 400596
rect 213184 399832 213236 399838
rect 213184 399774 213236 399780
rect 212448 334960 212500 334966
rect 212448 334902 212500 334908
rect 211804 266348 211856 266354
rect 211804 266290 211856 266296
rect 211068 4208 211120 4214
rect 211068 4150 211120 4156
rect 212460 3618 212488 334902
rect 213196 309126 213224 399774
rect 214564 399628 214616 399634
rect 214564 399570 214616 399576
rect 213828 325168 213880 325174
rect 213828 325110 213880 325116
rect 213184 309120 213236 309126
rect 213184 309062 213236 309068
rect 213840 3618 213868 325110
rect 214576 35902 214604 399570
rect 215208 319660 215260 319666
rect 215208 319602 215260 319608
rect 214564 35896 214616 35902
rect 214564 35838 214616 35844
rect 215220 3618 215248 319602
rect 215956 80034 215984 400590
rect 218704 399764 218756 399770
rect 218704 399706 218756 399712
rect 216588 336388 216640 336394
rect 216588 336330 216640 336336
rect 215944 80028 215996 80034
rect 215944 79970 215996 79976
rect 216600 3618 216628 336330
rect 217968 323808 218020 323814
rect 217968 323750 218020 323756
rect 217980 3618 218008 323750
rect 218716 122806 218744 399706
rect 220728 336456 220780 336462
rect 220728 336398 220780 336404
rect 219348 333668 219400 333674
rect 219348 333610 219400 333616
rect 218704 122800 218756 122806
rect 218704 122742 218756 122748
rect 219256 122120 219308 122126
rect 219256 122062 219308 122068
rect 219268 3618 219296 122062
rect 212276 3590 212488 3618
rect 213472 3590 213868 3618
rect 214668 3590 215248 3618
rect 215864 3590 216628 3618
rect 217060 3590 218008 3618
rect 218164 3590 219296 3618
rect 210988 3454 211108 3482
rect 211080 480 211108 3454
rect 212276 480 212304 3590
rect 213472 480 213500 3590
rect 214668 480 214696 3590
rect 215864 480 215892 3590
rect 217060 480 217088 3590
rect 218164 480 218192 3590
rect 219360 480 219388 333610
rect 220740 3346 220768 336398
rect 222108 328024 222160 328030
rect 222108 327966 222160 327972
rect 222120 3346 222148 327966
rect 222856 165578 222884 400998
rect 225604 400988 225656 400994
rect 225604 400930 225656 400936
rect 223488 335096 223540 335102
rect 223488 335038 223540 335044
rect 222844 165572 222896 165578
rect 222844 165514 222896 165520
rect 223500 3346 223528 335038
rect 224868 332240 224920 332246
rect 224868 332182 224920 332188
rect 224880 3346 224908 332182
rect 225616 51066 225644 400930
rect 225696 337272 225748 337278
rect 225696 337214 225748 337220
rect 225604 51060 225656 51066
rect 225604 51002 225656 51008
rect 225708 13122 225736 337214
rect 225800 252550 225828 401202
rect 227076 401192 227128 401198
rect 227076 401134 227128 401140
rect 226984 400104 227036 400110
rect 226984 400046 227036 400052
rect 226996 367062 227024 400046
rect 226984 367056 227036 367062
rect 226984 366998 227036 367004
rect 226984 329520 227036 329526
rect 226984 329462 227036 329468
rect 226248 326664 226300 326670
rect 226248 326606 226300 326612
rect 225788 252544 225840 252550
rect 225788 252486 225840 252492
rect 225696 13116 225748 13122
rect 225696 13058 225748 13064
rect 226260 3346 226288 326606
rect 226996 11762 227024 329462
rect 227088 136610 227116 401134
rect 227180 295322 227208 401270
rect 233332 401124 233384 401130
rect 233332 401066 233384 401072
rect 231768 400852 231820 400858
rect 231768 400794 231820 400800
rect 230664 400444 230716 400450
rect 230664 400386 230716 400392
rect 230676 399908 230704 400386
rect 231780 399908 231808 400794
rect 233344 399908 233372 401066
rect 234896 400920 234948 400926
rect 234896 400862 234948 400868
rect 233884 400376 233936 400382
rect 233884 400318 233936 400324
rect 233896 399908 233924 400318
rect 234908 399908 234936 400862
rect 235448 400512 235500 400518
rect 235448 400454 235500 400460
rect 235460 399908 235488 400454
rect 235828 399922 235856 401911
rect 235908 401882 235960 401888
rect 238024 400784 238076 400790
rect 238024 400726 238076 400732
rect 236736 399968 236788 399974
rect 235828 399894 235934 399922
rect 236486 399916 236736 399922
rect 236486 399910 236788 399916
rect 236486 399894 236776 399910
rect 238036 399908 238064 400726
rect 241704 400308 241756 400314
rect 241704 400250 241756 400256
rect 241244 400240 241296 400246
rect 241244 400182 241296 400188
rect 238576 400172 238628 400178
rect 238576 400114 238628 400120
rect 238588 399908 238616 400114
rect 239614 399906 239904 399922
rect 241256 399908 241284 400182
rect 241716 399908 241744 400250
rect 242268 399908 242296 401950
rect 243268 401872 243320 401878
rect 243268 401814 243320 401820
rect 242624 400036 242676 400042
rect 242624 399978 242676 399984
rect 242636 399922 242664 399978
rect 239614 399900 239916 399906
rect 239614 399894 239864 399900
rect 242636 399894 242834 399922
rect 243280 399908 243308 401814
rect 243832 399908 243860 404330
rect 244200 401878 244228 415414
rect 244924 402008 244976 402014
rect 244924 401950 244976 401956
rect 244188 401872 244240 401878
rect 244188 401814 244240 401820
rect 244372 401872 244424 401878
rect 244372 401814 244424 401820
rect 244384 399908 244412 401814
rect 244936 399908 244964 401950
rect 245396 401878 245424 438874
rect 245384 401872 245436 401878
rect 245384 401814 245436 401820
rect 245488 399922 245516 451250
rect 245580 402014 245608 462334
rect 245568 402008 245620 402014
rect 245568 401950 245620 401956
rect 246868 401878 246896 485794
rect 245936 401872 245988 401878
rect 245936 401814 245988 401820
rect 246856 401872 246908 401878
rect 246856 401814 246908 401820
rect 245410 399894 245516 399922
rect 245948 399908 245976 401814
rect 246960 399922 246988 509254
rect 248144 498228 248196 498234
rect 248144 498170 248196 498176
rect 248156 402014 248184 498170
rect 247040 402008 247092 402014
rect 247040 401950 247092 401956
rect 248144 402008 248196 402014
rect 248144 401950 248196 401956
rect 246514 399894 246988 399922
rect 247052 399908 247080 401950
rect 248248 401878 248276 532714
rect 247500 401872 247552 401878
rect 247500 401814 247552 401820
rect 248236 401872 248288 401878
rect 248236 401814 248288 401820
rect 247512 399908 247540 401814
rect 248340 399922 248368 556174
rect 249524 545148 249576 545154
rect 249524 545090 249576 545096
rect 249536 402014 249564 545090
rect 248604 402008 248656 402014
rect 248604 401950 248656 401956
rect 249524 402008 249576 402014
rect 249524 401950 249576 401956
rect 248078 399894 248368 399922
rect 248616 399908 248644 401950
rect 249628 400330 249656 579634
rect 249536 400302 249656 400330
rect 249536 399922 249564 400302
rect 249720 399922 249748 603094
rect 250996 592068 251048 592074
rect 250996 592010 251048 592016
rect 251008 402014 251036 592010
rect 250168 402008 250220 402014
rect 250168 401950 250220 401956
rect 250996 402008 251048 402014
rect 250996 401950 251048 401956
rect 249090 399894 249564 399922
rect 249642 399894 249748 399922
rect 250180 399908 250208 401950
rect 251100 399922 251128 626554
rect 251180 402008 251232 402014
rect 251180 401950 251232 401956
rect 250746 399894 251128 399922
rect 251192 399908 251220 401950
rect 252296 400330 252324 638930
rect 252388 402014 252416 650014
rect 252376 402008 252428 402014
rect 252376 401950 252428 401956
rect 252204 400302 252324 400330
rect 239864 399842 239916 399848
rect 252204 399786 252232 400302
rect 252480 399922 252508 673474
rect 252744 402008 252796 402014
rect 252744 401950 252796 401956
rect 252310 399894 252508 399922
rect 252756 399908 252784 401950
rect 253676 399922 253704 685850
rect 253768 402014 253796 696934
rect 253756 402008 253808 402014
rect 253756 401950 253808 401956
rect 253322 399894 253704 399922
rect 253860 399908 253888 700266
rect 254400 402756 254452 402762
rect 254400 402698 254452 402704
rect 254412 399908 254440 402698
rect 255148 399922 255176 700334
rect 255240 402762 255268 700402
rect 256436 402898 256464 700538
rect 255412 402892 255464 402898
rect 255412 402834 255464 402840
rect 256424 402892 256476 402898
rect 256424 402834 256476 402840
rect 255228 402756 255280 402762
rect 255228 402698 255280 402704
rect 254886 399894 255176 399922
rect 255424 399908 255452 402834
rect 256528 400058 256556 700674
rect 256608 700664 256660 700670
rect 256608 700606 256660 700612
rect 256344 400030 256556 400058
rect 256344 399922 256372 400030
rect 256620 399922 256648 700606
rect 256976 402892 257028 402898
rect 256976 402834 257028 402840
rect 255990 399894 256372 399922
rect 256450 399894 256648 399922
rect 256988 399908 257016 402834
rect 257908 399922 257936 700946
rect 259368 700936 259420 700942
rect 259368 700878 259420 700884
rect 257988 700868 258040 700874
rect 257988 700810 258040 700816
rect 258000 402898 258028 700810
rect 259276 700188 259328 700194
rect 259276 700130 259328 700136
rect 259184 700052 259236 700058
rect 259184 699994 259236 700000
rect 257988 402892 258040 402898
rect 257988 402834 258040 402840
rect 258540 402892 258592 402898
rect 258540 402834 258592 402840
rect 258080 402212 258132 402218
rect 258080 402154 258132 402160
rect 257554 399894 257936 399922
rect 258092 399908 258120 402154
rect 258552 399908 258580 402834
rect 259196 399922 259224 699994
rect 259288 402898 259316 700130
rect 259276 402892 259328 402898
rect 259276 402834 259328 402840
rect 259380 402218 259408 700878
rect 265072 700800 265124 700806
rect 265072 700742 265124 700748
rect 263784 700256 263836 700262
rect 263784 700198 263836 700204
rect 260656 700120 260708 700126
rect 260656 700062 260708 700068
rect 260668 402898 260696 700062
rect 262220 699984 262272 699990
rect 262220 699926 262272 699932
rect 262128 699916 262180 699922
rect 262128 699858 262180 699864
rect 260748 699712 260800 699718
rect 260748 699654 260800 699660
rect 259644 402892 259696 402898
rect 259644 402834 259696 402840
rect 260656 402892 260708 402898
rect 260656 402834 260708 402840
rect 259368 402212 259420 402218
rect 259368 402154 259420 402160
rect 259118 399894 259224 399922
rect 259656 399908 259684 402834
rect 260196 402008 260248 402014
rect 260196 401950 260248 401956
rect 260208 399908 260236 401950
rect 260760 399922 260788 699654
rect 262140 402898 262168 699858
rect 261208 402892 261260 402898
rect 261208 402834 261260 402840
rect 262128 402892 262180 402898
rect 262128 402834 262180 402840
rect 260682 399894 260788 399922
rect 261220 399908 261248 402834
rect 261760 402144 261812 402150
rect 261760 402086 261812 402092
rect 261772 399908 261800 402086
rect 262232 399908 262260 699926
rect 262864 552084 262916 552090
rect 262864 552026 262916 552032
rect 262772 402756 262824 402762
rect 262772 402698 262824 402704
rect 262784 399908 262812 402698
rect 262876 402150 262904 552026
rect 262864 402144 262916 402150
rect 262864 402086 262916 402092
rect 262956 401600 263008 401606
rect 262956 401542 263008 401548
rect 262968 399922 262996 401542
rect 263796 399922 263824 700198
rect 264244 495508 264296 495514
rect 264244 495450 264296 495456
rect 264256 402966 264284 495450
rect 264888 403028 264940 403034
rect 264888 402970 264940 402976
rect 264244 402960 264296 402966
rect 264244 402902 264296 402908
rect 264336 401940 264388 401946
rect 264336 401882 264388 401888
rect 262968 399894 263350 399922
rect 263796 399894 263902 399922
rect 264348 399908 264376 401882
rect 264900 399908 264928 402970
rect 264980 401940 265032 401946
rect 264980 401882 265032 401888
rect 251758 399758 252232 399786
rect 232504 399696 232556 399702
rect 232254 399644 232504 399650
rect 232254 399638 232556 399644
rect 232254 399622 232544 399638
rect 240322 399528 240378 399537
rect 240166 399486 240322 399514
rect 264992 399498 265020 401882
rect 265084 399922 265112 700742
rect 266544 700528 266596 700534
rect 266544 700470 266596 700476
rect 265624 437504 265676 437510
rect 265624 437446 265676 437452
rect 265636 402898 265664 437446
rect 265624 402892 265676 402898
rect 265624 402834 265676 402840
rect 265900 402824 265952 402830
rect 265900 402766 265952 402772
rect 265084 399894 265466 399922
rect 265912 399908 265940 402766
rect 266452 402620 266504 402626
rect 266452 402562 266504 402568
rect 266464 399908 266492 402562
rect 266556 399922 266584 700470
rect 267660 699718 267688 703520
rect 283852 699922 283880 703520
rect 283840 699916 283892 699922
rect 283840 699858 283892 699864
rect 267648 699712 267700 699718
rect 267648 699654 267700 699660
rect 300136 688634 300164 703520
rect 332520 700058 332548 703520
rect 348804 700126 348832 703520
rect 364996 700194 365024 703520
rect 397472 701010 397500 703520
rect 397460 701004 397512 701010
rect 397460 700946 397512 700952
rect 413664 700942 413692 703520
rect 413652 700936 413704 700942
rect 413652 700878 413704 700884
rect 429856 700874 429884 703520
rect 429844 700868 429896 700874
rect 429844 700810 429896 700816
rect 462332 700738 462360 703520
rect 462320 700732 462372 700738
rect 462320 700674 462372 700680
rect 478524 700670 478552 703520
rect 478512 700664 478564 700670
rect 478512 700606 478564 700612
rect 494808 700602 494836 703520
rect 494796 700596 494848 700602
rect 494796 700538 494848 700544
rect 527192 700466 527220 703520
rect 527180 700460 527232 700466
rect 527180 700402 527232 700408
rect 543476 700398 543504 703520
rect 543464 700392 543516 700398
rect 543464 700334 543516 700340
rect 559668 700330 559696 703520
rect 559656 700324 559708 700330
rect 559656 700266 559708 700272
rect 364984 700188 365036 700194
rect 364984 700130 365036 700136
rect 348792 700120 348844 700126
rect 348792 700062 348844 700068
rect 332508 700052 332560 700058
rect 332508 699994 332560 700000
rect 580170 698048 580226 698057
rect 580170 697983 580226 697992
rect 580184 696998 580212 697983
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 299664 688628 299716 688634
rect 299664 688570 299716 688576
rect 300124 688628 300176 688634
rect 300124 688570 300176 688576
rect 299676 685930 299704 688570
rect 580170 686352 580226 686361
rect 580170 686287 580226 686296
rect 299584 685902 299704 685930
rect 580184 685914 580212 686287
rect 580172 685908 580224 685914
rect 299584 684486 299612 685902
rect 580172 685850 580224 685856
rect 299572 684480 299624 684486
rect 299572 684422 299624 684428
rect 580170 674656 580226 674665
rect 580170 674591 580226 674600
rect 580184 673538 580212 674591
rect 580172 673532 580224 673538
rect 580172 673474 580224 673480
rect 299940 666596 299992 666602
rect 299940 666538 299992 666544
rect 299952 659682 299980 666538
rect 299768 659654 299980 659682
rect 267832 652792 267884 652798
rect 267832 652734 267884 652740
rect 267844 402778 267872 652734
rect 299768 647290 299796 659654
rect 580170 651128 580226 651137
rect 580170 651063 580226 651072
rect 580184 650078 580212 651063
rect 580172 650072 580224 650078
rect 580172 650014 580224 650020
rect 299664 647284 299716 647290
rect 299664 647226 299716 647232
rect 299756 647284 299808 647290
rect 299756 647226 299808 647232
rect 299676 640422 299704 647226
rect 299664 640416 299716 640422
rect 299664 640358 299716 640364
rect 299756 640416 299808 640422
rect 299756 640358 299808 640364
rect 299768 630698 299796 640358
rect 580170 639432 580226 639441
rect 580170 639367 580226 639376
rect 580184 638994 580212 639367
rect 580172 638988 580224 638994
rect 580172 638930 580224 638936
rect 299572 630692 299624 630698
rect 299572 630634 299624 630640
rect 299756 630692 299808 630698
rect 299756 630634 299808 630640
rect 299584 630578 299612 630634
rect 299584 630550 299704 630578
rect 299676 621058 299704 630550
rect 580170 627736 580226 627745
rect 580170 627671 580226 627680
rect 580184 626618 580212 627671
rect 580172 626612 580224 626618
rect 580172 626554 580224 626560
rect 299676 621030 299796 621058
rect 299768 611386 299796 621030
rect 299572 611380 299624 611386
rect 299572 611322 299624 611328
rect 299756 611380 299808 611386
rect 299756 611322 299808 611328
rect 299584 611266 299612 611322
rect 299584 611238 299704 611266
rect 299676 608598 299704 611238
rect 299664 608592 299716 608598
rect 299664 608534 299716 608540
rect 580170 604208 580226 604217
rect 580170 604143 580226 604152
rect 580184 603158 580212 604143
rect 580172 603152 580224 603158
rect 580172 603094 580224 603100
rect 299848 601724 299900 601730
rect 299848 601666 299900 601672
rect 299860 598942 299888 601666
rect 299848 598936 299900 598942
rect 299848 598878 299900 598884
rect 269304 594856 269356 594862
rect 269304 594798 269356 594804
rect 267844 402750 268148 402778
rect 268016 402688 268068 402694
rect 268016 402630 268068 402636
rect 267556 402076 267608 402082
rect 267556 402018 267608 402024
rect 266556 399894 267030 399922
rect 267568 399908 267596 402018
rect 268028 399908 268056 402630
rect 268120 399786 268148 402750
rect 269120 402552 269172 402558
rect 269120 402494 269172 402500
rect 269132 399908 269160 402494
rect 269316 402370 269344 594798
rect 580170 592512 580226 592521
rect 580170 592447 580226 592456
rect 580184 592074 580212 592447
rect 580172 592068 580224 592074
rect 580172 592010 580224 592016
rect 299940 589348 299992 589354
rect 299940 589290 299992 589296
rect 299952 582486 299980 589290
rect 299940 582480 299992 582486
rect 299940 582422 299992 582428
rect 299848 582344 299900 582350
rect 299848 582286 299900 582292
rect 299860 572642 299888 582286
rect 580170 580816 580226 580825
rect 580170 580751 580226 580760
rect 580184 579698 580212 580751
rect 580172 579692 580224 579698
rect 580172 579634 580224 579640
rect 299676 572614 299888 572642
rect 299676 569922 299704 572614
rect 299584 569894 299704 569922
rect 299584 563174 299612 569894
rect 299572 563168 299624 563174
rect 299572 563110 299624 563116
rect 299572 563032 299624 563038
rect 299572 562974 299624 562980
rect 299584 560561 299612 562974
rect 299570 560552 299626 560561
rect 299570 560487 299626 560496
rect 299570 560416 299626 560425
rect 299570 560351 299626 560360
rect 299584 553518 299612 560351
rect 580170 557288 580226 557297
rect 580170 557223 580226 557232
rect 580184 556238 580212 557223
rect 580172 556232 580224 556238
rect 580172 556174 580224 556180
rect 299572 553512 299624 553518
rect 299572 553454 299624 553460
rect 299480 553376 299532 553382
rect 299480 553318 299532 553324
rect 299492 549273 299520 553318
rect 299294 549264 299350 549273
rect 299294 549199 299350 549208
rect 299478 549264 299534 549273
rect 299478 549199 299534 549208
rect 299308 543726 299336 549199
rect 580170 545592 580226 545601
rect 580170 545527 580226 545536
rect 580184 545154 580212 545527
rect 580172 545148 580224 545154
rect 580172 545090 580224 545096
rect 299296 543720 299348 543726
rect 299296 543662 299348 543668
rect 299480 543720 299532 543726
rect 299480 543662 299532 543668
rect 299492 539594 299520 543662
rect 299492 539566 299612 539594
rect 270776 538280 270828 538286
rect 270776 538222 270828 538228
rect 270788 402642 270816 538222
rect 299584 531350 299612 539566
rect 580170 533896 580226 533905
rect 580170 533831 580226 533840
rect 580184 532778 580212 533831
rect 580172 532772 580224 532778
rect 580172 532714 580224 532720
rect 299572 531344 299624 531350
rect 299572 531286 299624 531292
rect 299756 531344 299808 531350
rect 299756 531286 299808 531292
rect 299768 524482 299796 531286
rect 299756 524476 299808 524482
rect 299756 524418 299808 524424
rect 299848 524408 299900 524414
rect 299848 524350 299900 524356
rect 299860 521665 299888 524350
rect 299662 521656 299718 521665
rect 299662 521591 299718 521600
rect 299846 521656 299902 521665
rect 299846 521591 299902 521600
rect 299676 512038 299704 521591
rect 299664 512032 299716 512038
rect 299664 511974 299716 511980
rect 299940 512032 299992 512038
rect 299940 511974 299992 511980
rect 299952 502382 299980 511974
rect 580170 510368 580226 510377
rect 580170 510303 580226 510312
rect 580184 509318 580212 510303
rect 580172 509312 580224 509318
rect 580172 509254 580224 509260
rect 299756 502376 299808 502382
rect 299478 502344 299534 502353
rect 299478 502279 299534 502288
rect 299754 502344 299756 502353
rect 299940 502376 299992 502382
rect 299808 502344 299810 502353
rect 299940 502318 299992 502324
rect 299754 502279 299810 502288
rect 299492 492697 299520 502279
rect 580170 498672 580226 498681
rect 580170 498607 580226 498616
rect 580184 498234 580212 498607
rect 580172 498228 580224 498234
rect 580172 498170 580224 498176
rect 299478 492688 299534 492697
rect 299478 492623 299534 492632
rect 299662 492688 299718 492697
rect 299662 492623 299664 492632
rect 299716 492623 299718 492632
rect 299664 492594 299716 492600
rect 580170 486840 580226 486849
rect 580170 486775 580226 486784
rect 580184 485858 580212 486775
rect 580172 485852 580224 485858
rect 580172 485794 580224 485800
rect 299664 485784 299716 485790
rect 299664 485726 299716 485732
rect 299676 483018 299704 485726
rect 299676 482990 299796 483018
rect 272524 480276 272576 480282
rect 272524 480218 272576 480224
rect 270788 402614 271552 402642
rect 271236 402484 271288 402490
rect 271236 402426 271288 402432
rect 270684 402416 270736 402422
rect 269316 402342 269896 402370
rect 270684 402358 270736 402364
rect 269580 402212 269632 402218
rect 269580 402154 269632 402160
rect 269592 399908 269620 402154
rect 269868 399922 269896 402342
rect 269868 399894 270158 399922
rect 270696 399908 270724 402358
rect 271248 399908 271276 402426
rect 271524 399922 271552 402614
rect 272248 402144 272300 402150
rect 272248 402086 272300 402092
rect 271524 399894 271722 399922
rect 272260 399908 272288 402086
rect 272536 401946 272564 480218
rect 299768 476134 299796 482990
rect 299572 476128 299624 476134
rect 299756 476128 299808 476134
rect 299624 476076 299704 476082
rect 299572 476070 299704 476076
rect 299756 476070 299808 476076
rect 299584 476054 299704 476070
rect 299676 473346 299704 476054
rect 299664 473340 299716 473346
rect 299664 473282 299716 473288
rect 299664 466404 299716 466410
rect 299664 466346 299716 466352
rect 299676 463706 299704 466346
rect 299676 463678 299796 463706
rect 299768 460902 299796 463678
rect 580170 463448 580226 463457
rect 580170 463383 580226 463392
rect 580184 462398 580212 463383
rect 580172 462392 580224 462398
rect 580172 462334 580224 462340
rect 299388 460896 299440 460902
rect 299388 460838 299440 460844
rect 299756 460896 299808 460902
rect 299756 460838 299808 460844
rect 299400 451330 299428 460838
rect 580170 451752 580226 451761
rect 580170 451687 580226 451696
rect 299400 451302 299520 451330
rect 580184 451314 580212 451687
rect 299492 449886 299520 451302
rect 580172 451308 580224 451314
rect 580172 451250 580224 451256
rect 299480 449880 299532 449886
rect 299480 449822 299532 449828
rect 299572 440292 299624 440298
rect 299572 440234 299624 440240
rect 299584 436830 299612 440234
rect 580170 439920 580226 439929
rect 580170 439855 580226 439864
rect 580184 438938 580212 439855
rect 580172 438932 580224 438938
rect 580172 438874 580224 438880
rect 299572 436824 299624 436830
rect 299572 436766 299624 436772
rect 299572 427780 299624 427786
rect 299572 427722 299624 427728
rect 273904 423700 273956 423706
rect 273904 423642 273956 423648
rect 273916 402966 273944 423642
rect 299584 418146 299612 427722
rect 299584 418118 299796 418146
rect 299768 415410 299796 418118
rect 580170 416528 580226 416537
rect 580170 416463 580226 416472
rect 580184 415478 580212 416463
rect 580172 415472 580224 415478
rect 580172 415414 580224 415420
rect 299756 415404 299808 415410
rect 299756 415346 299808 415352
rect 299664 405748 299716 405754
rect 299664 405690 299716 405696
rect 273812 402960 273864 402966
rect 273812 402902 273864 402908
rect 273904 402960 273956 402966
rect 273904 402902 273956 402908
rect 274916 402960 274968 402966
rect 274916 402902 274968 402908
rect 272800 402348 272852 402354
rect 272800 402290 272852 402296
rect 272524 401940 272576 401946
rect 272524 401882 272576 401888
rect 272812 399908 272840 402290
rect 273260 401940 273312 401946
rect 273260 401882 273312 401888
rect 273272 399908 273300 401882
rect 273824 399908 273852 402902
rect 274364 402280 274416 402286
rect 274364 402222 274416 402228
rect 274376 399908 274404 402222
rect 274928 399908 274956 402902
rect 275376 402892 275428 402898
rect 275376 402834 275428 402840
rect 275388 399908 275416 402834
rect 277032 402076 277084 402082
rect 277032 402018 277084 402024
rect 275928 401464 275980 401470
rect 275928 401406 275980 401412
rect 275940 399908 275968 401406
rect 276480 400104 276532 400110
rect 276480 400046 276532 400052
rect 276492 399908 276520 400046
rect 277044 399908 277072 402018
rect 299676 402014 299704 405690
rect 580170 404832 580226 404841
rect 580170 404767 580226 404776
rect 580184 404394 580212 404767
rect 580172 404388 580224 404394
rect 580172 404330 580224 404336
rect 299664 402008 299716 402014
rect 299664 401950 299716 401956
rect 485042 401976 485098 401985
rect 485042 401911 485098 401920
rect 289634 401840 289690 401849
rect 278596 401804 278648 401810
rect 289634 401775 289690 401784
rect 278596 401746 278648 401752
rect 277492 401396 277544 401402
rect 277492 401338 277544 401344
rect 277504 399908 277532 401338
rect 278608 399908 278636 401746
rect 280160 401736 280212 401742
rect 280160 401678 280212 401684
rect 279056 401328 279108 401334
rect 279056 401270 279108 401276
rect 279068 399908 279096 401270
rect 279608 400716 279660 400722
rect 279608 400658 279660 400664
rect 279620 399908 279648 400658
rect 280172 399908 280200 401678
rect 281724 401668 281776 401674
rect 281724 401610 281776 401616
rect 280712 401260 280764 401266
rect 280712 401202 280764 401208
rect 280724 399908 280752 401202
rect 281172 400580 281224 400586
rect 281172 400522 281224 400528
rect 281184 399908 281212 400522
rect 281736 399908 281764 401610
rect 284392 401192 284444 401198
rect 284392 401134 284444 401140
rect 283840 401056 283892 401062
rect 283840 400998 283892 401004
rect 283852 399908 283880 400998
rect 284404 399908 284432 401134
rect 287520 400988 287572 400994
rect 287520 400930 287572 400936
rect 286968 400648 287020 400654
rect 286968 400590 287020 400596
rect 286980 399908 287008 400590
rect 287532 399908 287560 400930
rect 289648 399908 289676 401775
rect 291936 401124 291988 401130
rect 291936 401066 291988 401072
rect 290556 400308 290608 400314
rect 290556 400250 290608 400256
rect 290464 400240 290516 400246
rect 290464 400182 290516 400188
rect 277676 399832 277728 399838
rect 268120 399758 268594 399786
rect 277728 399780 278070 399786
rect 277676 399774 278070 399780
rect 277688 399758 278070 399774
rect 285048 399770 285430 399786
rect 285036 399764 285430 399770
rect 285088 399758 285430 399764
rect 285036 399706 285088 399712
rect 288360 399634 288558 399650
rect 288348 399628 288558 399634
rect 288400 399622 288558 399628
rect 288348 399570 288400 399576
rect 282460 399560 282512 399566
rect 285588 399560 285640 399566
rect 282512 399508 282762 399514
rect 282460 399502 282762 399508
rect 285640 399508 285982 399514
rect 285588 399502 285982 399508
rect 240322 399463 240378 399472
rect 264980 399492 265032 399498
rect 282472 399486 282762 399502
rect 285600 399486 285982 399502
rect 264980 399434 265032 399440
rect 231582 399392 231638 399401
rect 231242 399350 231582 399378
rect 232962 399392 233018 399401
rect 232806 399350 232962 399378
rect 231582 399327 231638 399336
rect 232962 399327 233018 399336
rect 234066 399392 234122 399401
rect 237194 399392 237250 399401
rect 234122 399350 234370 399378
rect 237038 399350 237194 399378
rect 234066 399327 234122 399336
rect 237838 399392 237894 399401
rect 237590 399350 237838 399378
rect 237194 399327 237250 399336
rect 239402 399392 239458 399401
rect 239154 399350 239402 399378
rect 237838 399327 237894 399336
rect 240966 399392 241022 399401
rect 240718 399350 240966 399378
rect 239402 399327 239458 399336
rect 283010 399392 283066 399401
rect 281920 399362 282302 399378
rect 240966 399327 241022 399336
rect 281908 399356 282302 399362
rect 281960 399350 282302 399356
rect 284482 399392 284538 399401
rect 283066 399350 283314 399378
rect 283010 399327 283066 399336
rect 286138 399392 286194 399401
rect 284538 399350 284878 399378
rect 284482 399327 284538 399336
rect 287794 399392 287850 399401
rect 286194 399350 286442 399378
rect 286138 399327 286194 399336
rect 287850 399350 288098 399378
rect 288728 399362 289110 399378
rect 288716 399356 289110 399362
rect 287794 399327 287850 399336
rect 281908 399298 281960 399304
rect 288768 399350 289110 399356
rect 288716 399298 288768 399304
rect 229112 399214 230230 399242
rect 228364 337204 228416 337210
rect 228364 337146 228416 337152
rect 227628 336524 227680 336530
rect 227628 336466 227680 336472
rect 227168 295316 227220 295322
rect 227168 295258 227220 295264
rect 227076 136604 227128 136610
rect 227076 136546 227128 136552
rect 226984 11756 227036 11762
rect 226984 11698 227036 11704
rect 227640 3346 227668 336466
rect 228376 14482 228404 337146
rect 229008 335164 229060 335170
rect 229008 335106 229060 335112
rect 228364 14476 228416 14482
rect 228364 14418 228416 14424
rect 228916 11756 228968 11762
rect 228916 11698 228968 11704
rect 227720 4208 227772 4214
rect 227720 4150 227772 4156
rect 220556 3318 220768 3346
rect 221752 3318 222148 3346
rect 222948 3318 223528 3346
rect 224144 3318 224908 3346
rect 225340 3318 226288 3346
rect 226536 3318 227668 3346
rect 220556 480 220584 3318
rect 221752 480 221780 3318
rect 222948 480 222976 3318
rect 224144 480 224172 3318
rect 225340 480 225368 3318
rect 226536 480 226564 3318
rect 227732 480 227760 4150
rect 228928 480 228956 11698
rect 229020 4214 229048 335106
rect 229112 17950 229140 399214
rect 290476 346390 290504 400182
rect 290568 369850 290596 400250
rect 290648 400036 290700 400042
rect 290648 399978 290700 399984
rect 290660 393310 290688 399978
rect 290648 393304 290700 393310
rect 290648 393246 290700 393252
rect 290556 369844 290608 369850
rect 290556 369786 290608 369792
rect 290464 346384 290516 346390
rect 290464 346326 290516 346332
rect 270696 340190 270802 340218
rect 229204 340054 230046 340082
rect 229100 17944 229152 17950
rect 229100 17886 229152 17892
rect 229204 5030 229232 340054
rect 230124 335730 230152 340068
rect 229296 335702 230152 335730
rect 230216 335714 230244 340068
rect 230204 335708 230256 335714
rect 229192 5024 229244 5030
rect 229192 4966 229244 4972
rect 229296 4826 229324 335702
rect 230204 335650 230256 335656
rect 229376 335640 229428 335646
rect 229376 335582 229428 335588
rect 229388 4962 229416 335582
rect 230308 334218 230336 340068
rect 230492 337414 230520 340068
rect 230480 337408 230532 337414
rect 230480 337350 230532 337356
rect 230388 337000 230440 337006
rect 230388 336942 230440 336948
rect 230296 334212 230348 334218
rect 230296 334154 230348 334160
rect 230400 334098 230428 336942
rect 229756 334070 230428 334098
rect 229560 328500 229612 328506
rect 229560 328442 229612 328448
rect 229572 318782 229600 328442
rect 229756 319530 229784 334070
rect 230388 332308 230440 332314
rect 230388 332250 230440 332256
rect 229744 319524 229796 319530
rect 229744 319466 229796 319472
rect 229560 318776 229612 318782
rect 229560 318718 229612 318724
rect 229468 309256 229520 309262
rect 229468 309198 229520 309204
rect 229480 309126 229508 309198
rect 229468 309120 229520 309126
rect 229468 309062 229520 309068
rect 229560 299532 229612 299538
rect 229560 299474 229612 299480
rect 229572 294522 229600 299474
rect 229572 294494 229692 294522
rect 229664 282826 229692 294494
rect 229572 282798 229692 282826
rect 229572 280158 229600 282798
rect 229560 280152 229612 280158
rect 229560 280094 229612 280100
rect 229652 270564 229704 270570
rect 229652 270506 229704 270512
rect 229664 263514 229692 270506
rect 229572 263486 229692 263514
rect 229572 260846 229600 263486
rect 229560 260840 229612 260846
rect 229560 260782 229612 260788
rect 229652 251252 229704 251258
rect 229652 251194 229704 251200
rect 229664 244202 229692 251194
rect 229572 244174 229692 244202
rect 229572 241505 229600 244174
rect 229558 241496 229614 241505
rect 229558 241431 229614 241440
rect 229834 241496 229890 241505
rect 229834 241431 229890 241440
rect 229848 231878 229876 241431
rect 229652 231872 229704 231878
rect 229652 231814 229704 231820
rect 229836 231872 229888 231878
rect 229836 231814 229888 231820
rect 229664 224890 229692 231814
rect 229572 224862 229692 224890
rect 229572 222193 229600 224862
rect 229558 222184 229614 222193
rect 229558 222119 229614 222128
rect 229834 222184 229890 222193
rect 229834 222119 229890 222128
rect 229848 212566 229876 222119
rect 229652 212560 229704 212566
rect 229652 212502 229704 212508
rect 229836 212560 229888 212566
rect 229836 212502 229888 212508
rect 229664 205578 229692 212502
rect 229572 205550 229692 205578
rect 229572 202881 229600 205550
rect 229558 202872 229614 202881
rect 229558 202807 229614 202816
rect 229834 202872 229890 202881
rect 229834 202807 229890 202816
rect 229848 193254 229876 202807
rect 229652 193248 229704 193254
rect 229652 193190 229704 193196
rect 229836 193248 229888 193254
rect 229836 193190 229888 193196
rect 229664 186266 229692 193190
rect 229572 186238 229692 186266
rect 229572 183569 229600 186238
rect 229558 183560 229614 183569
rect 229558 183495 229614 183504
rect 229834 183560 229890 183569
rect 229834 183495 229890 183504
rect 229848 173942 229876 183495
rect 229652 173936 229704 173942
rect 229652 173878 229704 173884
rect 229836 173936 229888 173942
rect 229836 173878 229888 173884
rect 229664 166954 229692 173878
rect 229572 166926 229692 166954
rect 229572 164218 229600 166926
rect 229560 164212 229612 164218
rect 229560 164154 229612 164160
rect 229836 164212 229888 164218
rect 229836 164154 229888 164160
rect 229848 154601 229876 164154
rect 229650 154592 229706 154601
rect 229650 154527 229706 154536
rect 229834 154592 229890 154601
rect 229834 154527 229890 154536
rect 229664 147642 229692 154527
rect 229572 147614 229692 147642
rect 229572 138038 229600 147614
rect 229560 138032 229612 138038
rect 229560 137974 229612 137980
rect 229468 137964 229520 137970
rect 229468 137906 229520 137912
rect 229480 135289 229508 137906
rect 229466 135280 229522 135289
rect 229466 135215 229522 135224
rect 229650 135280 229706 135289
rect 229650 135215 229706 135224
rect 229664 128330 229692 135215
rect 229572 128302 229692 128330
rect 229572 118726 229600 128302
rect 229560 118720 229612 118726
rect 229560 118662 229612 118668
rect 229468 118652 229520 118658
rect 229468 118594 229520 118600
rect 229480 115977 229508 118594
rect 229466 115968 229522 115977
rect 229466 115903 229522 115912
rect 229650 115968 229706 115977
rect 229650 115903 229706 115912
rect 229664 109018 229692 115903
rect 229572 108990 229692 109018
rect 229572 99414 229600 108990
rect 229560 99408 229612 99414
rect 229560 99350 229612 99356
rect 229468 99340 229520 99346
rect 229468 99282 229520 99288
rect 229480 96665 229508 99282
rect 229466 96656 229522 96665
rect 229466 96591 229522 96600
rect 229650 96656 229706 96665
rect 229650 96591 229706 96600
rect 229664 89706 229692 96591
rect 229572 89678 229692 89706
rect 229572 80170 229600 89678
rect 229560 80164 229612 80170
rect 229560 80106 229612 80112
rect 229468 77376 229520 77382
rect 229520 77324 229600 77330
rect 229468 77318 229600 77324
rect 229480 77302 229600 77318
rect 229572 77246 229600 77302
rect 229560 77240 229612 77246
rect 229560 77182 229612 77188
rect 229652 67652 229704 67658
rect 229652 67594 229704 67600
rect 229664 67561 229692 67594
rect 229650 67552 229706 67561
rect 229650 67487 229706 67496
rect 229650 58032 229706 58041
rect 229650 57967 229706 57976
rect 229664 57934 229692 57967
rect 229652 57928 229704 57934
rect 229652 57870 229704 57876
rect 229560 48340 229612 48346
rect 229560 48282 229612 48288
rect 229572 41426 229600 48282
rect 229480 41410 229600 41426
rect 229468 41404 229600 41410
rect 229520 41398 229600 41404
rect 229652 41404 229704 41410
rect 229468 41346 229520 41352
rect 229652 41346 229704 41352
rect 229664 38622 229692 41346
rect 229652 38616 229704 38622
rect 229652 38558 229704 38564
rect 229560 29028 229612 29034
rect 229560 28970 229612 28976
rect 229572 22166 229600 28970
rect 229560 22160 229612 22166
rect 229560 22102 229612 22108
rect 229560 22024 229612 22030
rect 229560 21966 229612 21972
rect 229572 10334 229600 21966
rect 229560 10328 229612 10334
rect 229560 10270 229612 10276
rect 229376 4956 229428 4962
rect 229376 4898 229428 4904
rect 229284 4820 229336 4826
rect 229284 4762 229336 4768
rect 229008 4208 229060 4214
rect 229008 4150 229060 4156
rect 229100 3324 229152 3330
rect 229100 3266 229152 3272
rect 229112 3233 229140 3266
rect 229098 3224 229154 3233
rect 229098 3159 229154 3168
rect 230400 610 230428 332250
rect 230584 3369 230612 340068
rect 230690 340054 230796 340082
rect 230664 335640 230716 335646
rect 230664 335582 230716 335588
rect 230676 3505 230704 335582
rect 230768 4622 230796 340054
rect 230860 333282 230888 340068
rect 230952 337482 230980 340068
rect 231044 337550 231072 340068
rect 231136 340054 231242 340082
rect 231032 337544 231084 337550
rect 231032 337486 231084 337492
rect 230940 337476 230992 337482
rect 230940 337418 230992 337424
rect 231136 333282 231164 340054
rect 230860 333254 230980 333282
rect 230848 205692 230900 205698
rect 230848 205634 230900 205640
rect 230860 195974 230888 205634
rect 230848 195968 230900 195974
rect 230848 195910 230900 195916
rect 230848 186380 230900 186386
rect 230848 186322 230900 186328
rect 230860 176662 230888 186322
rect 230848 176656 230900 176662
rect 230848 176598 230900 176604
rect 230848 167068 230900 167074
rect 230848 167010 230900 167016
rect 230860 157350 230888 167010
rect 230848 157344 230900 157350
rect 230848 157286 230900 157292
rect 230848 51128 230900 51134
rect 230848 51070 230900 51076
rect 230860 41410 230888 51070
rect 230848 41404 230900 41410
rect 230848 41346 230900 41352
rect 230848 31816 230900 31822
rect 230848 31758 230900 31764
rect 230860 22098 230888 31758
rect 230848 22092 230900 22098
rect 230848 22034 230900 22040
rect 230848 12504 230900 12510
rect 230848 12446 230900 12452
rect 230860 6186 230888 12446
rect 230952 10402 230980 333254
rect 231044 333254 231164 333282
rect 231044 205698 231072 333254
rect 231320 331906 231348 340068
rect 231412 335646 231440 340068
rect 231504 340054 231610 340082
rect 231400 335640 231452 335646
rect 231400 335582 231452 335588
rect 231308 331900 231360 331906
rect 231308 331842 231360 331848
rect 231504 331786 231532 340054
rect 231688 333946 231716 340068
rect 231676 333940 231728 333946
rect 231676 333882 231728 333888
rect 231676 333804 231728 333810
rect 231676 333746 231728 333752
rect 231584 333192 231636 333198
rect 231584 333134 231636 333140
rect 231136 331758 231532 331786
rect 231032 205692 231084 205698
rect 231032 205634 231084 205640
rect 231032 195968 231084 195974
rect 231032 195910 231084 195916
rect 231044 186386 231072 195910
rect 231032 186380 231084 186386
rect 231032 186322 231084 186328
rect 231032 176656 231084 176662
rect 231032 176598 231084 176604
rect 231044 167074 231072 176598
rect 231032 167068 231084 167074
rect 231032 167010 231084 167016
rect 231032 157344 231084 157350
rect 231032 157286 231084 157292
rect 231044 51134 231072 157286
rect 231032 51128 231084 51134
rect 231032 51070 231084 51076
rect 231032 41404 231084 41410
rect 231032 41346 231084 41352
rect 231044 31822 231072 41346
rect 231032 31816 231084 31822
rect 231032 31758 231084 31764
rect 231032 22092 231084 22098
rect 231032 22034 231084 22040
rect 231044 12510 231072 22034
rect 231032 12504 231084 12510
rect 231032 12446 231084 12452
rect 230940 10396 230992 10402
rect 230940 10338 230992 10344
rect 230848 6180 230900 6186
rect 230848 6122 230900 6128
rect 230756 4616 230808 4622
rect 230756 4558 230808 4564
rect 231136 3641 231164 331758
rect 231596 328438 231624 333134
rect 231584 328432 231636 328438
rect 231584 328374 231636 328380
rect 231492 318844 231544 318850
rect 231492 318786 231544 318792
rect 231504 318730 231532 318786
rect 231504 318702 231624 318730
rect 231596 315314 231624 318702
rect 231584 315308 231636 315314
rect 231584 315250 231636 315256
rect 231688 8974 231716 333746
rect 231780 333198 231808 340068
rect 231964 337754 231992 340068
rect 231952 337748 232004 337754
rect 231952 337690 232004 337696
rect 232056 337618 232084 340068
rect 232044 337612 232096 337618
rect 232044 337554 232096 337560
rect 231952 337136 232004 337142
rect 231952 337078 232004 337084
rect 231768 333192 231820 333198
rect 231768 333134 231820 333140
rect 231964 331974 231992 337078
rect 232044 336048 232096 336054
rect 232044 335990 232096 335996
rect 232056 333962 232084 335990
rect 232148 334082 232176 340068
rect 232228 335980 232280 335986
rect 232228 335922 232280 335928
rect 232240 335458 232268 335922
rect 232332 335594 232360 340068
rect 232424 335730 232452 340068
rect 232530 340054 232636 340082
rect 232608 335866 232636 340054
rect 232700 336054 232728 340068
rect 232688 336048 232740 336054
rect 232688 335990 232740 335996
rect 232792 335986 232820 340068
rect 232884 337686 232912 340068
rect 232872 337680 232924 337686
rect 232872 337622 232924 337628
rect 232780 335980 232832 335986
rect 232780 335922 232832 335928
rect 232608 335838 233004 335866
rect 232424 335702 232820 335730
rect 232332 335566 232452 335594
rect 232240 335430 232360 335458
rect 232136 334076 232188 334082
rect 232136 334018 232188 334024
rect 232056 333934 232176 333962
rect 232044 333872 232096 333878
rect 232044 333814 232096 333820
rect 231952 331968 232004 331974
rect 231952 331910 232004 331916
rect 232056 10470 232084 333814
rect 232148 10538 232176 333934
rect 232228 333192 232280 333198
rect 232228 333134 232280 333140
rect 232240 10606 232268 333134
rect 232332 309806 232360 335430
rect 232424 313954 232452 335566
rect 232412 313948 232464 313954
rect 232412 313890 232464 313896
rect 232320 309800 232372 309806
rect 232320 309742 232372 309748
rect 232228 10600 232280 10606
rect 232228 10542 232280 10548
rect 232136 10532 232188 10538
rect 232136 10474 232188 10480
rect 232044 10464 232096 10470
rect 232044 10406 232096 10412
rect 231768 10328 231820 10334
rect 231768 10270 231820 10276
rect 231676 8968 231728 8974
rect 231676 8910 231728 8916
rect 231122 3632 231178 3641
rect 231122 3567 231178 3576
rect 231780 3534 231808 10270
rect 232792 3777 232820 335702
rect 232976 3913 233004 335838
rect 233068 333198 233096 340068
rect 233056 333192 233108 333198
rect 233056 333134 233108 333140
rect 233160 312594 233188 340068
rect 233252 336938 233280 340068
rect 233344 340054 233450 340082
rect 233240 336932 233292 336938
rect 233240 336874 233292 336880
rect 233240 336796 233292 336802
rect 233240 336738 233292 336744
rect 233252 335918 233280 336738
rect 233240 335912 233292 335918
rect 233240 335854 233292 335860
rect 233344 335594 233372 340054
rect 233528 335968 233556 340068
rect 233620 337822 233648 340068
rect 233712 340054 233818 340082
rect 233608 337816 233660 337822
rect 233608 337758 233660 337764
rect 233528 335940 233648 335968
rect 233516 335844 233568 335850
rect 233516 335786 233568 335792
rect 233252 335566 233372 335594
rect 233252 329118 233280 335566
rect 233332 335504 233384 335510
rect 233332 335446 233384 335452
rect 233240 329112 233292 329118
rect 233240 329054 233292 329060
rect 233344 324970 233372 335446
rect 233528 327758 233556 335786
rect 233620 335730 233648 335940
rect 233712 335850 233740 340054
rect 233700 335844 233752 335850
rect 233700 335786 233752 335792
rect 233620 335702 233740 335730
rect 233608 333736 233660 333742
rect 233608 333678 233660 333684
rect 233516 327752 233568 327758
rect 233516 327694 233568 327700
rect 233620 327078 233648 333678
rect 233608 327072 233660 327078
rect 233608 327014 233660 327020
rect 233332 324964 233384 324970
rect 233332 324906 233384 324912
rect 233516 317484 233568 317490
rect 233516 317426 233568 317432
rect 233148 312588 233200 312594
rect 233148 312530 233200 312536
rect 233528 309126 233556 317426
rect 233516 309120 233568 309126
rect 233516 309062 233568 309068
rect 233712 307086 233740 335702
rect 233896 333742 233924 340068
rect 234002 340054 234108 340082
rect 233884 333736 233936 333742
rect 233884 333678 233936 333684
rect 233884 333192 233936 333198
rect 233884 333134 233936 333140
rect 234080 333146 234108 340054
rect 234172 335510 234200 340068
rect 234160 335504 234212 335510
rect 234160 335446 234212 335452
rect 233896 320890 233924 333134
rect 234080 333118 234200 333146
rect 234068 332444 234120 332450
rect 234068 332386 234120 332392
rect 233884 320884 233936 320890
rect 233884 320826 233936 320832
rect 233700 307080 233752 307086
rect 233700 307022 233752 307028
rect 233148 10396 233200 10402
rect 233148 10338 233200 10344
rect 232962 3904 233018 3913
rect 232962 3839 233018 3848
rect 232778 3768 232834 3777
rect 232778 3703 232834 3712
rect 233160 3534 233188 10338
rect 233700 4820 233752 4826
rect 233700 4762 233752 4768
rect 231308 3528 231360 3534
rect 230662 3496 230718 3505
rect 230662 3431 230718 3440
rect 230938 3496 230994 3505
rect 231308 3470 231360 3476
rect 231768 3528 231820 3534
rect 231768 3470 231820 3476
rect 232504 3528 232556 3534
rect 232504 3470 232556 3476
rect 233148 3528 233200 3534
rect 233240 3528 233292 3534
rect 233148 3470 233200 3476
rect 233238 3496 233240 3505
rect 233292 3496 233294 3505
rect 230938 3431 230994 3440
rect 230952 3398 230980 3431
rect 230940 3392 230992 3398
rect 230570 3360 230626 3369
rect 230940 3334 230992 3340
rect 230570 3295 230626 3304
rect 230112 604 230164 610
rect 230112 546 230164 552
rect 230388 604 230440 610
rect 230388 546 230440 552
rect 230124 480 230152 546
rect 231320 480 231348 3470
rect 232516 480 232544 3470
rect 233238 3431 233294 3440
rect 233712 480 233740 4762
rect 234080 3602 234108 332386
rect 234068 3596 234120 3602
rect 234068 3538 234120 3544
rect 234172 3330 234200 333118
rect 234264 304298 234292 340068
rect 234356 332450 234384 340068
rect 234436 336932 234488 336938
rect 234436 336874 234488 336880
rect 234344 332444 234396 332450
rect 234344 332386 234396 332392
rect 234252 304292 234304 304298
rect 234252 304234 234304 304240
rect 234448 4049 234476 336874
rect 234540 323610 234568 340068
rect 234632 333130 234660 340068
rect 234738 340054 234844 340082
rect 234816 333282 234844 340054
rect 234908 337142 234936 340068
rect 234896 337136 234948 337142
rect 234896 337078 234948 337084
rect 234724 333254 234844 333282
rect 235000 333266 235028 340068
rect 234988 333260 235040 333266
rect 234620 333124 234672 333130
rect 234620 333066 234672 333072
rect 234528 323604 234580 323610
rect 234528 323546 234580 323552
rect 234434 4040 234490 4049
rect 234434 3975 234490 3984
rect 234724 3398 234752 333254
rect 234988 333202 235040 333208
rect 234988 333124 235040 333130
rect 234988 333066 235040 333072
rect 235000 319462 235028 333066
rect 234988 319456 235040 319462
rect 234988 319398 235040 319404
rect 235092 302938 235120 340068
rect 235276 336802 235304 340068
rect 235264 336796 235316 336802
rect 235264 336738 235316 336744
rect 235172 332988 235224 332994
rect 235172 332930 235224 332936
rect 235080 302932 235132 302938
rect 235080 302874 235132 302880
rect 234804 6180 234856 6186
rect 234804 6122 234856 6128
rect 234712 3392 234764 3398
rect 234712 3334 234764 3340
rect 234160 3324 234212 3330
rect 234160 3266 234212 3272
rect 233792 3256 233844 3262
rect 233790 3224 233792 3233
rect 233844 3224 233846 3233
rect 233790 3159 233846 3168
rect 234816 480 234844 6122
rect 235184 3670 235212 332930
rect 235368 326398 235396 340068
rect 235460 332994 235488 340068
rect 235644 334626 235672 340068
rect 235632 334620 235684 334626
rect 235632 334562 235684 334568
rect 235736 333282 235764 340068
rect 235644 333254 235764 333282
rect 235448 332988 235500 332994
rect 235448 332930 235500 332936
rect 235356 326392 235408 326398
rect 235356 326334 235408 326340
rect 235644 322250 235672 333254
rect 235632 322244 235684 322250
rect 235632 322186 235684 322192
rect 235828 4078 235856 340068
rect 236012 335510 236040 340068
rect 236104 335646 236132 340068
rect 236092 335640 236144 335646
rect 236092 335582 236144 335588
rect 236000 335504 236052 335510
rect 236000 335446 236052 335452
rect 236196 333962 236224 340068
rect 236276 336116 236328 336122
rect 236276 336058 236328 336064
rect 236104 333934 236224 333962
rect 236000 10464 236052 10470
rect 236000 10406 236052 10412
rect 235816 4072 235868 4078
rect 235816 4014 235868 4020
rect 235172 3664 235224 3670
rect 235172 3606 235224 3612
rect 236012 480 236040 10406
rect 236104 3806 236132 333934
rect 236288 333826 236316 336058
rect 236380 335714 236408 340068
rect 236472 335782 236500 340068
rect 236564 336122 236592 340068
rect 236656 340054 236762 340082
rect 236552 336116 236604 336122
rect 236552 336058 236604 336064
rect 236656 335866 236684 340054
rect 236840 337006 236868 340068
rect 236828 337000 236880 337006
rect 236828 336942 236880 336948
rect 236564 335838 236684 335866
rect 236460 335776 236512 335782
rect 236460 335718 236512 335724
rect 236368 335708 236420 335714
rect 236368 335650 236420 335656
rect 236564 335594 236592 335838
rect 236736 335776 236788 335782
rect 236736 335718 236788 335724
rect 236644 335708 236696 335714
rect 236644 335650 236696 335656
rect 236196 333798 236316 333826
rect 236380 335566 236592 335594
rect 236196 3874 236224 333798
rect 236276 333736 236328 333742
rect 236276 333678 236328 333684
rect 236288 3942 236316 333678
rect 236380 9178 236408 335566
rect 236460 335504 236512 335510
rect 236460 335446 236512 335452
rect 236368 9172 236420 9178
rect 236368 9114 236420 9120
rect 236472 9042 236500 335446
rect 236656 9110 236684 335650
rect 236748 10742 236776 335718
rect 236828 335640 236880 335646
rect 236828 335582 236880 335588
rect 236736 10736 236788 10742
rect 236736 10678 236788 10684
rect 236840 10674 236868 335582
rect 236932 333742 236960 340068
rect 236920 333736 236972 333742
rect 236920 333678 236972 333684
rect 237012 331288 237064 331294
rect 237012 331230 237064 331236
rect 236828 10668 236880 10674
rect 236828 10610 236880 10616
rect 236644 9104 236696 9110
rect 236644 9046 236696 9052
rect 236460 9036 236512 9042
rect 236460 8978 236512 8984
rect 237024 4010 237052 331230
rect 237116 9246 237144 340068
rect 237208 330546 237236 340068
rect 237300 331294 237328 340068
rect 237484 333010 237512 340068
rect 237576 333198 237604 340068
rect 237682 340054 237788 340082
rect 237760 335782 237788 340054
rect 237748 335776 237800 335782
rect 237748 335718 237800 335724
rect 237748 335640 237800 335646
rect 237748 335582 237800 335588
rect 237564 333192 237616 333198
rect 237564 333134 237616 333140
rect 237484 332982 237696 333010
rect 237288 331288 237340 331294
rect 237288 331230 237340 331236
rect 237196 330540 237248 330546
rect 237196 330482 237248 330488
rect 237668 327078 237696 332982
rect 237656 327072 237708 327078
rect 237656 327014 237708 327020
rect 237564 317484 237616 317490
rect 237564 317426 237616 317432
rect 237576 309126 237604 317426
rect 237564 309120 237616 309126
rect 237564 309062 237616 309068
rect 237656 309052 237708 309058
rect 237656 308994 237708 309000
rect 237668 298110 237696 308994
rect 237656 298104 237708 298110
rect 237656 298046 237708 298052
rect 237564 288448 237616 288454
rect 237564 288390 237616 288396
rect 237576 282826 237604 288390
rect 237576 282798 237696 282826
rect 237668 278769 237696 282798
rect 237654 278760 237710 278769
rect 237654 278695 237710 278704
rect 237654 264344 237710 264353
rect 237654 264279 237710 264288
rect 237668 259622 237696 264279
rect 237656 259616 237708 259622
rect 237656 259558 237708 259564
rect 237656 259480 237708 259486
rect 237656 259422 237708 259428
rect 237668 254046 237696 259422
rect 237656 254040 237708 254046
rect 237656 253982 237708 253988
rect 237564 253904 237616 253910
rect 237564 253846 237616 253852
rect 237576 248402 237604 253846
rect 237564 248396 237616 248402
rect 237564 248338 237616 248344
rect 237656 244180 237708 244186
rect 237656 244122 237708 244128
rect 237668 232014 237696 244122
rect 237656 232008 237708 232014
rect 237656 231950 237708 231956
rect 237472 227792 237524 227798
rect 237472 227734 237524 227740
rect 237484 219473 237512 227734
rect 237470 219464 237526 219473
rect 237470 219399 237526 219408
rect 237654 219464 237710 219473
rect 237654 219399 237710 219408
rect 237668 219366 237696 219399
rect 237656 219360 237708 219366
rect 237656 219302 237708 219308
rect 237656 214600 237708 214606
rect 237656 214542 237708 214548
rect 237668 201482 237696 214542
rect 237564 201476 237616 201482
rect 237564 201418 237616 201424
rect 237656 201476 237708 201482
rect 237656 201418 237708 201424
rect 237576 186386 237604 201418
rect 237564 186380 237616 186386
rect 237564 186322 237616 186328
rect 237656 186244 237708 186250
rect 237656 186186 237708 186192
rect 237668 174010 237696 186186
rect 237564 174004 237616 174010
rect 237564 173946 237616 173952
rect 237656 174004 237708 174010
rect 237656 173946 237708 173952
rect 237576 172514 237604 173946
rect 237564 172508 237616 172514
rect 237564 172450 237616 172456
rect 237564 167000 237616 167006
rect 237564 166942 237616 166948
rect 237576 162874 237604 166942
rect 237576 162858 237696 162874
rect 237564 162852 237708 162858
rect 237616 162846 237656 162852
rect 237564 162794 237616 162800
rect 237656 162794 237708 162800
rect 237576 153377 237604 162794
rect 237562 153368 237618 153377
rect 237562 153303 237618 153312
rect 237562 153232 237618 153241
rect 237562 153167 237564 153176
rect 237616 153167 237618 153176
rect 237564 153138 237616 153144
rect 237564 147620 237616 147626
rect 237564 147562 237616 147568
rect 237576 143562 237604 147562
rect 237576 143534 237696 143562
rect 237668 143478 237696 143534
rect 237656 143472 237708 143478
rect 237656 143414 237708 143420
rect 237564 134020 237616 134026
rect 237564 133962 237616 133968
rect 237576 124409 237604 133962
rect 237562 124400 237618 124409
rect 237562 124335 237618 124344
rect 237654 124264 237710 124273
rect 237654 124199 237710 124208
rect 237668 113218 237696 124199
rect 237564 113212 237616 113218
rect 237564 113154 237616 113160
rect 237656 113212 237708 113218
rect 237656 113154 237708 113160
rect 237576 113098 237604 113154
rect 237576 113070 237696 113098
rect 237668 99414 237696 113070
rect 237656 99408 237708 99414
rect 237656 99350 237708 99356
rect 237564 99340 237616 99346
rect 237564 99282 237616 99288
rect 237576 95198 237604 99282
rect 237564 95192 237616 95198
rect 237564 95134 237616 95140
rect 237656 85604 237708 85610
rect 237656 85546 237708 85552
rect 237668 82822 237696 85546
rect 237656 82816 237708 82822
rect 237656 82758 237708 82764
rect 237564 73228 237616 73234
rect 237564 73170 237616 73176
rect 237576 66366 237604 73170
rect 237564 66360 237616 66366
rect 237564 66302 237616 66308
rect 237472 66224 237524 66230
rect 237472 66166 237524 66172
rect 237484 64818 237512 66166
rect 237484 64790 237696 64818
rect 237668 56522 237696 64790
rect 237484 56494 237696 56522
rect 237484 46986 237512 56494
rect 237472 46980 237524 46986
rect 237472 46922 237524 46928
rect 237564 46980 237616 46986
rect 237564 46922 237616 46928
rect 237576 45558 237604 46922
rect 237564 45552 237616 45558
rect 237564 45494 237616 45500
rect 237656 35964 237708 35970
rect 237656 35906 237708 35912
rect 237668 19378 237696 35906
rect 237564 19372 237616 19378
rect 237564 19314 237616 19320
rect 237656 19372 237708 19378
rect 237656 19314 237708 19320
rect 237576 16590 237604 19314
rect 237564 16584 237616 16590
rect 237564 16526 237616 16532
rect 237760 9450 237788 335582
rect 237748 9444 237800 9450
rect 237748 9386 237800 9392
rect 237852 9382 237880 340068
rect 237944 329186 237972 340068
rect 237932 329180 237984 329186
rect 237932 329122 237984 329128
rect 237840 9376 237892 9382
rect 237840 9318 237892 9324
rect 237104 9240 237156 9246
rect 237104 9182 237156 9188
rect 237288 4888 237340 4894
rect 237288 4830 237340 4836
rect 237012 4004 237064 4010
rect 237012 3946 237064 3952
rect 236276 3936 236328 3942
rect 236276 3878 236328 3884
rect 236184 3868 236236 3874
rect 236184 3810 236236 3816
rect 236092 3800 236144 3806
rect 236092 3742 236144 3748
rect 237300 2530 237328 4830
rect 238036 4146 238064 340068
rect 238128 340054 238234 340082
rect 238128 335646 238156 340054
rect 238116 335640 238168 335646
rect 238116 335582 238168 335588
rect 238116 329792 238168 329798
rect 238116 329734 238168 329740
rect 238128 302326 238156 329734
rect 238312 327826 238340 340068
rect 238404 329798 238432 340068
rect 238484 335776 238536 335782
rect 238484 335718 238536 335724
rect 238392 329792 238444 329798
rect 238392 329734 238444 329740
rect 238300 327820 238352 327826
rect 238300 327762 238352 327768
rect 238116 302320 238168 302326
rect 238116 302262 238168 302268
rect 238208 302116 238260 302122
rect 238208 302058 238260 302064
rect 238220 289814 238248 302058
rect 238116 289808 238168 289814
rect 238116 289750 238168 289756
rect 238208 289808 238260 289814
rect 238208 289750 238260 289756
rect 238128 285002 238156 289750
rect 238128 284974 238248 285002
rect 238220 273306 238248 284974
rect 238128 273278 238248 273306
rect 238128 273170 238156 273278
rect 238128 273142 238248 273170
rect 238220 253994 238248 273142
rect 238128 253966 238248 253994
rect 238128 253858 238156 253966
rect 238128 253830 238248 253858
rect 238220 244338 238248 253830
rect 238220 244310 238340 244338
rect 238312 238921 238340 244310
rect 238298 238912 238354 238921
rect 238298 238847 238354 238856
rect 238114 238776 238170 238785
rect 238114 238711 238170 238720
rect 238128 237386 238156 238711
rect 238116 237380 238168 237386
rect 238116 237322 238168 237328
rect 238300 237380 238352 237386
rect 238300 237322 238352 237328
rect 238312 214554 238340 237322
rect 238220 214526 238340 214554
rect 238220 176610 238248 214526
rect 238128 176582 238248 176610
rect 238128 176338 238156 176582
rect 238128 176310 238248 176338
rect 238220 172514 238248 176310
rect 238208 172508 238260 172514
rect 238208 172450 238260 172456
rect 238208 162920 238260 162926
rect 238208 162862 238260 162868
rect 238220 153202 238248 162862
rect 238208 153196 238260 153202
rect 238208 153138 238260 153144
rect 238208 143608 238260 143614
rect 238208 143550 238260 143556
rect 238220 133906 238248 143550
rect 238128 133890 238248 133906
rect 238116 133884 238248 133890
rect 238168 133878 238248 133884
rect 238116 133826 238168 133832
rect 238128 133795 238156 133826
rect 238116 122868 238168 122874
rect 238116 122810 238168 122816
rect 238128 121446 238156 122810
rect 238116 121440 238168 121446
rect 238116 121382 238168 121388
rect 238116 113144 238168 113150
rect 238116 113086 238168 113092
rect 238128 103562 238156 113086
rect 238116 103556 238168 103562
rect 238116 103498 238168 103504
rect 238208 103556 238260 103562
rect 238208 103498 238260 103504
rect 238220 102134 238248 103498
rect 238208 102128 238260 102134
rect 238208 102070 238260 102076
rect 238116 92540 238168 92546
rect 238116 92482 238168 92488
rect 238128 85610 238156 92482
rect 238116 85604 238168 85610
rect 238116 85546 238168 85552
rect 238208 85604 238260 85610
rect 238208 85546 238260 85552
rect 238220 80186 238248 85546
rect 238128 80158 238248 80186
rect 238128 80050 238156 80158
rect 238128 80022 238248 80050
rect 238220 69034 238248 80022
rect 238128 69006 238248 69034
rect 238128 67640 238156 69006
rect 238128 67612 238248 67640
rect 238220 64870 238248 67612
rect 238208 64864 238260 64870
rect 238208 64806 238260 64812
rect 238208 55276 238260 55282
rect 238208 55218 238260 55224
rect 238220 51134 238248 55218
rect 238208 51128 238260 51134
rect 238208 51070 238260 51076
rect 238208 46980 238260 46986
rect 238208 46922 238260 46928
rect 238220 45558 238248 46922
rect 238208 45552 238260 45558
rect 238208 45494 238260 45500
rect 238208 36032 238260 36038
rect 238208 35974 238260 35980
rect 238220 35902 238248 35974
rect 238208 35896 238260 35902
rect 238208 35838 238260 35844
rect 238116 26308 238168 26314
rect 238116 26250 238168 26256
rect 238024 4140 238076 4146
rect 238024 4082 238076 4088
rect 238128 3602 238156 26250
rect 238392 6044 238444 6050
rect 238392 5986 238444 5992
rect 238116 3596 238168 3602
rect 238116 3538 238168 3544
rect 237208 2502 237328 2530
rect 237208 480 237236 2502
rect 238404 480 238432 5986
rect 238496 3466 238524 335718
rect 238588 9518 238616 340068
rect 238680 318102 238708 340068
rect 238668 318096 238720 318102
rect 238668 318038 238720 318044
rect 238668 133884 238720 133890
rect 238668 133826 238720 133832
rect 238680 124273 238708 133826
rect 238666 124264 238722 124273
rect 238666 124199 238722 124208
rect 238576 9512 238628 9518
rect 238576 9454 238628 9460
rect 238484 3460 238536 3466
rect 238484 3402 238536 3408
rect 238772 3262 238800 340068
rect 238852 335640 238904 335646
rect 238852 335582 238904 335588
rect 238864 326466 238892 335582
rect 238956 333418 238984 340068
rect 239048 336598 239076 340068
rect 239036 336592 239088 336598
rect 239036 336534 239088 336540
rect 238956 333390 239076 333418
rect 238944 333260 238996 333266
rect 238944 333202 238996 333208
rect 238852 326460 238904 326466
rect 238852 326402 238904 326408
rect 238956 319530 238984 333202
rect 238944 319524 238996 319530
rect 238944 319466 238996 319472
rect 238944 317484 238996 317490
rect 238944 317426 238996 317432
rect 238956 309126 238984 317426
rect 238944 309120 238996 309126
rect 238944 309062 238996 309068
rect 238944 299532 238996 299538
rect 238944 299474 238996 299480
rect 238956 263650 238984 299474
rect 238864 263622 238984 263650
rect 238864 263514 238892 263622
rect 238864 263486 238984 263514
rect 238956 244338 238984 263486
rect 238864 244310 238984 244338
rect 238864 244202 238892 244310
rect 238864 244174 238984 244202
rect 238956 229090 238984 244174
rect 238944 229084 238996 229090
rect 238944 229026 238996 229032
rect 238850 219464 238906 219473
rect 238850 219399 238906 219408
rect 238864 218890 238892 219399
rect 238852 218884 238904 218890
rect 238852 218826 238904 218832
rect 238944 205352 238996 205358
rect 238944 205294 238996 205300
rect 238956 186402 238984 205294
rect 238864 186374 238984 186402
rect 238864 186266 238892 186374
rect 238864 186238 238984 186266
rect 238956 167090 238984 186238
rect 238864 167062 238984 167090
rect 238864 166954 238892 167062
rect 238864 166926 238984 166954
rect 238956 162858 238984 166926
rect 238944 162852 238996 162858
rect 238944 162794 238996 162800
rect 238942 153232 238998 153241
rect 238942 153167 238944 153176
rect 238996 153167 238998 153176
rect 238944 153138 238996 153144
rect 238944 147212 238996 147218
rect 238944 147154 238996 147160
rect 238956 133890 238984 147154
rect 238944 133884 238996 133890
rect 238944 133826 238996 133832
rect 238942 124264 238998 124273
rect 238942 124199 238998 124208
rect 238956 122890 238984 124199
rect 238864 122862 238984 122890
rect 238864 121446 238892 122862
rect 238852 121440 238904 121446
rect 238852 121382 238904 121388
rect 238852 115388 238904 115394
rect 238852 115330 238904 115336
rect 238864 106350 238892 115330
rect 238852 106344 238904 106350
rect 238852 106286 238904 106292
rect 238852 106208 238904 106214
rect 238852 106150 238904 106156
rect 238864 95198 238892 106150
rect 238852 95192 238904 95198
rect 238852 95134 238904 95140
rect 238944 95124 238996 95130
rect 238944 95066 238996 95072
rect 238956 80186 238984 95066
rect 238864 80158 238984 80186
rect 238864 74610 238892 80158
rect 238864 74582 238984 74610
rect 238956 74526 238984 74582
rect 238944 74520 238996 74526
rect 238944 74462 238996 74468
rect 238944 64932 238996 64938
rect 238944 64874 238996 64880
rect 238956 55214 238984 64874
rect 238944 55208 238996 55214
rect 238944 55150 238996 55156
rect 238944 45620 238996 45626
rect 238944 45562 238996 45568
rect 238956 38690 238984 45562
rect 238944 38684 238996 38690
rect 238944 38626 238996 38632
rect 238852 38616 238904 38622
rect 238852 38558 238904 38564
rect 238864 29034 238892 38558
rect 238852 29028 238904 29034
rect 238852 28970 238904 28976
rect 238944 29028 238996 29034
rect 238944 28970 238996 28976
rect 238956 21486 238984 28970
rect 238944 21480 238996 21486
rect 238944 21422 238996 21428
rect 238852 16652 238904 16658
rect 238852 16594 238904 16600
rect 238760 3256 238812 3262
rect 238760 3198 238812 3204
rect 238864 3194 238892 16594
rect 239048 9586 239076 333390
rect 239140 333266 239168 340068
rect 239220 333804 239272 333810
rect 239220 333746 239272 333752
rect 239128 333260 239180 333266
rect 239128 333202 239180 333208
rect 239128 229084 239180 229090
rect 239128 229026 239180 229032
rect 239140 219473 239168 229026
rect 239126 219464 239182 219473
rect 239126 219399 239182 219408
rect 239128 162852 239180 162858
rect 239128 162794 239180 162800
rect 239140 153241 239168 162794
rect 239126 153232 239182 153241
rect 239126 153167 239182 153176
rect 239036 9580 239088 9586
rect 239036 9522 239088 9528
rect 239232 8906 239260 333746
rect 239324 9654 239352 340068
rect 239416 331294 239444 340068
rect 239404 331288 239456 331294
rect 239404 331230 239456 331236
rect 239312 9648 239364 9654
rect 239312 9590 239364 9596
rect 239220 8900 239272 8906
rect 239220 8842 239272 8848
rect 238852 3188 238904 3194
rect 238852 3130 238904 3136
rect 239508 3126 239536 340068
rect 239600 340054 239706 340082
rect 239600 333810 239628 340054
rect 239784 335646 239812 340068
rect 239772 335640 239824 335646
rect 239772 335582 239824 335588
rect 239588 333804 239640 333810
rect 239588 333746 239640 333752
rect 239588 331220 239640 331226
rect 239588 331162 239640 331168
rect 239600 325038 239628 331162
rect 239588 325032 239640 325038
rect 239588 324974 239640 324980
rect 239588 3460 239640 3466
rect 239588 3402 239640 3408
rect 239496 3120 239548 3126
rect 239496 3062 239548 3068
rect 239600 480 239628 3402
rect 239876 3058 239904 340068
rect 240060 8838 240088 340068
rect 240152 333180 240180 340068
rect 240244 338094 240272 340068
rect 240232 338088 240284 338094
rect 240232 338030 240284 338036
rect 240232 336796 240284 336802
rect 240232 336738 240284 336744
rect 240244 333334 240272 336738
rect 240324 335708 240376 335714
rect 240428 335696 240456 340068
rect 240520 335850 240548 340068
rect 240626 340054 240732 340082
rect 240508 335844 240560 335850
rect 240508 335786 240560 335792
rect 240428 335668 240548 335696
rect 240324 335650 240376 335656
rect 240232 333328 240284 333334
rect 240232 333270 240284 333276
rect 240152 333152 240272 333180
rect 240244 323678 240272 333152
rect 240232 323672 240284 323678
rect 240232 323614 240284 323620
rect 240048 8832 240100 8838
rect 240048 8774 240100 8780
rect 240336 8634 240364 335650
rect 240416 335572 240468 335578
rect 240416 335514 240468 335520
rect 240428 8702 240456 335514
rect 240520 331294 240548 335668
rect 240704 335646 240732 340054
rect 240692 335640 240744 335646
rect 240692 335582 240744 335588
rect 240796 335578 240824 340068
rect 240888 338094 240916 340068
rect 240876 338088 240928 338094
rect 240876 338030 240928 338036
rect 240980 337754 241008 340068
rect 241072 340054 241178 340082
rect 240968 337748 241020 337754
rect 240968 337690 241020 337696
rect 241072 335714 241100 340054
rect 241152 337544 241204 337550
rect 241152 337486 241204 337492
rect 241060 335708 241112 335714
rect 241060 335650 241112 335656
rect 240968 335640 241020 335646
rect 240968 335582 241020 335588
rect 240784 335572 240836 335578
rect 240784 335514 240836 335520
rect 240508 331288 240560 331294
rect 240508 331230 240560 331236
rect 240508 331152 240560 331158
rect 240508 331094 240560 331100
rect 240520 67590 240548 331094
rect 240692 328500 240744 328506
rect 240692 328442 240744 328448
rect 240704 316742 240732 328442
rect 240692 316736 240744 316742
rect 240692 316678 240744 316684
rect 240876 247036 240928 247042
rect 240876 246978 240928 246984
rect 240888 237425 240916 246978
rect 240874 237416 240930 237425
rect 240874 237351 240930 237360
rect 240876 229084 240928 229090
rect 240876 229026 240928 229032
rect 240888 219473 240916 229026
rect 240874 219464 240930 219473
rect 240874 219399 240930 219408
rect 240508 67584 240560 67590
rect 240508 67526 240560 67532
rect 240508 57996 240560 58002
rect 240508 57938 240560 57944
rect 240520 8770 240548 57938
rect 240874 27568 240930 27577
rect 240874 27503 240930 27512
rect 240888 18018 240916 27503
rect 240876 18012 240928 18018
rect 240876 17954 240928 17960
rect 240508 8764 240560 8770
rect 240508 8706 240560 8712
rect 240416 8696 240468 8702
rect 240416 8638 240468 8644
rect 240324 8628 240376 8634
rect 240324 8570 240376 8576
rect 240784 4956 240836 4962
rect 240784 4898 240836 4904
rect 239864 3052 239916 3058
rect 239864 2994 239916 3000
rect 240796 480 240824 4898
rect 240980 2990 241008 335582
rect 241164 334762 241192 337486
rect 241152 334756 241204 334762
rect 241152 334698 241204 334704
rect 241060 333328 241112 333334
rect 241060 333270 241112 333276
rect 241072 302002 241100 333270
rect 241256 312066 241284 340068
rect 241348 333334 241376 340068
rect 241428 335844 241480 335850
rect 241428 335786 241480 335792
rect 241336 333328 241388 333334
rect 241336 333270 241388 333276
rect 241440 322318 241468 335786
rect 241532 335646 241560 340068
rect 241624 336802 241652 340068
rect 241716 338026 241744 340068
rect 241808 340054 241914 340082
rect 241704 338020 241756 338026
rect 241704 337962 241756 337968
rect 241612 336796 241664 336802
rect 241612 336738 241664 336744
rect 241520 335640 241572 335646
rect 241520 335582 241572 335588
rect 241428 322312 241480 322318
rect 241428 322254 241480 322260
rect 241164 312038 241284 312066
rect 241164 311166 241192 312038
rect 241152 311160 241204 311166
rect 241152 311102 241204 311108
rect 241072 301974 241192 302002
rect 241164 289814 241192 301974
rect 241060 289808 241112 289814
rect 241060 289750 241112 289756
rect 241152 289808 241204 289814
rect 241152 289750 241204 289756
rect 241072 285002 241100 289750
rect 241072 284974 241192 285002
rect 241164 273306 241192 284974
rect 241072 273278 241192 273306
rect 241072 273170 241100 273278
rect 241072 273142 241192 273170
rect 241164 270502 241192 273142
rect 241152 270496 241204 270502
rect 241152 270438 241204 270444
rect 241152 260908 241204 260914
rect 241152 260850 241204 260856
rect 241164 253994 241192 260850
rect 241072 253966 241192 253994
rect 241072 253858 241100 253966
rect 241072 253830 241192 253858
rect 241164 247042 241192 253830
rect 241152 247036 241204 247042
rect 241152 246978 241204 246984
rect 241058 237416 241114 237425
rect 241058 237351 241114 237360
rect 241072 230466 241100 237351
rect 241072 230438 241192 230466
rect 241164 229090 241192 230438
rect 241152 229084 241204 229090
rect 241152 229026 241204 229032
rect 241058 219464 241114 219473
rect 241058 219399 241114 219408
rect 241072 215370 241100 219399
rect 241072 215342 241192 215370
rect 241164 201482 241192 215342
rect 241152 201476 241204 201482
rect 241152 201418 241204 201424
rect 241336 201476 241388 201482
rect 241336 201418 241388 201424
rect 241348 191865 241376 201418
rect 241150 191856 241206 191865
rect 241150 191791 241206 191800
rect 241334 191856 241390 191865
rect 241334 191791 241390 191800
rect 241164 182170 241192 191791
rect 241152 182164 241204 182170
rect 241152 182106 241204 182112
rect 241336 182164 241388 182170
rect 241336 182106 241388 182112
rect 241348 172553 241376 182106
rect 241150 172544 241206 172553
rect 241150 172479 241206 172488
rect 241334 172544 241390 172553
rect 241334 172479 241390 172488
rect 241164 162858 241192 172479
rect 241152 162852 241204 162858
rect 241152 162794 241204 162800
rect 241152 153264 241204 153270
rect 241152 153206 241204 153212
rect 241164 125769 241192 153206
rect 241150 125760 241206 125769
rect 241150 125695 241206 125704
rect 241058 125624 241114 125633
rect 241058 125559 241114 125568
rect 241072 124166 241100 125559
rect 241060 124160 241112 124166
rect 241060 124102 241112 124108
rect 241152 114572 241204 114578
rect 241152 114514 241204 114520
rect 241164 64870 241192 114514
rect 241152 64864 241204 64870
rect 241152 64806 241204 64812
rect 241152 55276 241204 55282
rect 241152 55218 241204 55224
rect 241164 51134 241192 55218
rect 241152 51128 241204 51134
rect 241152 51070 241204 51076
rect 241244 50992 241296 50998
rect 241244 50934 241296 50940
rect 241256 45558 241284 50934
rect 241244 45552 241296 45558
rect 241244 45494 241296 45500
rect 241244 35964 241296 35970
rect 241244 35906 241296 35912
rect 241256 29050 241284 35906
rect 241256 29022 241376 29050
rect 241348 28914 241376 29022
rect 241072 28886 241376 28914
rect 241072 27577 241100 28886
rect 241058 27568 241114 27577
rect 241058 27503 241114 27512
rect 241060 18012 241112 18018
rect 241060 17954 241112 17960
rect 241072 3738 241100 17954
rect 241808 8498 241836 340054
rect 241888 335640 241940 335646
rect 241888 335582 241940 335588
rect 241900 8566 241928 335582
rect 241992 334694 242020 340068
rect 241980 334688 242032 334694
rect 241980 334630 242032 334636
rect 241980 8968 242032 8974
rect 241980 8910 242032 8916
rect 241888 8560 241940 8566
rect 241888 8502 241940 8508
rect 241796 8492 241848 8498
rect 241796 8434 241848 8440
rect 241060 3732 241112 3738
rect 241060 3674 241112 3680
rect 240968 2984 241020 2990
rect 240968 2926 241020 2932
rect 241992 480 242020 8910
rect 242084 2922 242112 340068
rect 242164 335640 242216 335646
rect 242164 335582 242216 335588
rect 242072 2916 242124 2922
rect 242072 2858 242124 2864
rect 242176 2854 242204 335582
rect 242268 8430 242296 340068
rect 242360 330614 242388 340068
rect 242452 335646 242480 340068
rect 242440 335640 242492 335646
rect 242440 335582 242492 335588
rect 242532 335640 242584 335646
rect 242532 335582 242584 335588
rect 242348 330608 242400 330614
rect 242348 330550 242400 330556
rect 242544 320958 242572 335582
rect 242532 320952 242584 320958
rect 242532 320894 242584 320900
rect 242256 8424 242308 8430
rect 242256 8366 242308 8372
rect 242636 8362 242664 340068
rect 242728 335646 242756 340068
rect 242820 337822 242848 340068
rect 242808 337816 242860 337822
rect 242808 337758 242860 337764
rect 243004 337550 243032 340068
rect 243096 338094 243124 340068
rect 243084 338088 243136 338094
rect 243084 338030 243136 338036
rect 242992 337544 243044 337550
rect 242992 337486 243044 337492
rect 242900 337476 242952 337482
rect 242900 337418 242952 337424
rect 242912 336530 242940 337418
rect 242900 336524 242952 336530
rect 242900 336466 242952 336472
rect 242716 335640 242768 335646
rect 242716 335582 242768 335588
rect 243188 333402 243216 340068
rect 243176 333396 243228 333402
rect 243176 333338 243228 333344
rect 243372 332042 243400 340068
rect 243360 332036 243412 332042
rect 243360 331978 243412 331984
rect 243464 331922 243492 340068
rect 243188 331894 243492 331922
rect 242624 8356 242676 8362
rect 242624 8298 242676 8304
rect 243188 6254 243216 331894
rect 243268 331356 243320 331362
rect 243268 331298 243320 331304
rect 243280 6322 243308 331298
rect 243556 318850 243584 340068
rect 243636 332036 243688 332042
rect 243636 331978 243688 331984
rect 243360 318844 243412 318850
rect 243360 318786 243412 318792
rect 243544 318844 243596 318850
rect 243544 318786 243596 318792
rect 243372 309194 243400 318786
rect 243360 309188 243412 309194
rect 243360 309130 243412 309136
rect 243544 309188 243596 309194
rect 243544 309130 243596 309136
rect 243556 292618 243584 309130
rect 243464 292590 243584 292618
rect 243464 289814 243492 292590
rect 243452 289808 243504 289814
rect 243452 289750 243504 289756
rect 243544 280220 243596 280226
rect 243544 280162 243596 280168
rect 243556 278730 243584 280162
rect 243544 278724 243596 278730
rect 243544 278666 243596 278672
rect 243544 256760 243596 256766
rect 243544 256702 243596 256708
rect 243556 255270 243584 256702
rect 243544 255264 243596 255270
rect 243544 255206 243596 255212
rect 243544 240236 243596 240242
rect 243544 240178 243596 240184
rect 243556 237386 243584 240178
rect 243544 237380 243596 237386
rect 243544 237322 243596 237328
rect 243452 219496 243504 219502
rect 243452 219438 243504 219444
rect 243464 219366 243492 219438
rect 243452 219360 243504 219366
rect 243452 219302 243504 219308
rect 243544 202904 243596 202910
rect 243544 202846 243596 202852
rect 243556 196602 243584 202846
rect 243372 196574 243584 196602
rect 243372 191826 243400 196574
rect 243360 191820 243412 191826
rect 243360 191762 243412 191768
rect 243452 186312 243504 186318
rect 243452 186254 243504 186260
rect 243464 182186 243492 186254
rect 243464 182158 243584 182186
rect 243556 182102 243584 182158
rect 243544 182096 243596 182102
rect 243544 182038 243596 182044
rect 243452 174412 243504 174418
rect 243452 174354 243504 174360
rect 243464 167074 243492 174354
rect 243452 167068 243504 167074
rect 243452 167010 243504 167016
rect 243544 166932 243596 166938
rect 243544 166874 243596 166880
rect 243556 157418 243584 166874
rect 243544 157412 243596 157418
rect 243544 157354 243596 157360
rect 243452 153332 243504 153338
rect 243452 153274 243504 153280
rect 243464 147762 243492 153274
rect 243452 147756 243504 147762
rect 243452 147698 243504 147704
rect 243452 147620 243504 147626
rect 243452 147562 243504 147568
rect 243464 143562 243492 147562
rect 243464 143534 243584 143562
rect 243556 142118 243584 143534
rect 243544 142112 243596 142118
rect 243544 142054 243596 142060
rect 243452 124228 243504 124234
rect 243452 124170 243504 124176
rect 243464 118930 243492 124170
rect 243452 118924 243504 118930
rect 243452 118866 243504 118872
rect 243544 108996 243596 109002
rect 243544 108938 243596 108944
rect 243556 101454 243584 108938
rect 243544 101448 243596 101454
rect 243544 101390 243596 101396
rect 243544 101312 243596 101318
rect 243544 101254 243596 101260
rect 243556 86970 243584 101254
rect 243544 86964 243596 86970
rect 243544 86906 243596 86912
rect 243544 77308 243596 77314
rect 243544 77250 243596 77256
rect 243556 60738 243584 77250
rect 243464 60710 243584 60738
rect 243464 51202 243492 60710
rect 243452 51196 243504 51202
rect 243452 51138 243504 51144
rect 243452 51060 243504 51066
rect 243452 51002 243504 51008
rect 243464 48362 243492 51002
rect 243464 48334 243584 48362
rect 243556 48278 243584 48334
rect 243544 48272 243596 48278
rect 243544 48214 243596 48220
rect 243544 27668 243596 27674
rect 243544 27610 243596 27616
rect 243556 27538 243584 27610
rect 243544 27532 243596 27538
rect 243544 27474 243596 27480
rect 243452 22092 243504 22098
rect 243452 22034 243504 22040
rect 243464 12510 243492 22034
rect 243452 12504 243504 12510
rect 243452 12446 243504 12452
rect 243360 12436 243412 12442
rect 243360 12378 243412 12384
rect 243372 7614 243400 12378
rect 243360 7608 243412 7614
rect 243360 7550 243412 7556
rect 243268 6316 243320 6322
rect 243268 6258 243320 6264
rect 243176 6248 243228 6254
rect 243176 6190 243228 6196
rect 243648 5098 243676 331978
rect 243740 5166 243768 340068
rect 243832 331362 243860 340068
rect 243820 331356 243872 331362
rect 243820 331298 243872 331304
rect 243924 321026 243952 340068
rect 244016 340054 244122 340082
rect 243912 321020 243964 321026
rect 243912 320962 243964 320968
rect 244016 5234 244044 340054
rect 244200 331974 244228 340068
rect 244306 340054 244412 340082
rect 244280 335844 244332 335850
rect 244280 335786 244332 335792
rect 244292 335458 244320 335786
rect 244384 335594 244412 340054
rect 244476 335714 244504 340068
rect 244568 335730 244596 340068
rect 244660 335918 244688 340068
rect 244752 340054 244858 340082
rect 244648 335912 244700 335918
rect 244648 335854 244700 335860
rect 244752 335850 244780 340054
rect 244740 335844 244792 335850
rect 244740 335786 244792 335792
rect 244464 335708 244516 335714
rect 244568 335702 244872 335730
rect 244464 335650 244516 335656
rect 244648 335640 244700 335646
rect 244384 335566 244596 335594
rect 244648 335582 244700 335588
rect 244292 335430 244504 335458
rect 244280 335368 244332 335374
rect 244280 335310 244332 335316
rect 244372 335368 244424 335374
rect 244372 335310 244424 335316
rect 244292 332110 244320 335310
rect 244280 332104 244332 332110
rect 244280 332046 244332 332052
rect 244188 331968 244240 331974
rect 244188 331910 244240 331916
rect 244384 327894 244412 335310
rect 244476 330750 244504 335430
rect 244464 330744 244516 330750
rect 244464 330686 244516 330692
rect 244372 327888 244424 327894
rect 244372 327830 244424 327836
rect 244568 318170 244596 335566
rect 244660 322386 244688 335582
rect 244740 331900 244792 331906
rect 244740 331842 244792 331848
rect 244752 329254 244780 331842
rect 244740 329248 244792 329254
rect 244740 329190 244792 329196
rect 244844 325106 244872 335702
rect 244936 335646 244964 340068
rect 245028 335646 245056 340068
rect 245120 337890 245148 340068
rect 245212 340054 245318 340082
rect 245108 337884 245160 337890
rect 245108 337826 245160 337832
rect 245108 335912 245160 335918
rect 245108 335854 245160 335860
rect 244924 335640 244976 335646
rect 244924 335582 244976 335588
rect 245016 335640 245068 335646
rect 245016 335582 245068 335588
rect 244832 325100 244884 325106
rect 244832 325042 244884 325048
rect 244648 322380 244700 322386
rect 244648 322322 244700 322328
rect 244556 318164 244608 318170
rect 244556 318106 244608 318112
rect 245120 316810 245148 335854
rect 245212 335374 245240 340054
rect 245292 336796 245344 336802
rect 245292 336738 245344 336744
rect 245200 335368 245252 335374
rect 245200 335310 245252 335316
rect 245304 333470 245332 336738
rect 245292 333464 245344 333470
rect 245292 333406 245344 333412
rect 245396 333282 245424 340068
rect 245212 333254 245424 333282
rect 245108 316804 245160 316810
rect 245108 316746 245160 316752
rect 244186 228168 244242 228177
rect 244186 228103 244242 228112
rect 244200 228018 244228 228103
rect 244370 228032 244426 228041
rect 244200 227990 244370 228018
rect 244370 227967 244426 227976
rect 244278 75984 244334 75993
rect 244462 75984 244518 75993
rect 244334 75942 244462 75970
rect 244278 75919 244334 75928
rect 244462 75919 244518 75928
rect 245212 15910 245240 333254
rect 245488 331906 245516 340068
rect 245568 337408 245620 337414
rect 245568 337350 245620 337356
rect 245580 335782 245608 337350
rect 245568 335776 245620 335782
rect 245568 335718 245620 335724
rect 245568 335640 245620 335646
rect 245568 335582 245620 335588
rect 245672 335594 245700 340068
rect 245764 335714 245792 340068
rect 245856 336802 245884 340068
rect 245844 336796 245896 336802
rect 245844 336738 245896 336744
rect 246040 335714 246068 340068
rect 245752 335708 245804 335714
rect 245752 335650 245804 335656
rect 246028 335708 246080 335714
rect 246028 335650 246080 335656
rect 245476 331900 245528 331906
rect 245476 331842 245528 331848
rect 245580 315382 245608 335582
rect 245672 335566 246068 335594
rect 245936 335504 245988 335510
rect 245936 335446 245988 335452
rect 245948 323746 245976 335446
rect 246040 329322 246068 335566
rect 246028 329316 246080 329322
rect 246028 329258 246080 329264
rect 245936 323740 245988 323746
rect 245936 323682 245988 323688
rect 245568 315376 245620 315382
rect 245568 315318 245620 315324
rect 246132 314022 246160 340068
rect 246224 335850 246252 340068
rect 246316 340054 246422 340082
rect 246212 335844 246264 335850
rect 246212 335786 246264 335792
rect 246316 335730 246344 340054
rect 246224 335702 246344 335730
rect 246224 335510 246252 335702
rect 246500 335594 246528 340068
rect 246592 337686 246620 340068
rect 246580 337680 246632 337686
rect 246580 337622 246632 337628
rect 246776 337142 246804 340068
rect 246764 337136 246816 337142
rect 246764 337078 246816 337084
rect 246672 335708 246724 335714
rect 246672 335650 246724 335656
rect 246316 335566 246528 335594
rect 246212 335504 246264 335510
rect 246212 335446 246264 335452
rect 246120 314016 246172 314022
rect 246120 313958 246172 313964
rect 246316 312662 246344 335566
rect 246396 335504 246448 335510
rect 246396 335446 246448 335452
rect 246408 319598 246436 335446
rect 246684 326534 246712 335650
rect 246868 330818 246896 340068
rect 246960 337754 246988 340068
rect 246948 337748 247000 337754
rect 246948 337690 247000 337696
rect 247040 336796 247092 336802
rect 247040 336738 247092 336744
rect 247052 332178 247080 336738
rect 247040 332172 247092 332178
rect 247040 332114 247092 332120
rect 246856 330812 246908 330818
rect 246856 330754 246908 330760
rect 247144 327962 247172 340068
rect 247236 334778 247264 340068
rect 247328 334898 247356 340068
rect 247408 335640 247460 335646
rect 247408 335582 247460 335588
rect 247316 334892 247368 334898
rect 247316 334834 247368 334840
rect 247236 334750 247356 334778
rect 247132 327956 247184 327962
rect 247132 327898 247184 327904
rect 246672 326528 246724 326534
rect 246672 326470 246724 326476
rect 246396 319592 246448 319598
rect 246396 319534 246448 319540
rect 246304 312656 246356 312662
rect 246304 312598 246356 312604
rect 245200 15904 245252 15910
rect 245200 15846 245252 15852
rect 247328 7682 247356 334750
rect 247420 7750 247448 335582
rect 247512 335458 247540 340068
rect 247604 335646 247632 340068
rect 247710 340054 247816 340082
rect 247684 337068 247736 337074
rect 247684 337010 247736 337016
rect 247592 335640 247644 335646
rect 247592 335582 247644 335588
rect 247512 335430 247632 335458
rect 247604 326602 247632 335430
rect 247592 326596 247644 326602
rect 247592 326538 247644 326544
rect 247408 7744 247460 7750
rect 247408 7686 247460 7692
rect 247316 7676 247368 7682
rect 247316 7618 247368 7624
rect 247696 5506 247724 337010
rect 247788 333538 247816 340054
rect 247776 333532 247828 333538
rect 247776 333474 247828 333480
rect 247880 6390 247908 340068
rect 247972 7818 248000 340068
rect 248064 336190 248092 340068
rect 248156 340054 248262 340082
rect 248052 336184 248104 336190
rect 248052 336126 248104 336132
rect 247960 7812 248012 7818
rect 247960 7754 248012 7760
rect 248156 6458 248184 340054
rect 248340 7886 248368 340068
rect 248432 336802 248460 340068
rect 248512 337000 248564 337006
rect 248512 336942 248564 336948
rect 248420 336796 248472 336802
rect 248420 336738 248472 336744
rect 248524 336326 248552 336942
rect 248512 336320 248564 336326
rect 248512 336262 248564 336268
rect 248512 335844 248564 335850
rect 248512 335786 248564 335792
rect 248420 335708 248472 335714
rect 248420 335650 248472 335656
rect 248432 333606 248460 335650
rect 248420 333600 248472 333606
rect 248420 333542 248472 333548
rect 248418 228032 248474 228041
rect 248418 227967 248474 227976
rect 248432 227633 248460 227967
rect 248418 227624 248474 227633
rect 248418 227559 248474 227568
rect 248328 7880 248380 7886
rect 248328 7822 248380 7828
rect 248144 6452 248196 6458
rect 248144 6394 248196 6400
rect 247868 6384 247920 6390
rect 247868 6326 247920 6332
rect 244372 5500 244424 5506
rect 244372 5442 244424 5448
rect 247684 5500 247736 5506
rect 247684 5442 247736 5448
rect 244004 5228 244056 5234
rect 244004 5170 244056 5176
rect 243728 5160 243780 5166
rect 243728 5102 243780 5108
rect 243636 5092 243688 5098
rect 243636 5034 243688 5040
rect 243176 3528 243228 3534
rect 243176 3470 243228 3476
rect 242164 2848 242216 2854
rect 242164 2790 242216 2796
rect 243188 480 243216 3470
rect 244384 480 244412 5442
rect 248524 5370 248552 335786
rect 248616 6526 248644 340068
rect 248708 336122 248736 340068
rect 248696 336116 248748 336122
rect 248696 336058 248748 336064
rect 248800 335714 248828 340068
rect 248892 340054 248998 340082
rect 248788 335708 248840 335714
rect 248788 335650 248840 335656
rect 248892 335594 248920 340054
rect 248972 335708 249024 335714
rect 248972 335650 249024 335656
rect 248708 335566 248920 335594
rect 248708 6594 248736 335566
rect 248984 335458 249012 335650
rect 248800 335430 249012 335458
rect 248800 6662 248828 335430
rect 248880 335368 248932 335374
rect 248880 335310 248932 335316
rect 248892 106185 248920 335310
rect 249076 333690 249104 340068
rect 249182 340054 249288 340082
rect 249260 335646 249288 340054
rect 249352 335714 249380 340068
rect 249340 335708 249392 335714
rect 249340 335650 249392 335656
rect 249248 335640 249300 335646
rect 249248 335582 249300 335588
rect 248984 333662 249104 333690
rect 248984 106214 249012 333662
rect 249444 329050 249472 340068
rect 249536 335850 249564 340068
rect 249616 336932 249668 336938
rect 249616 336874 249668 336880
rect 249524 335844 249576 335850
rect 249524 335786 249576 335792
rect 249628 335730 249656 336874
rect 249536 335702 249656 335730
rect 249536 335102 249564 335702
rect 249616 335640 249668 335646
rect 249616 335582 249668 335588
rect 249524 335096 249576 335102
rect 249524 335038 249576 335044
rect 249064 329044 249116 329050
rect 249064 328986 249116 328992
rect 249432 329044 249484 329050
rect 249432 328986 249484 328992
rect 249076 106282 249104 328986
rect 249156 328500 249208 328506
rect 249156 328442 249208 328448
rect 249168 318782 249196 328442
rect 249156 318776 249208 318782
rect 249156 318718 249208 318724
rect 249156 309188 249208 309194
rect 249156 309130 249208 309136
rect 249064 106276 249116 106282
rect 249064 106218 249116 106224
rect 249168 106214 249196 309130
rect 248972 106208 249024 106214
rect 248878 106176 248934 106185
rect 248972 106150 249024 106156
rect 249156 106208 249208 106214
rect 249156 106150 249208 106156
rect 248878 106111 248934 106120
rect 249064 106140 249116 106146
rect 249064 106082 249116 106088
rect 248970 105904 249026 105913
rect 248970 105839 249026 105848
rect 248984 101402 249012 105839
rect 248892 101374 249012 101402
rect 248892 86970 248920 101374
rect 248972 97844 249024 97850
rect 248972 97786 249024 97792
rect 248880 86964 248932 86970
rect 248880 86906 248932 86912
rect 248984 86902 249012 97786
rect 249076 86902 249104 106082
rect 249156 106072 249208 106078
rect 249156 106014 249208 106020
rect 249168 86970 249196 106014
rect 249156 86964 249208 86970
rect 249156 86906 249208 86912
rect 248972 86896 249024 86902
rect 248972 86838 249024 86844
rect 249064 86896 249116 86902
rect 249064 86838 249116 86844
rect 249064 86760 249116 86766
rect 249064 86702 249116 86708
rect 248880 82136 248932 82142
rect 248880 82078 248932 82084
rect 248892 6730 248920 82078
rect 248972 78464 249024 78470
rect 248972 78406 249024 78412
rect 248984 8022 249012 78406
rect 249076 8090 249104 86702
rect 249156 77308 249208 77314
rect 249156 77250 249208 77256
rect 249168 48226 249196 77250
rect 249168 48198 249288 48226
rect 249260 38690 249288 48198
rect 249156 38684 249208 38690
rect 249156 38626 249208 38632
rect 249248 38684 249300 38690
rect 249248 38626 249300 38632
rect 249064 8084 249116 8090
rect 249064 8026 249116 8032
rect 248972 8016 249024 8022
rect 248972 7958 249024 7964
rect 249168 7954 249196 38626
rect 249156 7948 249208 7954
rect 249156 7890 249208 7896
rect 248880 6724 248932 6730
rect 248880 6666 248932 6672
rect 248788 6656 248840 6662
rect 248788 6598 248840 6604
rect 248696 6588 248748 6594
rect 248696 6530 248748 6536
rect 248604 6520 248656 6526
rect 248604 6462 248656 6468
rect 248512 5364 248564 5370
rect 248512 5306 248564 5312
rect 249628 5302 249656 335582
rect 249720 335374 249748 340068
rect 249812 335510 249840 340068
rect 249918 340054 250024 340082
rect 249800 335504 249852 335510
rect 249800 335446 249852 335452
rect 249708 335368 249760 335374
rect 249708 335310 249760 335316
rect 249800 335368 249852 335374
rect 249800 335310 249852 335316
rect 249812 6866 249840 335310
rect 249892 335300 249944 335306
rect 249892 335242 249944 335248
rect 249800 6860 249852 6866
rect 249800 6802 249852 6808
rect 249616 5296 249668 5302
rect 249616 5238 249668 5244
rect 249904 4758 249932 335242
rect 249996 5438 250024 340054
rect 250088 335594 250116 340068
rect 250180 335714 250208 340068
rect 250286 340054 250392 340082
rect 250364 335782 250392 340054
rect 250352 335776 250404 335782
rect 250352 335718 250404 335724
rect 250168 335708 250220 335714
rect 250168 335650 250220 335656
rect 250088 335566 250392 335594
rect 250076 335504 250128 335510
rect 250076 335446 250128 335452
rect 250088 8158 250116 335446
rect 250076 8152 250128 8158
rect 250076 8094 250128 8100
rect 250364 6798 250392 335566
rect 250456 335374 250484 340068
rect 250444 335368 250496 335374
rect 250444 335310 250496 335316
rect 250548 8294 250576 340068
rect 250640 335306 250668 340068
rect 250720 335708 250772 335714
rect 250720 335650 250772 335656
rect 250628 335300 250680 335306
rect 250628 335242 250680 335248
rect 250536 8288 250588 8294
rect 250536 8230 250588 8236
rect 250732 8226 250760 335650
rect 250720 8220 250772 8226
rect 250720 8162 250772 8168
rect 250352 6792 250404 6798
rect 250352 6734 250404 6740
rect 250824 6118 250852 340068
rect 250916 7546 250944 340068
rect 250904 7540 250956 7546
rect 250904 7482 250956 7488
rect 250812 6112 250864 6118
rect 250812 6054 250864 6060
rect 249984 5432 250036 5438
rect 249984 5374 250036 5380
rect 249892 4752 249944 4758
rect 249892 4694 249944 4700
rect 251008 4690 251036 340068
rect 251088 335776 251140 335782
rect 251088 335718 251140 335724
rect 251100 5234 251128 335718
rect 251192 329390 251220 340068
rect 251284 337414 251312 340068
rect 251272 337408 251324 337414
rect 251272 337350 251324 337356
rect 251272 337204 251324 337210
rect 251272 337146 251324 337152
rect 251180 329384 251232 329390
rect 251180 329326 251232 329332
rect 251284 326398 251312 337146
rect 251376 337006 251404 340068
rect 251364 337000 251416 337006
rect 251364 336942 251416 336948
rect 251364 335912 251416 335918
rect 251364 335854 251416 335860
rect 251376 334966 251404 335854
rect 251456 335776 251508 335782
rect 251456 335718 251508 335724
rect 251364 334960 251416 334966
rect 251364 334902 251416 334908
rect 251272 326392 251324 326398
rect 251272 326334 251324 326340
rect 251468 323814 251496 335718
rect 251560 335714 251588 340068
rect 251652 335714 251680 340068
rect 251744 335918 251772 340068
rect 251836 340054 251942 340082
rect 251732 335912 251784 335918
rect 251732 335854 251784 335860
rect 251548 335708 251600 335714
rect 251548 335650 251600 335656
rect 251640 335708 251692 335714
rect 251640 335650 251692 335656
rect 251836 335594 251864 340054
rect 251916 336796 251968 336802
rect 251916 336738 251968 336744
rect 251560 335566 251864 335594
rect 251928 335594 251956 336738
rect 252020 335753 252048 340068
rect 252112 336394 252140 340068
rect 252204 340054 252310 340082
rect 252100 336388 252152 336394
rect 252100 336330 252152 336336
rect 252204 335782 252232 340054
rect 252284 336864 252336 336870
rect 252284 336806 252336 336812
rect 252192 335776 252244 335782
rect 252006 335744 252062 335753
rect 252192 335718 252244 335724
rect 252296 335714 252324 336806
rect 252006 335679 252062 335688
rect 252100 335708 252152 335714
rect 252100 335650 252152 335656
rect 252284 335708 252336 335714
rect 252284 335650 252336 335656
rect 251928 335566 252048 335594
rect 251560 325174 251588 335566
rect 251916 335504 251968 335510
rect 251638 335472 251694 335481
rect 251916 335446 251968 335452
rect 251638 335407 251694 335416
rect 251548 325168 251600 325174
rect 251548 325110 251600 325116
rect 251456 323808 251508 323814
rect 251456 323750 251508 323756
rect 251652 319666 251680 335407
rect 251732 335368 251784 335374
rect 251732 335310 251784 335316
rect 251744 332314 251772 335310
rect 251732 332308 251784 332314
rect 251732 332250 251784 332256
rect 251732 326392 251784 326398
rect 251732 326334 251784 326340
rect 251640 319660 251692 319666
rect 251640 319602 251692 319608
rect 251744 313970 251772 326334
rect 251744 313942 251864 313970
rect 251836 307766 251864 313942
rect 251824 307760 251876 307766
rect 251824 307702 251876 307708
rect 251732 298172 251784 298178
rect 251732 298114 251784 298120
rect 251744 292534 251772 298114
rect 251732 292528 251784 292534
rect 251732 292470 251784 292476
rect 251640 287088 251692 287094
rect 251640 287030 251692 287036
rect 251652 260846 251680 287030
rect 251364 260840 251416 260846
rect 251364 260782 251416 260788
rect 251640 260840 251692 260846
rect 251640 260782 251692 260788
rect 251376 258097 251404 260782
rect 251362 258088 251418 258097
rect 251362 258023 251418 258032
rect 251362 257952 251418 257961
rect 251362 257887 251418 257896
rect 251376 253230 251404 257887
rect 251364 253224 251416 253230
rect 251364 253166 251416 253172
rect 251548 253224 251600 253230
rect 251548 253166 251600 253172
rect 251560 245002 251588 253166
rect 251548 244996 251600 245002
rect 251548 244938 251600 244944
rect 251732 244996 251784 245002
rect 251732 244938 251784 244944
rect 251744 237538 251772 244938
rect 251744 237510 251864 237538
rect 251836 225010 251864 237510
rect 251824 225004 251876 225010
rect 251824 224946 251876 224952
rect 251824 222216 251876 222222
rect 251824 222158 251876 222164
rect 251836 217410 251864 222158
rect 251560 217382 251864 217410
rect 251560 205698 251588 217382
rect 251548 205692 251600 205698
rect 251548 205634 251600 205640
rect 251548 205556 251600 205562
rect 251548 205498 251600 205504
rect 251560 202881 251588 205498
rect 251546 202872 251602 202881
rect 251546 202807 251602 202816
rect 251730 202872 251786 202881
rect 251730 202807 251786 202816
rect 251744 197946 251772 202807
rect 251640 197940 251692 197946
rect 251640 197882 251692 197888
rect 251732 197940 251784 197946
rect 251732 197882 251784 197888
rect 251652 171086 251680 197882
rect 251640 171080 251692 171086
rect 251640 171022 251692 171028
rect 251824 171080 251876 171086
rect 251824 171022 251876 171028
rect 251836 151842 251864 171022
rect 251732 151836 251784 151842
rect 251732 151778 251784 151784
rect 251824 151836 251876 151842
rect 251824 151778 251876 151784
rect 251744 137154 251772 151778
rect 251732 137148 251784 137154
rect 251732 137090 251784 137096
rect 251640 132524 251692 132530
rect 251640 132466 251692 132472
rect 251652 124302 251680 132466
rect 251640 124296 251692 124302
rect 251640 124238 251692 124244
rect 251732 124092 251784 124098
rect 251732 124034 251784 124040
rect 251744 110514 251772 124034
rect 251744 110486 251864 110514
rect 251836 110430 251864 110486
rect 251824 110424 251876 110430
rect 251824 110366 251876 110372
rect 251744 100774 251772 100805
rect 251732 100768 251784 100774
rect 251784 100716 251864 100722
rect 251732 100710 251864 100716
rect 251744 100694 251864 100710
rect 251836 95962 251864 100694
rect 251744 95934 251864 95962
rect 251744 84182 251772 95934
rect 251732 84176 251784 84182
rect 251732 84118 251784 84124
rect 251824 74588 251876 74594
rect 251824 74530 251876 74536
rect 251836 66298 251864 74530
rect 251640 66292 251692 66298
rect 251640 66234 251692 66240
rect 251824 66292 251876 66298
rect 251824 66234 251876 66240
rect 251652 48346 251680 66234
rect 251548 48340 251600 48346
rect 251548 48282 251600 48288
rect 251640 48340 251692 48346
rect 251640 48282 251692 48288
rect 251560 45014 251588 48282
rect 251548 45008 251600 45014
rect 251548 44950 251600 44956
rect 251732 45008 251784 45014
rect 251732 44950 251784 44956
rect 251744 18018 251772 44950
rect 251640 18012 251692 18018
rect 251640 17954 251692 17960
rect 251732 18012 251784 18018
rect 251732 17954 251784 17960
rect 251652 8974 251680 17954
rect 251928 10334 251956 335446
rect 252020 11762 252048 335566
rect 252112 326398 252140 335650
rect 252388 335594 252416 340068
rect 252480 336002 252508 340068
rect 252664 336462 252692 340068
rect 252652 336456 252704 336462
rect 252652 336398 252704 336404
rect 252480 335974 252600 336002
rect 252204 335566 252416 335594
rect 252100 326392 252152 326398
rect 252100 326334 252152 326340
rect 252204 122126 252232 335566
rect 252572 335458 252600 335974
rect 252388 335430 252600 335458
rect 252388 333674 252416 335430
rect 252376 333668 252428 333674
rect 252376 333610 252428 333616
rect 252756 328030 252784 340068
rect 252848 336938 252876 340068
rect 252836 336932 252888 336938
rect 252836 336874 252888 336880
rect 252928 335640 252980 335646
rect 252928 335582 252980 335588
rect 252744 328024 252796 328030
rect 252744 327966 252796 327972
rect 252284 326392 252336 326398
rect 252284 326334 252336 326340
rect 252296 321094 252324 326334
rect 252284 321088 252336 321094
rect 252284 321030 252336 321036
rect 252192 122120 252244 122126
rect 252192 122062 252244 122068
rect 252008 11756 252060 11762
rect 252008 11698 252060 11704
rect 252940 10402 252968 335582
rect 253032 332246 253060 340068
rect 253020 332240 253072 332246
rect 253020 332182 253072 332188
rect 253124 326670 253152 340068
rect 253230 340054 253336 340082
rect 253204 337952 253256 337958
rect 253204 337894 253256 337900
rect 253112 326664 253164 326670
rect 253112 326606 253164 326612
rect 253216 10470 253244 337894
rect 253308 337482 253336 340054
rect 253296 337476 253348 337482
rect 253296 337418 253348 337424
rect 253400 335170 253428 340068
rect 253492 336802 253520 340068
rect 253584 337006 253612 340068
rect 253572 337000 253624 337006
rect 253572 336942 253624 336948
rect 253768 336870 253796 340068
rect 253756 336864 253808 336870
rect 253756 336806 253808 336812
rect 253480 336796 253532 336802
rect 253480 336738 253532 336744
rect 253860 335646 253888 340068
rect 253966 340054 254072 340082
rect 254044 335714 254072 340054
rect 254032 335708 254084 335714
rect 254032 335650 254084 335656
rect 253848 335640 253900 335646
rect 253848 335582 253900 335588
rect 254136 335578 254164 340068
rect 254228 337958 254256 340068
rect 254216 337952 254268 337958
rect 254216 337894 254268 337900
rect 254320 335628 254348 340068
rect 254400 335708 254452 335714
rect 254400 335650 254452 335656
rect 254228 335600 254348 335628
rect 254124 335572 254176 335578
rect 254124 335514 254176 335520
rect 254122 335472 254178 335481
rect 254122 335407 254178 335416
rect 253388 335164 253440 335170
rect 253388 335106 253440 335112
rect 254136 318850 254164 335407
rect 254032 318844 254084 318850
rect 254032 318786 254084 318792
rect 254124 318844 254176 318850
rect 254124 318786 254176 318792
rect 254044 298314 254072 318786
rect 254032 298308 254084 298314
rect 254032 298250 254084 298256
rect 254032 298172 254084 298178
rect 254032 298114 254084 298120
rect 254044 296721 254072 298114
rect 253846 296712 253902 296721
rect 253846 296647 253902 296656
rect 254030 296712 254086 296721
rect 254030 296647 254086 296656
rect 253860 287094 253888 296647
rect 253848 287088 253900 287094
rect 253848 287030 253900 287036
rect 254032 287088 254084 287094
rect 254032 287030 254084 287036
rect 254044 260914 254072 287030
rect 254032 260908 254084 260914
rect 254032 260850 254084 260856
rect 253940 258120 253992 258126
rect 253940 258062 253992 258068
rect 253952 238762 253980 258062
rect 253952 238746 254072 238762
rect 253952 238740 254084 238746
rect 253952 238734 254032 238740
rect 254032 238682 254084 238688
rect 254032 230308 254084 230314
rect 254032 230250 254084 230256
rect 254044 225706 254072 230250
rect 253952 225678 254072 225706
rect 253952 201521 253980 225678
rect 253938 201512 253994 201521
rect 253938 201447 253994 201456
rect 254122 201512 254178 201521
rect 254122 201447 254178 201456
rect 254136 197962 254164 201447
rect 254044 197934 254164 197962
rect 254044 186402 254072 197934
rect 254044 186374 254164 186402
rect 254136 186266 254164 186374
rect 253952 186238 254164 186266
rect 253952 173942 253980 186238
rect 253940 173936 253992 173942
rect 253940 173878 253992 173884
rect 254124 173868 254176 173874
rect 254124 173810 254176 173816
rect 254136 151842 254164 173810
rect 253940 151836 253992 151842
rect 253940 151778 253992 151784
rect 254124 151836 254176 151842
rect 254124 151778 254176 151784
rect 253952 144945 253980 151778
rect 253938 144936 253994 144945
rect 253938 144871 253994 144880
rect 254122 144936 254178 144945
rect 254122 144871 254178 144880
rect 254136 142118 254164 144871
rect 254124 142112 254176 142118
rect 254124 142054 254176 142060
rect 254032 132524 254084 132530
rect 254032 132466 254084 132472
rect 254044 124234 254072 132466
rect 253940 124228 253992 124234
rect 253940 124170 253992 124176
rect 254032 124228 254084 124234
rect 254032 124170 254084 124176
rect 253952 122806 253980 124170
rect 253940 122800 253992 122806
rect 253940 122742 253992 122748
rect 254124 111852 254176 111858
rect 254124 111794 254176 111800
rect 254136 103630 254164 111794
rect 253940 103624 253992 103630
rect 253940 103566 253992 103572
rect 254124 103624 254176 103630
rect 254124 103566 254176 103572
rect 253952 100722 253980 103566
rect 253860 100694 253980 100722
rect 253860 95266 253888 100694
rect 253848 95260 253900 95266
rect 253848 95202 253900 95208
rect 253848 91112 253900 91118
rect 253848 91054 253900 91060
rect 253860 85610 253888 91054
rect 253848 85604 253900 85610
rect 253848 85546 253900 85552
rect 253940 85604 253992 85610
rect 253940 85546 253992 85552
rect 253952 80170 253980 85546
rect 253940 80164 253992 80170
rect 253940 80106 253992 80112
rect 253940 75880 253992 75886
rect 253940 75822 253992 75828
rect 253952 43518 253980 75822
rect 253940 43512 253992 43518
rect 253940 43454 253992 43460
rect 254124 43512 254176 43518
rect 254124 43454 254176 43460
rect 254136 29102 254164 43454
rect 254124 29096 254176 29102
rect 254124 29038 254176 29044
rect 253940 28960 253992 28966
rect 253940 28902 253992 28908
rect 253952 18086 253980 28902
rect 253940 18080 253992 18086
rect 253940 18022 253992 18028
rect 253940 16652 253992 16658
rect 253940 16594 253992 16600
rect 253204 10464 253256 10470
rect 253204 10406 253256 10412
rect 252928 10396 252980 10402
rect 252928 10338 252980 10344
rect 251916 10328 251968 10334
rect 251916 10270 251968 10276
rect 251640 8968 251692 8974
rect 251640 8910 251692 8916
rect 251088 5228 251140 5234
rect 251088 5170 251140 5176
rect 250996 4684 251048 4690
rect 250996 4626 251048 4632
rect 246764 3868 246816 3874
rect 246764 3810 246816 3816
rect 245568 3664 245620 3670
rect 245568 3606 245620 3612
rect 245580 480 245608 3606
rect 246776 480 246804 3810
rect 247960 3732 248012 3738
rect 247960 3674 248012 3680
rect 247972 480 248000 3674
rect 252652 3596 252704 3602
rect 252652 3538 252704 3544
rect 249156 3392 249208 3398
rect 249156 3334 249208 3340
rect 249168 480 249196 3334
rect 251456 3324 251508 3330
rect 251456 3266 251508 3272
rect 250352 2916 250404 2922
rect 250352 2858 250404 2864
rect 250364 480 250392 2858
rect 251468 480 251496 3266
rect 252664 480 252692 3538
rect 253952 3534 253980 16594
rect 254228 4894 254256 335600
rect 254308 335368 254360 335374
rect 254308 335310 254360 335316
rect 254320 4962 254348 335310
rect 254308 4956 254360 4962
rect 254308 4898 254360 4904
rect 254216 4888 254268 4894
rect 254216 4830 254268 4836
rect 254412 4826 254440 335650
rect 254504 335322 254532 340068
rect 254596 335481 254624 340068
rect 254582 335472 254638 335481
rect 254582 335407 254638 335416
rect 254688 335374 254716 340068
rect 254872 337210 254900 340068
rect 254860 337204 254912 337210
rect 254860 337146 254912 337152
rect 254860 336864 254912 336870
rect 254860 336806 254912 336812
rect 254768 336796 254820 336802
rect 254768 336738 254820 336744
rect 254676 335368 254728 335374
rect 254504 335294 254624 335322
rect 254676 335310 254728 335316
rect 254492 335232 254544 335238
rect 254492 335174 254544 335180
rect 254504 6186 254532 335174
rect 254492 6180 254544 6186
rect 254492 6122 254544 6128
rect 254596 6050 254624 335294
rect 254780 335186 254808 336738
rect 254688 335158 254808 335186
rect 254584 6044 254636 6050
rect 254584 5986 254636 5992
rect 254400 4820 254452 4826
rect 254400 4762 254452 4768
rect 254688 3738 254716 335158
rect 254872 335050 254900 336806
rect 254780 335022 254900 335050
rect 254676 3732 254728 3738
rect 254676 3674 254728 3680
rect 253940 3528 253992 3534
rect 253940 3470 253992 3476
rect 253848 3460 253900 3466
rect 253848 3402 253900 3408
rect 253860 480 253888 3402
rect 254780 3330 254808 335022
rect 254964 3942 254992 340068
rect 255056 337074 255084 340068
rect 255148 340054 255254 340082
rect 255044 337068 255096 337074
rect 255044 337010 255096 337016
rect 255044 4072 255096 4078
rect 255044 4014 255096 4020
rect 254952 3936 255004 3942
rect 254952 3878 255004 3884
rect 254768 3324 254820 3330
rect 254768 3266 254820 3272
rect 255056 480 255084 4014
rect 255148 3670 255176 340054
rect 255332 3874 255360 340068
rect 255424 336802 255452 340068
rect 255412 336796 255464 336802
rect 255412 336738 255464 336744
rect 255504 335640 255556 335646
rect 255504 335582 255556 335588
rect 255516 4146 255544 335582
rect 255504 4140 255556 4146
rect 255504 4082 255556 4088
rect 255320 3868 255372 3874
rect 255320 3810 255372 3816
rect 255136 3664 255188 3670
rect 255136 3606 255188 3612
rect 255608 3398 255636 340068
rect 255700 335374 255728 340068
rect 255792 336870 255820 340068
rect 255884 340054 255990 340082
rect 255780 336864 255832 336870
rect 255780 336806 255832 336812
rect 255884 335628 255912 340054
rect 255792 335600 255912 335628
rect 255688 335368 255740 335374
rect 255688 335310 255740 335316
rect 255688 335232 255740 335238
rect 255688 335174 255740 335180
rect 255700 3466 255728 335174
rect 255792 3602 255820 335600
rect 256068 335578 256096 340068
rect 256056 335572 256108 335578
rect 256056 335514 256108 335520
rect 256160 335458 256188 340068
rect 256252 340054 256358 340082
rect 256252 335646 256280 340054
rect 256240 335640 256292 335646
rect 256240 335582 256292 335588
rect 255884 335430 256188 335458
rect 255884 4078 255912 335430
rect 256056 335368 256108 335374
rect 256056 335310 256108 335316
rect 255872 4072 255924 4078
rect 255872 4014 255924 4020
rect 255780 3596 255832 3602
rect 255780 3538 255832 3544
rect 255688 3460 255740 3466
rect 255688 3402 255740 3408
rect 255596 3392 255648 3398
rect 255596 3334 255648 3340
rect 256068 2922 256096 335310
rect 256436 335306 256464 340068
rect 256528 336802 256556 340068
rect 256712 337142 256740 340068
rect 256700 337136 256752 337142
rect 256700 337078 256752 337084
rect 256516 336796 256568 336802
rect 256516 336738 256568 336744
rect 256804 335510 256832 340068
rect 256896 337074 256924 340068
rect 256884 337068 256936 337074
rect 256884 337010 256936 337016
rect 257080 337006 257108 340068
rect 257172 337890 257200 340068
rect 257160 337884 257212 337890
rect 257160 337826 257212 337832
rect 257264 337686 257292 340068
rect 257252 337680 257304 337686
rect 257252 337622 257304 337628
rect 257448 337278 257476 340068
rect 257540 337754 257568 340068
rect 257528 337748 257580 337754
rect 257528 337690 257580 337696
rect 257436 337272 257488 337278
rect 257436 337214 257488 337220
rect 257068 337000 257120 337006
rect 257068 336942 257120 336948
rect 257160 336932 257212 336938
rect 257160 336874 257212 336880
rect 257068 336864 257120 336870
rect 257068 336806 257120 336812
rect 256792 335504 256844 335510
rect 256792 335446 256844 335452
rect 256424 335300 256476 335306
rect 256424 335242 256476 335248
rect 256608 331764 256660 331770
rect 256608 331706 256660 331712
rect 256620 325689 256648 331706
rect 256422 325680 256478 325689
rect 256422 325615 256478 325624
rect 256606 325680 256662 325689
rect 256606 325615 256662 325624
rect 256436 316062 256464 325615
rect 256424 316056 256476 316062
rect 256422 316024 256424 316033
rect 256608 316056 256660 316062
rect 256476 316024 256478 316033
rect 256422 315959 256478 315968
rect 256606 316024 256608 316033
rect 256660 316024 256662 316033
rect 256606 315959 256662 315968
rect 256436 306406 256464 315959
rect 256424 306400 256476 306406
rect 256424 306342 256476 306348
rect 256700 306400 256752 306406
rect 256700 306342 256752 306348
rect 256712 302122 256740 306342
rect 256516 302116 256568 302122
rect 256516 302058 256568 302064
rect 256700 302116 256752 302122
rect 256700 302058 256752 302064
rect 256528 289882 256556 302058
rect 256516 289876 256568 289882
rect 256516 289818 256568 289824
rect 256608 289740 256660 289746
rect 256608 289682 256660 289688
rect 256620 244338 256648 289682
rect 256528 244310 256648 244338
rect 256528 244202 256556 244310
rect 256528 244174 256648 244202
rect 256620 222222 256648 244174
rect 256516 222216 256568 222222
rect 256516 222158 256568 222164
rect 256608 222216 256660 222222
rect 256608 222158 256660 222164
rect 256528 217274 256556 222158
rect 256528 217246 256648 217274
rect 256620 186402 256648 217246
rect 256528 186374 256648 186402
rect 256528 186266 256556 186374
rect 256528 186238 256648 186266
rect 256620 174010 256648 186238
rect 256608 174004 256660 174010
rect 256608 173946 256660 173952
rect 256516 169788 256568 169794
rect 256516 169730 256568 169736
rect 256528 166410 256556 169730
rect 256528 166382 256648 166410
rect 256620 151842 256648 166382
rect 256608 151836 256660 151842
rect 256608 151778 256660 151784
rect 256884 151836 256936 151842
rect 256884 151778 256936 151784
rect 256896 150498 256924 151778
rect 256804 150470 256924 150498
rect 256804 149054 256832 150470
rect 256792 149048 256844 149054
rect 256792 148990 256844 148996
rect 256424 139460 256476 139466
rect 256424 139402 256476 139408
rect 256436 132433 256464 139402
rect 256422 132424 256478 132433
rect 256422 132359 256478 132368
rect 256606 132424 256662 132433
rect 256606 132359 256662 132368
rect 256620 127514 256648 132359
rect 256528 127486 256648 127514
rect 256528 122806 256556 127486
rect 256516 122800 256568 122806
rect 256516 122742 256568 122748
rect 256608 113212 256660 113218
rect 256608 113154 256660 113160
rect 256620 104802 256648 113154
rect 256620 104774 256740 104802
rect 256712 85610 256740 104774
rect 256516 85604 256568 85610
rect 256516 85546 256568 85552
rect 256700 85604 256752 85610
rect 256700 85546 256752 85552
rect 256528 80102 256556 85546
rect 256516 80096 256568 80102
rect 256516 80038 256568 80044
rect 256608 79960 256660 79966
rect 256608 79902 256660 79908
rect 256620 66298 256648 79902
rect 256516 66292 256568 66298
rect 256516 66234 256568 66240
rect 256608 66292 256660 66298
rect 256608 66234 256660 66240
rect 256528 56642 256556 66234
rect 256516 56636 256568 56642
rect 256516 56578 256568 56584
rect 256608 56636 256660 56642
rect 256608 56578 256660 56584
rect 256620 37262 256648 56578
rect 256608 37256 256660 37262
rect 256608 37198 256660 37204
rect 256700 37256 256752 37262
rect 256700 37198 256752 37204
rect 256712 35902 256740 37198
rect 256700 35896 256752 35902
rect 256700 35838 256752 35844
rect 256608 26308 256660 26314
rect 256608 26250 256660 26256
rect 256620 26194 256648 26250
rect 256528 26166 256648 26194
rect 256528 16726 256556 26166
rect 256516 16720 256568 16726
rect 256516 16662 256568 16668
rect 256608 16652 256660 16658
rect 256608 16594 256660 16600
rect 256620 9738 256648 16594
rect 256620 9710 256740 9738
rect 256712 9466 256740 9710
rect 256528 9438 256740 9466
rect 256528 8294 256556 9438
rect 256516 8288 256568 8294
rect 256516 8230 256568 8236
rect 257080 4758 257108 336806
rect 257172 316742 257200 336874
rect 257632 336870 257660 340068
rect 257724 340054 257830 340082
rect 257620 336864 257672 336870
rect 257620 336806 257672 336812
rect 257344 336796 257396 336802
rect 257344 336738 257396 336744
rect 257528 336796 257580 336802
rect 257528 336738 257580 336744
rect 257160 316736 257212 316742
rect 257160 316678 257212 316684
rect 257068 4752 257120 4758
rect 257068 4694 257120 4700
rect 256240 4140 256292 4146
rect 256240 4082 256292 4088
rect 256056 2916 256108 2922
rect 256056 2858 256108 2864
rect 256252 480 256280 4082
rect 257356 4078 257384 336738
rect 257436 8288 257488 8294
rect 257436 8230 257488 8236
rect 257344 4072 257396 4078
rect 257344 4014 257396 4020
rect 257448 480 257476 8230
rect 257540 5370 257568 336738
rect 257724 5506 257752 340054
rect 257804 337000 257856 337006
rect 257804 336942 257856 336948
rect 257816 335628 257844 336942
rect 257908 336938 257936 340068
rect 257896 336932 257948 336938
rect 257896 336874 257948 336880
rect 258000 336802 258028 340068
rect 258080 337068 258132 337074
rect 258080 337010 258132 337016
rect 257988 336796 258040 336802
rect 257988 336738 258040 336744
rect 258092 336682 258120 337010
rect 258000 336654 258120 336682
rect 257816 335600 257936 335628
rect 257804 335504 257856 335510
rect 257804 335446 257856 335452
rect 257712 5500 257764 5506
rect 257712 5442 257764 5448
rect 257528 5364 257580 5370
rect 257528 5306 257580 5312
rect 257816 4010 257844 335446
rect 257804 4004 257856 4010
rect 257804 3946 257856 3952
rect 257908 3874 257936 335600
rect 258000 3942 258028 336654
rect 258184 5438 258212 340068
rect 258276 337618 258304 340068
rect 258264 337612 258316 337618
rect 258264 337554 258316 337560
rect 258368 337006 258396 340068
rect 258448 337136 258500 337142
rect 258448 337078 258500 337084
rect 258356 337000 258408 337006
rect 258356 336942 258408 336948
rect 258264 336932 258316 336938
rect 258264 336874 258316 336880
rect 258172 5432 258224 5438
rect 258172 5374 258224 5380
rect 258276 4962 258304 336874
rect 258356 336864 258408 336870
rect 258356 336806 258408 336812
rect 258368 5030 258396 336806
rect 258356 5024 258408 5030
rect 258356 4966 258408 4972
rect 258264 4956 258316 4962
rect 258264 4898 258316 4904
rect 258460 4146 258488 337078
rect 258552 336802 258580 340068
rect 258644 337142 258672 340068
rect 258632 337136 258684 337142
rect 258632 337078 258684 337084
rect 258540 336796 258592 336802
rect 258540 336738 258592 336744
rect 258736 333146 258764 340068
rect 258552 333118 258764 333146
rect 258828 340054 258934 340082
rect 258552 328438 258580 333118
rect 258540 328432 258592 328438
rect 258540 328374 258592 328380
rect 258632 328432 258684 328438
rect 258632 328374 258684 328380
rect 258644 253994 258672 328374
rect 258552 253966 258672 253994
rect 258552 253858 258580 253966
rect 258552 253830 258672 253858
rect 258644 244458 258672 253830
rect 258632 244452 258684 244458
rect 258632 244394 258684 244400
rect 258540 240168 258592 240174
rect 258540 240110 258592 240116
rect 258552 230518 258580 240110
rect 258540 230512 258592 230518
rect 258540 230454 258592 230460
rect 258632 230512 258684 230518
rect 258632 230454 258684 230460
rect 258644 225706 258672 230454
rect 258552 225678 258672 225706
rect 258552 218090 258580 225678
rect 258552 218062 258764 218090
rect 258736 202910 258764 218062
rect 258632 202904 258684 202910
rect 258632 202846 258684 202852
rect 258724 202904 258776 202910
rect 258724 202846 258776 202852
rect 258644 180810 258672 202846
rect 258632 180804 258684 180810
rect 258632 180746 258684 180752
rect 258632 171216 258684 171222
rect 258632 171158 258684 171164
rect 258644 171086 258672 171158
rect 258632 171080 258684 171086
rect 258632 171022 258684 171028
rect 258632 161492 258684 161498
rect 258632 161434 258684 161440
rect 258644 151774 258672 161434
rect 258632 151768 258684 151774
rect 258632 151710 258684 151716
rect 258632 142180 258684 142186
rect 258632 142122 258684 142128
rect 258644 132546 258672 142122
rect 258552 132518 258672 132546
rect 258552 131102 258580 132518
rect 258540 131096 258592 131102
rect 258540 131038 258592 131044
rect 258632 121508 258684 121514
rect 258632 121450 258684 121456
rect 258644 111790 258672 121450
rect 258632 111784 258684 111790
rect 258632 111726 258684 111732
rect 258632 102196 258684 102202
rect 258632 102138 258684 102144
rect 258644 97306 258672 102138
rect 258632 97300 258684 97306
rect 258632 97242 258684 97248
rect 258540 84244 258592 84250
rect 258540 84186 258592 84192
rect 258552 84153 258580 84186
rect 258538 84144 258594 84153
rect 258538 84079 258594 84088
rect 258722 84008 258778 84017
rect 258722 83943 258778 83952
rect 258736 80050 258764 83943
rect 258644 80022 258764 80050
rect 258644 74526 258672 80022
rect 258632 74520 258684 74526
rect 258632 74462 258684 74468
rect 258540 65000 258592 65006
rect 258540 64942 258592 64948
rect 258552 64870 258580 64942
rect 258540 64864 258592 64870
rect 258540 64806 258592 64812
rect 258632 64864 258684 64870
rect 258632 64806 258684 64812
rect 258644 63510 258672 64806
rect 258632 63504 258684 63510
rect 258632 63446 258684 63452
rect 258632 45620 258684 45626
rect 258632 45562 258684 45568
rect 258644 30410 258672 45562
rect 258552 30382 258672 30410
rect 258552 18018 258580 30382
rect 258540 18012 258592 18018
rect 258540 17954 258592 17960
rect 258632 18012 258684 18018
rect 258632 17954 258684 17960
rect 258644 9738 258672 17954
rect 258644 9710 258764 9738
rect 258736 9602 258764 9710
rect 258552 9574 258764 9602
rect 258552 5166 258580 9574
rect 258540 5160 258592 5166
rect 258540 5102 258592 5108
rect 258828 5098 258856 340054
rect 258908 336796 258960 336802
rect 258908 336738 258960 336744
rect 258920 5234 258948 336738
rect 259012 318102 259040 340068
rect 259104 336870 259132 340068
rect 259184 337000 259236 337006
rect 259184 336942 259236 336948
rect 259092 336864 259144 336870
rect 259092 336806 259144 336812
rect 259196 323474 259224 336942
rect 259288 336938 259316 340068
rect 259276 336932 259328 336938
rect 259276 336874 259328 336880
rect 259380 323610 259408 340068
rect 259472 334082 259500 340068
rect 259656 337482 259684 340068
rect 259644 337476 259696 337482
rect 259644 337418 259696 337424
rect 259460 334076 259512 334082
rect 259460 334018 259512 334024
rect 259748 330478 259776 340068
rect 259854 340054 259960 340082
rect 259828 336932 259880 336938
rect 259828 336874 259880 336880
rect 259736 330472 259788 330478
rect 259736 330414 259788 330420
rect 259368 323604 259420 323610
rect 259368 323546 259420 323552
rect 259184 323468 259236 323474
rect 259184 323410 259236 323416
rect 259368 323468 259420 323474
rect 259368 323410 259420 323416
rect 259000 318096 259052 318102
rect 259000 318038 259052 318044
rect 259380 253994 259408 323410
rect 259288 253966 259408 253994
rect 259288 253858 259316 253966
rect 259288 253830 259408 253858
rect 259380 244322 259408 253830
rect 259368 244316 259420 244322
rect 259368 244258 259420 244264
rect 259276 244248 259328 244254
rect 259276 244190 259328 244196
rect 259288 240106 259316 244190
rect 259184 240100 259236 240106
rect 259184 240042 259236 240048
rect 259276 240100 259328 240106
rect 259276 240042 259328 240048
rect 259196 231826 259224 240042
rect 259196 231798 259500 231826
rect 259472 228154 259500 231798
rect 259472 228126 259592 228154
rect 259458 228032 259514 228041
rect 259458 227967 259460 227976
rect 259512 227967 259514 227976
rect 259460 227938 259512 227944
rect 259564 220862 259592 228126
rect 259552 220856 259604 220862
rect 259552 220798 259604 220804
rect 259644 220856 259696 220862
rect 259644 220798 259696 220804
rect 259734 220824 259790 220833
rect 259656 212566 259684 220798
rect 259734 220759 259790 220768
rect 259368 212560 259420 212566
rect 259368 212502 259420 212508
rect 259644 212560 259696 212566
rect 259644 212502 259696 212508
rect 259380 180810 259408 212502
rect 259748 211177 259776 220759
rect 259734 211168 259790 211177
rect 259734 211103 259790 211112
rect 259736 201476 259788 201482
rect 259736 201418 259788 201424
rect 259748 191865 259776 201418
rect 259734 191856 259790 191865
rect 259734 191791 259790 191800
rect 259276 180804 259328 180810
rect 259276 180746 259328 180752
rect 259368 180804 259420 180810
rect 259368 180746 259420 180752
rect 259288 171170 259316 180746
rect 259288 171142 259408 171170
rect 259380 171086 259408 171142
rect 259368 171080 259420 171086
rect 259368 171022 259420 171028
rect 259368 161560 259420 161566
rect 259368 161502 259420 161508
rect 259380 160070 259408 161502
rect 259368 160064 259420 160070
rect 259368 160006 259420 160012
rect 259276 142180 259328 142186
rect 259276 142122 259328 142128
rect 259288 122806 259316 142122
rect 259276 122800 259328 122806
rect 259276 122742 259328 122748
rect 259368 122732 259420 122738
rect 259368 122674 259420 122680
rect 259380 85814 259408 122674
rect 259368 85808 259420 85814
rect 259368 85750 259420 85756
rect 259276 85740 259328 85746
rect 259276 85682 259328 85688
rect 259288 84182 259316 85682
rect 259276 84176 259328 84182
rect 259276 84118 259328 84124
rect 259368 74588 259420 74594
rect 259368 74530 259420 74536
rect 259380 66298 259408 74530
rect 259276 66292 259328 66298
rect 259276 66234 259328 66240
rect 259368 66292 259420 66298
rect 259368 66234 259420 66240
rect 259288 43518 259316 66234
rect 259276 43512 259328 43518
rect 259276 43454 259328 43460
rect 259460 43512 259512 43518
rect 259460 43454 259512 43460
rect 259472 35902 259500 43454
rect 259460 35896 259512 35902
rect 259460 35838 259512 35844
rect 259276 26308 259328 26314
rect 259276 26250 259328 26256
rect 259288 11234 259316 26250
rect 259196 11206 259316 11234
rect 259196 7426 259224 11206
rect 259840 9178 259868 336874
rect 259932 334830 259960 340054
rect 260024 336802 260052 340068
rect 260116 337074 260144 340068
rect 260208 337414 260236 340068
rect 260196 337408 260248 337414
rect 260196 337350 260248 337356
rect 260104 337068 260156 337074
rect 260104 337010 260156 337016
rect 260012 336796 260064 336802
rect 260012 336738 260064 336744
rect 260300 335730 260328 340068
rect 260484 337210 260512 340068
rect 260576 337346 260604 340068
rect 260564 337340 260616 337346
rect 260564 337282 260616 337288
rect 260472 337204 260524 337210
rect 260472 337146 260524 337152
rect 260564 337068 260616 337074
rect 260564 337010 260616 337016
rect 260472 336796 260524 336802
rect 260472 336738 260524 336744
rect 260024 335702 260328 335730
rect 259920 334824 259972 334830
rect 259920 334766 259972 334772
rect 259920 280152 259972 280158
rect 259920 280094 259972 280100
rect 259932 278730 259960 280094
rect 259920 278724 259972 278730
rect 259920 278666 259972 278672
rect 259920 244996 259972 245002
rect 259920 244938 259972 244944
rect 259932 235346 259960 244938
rect 259920 235340 259972 235346
rect 259920 235282 259972 235288
rect 260024 212634 260052 335702
rect 260196 334824 260248 334830
rect 260196 334766 260248 334772
rect 260208 307766 260236 334766
rect 260380 334076 260432 334082
rect 260380 334018 260432 334024
rect 260392 307766 260420 334018
rect 260196 307760 260248 307766
rect 260196 307702 260248 307708
rect 260380 307760 260432 307766
rect 260380 307702 260432 307708
rect 260288 299396 260340 299402
rect 260288 299338 260340 299344
rect 260300 281994 260328 299338
rect 260104 281988 260156 281994
rect 260104 281930 260156 281936
rect 260288 281988 260340 281994
rect 260288 281930 260340 281936
rect 260116 280158 260144 281930
rect 260288 280220 260340 280226
rect 260288 280162 260340 280168
rect 260104 280152 260156 280158
rect 260104 280094 260156 280100
rect 260300 275330 260328 280162
rect 260288 275324 260340 275330
rect 260288 275266 260340 275272
rect 260104 267776 260156 267782
rect 260104 267718 260156 267724
rect 260116 258058 260144 267718
rect 260380 259480 260432 259486
rect 260380 259422 260432 259428
rect 260392 258058 260420 259422
rect 260104 258052 260156 258058
rect 260104 257994 260156 258000
rect 260380 258052 260432 258058
rect 260380 257994 260432 258000
rect 260104 249756 260156 249762
rect 260104 249698 260156 249704
rect 260116 245002 260144 249698
rect 260196 248464 260248 248470
rect 260196 248406 260248 248412
rect 260104 244996 260156 245002
rect 260104 244938 260156 244944
rect 260208 240106 260236 248406
rect 260196 240100 260248 240106
rect 260196 240042 260248 240048
rect 260196 235340 260248 235346
rect 260196 235282 260248 235288
rect 260208 222222 260236 235282
rect 260288 230512 260340 230518
rect 260288 230454 260340 230460
rect 260300 222358 260328 230454
rect 260288 222352 260340 222358
rect 260288 222294 260340 222300
rect 260104 222216 260156 222222
rect 260104 222158 260156 222164
rect 260196 222216 260248 222222
rect 260196 222158 260248 222164
rect 260288 222216 260340 222222
rect 260288 222158 260340 222164
rect 260116 220833 260144 222158
rect 260300 220833 260328 222158
rect 260102 220824 260158 220833
rect 260102 220759 260158 220768
rect 260286 220824 260342 220833
rect 260286 220759 260342 220768
rect 260012 212628 260064 212634
rect 260012 212570 260064 212576
rect 260012 212492 260064 212498
rect 260012 212434 260064 212440
rect 259918 211168 259974 211177
rect 259918 211103 259974 211112
rect 259932 202910 259960 211103
rect 259920 202904 259972 202910
rect 259920 202846 259972 202852
rect 259918 191856 259974 191865
rect 259918 191791 259974 191800
rect 259932 186318 259960 191791
rect 259920 186312 259972 186318
rect 259920 186254 259972 186260
rect 259918 183560 259974 183569
rect 259918 183495 259974 183504
rect 259932 178770 259960 183495
rect 259920 178764 259972 178770
rect 259920 178706 259972 178712
rect 260024 19446 260052 212434
rect 260194 211168 260250 211177
rect 260194 211103 260250 211112
rect 260208 202910 260236 211103
rect 260104 202904 260156 202910
rect 260104 202846 260156 202852
rect 260196 202904 260248 202910
rect 260196 202846 260248 202852
rect 260288 202904 260340 202910
rect 260288 202846 260340 202852
rect 260116 201482 260144 202846
rect 260300 201482 260328 202846
rect 260104 201476 260156 201482
rect 260104 201418 260156 201424
rect 260288 201476 260340 201482
rect 260288 201418 260340 201424
rect 260196 191888 260248 191894
rect 260196 191830 260248 191836
rect 260208 188442 260236 191830
rect 260208 188414 260328 188442
rect 260104 186312 260156 186318
rect 260104 186254 260156 186260
rect 260116 183569 260144 186254
rect 260102 183560 260158 183569
rect 260300 183530 260328 188414
rect 260102 183495 260158 183504
rect 260288 183524 260340 183530
rect 260288 183466 260340 183472
rect 260104 178764 260156 178770
rect 260104 178706 260156 178712
rect 260288 178764 260340 178770
rect 260288 178706 260340 178712
rect 260116 164218 260144 178706
rect 260300 164218 260328 178706
rect 260104 164212 260156 164218
rect 260104 164154 260156 164160
rect 260196 164212 260248 164218
rect 260196 164154 260248 164160
rect 260288 164212 260340 164218
rect 260288 164154 260340 164160
rect 260380 164212 260432 164218
rect 260380 164154 260432 164160
rect 260208 162858 260236 164154
rect 260196 162852 260248 162858
rect 260196 162794 260248 162800
rect 260392 154698 260420 164154
rect 260380 154692 260432 154698
rect 260380 154634 260432 154640
rect 260288 154556 260340 154562
rect 260288 154498 260340 154504
rect 260196 153332 260248 153338
rect 260196 153274 260248 153280
rect 260208 145081 260236 153274
rect 260194 145072 260250 145081
rect 260194 145007 260250 145016
rect 260102 144936 260158 144945
rect 260300 144906 260328 154498
rect 260102 144871 260104 144880
rect 260156 144871 260158 144880
rect 260196 144900 260248 144906
rect 260104 144842 260156 144848
rect 260196 144842 260248 144848
rect 260288 144900 260340 144906
rect 260288 144842 260340 144848
rect 260380 144900 260432 144906
rect 260380 144842 260432 144848
rect 260104 138712 260156 138718
rect 260104 138654 260156 138660
rect 260116 134065 260144 138654
rect 260102 134056 260158 134065
rect 260102 133991 260158 134000
rect 260208 125662 260236 144842
rect 260392 138718 260420 144842
rect 260380 138712 260432 138718
rect 260380 138654 260432 138660
rect 260286 133920 260342 133929
rect 260286 133855 260288 133864
rect 260340 133855 260342 133864
rect 260288 133826 260340 133832
rect 260104 125656 260156 125662
rect 260104 125598 260156 125604
rect 260196 125656 260248 125662
rect 260196 125598 260248 125604
rect 260116 124166 260144 125598
rect 260288 124296 260340 124302
rect 260288 124238 260340 124244
rect 260300 124166 260328 124238
rect 260104 124160 260156 124166
rect 260104 124102 260156 124108
rect 260288 124160 260340 124166
rect 260288 124102 260340 124108
rect 260196 114572 260248 114578
rect 260196 114514 260248 114520
rect 260380 114572 260432 114578
rect 260380 114514 260432 114520
rect 260208 104938 260236 114514
rect 260392 104938 260420 114514
rect 260116 104910 260236 104938
rect 260300 104910 260420 104938
rect 260116 102134 260144 104910
rect 260104 102128 260156 102134
rect 260104 102070 260156 102076
rect 260300 99414 260328 104910
rect 260288 99408 260340 99414
rect 260288 99350 260340 99356
rect 260380 99340 260432 99346
rect 260380 99282 260432 99288
rect 260196 92540 260248 92546
rect 260196 92482 260248 92488
rect 260208 72570 260236 92482
rect 260392 86562 260420 99282
rect 260380 86556 260432 86562
rect 260380 86498 260432 86504
rect 260380 75948 260432 75954
rect 260380 75890 260432 75896
rect 260116 72542 260236 72570
rect 260116 67590 260144 72542
rect 260392 72434 260420 75890
rect 260208 72406 260420 72434
rect 260104 67584 260156 67590
rect 260104 67526 260156 67532
rect 260208 67538 260236 72406
rect 260208 67510 260328 67538
rect 260196 67448 260248 67454
rect 260196 67390 260248 67396
rect 260208 48414 260236 67390
rect 260300 58002 260328 67510
rect 260288 57996 260340 58002
rect 260288 57938 260340 57944
rect 260380 57996 260432 58002
rect 260380 57938 260432 57944
rect 260392 48414 260420 57938
rect 260196 48408 260248 48414
rect 260196 48350 260248 48356
rect 260380 48408 260432 48414
rect 260380 48350 260432 48356
rect 260104 46980 260156 46986
rect 260104 46922 260156 46928
rect 260288 46980 260340 46986
rect 260288 46922 260340 46928
rect 260116 19514 260144 46922
rect 260104 19508 260156 19514
rect 260104 19450 260156 19456
rect 260012 19440 260064 19446
rect 260012 19382 260064 19388
rect 260300 19378 260328 46922
rect 260104 19372 260156 19378
rect 260104 19314 260156 19320
rect 260288 19372 260340 19378
rect 260288 19314 260340 19320
rect 260012 19304 260064 19310
rect 260012 19246 260064 19252
rect 259920 18012 259972 18018
rect 259920 17954 259972 17960
rect 259932 17882 259960 17954
rect 259920 17876 259972 17882
rect 259920 17818 259972 17824
rect 260024 9246 260052 19246
rect 260116 18057 260144 19314
rect 260102 18048 260158 18057
rect 260102 17983 260158 17992
rect 260378 18048 260434 18057
rect 260378 17983 260434 17992
rect 260392 17882 260420 17983
rect 260104 17876 260156 17882
rect 260104 17818 260156 17824
rect 260380 17876 260432 17882
rect 260380 17818 260432 17824
rect 260012 9240 260064 9246
rect 260012 9182 260064 9188
rect 259828 9172 259880 9178
rect 259828 9114 259880 9120
rect 259196 7398 259316 7426
rect 259288 5302 259316 7398
rect 259276 5296 259328 5302
rect 259276 5238 259328 5244
rect 258908 5228 258960 5234
rect 258908 5170 258960 5176
rect 258816 5092 258868 5098
rect 258816 5034 258868 5040
rect 260116 4826 260144 17818
rect 260484 9314 260512 336738
rect 260576 333742 260604 337010
rect 260668 336938 260696 340068
rect 260852 337074 260880 340068
rect 260944 337550 260972 340068
rect 261050 340054 261156 340082
rect 260932 337544 260984 337550
rect 260932 337486 260984 337492
rect 260932 337136 260984 337142
rect 260932 337078 260984 337084
rect 260840 337068 260892 337074
rect 260840 337010 260892 337016
rect 260656 336932 260708 336938
rect 260656 336874 260708 336880
rect 260840 336864 260892 336870
rect 260840 336806 260892 336812
rect 260656 336796 260708 336802
rect 260656 336738 260708 336744
rect 260564 333736 260616 333742
rect 260564 333678 260616 333684
rect 260668 332382 260696 336738
rect 260656 332376 260708 332382
rect 260656 332318 260708 332324
rect 260852 322522 260880 336806
rect 260944 336802 260972 337078
rect 261024 337000 261076 337006
rect 261024 336942 261076 336948
rect 260932 336796 260984 336802
rect 260932 336738 260984 336744
rect 260840 322516 260892 322522
rect 260840 322458 260892 322464
rect 261036 310010 261064 336942
rect 261128 333418 261156 340054
rect 261220 336938 261248 340068
rect 261312 337142 261340 340068
rect 261300 337136 261352 337142
rect 261300 337078 261352 337084
rect 261208 336932 261260 336938
rect 261208 336874 261260 336880
rect 261300 336796 261352 336802
rect 261300 336738 261352 336744
rect 261208 336660 261260 336666
rect 261208 336602 261260 336608
rect 261220 333538 261248 336602
rect 261208 333532 261260 333538
rect 261208 333474 261260 333480
rect 261128 333390 261248 333418
rect 261024 310004 261076 310010
rect 261024 309946 261076 309952
rect 260564 307760 260616 307766
rect 260564 307702 260616 307708
rect 260576 280226 260604 307702
rect 260564 280220 260616 280226
rect 260564 280162 260616 280168
rect 260564 275324 260616 275330
rect 260564 275266 260616 275272
rect 260576 259486 260604 275266
rect 260564 259480 260616 259486
rect 260564 259422 260616 259428
rect 260562 220824 260618 220833
rect 260562 220759 260618 220768
rect 260576 211177 260604 220759
rect 260562 211168 260618 211177
rect 260562 211103 260618 211112
rect 260472 9308 260524 9314
rect 260472 9250 260524 9256
rect 261220 8974 261248 333390
rect 261312 9042 261340 336738
rect 261404 9110 261432 340068
rect 261484 337272 261536 337278
rect 261484 337214 261536 337220
rect 261496 333674 261524 337214
rect 261588 336870 261616 340068
rect 261680 337278 261708 340068
rect 261668 337272 261720 337278
rect 261668 337214 261720 337220
rect 261668 337136 261720 337142
rect 261668 337078 261720 337084
rect 261576 336864 261628 336870
rect 261576 336806 261628 336812
rect 261576 336728 261628 336734
rect 261576 336670 261628 336676
rect 261484 333668 261536 333674
rect 261484 333610 261536 333616
rect 261484 333532 261536 333538
rect 261484 333474 261536 333480
rect 261392 9104 261444 9110
rect 261392 9046 261444 9052
rect 261300 9036 261352 9042
rect 261300 8978 261352 8984
rect 261208 8968 261260 8974
rect 261208 8910 261260 8916
rect 260196 8356 260248 8362
rect 260196 8298 260248 8304
rect 260208 4894 260236 8298
rect 261496 8294 261524 333474
rect 261588 319462 261616 336670
rect 261680 336530 261708 337078
rect 261772 336802 261800 340068
rect 261852 337068 261904 337074
rect 261852 337010 261904 337016
rect 261760 336796 261812 336802
rect 261760 336738 261812 336744
rect 261668 336524 261720 336530
rect 261668 336466 261720 336472
rect 261864 328098 261892 337010
rect 261956 337006 261984 340068
rect 262048 337090 262076 340068
rect 262140 337210 262168 340068
rect 262324 337754 262352 340068
rect 262416 337822 262444 340068
rect 262404 337816 262456 337822
rect 262404 337758 262456 337764
rect 262220 337748 262272 337754
rect 262220 337690 262272 337696
rect 262312 337748 262364 337754
rect 262312 337690 262364 337696
rect 262128 337204 262180 337210
rect 262128 337146 262180 337152
rect 262048 337062 262168 337090
rect 261944 337000 261996 337006
rect 261944 336942 261996 336948
rect 262036 336932 262088 336938
rect 262036 336874 262088 336880
rect 261944 336864 261996 336870
rect 261944 336806 261996 336812
rect 261956 332314 261984 336806
rect 261944 332308 261996 332314
rect 261944 332250 261996 332256
rect 262048 329526 262076 336874
rect 262140 335034 262168 337062
rect 262232 336802 262260 337690
rect 262508 337260 262536 340068
rect 262324 337232 262536 337260
rect 262600 340054 262706 340082
rect 262220 336796 262272 336802
rect 262220 336738 262272 336744
rect 262128 335028 262180 335034
rect 262128 334970 262180 334976
rect 262324 334966 262352 337232
rect 262404 337000 262456 337006
rect 262404 336942 262456 336948
rect 262312 334960 262364 334966
rect 262312 334902 262364 334908
rect 262036 329520 262088 329526
rect 262036 329462 262088 329468
rect 261852 328092 261904 328098
rect 261852 328034 261904 328040
rect 261576 319456 261628 319462
rect 261576 319398 261628 319404
rect 262416 318306 262444 336942
rect 262496 336796 262548 336802
rect 262496 336738 262548 336744
rect 262508 330954 262536 336738
rect 262496 330948 262548 330954
rect 262496 330890 262548 330896
rect 262600 319734 262628 340054
rect 262784 337074 262812 340068
rect 262772 337068 262824 337074
rect 262772 337010 262824 337016
rect 262772 336932 262824 336938
rect 262772 336874 262824 336880
rect 262680 336864 262732 336870
rect 262680 336806 262732 336812
rect 262588 319728 262640 319734
rect 262588 319670 262640 319676
rect 262404 318300 262456 318306
rect 262404 318242 262456 318248
rect 261484 8288 261536 8294
rect 261484 8230 261536 8236
rect 262692 5574 262720 336806
rect 262784 5642 262812 336874
rect 262876 336802 262904 340068
rect 262956 337068 263008 337074
rect 262956 337010 263008 337016
rect 262864 336796 262916 336802
rect 262864 336738 262916 336744
rect 262864 336660 262916 336666
rect 262864 336602 262916 336608
rect 262876 333418 262904 336602
rect 262968 333606 262996 337010
rect 263060 337006 263088 340068
rect 263048 337000 263100 337006
rect 263048 336942 263100 336948
rect 263152 336870 263180 340068
rect 263140 336864 263192 336870
rect 263140 336806 263192 336812
rect 262956 333600 263008 333606
rect 262956 333542 263008 333548
rect 262876 333390 262996 333418
rect 262864 333328 262916 333334
rect 262864 333270 262916 333276
rect 262772 5636 262824 5642
rect 262772 5578 262824 5584
rect 262680 5568 262732 5574
rect 262680 5510 262732 5516
rect 260196 4888 260248 4894
rect 260196 4830 260248 4836
rect 260104 4820 260156 4826
rect 260104 4762 260156 4768
rect 262876 4146 262904 333270
rect 262968 6934 262996 333390
rect 263244 326738 263272 340068
rect 263336 340054 263442 340082
rect 263232 326732 263284 326738
rect 263232 326674 263284 326680
rect 263336 293350 263364 340054
rect 263416 337884 263468 337890
rect 263416 337826 263468 337832
rect 263428 333334 263456 337826
rect 263520 336938 263548 340068
rect 263612 337958 263640 340068
rect 263600 337952 263652 337958
rect 263600 337894 263652 337900
rect 263508 336932 263560 336938
rect 263796 336920 263824 340068
rect 263888 336954 263916 340068
rect 263980 337346 264008 340068
rect 263968 337340 264020 337346
rect 263968 337282 264020 337288
rect 263888 336926 264100 336954
rect 263508 336874 263560 336880
rect 263704 336892 263824 336920
rect 263416 333328 263468 333334
rect 263416 333270 263468 333276
rect 263704 330886 263732 336892
rect 263968 336864 264020 336870
rect 263968 336806 264020 336812
rect 263784 336796 263836 336802
rect 263784 336738 263836 336744
rect 263692 330880 263744 330886
rect 263692 330822 263744 330828
rect 263796 325242 263824 336738
rect 263784 325236 263836 325242
rect 263784 325178 263836 325184
rect 263980 308582 264008 336806
rect 263968 308576 264020 308582
rect 263968 308518 264020 308524
rect 263324 293344 263376 293350
rect 263324 293286 263376 293292
rect 262956 6928 263008 6934
rect 262956 6870 263008 6876
rect 264072 5710 264100 336926
rect 264164 336802 264192 340068
rect 264152 336796 264204 336802
rect 264152 336738 264204 336744
rect 264256 5778 264284 340068
rect 264362 340054 264468 340082
rect 264336 336796 264388 336802
rect 264336 336738 264388 336744
rect 264348 5846 264376 336738
rect 264440 334898 264468 340054
rect 264428 334892 264480 334898
rect 264428 334834 264480 334840
rect 264532 322454 264560 340068
rect 264624 336802 264652 340068
rect 264730 340054 264836 340082
rect 264612 336796 264664 336802
rect 264612 336738 264664 336744
rect 264808 335594 264836 340054
rect 264900 336870 264928 340068
rect 264992 337142 265020 340068
rect 264980 337136 265032 337142
rect 264980 337078 265032 337084
rect 264980 337000 265032 337006
rect 264980 336942 265032 336948
rect 264888 336864 264940 336870
rect 264888 336806 264940 336812
rect 264808 335566 264928 335594
rect 264900 329458 264928 335566
rect 264888 329452 264940 329458
rect 264888 329394 264940 329400
rect 264520 322448 264572 322454
rect 264520 322390 264572 322396
rect 264336 5840 264388 5846
rect 264336 5782 264388 5788
rect 264992 5794 265020 336942
rect 265084 10062 265112 340068
rect 265268 337278 265296 340068
rect 265256 337272 265308 337278
rect 265256 337214 265308 337220
rect 265164 337068 265216 337074
rect 265164 337010 265216 337016
rect 265176 323882 265204 337010
rect 265256 337000 265308 337006
rect 265256 336942 265308 336948
rect 265164 323876 265216 323882
rect 265164 323818 265216 323824
rect 265268 311794 265296 336942
rect 265360 336326 265388 340068
rect 265452 336938 265480 340068
rect 265532 337816 265584 337822
rect 265532 337758 265584 337764
rect 265440 336932 265492 336938
rect 265440 336874 265492 336880
rect 265544 336462 265572 337758
rect 265636 337482 265664 340068
rect 265624 337476 265676 337482
rect 265624 337418 265676 337424
rect 265624 336864 265676 336870
rect 265624 336806 265676 336812
rect 265532 336456 265584 336462
rect 265532 336398 265584 336404
rect 265348 336320 265400 336326
rect 265348 336262 265400 336268
rect 265532 336320 265584 336326
rect 265532 336262 265584 336268
rect 265544 318850 265572 336262
rect 265348 318844 265400 318850
rect 265348 318786 265400 318792
rect 265532 318844 265584 318850
rect 265532 318786 265584 318792
rect 265360 318730 265388 318786
rect 265360 318702 265572 318730
rect 265268 311766 265388 311794
rect 265072 10056 265124 10062
rect 265072 9998 265124 10004
rect 265360 6118 265388 311766
rect 265348 6112 265400 6118
rect 265348 6054 265400 6060
rect 265544 5982 265572 318702
rect 265636 10266 265664 336806
rect 265728 336802 265756 340068
rect 265716 336796 265768 336802
rect 265716 336738 265768 336744
rect 265820 333282 265848 340068
rect 265900 337136 265952 337142
rect 265900 337078 265952 337084
rect 265912 336954 265940 337078
rect 266004 337074 266032 340068
rect 265992 337068 266044 337074
rect 265992 337010 266044 337016
rect 266096 337006 266124 340068
rect 266084 337000 266136 337006
rect 265912 336926 266032 336954
rect 266084 336942 266136 336948
rect 265900 336796 265952 336802
rect 265900 336738 265952 336744
rect 265728 333254 265848 333282
rect 265624 10260 265676 10266
rect 265624 10202 265676 10208
rect 265728 10198 265756 333254
rect 265912 326398 265940 336738
rect 265900 326392 265952 326398
rect 265900 326334 265952 326340
rect 265900 326256 265952 326262
rect 265900 326198 265952 326204
rect 265716 10192 265768 10198
rect 265716 10134 265768 10140
rect 265912 10130 265940 326198
rect 265900 10124 265952 10130
rect 265900 10066 265952 10072
rect 265532 5976 265584 5982
rect 265532 5918 265584 5924
rect 266004 5914 266032 336926
rect 266188 336870 266216 340068
rect 266372 337822 266400 340068
rect 266360 337816 266412 337822
rect 266360 337758 266412 337764
rect 266360 337000 266412 337006
rect 266360 336942 266412 336948
rect 266268 336932 266320 336938
rect 266268 336874 266320 336880
rect 266176 336864 266228 336870
rect 266176 336806 266228 336812
rect 266084 336796 266136 336802
rect 266084 336738 266136 336744
rect 266096 333538 266124 336738
rect 266084 333532 266136 333538
rect 266084 333474 266136 333480
rect 266084 326392 266136 326398
rect 266084 326334 266136 326340
rect 266096 6050 266124 326334
rect 266280 326262 266308 336874
rect 266268 326256 266320 326262
rect 266268 326198 266320 326204
rect 266372 10810 266400 336942
rect 266360 10804 266412 10810
rect 266360 10746 266412 10752
rect 266464 6866 266492 340068
rect 266556 11014 266584 340068
rect 266740 337074 266768 340068
rect 266728 337068 266780 337074
rect 266728 337010 266780 337016
rect 266728 336932 266780 336938
rect 266728 336874 266780 336880
rect 266636 336796 266688 336802
rect 266636 336738 266688 336744
rect 266648 326670 266676 336738
rect 266636 326664 266688 326670
rect 266636 326606 266688 326612
rect 266544 11008 266596 11014
rect 266544 10950 266596 10956
rect 266452 6860 266504 6866
rect 266452 6802 266504 6808
rect 266740 6730 266768 336874
rect 266832 6798 266860 340068
rect 266924 336870 266952 340068
rect 267004 337816 267056 337822
rect 267004 337758 267056 337764
rect 266912 336864 266964 336870
rect 266912 336806 266964 336812
rect 267016 336326 267044 337758
rect 267108 336802 267136 340068
rect 267200 336938 267228 340068
rect 267188 336932 267240 336938
rect 267188 336874 267240 336880
rect 267096 336796 267148 336802
rect 267096 336738 267148 336744
rect 267188 336796 267240 336802
rect 267188 336738 267240 336744
rect 267004 336320 267056 336326
rect 267004 336262 267056 336268
rect 267200 316946 267228 336738
rect 267188 316940 267240 316946
rect 267188 316882 267240 316888
rect 267292 10878 267320 340068
rect 267372 336864 267424 336870
rect 267372 336806 267424 336812
rect 267384 10946 267412 336806
rect 267476 336802 267504 340068
rect 267568 338094 267596 340068
rect 267556 338088 267608 338094
rect 267556 338030 267608 338036
rect 267660 337006 267688 340068
rect 267740 337952 267792 337958
rect 267740 337894 267792 337900
rect 267648 337000 267700 337006
rect 267648 336942 267700 336948
rect 267648 336864 267700 336870
rect 267648 336806 267700 336812
rect 267464 336796 267516 336802
rect 267464 336738 267516 336744
rect 267660 332178 267688 336806
rect 267752 336394 267780 337894
rect 267740 336388 267792 336394
rect 267740 336330 267792 336336
rect 267648 332172 267700 332178
rect 267648 332114 267700 332120
rect 267844 329390 267872 340068
rect 267936 337822 267964 340068
rect 267924 337816 267976 337822
rect 267924 337758 267976 337764
rect 267924 337000 267976 337006
rect 267924 336942 267976 336948
rect 267832 329384 267884 329390
rect 267832 329326 267884 329332
rect 267464 328500 267516 328506
rect 267464 328442 267516 328448
rect 267372 10940 267424 10946
rect 267372 10882 267424 10888
rect 267280 10872 267332 10878
rect 267280 10814 267332 10820
rect 267004 8288 267056 8294
rect 267004 8230 267056 8236
rect 266820 6792 266872 6798
rect 266820 6734 266872 6740
rect 266728 6724 266780 6730
rect 266728 6666 266780 6672
rect 266084 6044 266136 6050
rect 266084 5986 266136 5992
rect 265992 5908 266044 5914
rect 265992 5850 266044 5856
rect 264244 5772 264296 5778
rect 264992 5766 265848 5794
rect 264244 5714 264296 5720
rect 264060 5704 264112 5710
rect 264060 5646 264112 5652
rect 258448 4140 258500 4146
rect 258448 4082 258500 4088
rect 259828 4140 259880 4146
rect 259828 4082 259880 4088
rect 262864 4140 262916 4146
rect 262864 4082 262916 4088
rect 264612 4140 264664 4146
rect 264612 4082 264664 4088
rect 258632 4072 258684 4078
rect 258632 4014 258684 4020
rect 257988 3936 258040 3942
rect 257988 3878 258040 3884
rect 257896 3868 257948 3874
rect 257896 3810 257948 3816
rect 258644 480 258672 4014
rect 259840 480 259868 4082
rect 261024 4004 261076 4010
rect 261024 3946 261076 3952
rect 261036 480 261064 3946
rect 262220 3936 262272 3942
rect 262220 3878 262272 3884
rect 262232 480 262260 3878
rect 263416 3868 263468 3874
rect 263416 3810 263468 3816
rect 263428 480 263456 3810
rect 264624 480 264652 4082
rect 265820 480 265848 5766
rect 267016 480 267044 8230
rect 267476 6662 267504 328442
rect 267646 310992 267702 311001
rect 267646 310927 267702 310936
rect 267660 310593 267688 310927
rect 267646 310584 267702 310593
rect 267646 310519 267702 310528
rect 267464 6656 267516 6662
rect 267464 6598 267516 6604
rect 267936 6458 267964 336942
rect 268028 331294 268056 340068
rect 268016 331288 268068 331294
rect 268016 331230 268068 331236
rect 268016 329180 268068 329186
rect 268016 329122 268068 329128
rect 268028 318730 268056 329122
rect 268212 319666 268240 340068
rect 268304 336938 268332 340068
rect 268410 340054 268516 340082
rect 268292 336932 268344 336938
rect 268292 336874 268344 336880
rect 268292 336796 268344 336802
rect 268292 336738 268344 336744
rect 268200 319660 268252 319666
rect 268200 319602 268252 319608
rect 268028 318702 268148 318730
rect 268120 9466 268148 318702
rect 268304 315518 268332 336738
rect 268488 335594 268516 340054
rect 268580 336802 268608 340068
rect 268672 337006 268700 340068
rect 268660 337000 268712 337006
rect 268660 336942 268712 336948
rect 268568 336796 268620 336802
rect 268568 336738 268620 336744
rect 268660 336796 268712 336802
rect 268660 336738 268712 336744
rect 268488 335566 268608 335594
rect 268476 331220 268528 331226
rect 268476 331162 268528 331168
rect 268292 315512 268344 315518
rect 268292 315454 268344 315460
rect 268488 10742 268516 331162
rect 268476 10736 268528 10742
rect 268476 10678 268528 10684
rect 268580 10674 268608 335566
rect 268672 309942 268700 336738
rect 268660 309936 268712 309942
rect 268660 309878 268712 309884
rect 268568 10668 268620 10674
rect 268568 10610 268620 10616
rect 268764 10606 268792 340068
rect 268844 336932 268896 336938
rect 268844 336874 268896 336880
rect 268752 10600 268804 10606
rect 268752 10542 268804 10548
rect 268120 9438 268240 9466
rect 268108 6928 268160 6934
rect 268108 6870 268160 6876
rect 267924 6452 267976 6458
rect 267924 6394 267976 6400
rect 268120 480 268148 6870
rect 268212 6390 268240 9438
rect 268856 6526 268884 336874
rect 268948 336802 268976 340068
rect 268936 336796 268988 336802
rect 268936 336738 268988 336744
rect 269040 329186 269068 340068
rect 269028 329180 269080 329186
rect 269028 329122 269080 329128
rect 269132 325938 269160 340068
rect 269316 336954 269344 340068
rect 269224 336926 269344 336954
rect 269224 330818 269252 336926
rect 269304 335708 269356 335714
rect 269304 335650 269356 335656
rect 269212 330812 269264 330818
rect 269212 330754 269264 330760
rect 269132 325910 269252 325938
rect 269224 325718 269252 325910
rect 269028 325712 269080 325718
rect 269026 325680 269028 325689
rect 269120 325712 269172 325718
rect 269080 325680 269082 325689
rect 269120 325654 269172 325660
rect 269212 325712 269264 325718
rect 269212 325654 269264 325660
rect 269026 325615 269082 325624
rect 269028 318708 269080 318714
rect 269028 318650 269080 318656
rect 269040 6594 269068 318650
rect 269132 10538 269160 325654
rect 269210 325544 269266 325553
rect 269210 325479 269266 325488
rect 269224 318714 269252 325479
rect 269212 318708 269264 318714
rect 269212 318650 269264 318656
rect 269120 10532 269172 10538
rect 269120 10474 269172 10480
rect 269316 10402 269344 335650
rect 269408 335442 269436 340068
rect 269514 340054 269620 340082
rect 269488 336796 269540 336802
rect 269488 336738 269540 336744
rect 269396 335436 269448 335442
rect 269396 335378 269448 335384
rect 269304 10396 269356 10402
rect 269304 10338 269356 10344
rect 269028 6588 269080 6594
rect 269028 6530 269080 6536
rect 268844 6520 268896 6526
rect 268844 6462 268896 6468
rect 268200 6384 268252 6390
rect 268200 6326 268252 6332
rect 269500 6254 269528 336738
rect 269592 335510 269620 340054
rect 269580 335504 269632 335510
rect 269580 335446 269632 335452
rect 269580 335368 269632 335374
rect 269580 335310 269632 335316
rect 269488 6248 269540 6254
rect 269488 6190 269540 6196
rect 269304 4752 269356 4758
rect 269304 4694 269356 4700
rect 269316 480 269344 4694
rect 269592 2854 269620 335310
rect 269684 322386 269712 340068
rect 269776 336802 269804 340068
rect 269764 336796 269816 336802
rect 269764 336738 269816 336744
rect 269868 335714 269896 340068
rect 269960 340054 270066 340082
rect 269856 335708 269908 335714
rect 269856 335650 269908 335656
rect 269960 335594 269988 340054
rect 270040 336796 270092 336802
rect 270040 336738 270092 336744
rect 269868 335566 269988 335594
rect 269672 322380 269724 322386
rect 269672 322322 269724 322328
rect 269868 314158 269896 335566
rect 269948 335504 270000 335510
rect 269948 335446 270000 335452
rect 269856 314152 269908 314158
rect 269856 314094 269908 314100
rect 269960 10470 269988 335446
rect 269948 10464 270000 10470
rect 269948 10406 270000 10412
rect 270052 10334 270080 336738
rect 270144 335594 270172 340068
rect 270236 336802 270264 340068
rect 270328 340054 270434 340082
rect 270224 336796 270276 336802
rect 270224 336738 270276 336744
rect 270144 335566 270264 335594
rect 270132 335436 270184 335442
rect 270132 335378 270184 335384
rect 270040 10328 270092 10334
rect 270040 10270 270092 10276
rect 270144 6322 270172 335378
rect 270132 6316 270184 6322
rect 270132 6258 270184 6264
rect 270236 6186 270264 335566
rect 270328 335374 270356 340054
rect 270512 337142 270540 340068
rect 270500 337136 270552 337142
rect 270500 337078 270552 337084
rect 270604 336938 270632 340068
rect 270696 337113 270724 340190
rect 270880 337521 270908 340068
rect 270866 337512 270922 337521
rect 270866 337447 270922 337456
rect 270682 337104 270738 337113
rect 270682 337039 270738 337048
rect 270592 336932 270644 336938
rect 270592 336874 270644 336880
rect 270684 336796 270736 336802
rect 270684 336738 270736 336744
rect 270774 336798 270830 336807
rect 270316 335368 270368 335374
rect 270316 335310 270368 335316
rect 270500 316736 270552 316742
rect 270500 316678 270552 316684
rect 270408 227996 270460 228002
rect 270408 227938 270460 227944
rect 270420 227905 270448 227938
rect 270406 227896 270462 227905
rect 270406 227831 270462 227840
rect 270512 7614 270540 316678
rect 270500 7608 270552 7614
rect 270500 7550 270552 7556
rect 270224 6180 270276 6186
rect 270224 6122 270276 6128
rect 270500 5500 270552 5506
rect 270500 5442 270552 5448
rect 269580 2848 269632 2854
rect 269580 2790 269632 2796
rect 270512 480 270540 5442
rect 270696 2990 270724 336738
rect 270774 336733 270830 336742
rect 270788 322266 270816 336733
rect 270972 323814 271000 340068
rect 271156 337550 271184 340068
rect 271144 337544 271196 337550
rect 271144 337486 271196 337492
rect 271248 337278 271276 340068
rect 271354 340054 271460 340082
rect 271328 337340 271380 337346
rect 271328 337282 271380 337288
rect 271236 337272 271288 337278
rect 271236 337214 271288 337220
rect 271236 336932 271288 336938
rect 271236 336874 271288 336880
rect 271052 336796 271104 336802
rect 271052 336738 271104 336744
rect 270960 323808 271012 323814
rect 270960 323750 271012 323756
rect 270788 322238 271000 322266
rect 270972 278746 271000 322238
rect 270880 278718 271000 278746
rect 270880 269142 270908 278718
rect 270868 269136 270920 269142
rect 270774 269104 270830 269113
rect 270960 269136 271012 269142
rect 270868 269078 270920 269084
rect 270958 269104 270960 269113
rect 271012 269104 271014 269113
rect 270774 269039 270830 269048
rect 270958 269039 271014 269048
rect 270788 259486 270816 269039
rect 270776 259480 270828 259486
rect 270776 259422 270828 259428
rect 270960 259480 271012 259486
rect 270960 259422 271012 259428
rect 270972 249801 271000 259422
rect 270774 249792 270830 249801
rect 270774 249727 270830 249736
rect 270958 249792 271014 249801
rect 270958 249727 271014 249736
rect 270788 240174 270816 249727
rect 270776 240168 270828 240174
rect 270776 240110 270828 240116
rect 270960 240168 271012 240174
rect 270960 240110 271012 240116
rect 270972 220794 271000 240110
rect 270960 220788 271012 220794
rect 270960 220730 271012 220736
rect 270960 211200 271012 211206
rect 270960 211142 271012 211148
rect 270972 191826 271000 211142
rect 270960 191820 271012 191826
rect 270960 191762 271012 191768
rect 270960 182232 271012 182238
rect 270960 182174 271012 182180
rect 270972 180810 271000 182174
rect 270960 180804 271012 180810
rect 270960 180746 271012 180752
rect 270776 171148 270828 171154
rect 270776 171090 270828 171096
rect 270788 162897 270816 171090
rect 270774 162888 270830 162897
rect 270774 162823 270830 162832
rect 270774 162616 270830 162625
rect 270774 162551 270830 162560
rect 270788 153241 270816 162551
rect 270774 153232 270830 153241
rect 270774 153167 270830 153176
rect 270958 153232 271014 153241
rect 270958 153167 271014 153176
rect 270972 118726 271000 153167
rect 270960 118720 271012 118726
rect 270960 118662 271012 118668
rect 270960 118584 271012 118590
rect 270960 118526 271012 118532
rect 270684 2984 270736 2990
rect 270684 2926 270736 2932
rect 270972 2922 271000 118526
rect 271064 3058 271092 336738
rect 271248 325174 271276 336874
rect 271340 332246 271368 337282
rect 271328 332240 271380 332246
rect 271328 332182 271380 332188
rect 271236 325168 271288 325174
rect 271236 325110 271288 325116
rect 271432 311234 271460 340054
rect 271524 336802 271552 340068
rect 271512 336796 271564 336802
rect 271512 336738 271564 336744
rect 271616 333470 271644 340068
rect 271604 333464 271656 333470
rect 271604 333406 271656 333412
rect 271708 316878 271736 340068
rect 271892 336870 271920 340068
rect 271984 337958 272012 340068
rect 271972 337952 272024 337958
rect 271972 337894 272024 337900
rect 271880 336864 271932 336870
rect 271880 336806 271932 336812
rect 271972 336796 272024 336802
rect 271972 336738 272024 336744
rect 271696 316872 271748 316878
rect 271696 316814 271748 316820
rect 271420 311228 271472 311234
rect 271420 311170 271472 311176
rect 271696 7608 271748 7614
rect 271696 7550 271748 7556
rect 271052 3052 271104 3058
rect 271052 2994 271104 3000
rect 270960 2916 271012 2922
rect 270960 2858 271012 2864
rect 271708 480 271736 7550
rect 271984 3194 272012 336738
rect 272076 315450 272104 340068
rect 272156 336864 272208 336870
rect 272156 336806 272208 336812
rect 272168 335594 272196 336806
rect 272260 336802 272288 340068
rect 272352 337074 272380 340068
rect 272340 337068 272392 337074
rect 272340 337010 272392 337016
rect 272340 336932 272392 336938
rect 272340 336874 272392 336880
rect 272248 336796 272300 336802
rect 272248 336738 272300 336744
rect 272168 335566 272288 335594
rect 272156 335504 272208 335510
rect 272156 335446 272208 335452
rect 272168 321094 272196 335446
rect 272156 321088 272208 321094
rect 272156 321030 272208 321036
rect 272064 315444 272116 315450
rect 272064 315386 272116 315392
rect 272154 173904 272210 173913
rect 272154 173839 272210 173848
rect 272168 164257 272196 173839
rect 272154 164248 272210 164257
rect 272154 164183 272210 164192
rect 272154 74488 272210 74497
rect 272154 74423 272210 74432
rect 272168 64977 272196 74423
rect 272154 64968 272210 64977
rect 272154 64903 272210 64912
rect 271972 3188 272024 3194
rect 271972 3130 272024 3136
rect 272260 3126 272288 335566
rect 272352 329254 272380 336874
rect 272444 336802 272472 340068
rect 272524 337204 272576 337210
rect 272524 337146 272576 337152
rect 272432 336796 272484 336802
rect 272432 336738 272484 336744
rect 272536 335510 272564 337146
rect 272524 335504 272576 335510
rect 272524 335446 272576 335452
rect 272524 331220 272576 331226
rect 272524 331162 272576 331168
rect 272340 329248 272392 329254
rect 272340 329190 272392 329196
rect 272536 326466 272564 331162
rect 272524 326460 272576 326466
rect 272524 326402 272576 326408
rect 272524 326256 272576 326262
rect 272524 326198 272576 326204
rect 272432 317484 272484 317490
rect 272432 317426 272484 317432
rect 272444 273358 272472 317426
rect 272432 273352 272484 273358
rect 272432 273294 272484 273300
rect 272340 273216 272392 273222
rect 272340 273158 272392 273164
rect 272352 241534 272380 273158
rect 272340 241528 272392 241534
rect 272340 241470 272392 241476
rect 272432 241528 272484 241534
rect 272432 241470 272484 241476
rect 272444 215422 272472 241470
rect 272432 215416 272484 215422
rect 272432 215358 272484 215364
rect 272340 215280 272392 215286
rect 272340 215222 272392 215228
rect 272352 173913 272380 215222
rect 272338 173904 272394 173913
rect 272338 173839 272394 173848
rect 272338 164248 272394 164257
rect 272338 164183 272394 164192
rect 272352 157298 272380 164183
rect 272352 157270 272472 157298
rect 272444 130370 272472 157270
rect 272352 130342 272472 130370
rect 272352 125594 272380 130342
rect 272340 125588 272392 125594
rect 272340 125530 272392 125536
rect 272432 125588 272484 125594
rect 272432 125530 272484 125536
rect 272444 124166 272472 125530
rect 272432 124160 272484 124166
rect 272432 124102 272484 124108
rect 272432 111852 272484 111858
rect 272432 111794 272484 111800
rect 272444 111722 272472 111794
rect 272432 111716 272484 111722
rect 272432 111658 272484 111664
rect 272340 102196 272392 102202
rect 272340 102138 272392 102144
rect 272352 102082 272380 102138
rect 272352 102054 272472 102082
rect 272444 97306 272472 102054
rect 272432 97300 272484 97306
rect 272432 97242 272484 97248
rect 272340 74588 272392 74594
rect 272340 74530 272392 74536
rect 272352 74497 272380 74530
rect 272338 74488 272394 74497
rect 272338 74423 272394 74432
rect 272430 64968 272486 64977
rect 272430 64903 272486 64912
rect 272444 64870 272472 64903
rect 272432 64864 272484 64870
rect 272432 64806 272484 64812
rect 272340 64796 272392 64802
rect 272340 64738 272392 64744
rect 272352 3262 272380 64738
rect 272536 4214 272564 326198
rect 272628 317490 272656 340068
rect 272720 336938 272748 340068
rect 272708 336932 272760 336938
rect 272708 336874 272760 336880
rect 272708 336796 272760 336802
rect 272708 336738 272760 336744
rect 272616 317484 272668 317490
rect 272616 317426 272668 317432
rect 272720 307222 272748 336738
rect 272708 307216 272760 307222
rect 272708 307158 272760 307164
rect 272812 305726 272840 340068
rect 272892 336796 272944 336802
rect 272892 336738 272944 336744
rect 272800 305720 272852 305726
rect 272800 305662 272852 305668
rect 272904 291922 272932 336738
rect 272892 291916 272944 291922
rect 272892 291858 272944 291864
rect 272616 124160 272668 124166
rect 272616 124102 272668 124108
rect 272628 121446 272656 124102
rect 272616 121440 272668 121446
rect 272616 121382 272668 121388
rect 272892 5364 272944 5370
rect 272892 5306 272944 5312
rect 272524 4208 272576 4214
rect 272524 4150 272576 4156
rect 272340 3256 272392 3262
rect 272340 3198 272392 3204
rect 272248 3120 272300 3126
rect 272248 3062 272300 3068
rect 272904 480 272932 5306
rect 272996 3330 273024 340068
rect 273088 337210 273116 340068
rect 273076 337204 273128 337210
rect 273076 337146 273128 337152
rect 273076 337068 273128 337074
rect 273076 337010 273128 337016
rect 273088 330750 273116 337010
rect 273180 336802 273208 340068
rect 273364 337074 273392 340068
rect 273456 337346 273484 340068
rect 273444 337340 273496 337346
rect 273444 337282 273496 337288
rect 273352 337068 273404 337074
rect 273352 337010 273404 337016
rect 273444 337000 273496 337006
rect 273444 336942 273496 336948
rect 273260 336932 273312 336938
rect 273260 336874 273312 336880
rect 273168 336796 273220 336802
rect 273168 336738 273220 336744
rect 273076 330744 273128 330750
rect 273076 330686 273128 330692
rect 273272 326398 273300 336874
rect 273352 336864 273404 336870
rect 273352 336806 273404 336812
rect 273364 327962 273392 336806
rect 273352 327956 273404 327962
rect 273352 327898 273404 327904
rect 273260 326392 273312 326398
rect 273260 326334 273312 326340
rect 273456 4010 273484 336942
rect 273548 314090 273576 340068
rect 273628 336796 273680 336802
rect 273628 336738 273680 336744
rect 273640 325106 273668 336738
rect 273732 327162 273760 340068
rect 273824 336870 273852 340068
rect 273930 340054 274036 340082
rect 273904 337816 273956 337822
rect 273904 337758 273956 337764
rect 273812 336864 273864 336870
rect 273812 336806 273864 336812
rect 273916 332042 273944 337758
rect 273904 332036 273956 332042
rect 273904 331978 273956 331984
rect 273732 327134 273944 327162
rect 273720 326392 273772 326398
rect 273720 326334 273772 326340
rect 273812 326392 273864 326398
rect 273812 326334 273864 326340
rect 273628 325100 273680 325106
rect 273628 325042 273680 325048
rect 273536 314084 273588 314090
rect 273536 314026 273588 314032
rect 273732 4078 273760 326334
rect 273720 4072 273772 4078
rect 273720 4014 273772 4020
rect 273444 4004 273496 4010
rect 273444 3946 273496 3952
rect 273824 3398 273852 326334
rect 273916 4146 273944 327134
rect 274008 323626 274036 340054
rect 274100 336938 274128 340068
rect 274088 336932 274140 336938
rect 274088 336874 274140 336880
rect 274192 336802 274220 340068
rect 274180 336796 274232 336802
rect 274180 336738 274232 336744
rect 274284 333282 274312 340068
rect 274364 337068 274416 337074
rect 274364 337010 274416 337016
rect 274192 333254 274312 333282
rect 274008 323598 274128 323626
rect 274100 304366 274128 323598
rect 274088 304360 274140 304366
rect 274088 304302 274140 304308
rect 274192 290562 274220 333254
rect 274376 326398 274404 337010
rect 274468 337006 274496 340068
rect 274560 337822 274588 340068
rect 274548 337816 274600 337822
rect 274548 337758 274600 337764
rect 274548 337340 274600 337346
rect 274548 337282 274600 337288
rect 274456 337000 274508 337006
rect 274456 336942 274508 336948
rect 274560 334830 274588 337282
rect 274548 334824 274600 334830
rect 274548 334766 274600 334772
rect 274652 326806 274680 340068
rect 274836 337142 274864 340068
rect 274928 338094 274956 340068
rect 274916 338088 274968 338094
rect 274916 338030 274968 338036
rect 274824 337136 274876 337142
rect 274824 337078 274876 337084
rect 274732 337068 274784 337074
rect 274732 337010 274784 337016
rect 274640 326800 274692 326806
rect 274640 326742 274692 326748
rect 274744 326602 274772 337010
rect 274824 336932 274876 336938
rect 274824 336874 274876 336880
rect 274836 333282 274864 336874
rect 274916 336864 274968 336870
rect 274916 336806 274968 336812
rect 274928 335594 274956 336806
rect 275020 336802 275048 340068
rect 275008 336796 275060 336802
rect 275008 336738 275060 336744
rect 274928 335566 275048 335594
rect 274836 333254 274956 333282
rect 274732 326596 274784 326602
rect 274732 326538 274784 326544
rect 274364 326392 274416 326398
rect 274364 326334 274416 326340
rect 274928 311166 274956 333254
rect 274916 311160 274968 311166
rect 274916 311102 274968 311108
rect 274180 290556 274232 290562
rect 274180 290498 274232 290504
rect 274916 27600 274968 27606
rect 274916 27542 274968 27548
rect 274928 26246 274956 27542
rect 274916 26240 274968 26246
rect 274916 26182 274968 26188
rect 274916 16652 274968 16658
rect 274916 16594 274968 16600
rect 274928 9586 274956 16594
rect 274916 9580 274968 9586
rect 274916 9522 274968 9528
rect 274088 5432 274140 5438
rect 274088 5374 274140 5380
rect 273904 4140 273956 4146
rect 273904 4082 273956 4088
rect 273812 3392 273864 3398
rect 273812 3334 273864 3340
rect 272984 3324 273036 3330
rect 272984 3266 273036 3272
rect 274100 480 274128 5374
rect 275020 3806 275048 335566
rect 275112 3874 275140 340068
rect 275190 337784 275246 337793
rect 275190 337719 275246 337728
rect 275204 337686 275232 337719
rect 275192 337680 275244 337686
rect 275192 337622 275244 337628
rect 275296 336258 275324 340068
rect 275388 336938 275416 340068
rect 275376 336932 275428 336938
rect 275376 336874 275428 336880
rect 275480 336870 275508 340068
rect 275664 337074 275692 340068
rect 275652 337068 275704 337074
rect 275652 337010 275704 337016
rect 275468 336864 275520 336870
rect 275468 336806 275520 336812
rect 275376 336796 275428 336802
rect 275376 336738 275428 336744
rect 275284 336252 275336 336258
rect 275284 336194 275336 336200
rect 275282 314800 275338 314809
rect 275282 314735 275338 314744
rect 275296 314650 275324 314735
rect 275204 314622 275324 314650
rect 275204 305046 275232 314622
rect 275388 312730 275416 336738
rect 275756 334914 275784 340068
rect 275572 334886 275784 334914
rect 275376 312724 275428 312730
rect 275376 312666 275428 312672
rect 275192 305040 275244 305046
rect 275192 304982 275244 304988
rect 275284 305040 275336 305046
rect 275284 304982 275336 304988
rect 275296 302326 275324 304982
rect 275572 303006 275600 334886
rect 275744 331152 275796 331158
rect 275744 331094 275796 331100
rect 275560 303000 275612 303006
rect 275560 302942 275612 302948
rect 275284 302320 275336 302326
rect 275284 302262 275336 302268
rect 275376 302116 275428 302122
rect 275376 302058 275428 302064
rect 275388 292670 275416 302058
rect 275376 292664 275428 292670
rect 275376 292606 275428 292612
rect 275284 292528 275336 292534
rect 275284 292470 275336 292476
rect 275296 287042 275324 292470
rect 275296 287014 275416 287042
rect 275388 282946 275416 287014
rect 275376 282940 275428 282946
rect 275376 282882 275428 282888
rect 275284 282872 275336 282878
rect 275284 282814 275336 282820
rect 275296 273850 275324 282814
rect 275296 273822 275416 273850
rect 275388 260982 275416 273822
rect 275376 260976 275428 260982
rect 275376 260918 275428 260924
rect 275284 260772 275336 260778
rect 275284 260714 275336 260720
rect 275296 249830 275324 260714
rect 275284 249824 275336 249830
rect 275284 249766 275336 249772
rect 275284 248464 275336 248470
rect 275284 248406 275336 248412
rect 275296 240174 275324 248406
rect 275284 240168 275336 240174
rect 275284 240110 275336 240116
rect 275376 240168 275428 240174
rect 275376 240110 275428 240116
rect 275388 238746 275416 240110
rect 275376 238740 275428 238746
rect 275376 238682 275428 238688
rect 275560 238740 275612 238746
rect 275560 238682 275612 238688
rect 275572 229129 275600 238682
rect 275374 229120 275430 229129
rect 275374 229055 275430 229064
rect 275558 229120 275614 229129
rect 275558 229055 275614 229064
rect 275388 225706 275416 229055
rect 275296 225678 275416 225706
rect 275296 209778 275324 225678
rect 275284 209772 275336 209778
rect 275284 209714 275336 209720
rect 275284 205624 275336 205630
rect 275284 205566 275336 205572
rect 275296 200138 275324 205566
rect 275296 200110 275416 200138
rect 275388 190670 275416 200110
rect 275376 190664 275428 190670
rect 275376 190606 275428 190612
rect 275284 190528 275336 190534
rect 275284 190470 275336 190476
rect 275296 186386 275324 190470
rect 275284 186380 275336 186386
rect 275284 186322 275336 186328
rect 275376 186244 275428 186250
rect 275376 186186 275428 186192
rect 275388 180810 275416 186186
rect 275376 180804 275428 180810
rect 275376 180746 275428 180752
rect 275192 171148 275244 171154
rect 275192 171090 275244 171096
rect 275204 171018 275232 171090
rect 275192 171012 275244 171018
rect 275192 170954 275244 170960
rect 275376 161492 275428 161498
rect 275376 161434 275428 161440
rect 275388 142186 275416 161434
rect 275376 142180 275428 142186
rect 275376 142122 275428 142128
rect 275468 142180 275520 142186
rect 275468 142122 275520 142128
rect 275480 135318 275508 142122
rect 275468 135312 275520 135318
rect 275468 135254 275520 135260
rect 275376 135244 275428 135250
rect 275376 135186 275428 135192
rect 275388 133890 275416 135186
rect 275376 133884 275428 133890
rect 275376 133826 275428 133832
rect 275376 124228 275428 124234
rect 275376 124170 275428 124176
rect 275388 119354 275416 124170
rect 275296 119326 275416 119354
rect 275296 93838 275324 119326
rect 275284 93832 275336 93838
rect 275284 93774 275336 93780
rect 275284 84244 275336 84250
rect 275284 84186 275336 84192
rect 275296 56574 275324 84186
rect 275284 56568 275336 56574
rect 275284 56510 275336 56516
rect 275284 51060 275336 51066
rect 275284 51002 275336 51008
rect 275296 37210 275324 51002
rect 275296 37182 275416 37210
rect 275388 27606 275416 37182
rect 275376 27600 275428 27606
rect 275376 27542 275428 27548
rect 275376 9580 275428 9586
rect 275376 9522 275428 9528
rect 275388 8294 275416 9522
rect 275376 8288 275428 8294
rect 275376 8230 275428 8236
rect 275284 4208 275336 4214
rect 275284 4150 275336 4156
rect 275100 3868 275152 3874
rect 275100 3810 275152 3816
rect 275008 3800 275060 3806
rect 275008 3742 275060 3748
rect 275296 480 275324 4150
rect 275756 3942 275784 331094
rect 275848 325825 275876 340068
rect 276032 337822 276060 340068
rect 276020 337816 276072 337822
rect 276020 337758 276072 337764
rect 276124 337006 276152 340068
rect 276112 337000 276164 337006
rect 276112 336942 276164 336948
rect 276020 336864 276072 336870
rect 276020 336806 276072 336812
rect 275834 325816 275890 325825
rect 275834 325751 275890 325760
rect 276032 289202 276060 336806
rect 276112 336728 276164 336734
rect 276112 336670 276164 336676
rect 276020 289196 276072 289202
rect 276020 289138 276072 289144
rect 275744 3936 275796 3942
rect 275744 3878 275796 3884
rect 276124 3466 276152 336670
rect 276216 334558 276244 340068
rect 276400 336802 276428 340068
rect 276492 336870 276520 340068
rect 276480 336864 276532 336870
rect 276480 336806 276532 336812
rect 276388 336796 276440 336802
rect 276388 336738 276440 336744
rect 276204 334552 276256 334558
rect 276204 334494 276256 334500
rect 276584 330052 276612 340068
rect 276664 336796 276716 336802
rect 276664 336738 276716 336744
rect 276676 330682 276704 336738
rect 276664 330676 276716 330682
rect 276664 330618 276716 330624
rect 276492 330024 276612 330052
rect 276388 329316 276440 329322
rect 276388 329258 276440 329264
rect 276296 326392 276348 326398
rect 276296 326334 276348 326340
rect 276308 287774 276336 326334
rect 276296 287768 276348 287774
rect 276296 287710 276348 287716
rect 276400 3534 276428 329258
rect 276492 144906 276520 330024
rect 276768 318238 276796 340068
rect 276756 318232 276808 318238
rect 276756 318174 276808 318180
rect 276860 300218 276888 340068
rect 276952 336938 276980 340068
rect 277032 337000 277084 337006
rect 277032 336942 277084 336948
rect 276940 336932 276992 336938
rect 276940 336874 276992 336880
rect 276940 336796 276992 336802
rect 276940 336738 276992 336744
rect 276952 326398 276980 336738
rect 276940 326392 276992 326398
rect 276940 326334 276992 326340
rect 277044 301578 277072 336942
rect 277136 334642 277164 340068
rect 277228 336802 277256 340068
rect 277320 336870 277348 340068
rect 277504 338026 277532 340068
rect 277492 338020 277544 338026
rect 277492 337962 277544 337968
rect 277596 337770 277624 340068
rect 277412 337742 277624 337770
rect 277308 336864 277360 336870
rect 277308 336806 277360 336812
rect 277216 336796 277268 336802
rect 277216 336738 277268 336744
rect 277136 334614 277348 334642
rect 277124 334552 277176 334558
rect 277124 334494 277176 334500
rect 277032 301572 277084 301578
rect 277032 301514 277084 301520
rect 276848 300212 276900 300218
rect 276848 300154 276900 300160
rect 276480 144900 276532 144906
rect 276480 144842 276532 144848
rect 276480 135312 276532 135318
rect 276480 135254 276532 135260
rect 276492 125610 276520 135254
rect 276492 125582 276612 125610
rect 276584 119406 276612 125582
rect 276572 119400 276624 119406
rect 276572 119342 276624 119348
rect 276480 107636 276532 107642
rect 276480 107578 276532 107584
rect 276492 19310 276520 107578
rect 276480 19304 276532 19310
rect 276480 19246 276532 19252
rect 276480 9716 276532 9722
rect 276480 9658 276532 9664
rect 276492 7970 276520 9658
rect 276492 7942 276612 7970
rect 276480 5296 276532 5302
rect 276480 5238 276532 5244
rect 276388 3528 276440 3534
rect 276388 3470 276440 3476
rect 276112 3460 276164 3466
rect 276112 3402 276164 3408
rect 276492 480 276520 5238
rect 276584 3602 276612 7942
rect 277136 3670 277164 334494
rect 277320 322318 277348 334614
rect 277412 327894 277440 337742
rect 277492 337612 277544 337618
rect 277492 337554 277544 337560
rect 277400 327888 277452 327894
rect 277400 327830 277452 327836
rect 277308 322312 277360 322318
rect 277308 322254 277360 322260
rect 277504 307154 277532 337554
rect 277584 336796 277636 336802
rect 277584 336738 277636 336744
rect 277492 307148 277544 307154
rect 277492 307090 277544 307096
rect 277596 298790 277624 336738
rect 277688 335578 277716 340068
rect 277872 338162 277900 340068
rect 277860 338156 277912 338162
rect 277860 338098 277912 338104
rect 277768 337408 277820 337414
rect 277768 337350 277820 337356
rect 277780 336802 277808 337350
rect 277860 337340 277912 337346
rect 277860 337282 277912 337288
rect 277768 336796 277820 336802
rect 277768 336738 277820 336744
rect 277676 335572 277728 335578
rect 277676 335514 277728 335520
rect 277676 335368 277728 335374
rect 277676 335310 277728 335316
rect 277584 298784 277636 298790
rect 277584 298726 277636 298732
rect 277688 8242 277716 335310
rect 277872 325038 277900 337282
rect 277964 336802 277992 340068
rect 277952 336796 278004 336802
rect 277952 336738 278004 336744
rect 278056 333198 278084 340068
rect 278136 338156 278188 338162
rect 278136 338098 278188 338104
rect 278148 337074 278176 338098
rect 278240 337074 278268 340068
rect 278332 337414 278360 340068
rect 278320 337408 278372 337414
rect 278320 337350 278372 337356
rect 278136 337068 278188 337074
rect 278136 337010 278188 337016
rect 278228 337068 278280 337074
rect 278228 337010 278280 337016
rect 278228 336796 278280 336802
rect 278228 336738 278280 336744
rect 278044 333192 278096 333198
rect 278044 333134 278096 333140
rect 277952 333124 278004 333130
rect 277952 333066 278004 333072
rect 277860 325032 277912 325038
rect 277860 324974 277912 324980
rect 277964 317490 277992 333066
rect 278044 333056 278096 333062
rect 278044 332998 278096 333004
rect 278056 323626 278084 332998
rect 278056 323598 278176 323626
rect 277860 317484 277912 317490
rect 277860 317426 277912 317432
rect 277952 317484 278004 317490
rect 277952 317426 278004 317432
rect 277872 304978 277900 317426
rect 278148 307834 278176 323598
rect 278240 321026 278268 336738
rect 278424 333062 278452 340068
rect 278504 338020 278556 338026
rect 278504 337962 278556 337968
rect 278516 336802 278544 337962
rect 278608 337346 278636 340068
rect 278700 337618 278728 340068
rect 278806 340054 278912 340082
rect 278780 338088 278832 338094
rect 278780 338030 278832 338036
rect 278688 337612 278740 337618
rect 278688 337554 278740 337560
rect 278686 337512 278742 337521
rect 278686 337447 278742 337456
rect 278596 337340 278648 337346
rect 278596 337282 278648 337288
rect 278596 337000 278648 337006
rect 278596 336942 278648 336948
rect 278504 336796 278556 336802
rect 278504 336738 278556 336744
rect 278608 333402 278636 336942
rect 278700 335186 278728 337447
rect 278792 337278 278820 338030
rect 278780 337272 278832 337278
rect 278780 337214 278832 337220
rect 278780 337068 278832 337074
rect 278780 337010 278832 337016
rect 278792 335322 278820 337010
rect 278884 335458 278912 340054
rect 278976 335594 279004 340068
rect 279068 337006 279096 340068
rect 279160 337074 279188 340068
rect 279240 337952 279292 337958
rect 279240 337894 279292 337900
rect 279252 337793 279280 337894
rect 279238 337784 279294 337793
rect 279238 337719 279294 337728
rect 279240 337136 279292 337142
rect 279240 337078 279292 337084
rect 279148 337068 279200 337074
rect 279148 337010 279200 337016
rect 279056 337000 279108 337006
rect 279056 336942 279108 336948
rect 279252 335730 279280 337078
rect 279344 336938 279372 340068
rect 279332 336932 279384 336938
rect 279332 336874 279384 336880
rect 279252 335702 279372 335730
rect 278976 335566 279280 335594
rect 278884 335430 279188 335458
rect 278792 335294 279096 335322
rect 278872 335232 278924 335238
rect 278700 335158 278820 335186
rect 278872 335174 278924 335180
rect 278596 333396 278648 333402
rect 278596 333338 278648 333344
rect 278412 333056 278464 333062
rect 278412 332998 278464 333004
rect 278792 332450 278820 335158
rect 278780 332444 278832 332450
rect 278780 332386 278832 332392
rect 278228 321020 278280 321026
rect 278228 320962 278280 320968
rect 278780 319456 278832 319462
rect 278780 319398 278832 319404
rect 278044 307828 278096 307834
rect 278044 307770 278096 307776
rect 278136 307828 278188 307834
rect 278136 307770 278188 307776
rect 278056 306377 278084 307770
rect 278042 306368 278098 306377
rect 278042 306303 278098 306312
rect 278318 306368 278374 306377
rect 278318 306303 278374 306312
rect 277860 304972 277912 304978
rect 277860 304914 277912 304920
rect 278228 304972 278280 304978
rect 278228 304914 278280 304920
rect 278136 296744 278188 296750
rect 278136 296686 278188 296692
rect 277950 295352 278006 295361
rect 277950 295287 278006 295296
rect 277964 289610 277992 295287
rect 277952 289604 278004 289610
rect 277952 289546 278004 289552
rect 277860 277432 277912 277438
rect 277860 277374 277912 277380
rect 278042 277400 278098 277409
rect 277872 254590 277900 277374
rect 278148 277386 278176 296686
rect 278240 295361 278268 304914
rect 278332 296750 278360 306303
rect 278320 296744 278372 296750
rect 278320 296686 278372 296692
rect 278226 295352 278282 295361
rect 278226 295287 278282 295296
rect 278098 277358 278176 277386
rect 278042 277335 278098 277344
rect 278318 277264 278374 277273
rect 278318 277199 278374 277208
rect 277860 254584 277912 254590
rect 277860 254526 277912 254532
rect 278044 254584 278096 254590
rect 278044 254526 278096 254532
rect 278056 248402 278084 254526
rect 277860 248396 277912 248402
rect 277860 248338 277912 248344
rect 278044 248396 278096 248402
rect 278044 248338 278096 248344
rect 277872 238785 277900 248338
rect 278332 241534 278360 277199
rect 278228 241528 278280 241534
rect 278228 241470 278280 241476
rect 278320 241528 278372 241534
rect 278320 241470 278372 241476
rect 277858 238776 277914 238785
rect 277768 238740 277820 238746
rect 277858 238711 277914 238720
rect 278042 238776 278098 238785
rect 278042 238711 278044 238720
rect 277768 238682 277820 238688
rect 278096 238711 278098 238720
rect 278044 238682 278096 238688
rect 277780 229129 277808 238682
rect 277766 229120 277822 229129
rect 277766 229055 277822 229064
rect 277950 229120 278006 229129
rect 277950 229055 278006 229064
rect 277964 225214 277992 229055
rect 277952 225208 278004 225214
rect 277952 225150 278004 225156
rect 277952 220856 278004 220862
rect 277952 220798 278004 220804
rect 277964 219434 277992 220798
rect 277952 219428 278004 219434
rect 277952 219370 278004 219376
rect 277860 209840 277912 209846
rect 277860 209782 277912 209788
rect 277872 205578 277900 209782
rect 278240 205714 278268 241470
rect 278056 205686 278268 205714
rect 277872 205550 277992 205578
rect 277964 191894 277992 205550
rect 278056 202881 278084 205686
rect 278042 202872 278098 202881
rect 278042 202807 278098 202816
rect 278226 202872 278282 202881
rect 278226 202807 278282 202816
rect 277952 191888 278004 191894
rect 277952 191830 278004 191836
rect 278044 191752 278096 191758
rect 278044 191694 278096 191700
rect 278056 190466 278084 191694
rect 277768 190460 277820 190466
rect 277768 190402 277820 190408
rect 278044 190460 278096 190466
rect 278044 190402 278096 190408
rect 277780 180849 277808 190402
rect 278240 186318 278268 202807
rect 278228 186312 278280 186318
rect 278228 186254 278280 186260
rect 278412 186312 278464 186318
rect 278412 186254 278464 186260
rect 277766 180840 277822 180849
rect 277766 180775 277822 180784
rect 277950 180840 278006 180849
rect 277950 180775 278006 180784
rect 277964 171154 277992 180775
rect 278424 178786 278452 186254
rect 278332 178758 278452 178786
rect 277860 171148 277912 171154
rect 277860 171090 277912 171096
rect 277952 171148 278004 171154
rect 277952 171090 278004 171096
rect 277872 161498 277900 171090
rect 277860 161492 277912 161498
rect 277860 161434 277912 161440
rect 278136 161492 278188 161498
rect 278136 161434 278188 161440
rect 278148 153218 278176 161434
rect 278056 153190 278176 153218
rect 278056 144888 278084 153190
rect 278332 147694 278360 178758
rect 278136 147688 278188 147694
rect 278136 147630 278188 147636
rect 278320 147688 278372 147694
rect 278320 147630 278372 147636
rect 277872 144860 278084 144888
rect 277872 128330 277900 144860
rect 278148 142882 278176 147630
rect 278056 142854 278176 142882
rect 278056 137986 278084 142854
rect 278056 137958 278176 137986
rect 278148 135250 278176 137958
rect 278136 135244 278188 135250
rect 278136 135186 278188 135192
rect 277872 128302 278084 128330
rect 278056 120714 278084 128302
rect 278228 128308 278280 128314
rect 278228 128250 278280 128256
rect 277964 120686 278084 120714
rect 277964 109154 277992 120686
rect 278240 114578 278268 128250
rect 278228 114572 278280 114578
rect 278228 114514 278280 114520
rect 277872 109126 277992 109154
rect 277872 109018 277900 109126
rect 277872 108990 278084 109018
rect 278056 101402 278084 108990
rect 278320 104916 278372 104922
rect 278320 104858 278372 104864
rect 277872 101374 278084 101402
rect 277872 99226 277900 101374
rect 277872 99198 277992 99226
rect 277964 89706 277992 99198
rect 278332 96665 278360 104858
rect 278134 96656 278190 96665
rect 278134 96591 278190 96600
rect 278318 96656 278374 96665
rect 278318 96591 278374 96600
rect 277780 89678 277992 89706
rect 277780 62778 277808 89678
rect 278148 80186 278176 96591
rect 278056 80158 278176 80186
rect 278056 80050 278084 80158
rect 278056 80022 278176 80050
rect 278148 67658 278176 80022
rect 278044 67652 278096 67658
rect 278044 67594 278096 67600
rect 278136 67652 278188 67658
rect 278136 67594 278188 67600
rect 277780 62750 277992 62778
rect 277964 26874 277992 62750
rect 278056 51066 278084 67594
rect 278044 51060 278096 51066
rect 278044 51002 278096 51008
rect 278228 51060 278280 51066
rect 278228 51002 278280 51008
rect 278240 46918 278268 51002
rect 278228 46912 278280 46918
rect 278228 46854 278280 46860
rect 278044 37324 278096 37330
rect 278044 37266 278096 37272
rect 278056 27538 278084 37266
rect 278044 27532 278096 27538
rect 278044 27474 278096 27480
rect 277964 26846 278084 26874
rect 278056 12458 278084 26846
rect 277596 8214 277716 8242
rect 277872 12430 278084 12458
rect 277596 4049 277624 8214
rect 277676 5228 277728 5234
rect 277676 5170 277728 5176
rect 277582 4040 277638 4049
rect 277582 3975 277638 3984
rect 277124 3664 277176 3670
rect 277124 3606 277176 3612
rect 276572 3596 276624 3602
rect 276572 3538 276624 3544
rect 277688 480 277716 5170
rect 277872 3913 277900 12430
rect 278228 9716 278280 9722
rect 278228 9658 278280 9664
rect 277858 3904 277914 3913
rect 277858 3839 277914 3848
rect 278240 3777 278268 9658
rect 278226 3768 278282 3777
rect 278226 3703 278282 3712
rect 278792 626 278820 319398
rect 278884 283626 278912 335174
rect 278964 335164 279016 335170
rect 278964 335106 279016 335112
rect 278976 323746 279004 335106
rect 279068 329186 279096 335294
rect 279160 330070 279188 335430
rect 279148 330064 279200 330070
rect 279148 330006 279200 330012
rect 279056 329180 279108 329186
rect 279056 329122 279108 329128
rect 278964 323740 279016 323746
rect 278964 323682 279016 323688
rect 279252 320958 279280 335566
rect 279344 335238 279372 335702
rect 279436 335594 279464 340068
rect 279528 336802 279556 340068
rect 279712 338094 279740 340068
rect 279700 338088 279752 338094
rect 279700 338030 279752 338036
rect 279608 337748 279660 337754
rect 279608 337690 279660 337696
rect 279516 336796 279568 336802
rect 279516 336738 279568 336744
rect 279620 336598 279648 337690
rect 279700 337000 279752 337006
rect 279700 336942 279752 336948
rect 279608 336592 279660 336598
rect 279608 336534 279660 336540
rect 279436 335566 279648 335594
rect 279516 335504 279568 335510
rect 279516 335446 279568 335452
rect 279332 335232 279384 335238
rect 279332 335174 279384 335180
rect 279240 320952 279292 320958
rect 279240 320894 279292 320900
rect 279528 314022 279556 335446
rect 279620 326466 279648 335566
rect 279608 326460 279660 326466
rect 279608 326402 279660 326408
rect 279712 326346 279740 336942
rect 279804 335510 279832 340068
rect 279896 337142 279924 340068
rect 280080 337278 280108 340068
rect 280068 337272 280120 337278
rect 280068 337214 280120 337220
rect 279884 337136 279936 337142
rect 279884 337078 279936 337084
rect 280068 337068 280120 337074
rect 280068 337010 280120 337016
rect 279884 336932 279936 336938
rect 279884 336874 279936 336880
rect 279792 335504 279844 335510
rect 279792 335446 279844 335452
rect 279896 330154 279924 336874
rect 279976 336796 280028 336802
rect 279976 336738 280028 336744
rect 279620 326318 279740 326346
rect 279804 330126 279924 330154
rect 279516 314016 279568 314022
rect 279516 313958 279568 313964
rect 279620 286346 279648 326318
rect 279700 326256 279752 326262
rect 279700 326198 279752 326204
rect 279608 286340 279660 286346
rect 279608 286282 279660 286288
rect 279712 284986 279740 326198
rect 279804 315382 279832 330126
rect 279884 330064 279936 330070
rect 279884 330006 279936 330012
rect 279792 315376 279844 315382
rect 279792 315318 279844 315324
rect 279700 284980 279752 284986
rect 279700 284922 279752 284928
rect 278872 283620 278924 283626
rect 278872 283562 278924 283568
rect 279792 8084 279844 8090
rect 279792 8026 279844 8032
rect 279804 3369 279832 8026
rect 279896 3641 279924 330006
rect 279988 8090 280016 336738
rect 279976 8084 280028 8090
rect 279976 8026 280028 8032
rect 280080 7970 280108 337010
rect 280172 336802 280200 340068
rect 280160 336796 280212 336802
rect 280160 336738 280212 336744
rect 280160 336660 280212 336666
rect 280160 336602 280212 336608
rect 280172 335374 280200 336602
rect 280160 335368 280212 335374
rect 280160 335310 280212 335316
rect 280160 335232 280212 335238
rect 280160 335174 280212 335180
rect 280172 329322 280200 335174
rect 280160 329316 280212 329322
rect 280160 329258 280212 329264
rect 280264 282198 280292 340068
rect 280448 337074 280476 340068
rect 280436 337068 280488 337074
rect 280436 337010 280488 337016
rect 280344 337000 280396 337006
rect 280344 336942 280396 336948
rect 280356 326398 280384 336942
rect 280540 336802 280568 340068
rect 280632 336938 280660 340068
rect 280712 337544 280764 337550
rect 280712 337486 280764 337492
rect 280620 336932 280672 336938
rect 280620 336874 280672 336880
rect 280436 336796 280488 336802
rect 280436 336738 280488 336744
rect 280528 336796 280580 336802
rect 280528 336738 280580 336744
rect 280448 335458 280476 336738
rect 280724 336666 280752 337486
rect 280816 337142 280844 340068
rect 280804 337136 280856 337142
rect 280804 337078 280856 337084
rect 280908 337006 280936 340068
rect 280896 337000 280948 337006
rect 280896 336942 280948 336948
rect 281000 336802 281028 340068
rect 281184 337618 281212 340068
rect 281172 337612 281224 337618
rect 281172 337554 281224 337560
rect 281172 336932 281224 336938
rect 281172 336874 281224 336880
rect 280804 336796 280856 336802
rect 280804 336738 280856 336744
rect 280988 336796 281040 336802
rect 280988 336738 281040 336744
rect 280712 336660 280764 336666
rect 280712 336602 280764 336608
rect 280816 336546 280844 336738
rect 280896 336728 280948 336734
rect 280896 336670 280948 336676
rect 280724 336518 280844 336546
rect 280448 335430 280660 335458
rect 280528 335368 280580 335374
rect 280528 335310 280580 335316
rect 280436 335300 280488 335306
rect 280436 335242 280488 335248
rect 280448 326602 280476 335242
rect 280436 326596 280488 326602
rect 280436 326538 280488 326544
rect 280344 326392 280396 326398
rect 280344 326334 280396 326340
rect 280540 326210 280568 335310
rect 280632 326346 280660 335430
rect 280724 326482 280752 336518
rect 280724 326454 280844 326482
rect 280632 326318 280752 326346
rect 280540 326182 280660 326210
rect 280632 316810 280660 326182
rect 280724 319530 280752 326318
rect 280712 319524 280764 319530
rect 280712 319466 280764 319472
rect 280620 316804 280672 316810
rect 280620 316746 280672 316752
rect 280252 282192 280304 282198
rect 280252 282134 280304 282140
rect 280250 76120 280306 76129
rect 280250 76055 280252 76064
rect 280304 76055 280306 76064
rect 280252 76026 280304 76032
rect 279988 7942 280108 7970
rect 279882 3632 279938 3641
rect 279882 3567 279938 3576
rect 279988 3505 280016 7942
rect 280816 7614 280844 326454
rect 280908 312662 280936 336670
rect 280988 326392 281040 326398
rect 280988 326334 281040 326340
rect 281080 326392 281132 326398
rect 281080 326334 281132 326340
rect 280896 312656 280948 312662
rect 280896 312598 280948 312604
rect 281000 309874 281028 326334
rect 280988 309868 281040 309874
rect 280988 309810 281040 309816
rect 281092 308514 281120 326334
rect 281184 326210 281212 336874
rect 281276 326398 281304 340068
rect 281264 326392 281316 326398
rect 281264 326334 281316 326340
rect 281184 326182 281304 326210
rect 281080 308508 281132 308514
rect 281080 308450 281132 308456
rect 281276 280838 281304 326182
rect 281264 280832 281316 280838
rect 281264 280774 281316 280780
rect 281368 279478 281396 340068
rect 281552 337006 281580 340068
rect 281540 337000 281592 337006
rect 281540 336942 281592 336948
rect 281644 336802 281672 340068
rect 281448 336796 281500 336802
rect 281448 336738 281500 336744
rect 281632 336796 281684 336802
rect 281632 336738 281684 336744
rect 281356 279472 281408 279478
rect 281356 279414 281408 279420
rect 281460 134570 281488 336738
rect 281736 335730 281764 340068
rect 281920 337414 281948 340068
rect 281908 337408 281960 337414
rect 281908 337350 281960 337356
rect 281644 335702 281764 335730
rect 281644 335102 281672 335702
rect 282012 335594 282040 340068
rect 282104 336802 282132 340068
rect 282288 337278 282316 340068
rect 282276 337272 282328 337278
rect 282276 337214 282328 337220
rect 282092 336796 282144 336802
rect 282092 336738 282144 336744
rect 281736 335566 282040 335594
rect 281632 335096 281684 335102
rect 281632 335038 281684 335044
rect 281736 318170 281764 335566
rect 282380 335458 282408 340068
rect 281828 335430 282408 335458
rect 281828 323678 281856 335430
rect 282472 335322 282500 340068
rect 282656 337890 282684 340068
rect 282644 337884 282696 337890
rect 282644 337826 282696 337832
rect 282552 337204 282604 337210
rect 282552 337146 282604 337152
rect 281920 335294 282500 335322
rect 281816 323672 281868 323678
rect 281816 323614 281868 323620
rect 281724 318164 281776 318170
rect 281724 318106 281776 318112
rect 281540 318096 281592 318102
rect 281540 318038 281592 318044
rect 281448 134564 281500 134570
rect 281448 134506 281500 134512
rect 280804 7608 280856 7614
rect 280804 7550 280856 7556
rect 280068 5160 280120 5166
rect 280068 5102 280120 5108
rect 279974 3496 280030 3505
rect 279974 3431 280030 3440
rect 279790 3360 279846 3369
rect 279790 3295 279846 3304
rect 278792 598 278912 626
rect 278884 480 278912 598
rect 280080 480 280108 5102
rect 281264 5092 281316 5098
rect 281264 5034 281316 5040
rect 281276 480 281304 5034
rect 281552 610 281580 318038
rect 281920 278050 281948 335294
rect 282564 335186 282592 337146
rect 282644 336796 282696 336802
rect 282644 336738 282696 336744
rect 282104 335158 282592 335186
rect 281908 278044 281960 278050
rect 281908 277986 281960 277992
rect 282104 276690 282132 335158
rect 282552 335096 282604 335102
rect 282552 335038 282604 335044
rect 282564 297498 282592 335038
rect 282552 297492 282604 297498
rect 282552 297434 282604 297440
rect 282656 291854 282684 336738
rect 282748 307086 282776 340068
rect 282840 337210 282868 340068
rect 283024 337822 283052 340068
rect 283012 337816 283064 337822
rect 283012 337758 283064 337764
rect 283012 337272 283064 337278
rect 283012 337214 283064 337220
rect 282828 337204 282880 337210
rect 282828 337146 282880 337152
rect 282920 337204 282972 337210
rect 282920 337146 282972 337152
rect 282828 336728 282880 336734
rect 282828 336670 282880 336676
rect 282840 327826 282868 336670
rect 282828 327820 282880 327826
rect 282828 327762 282880 327768
rect 282736 307080 282788 307086
rect 282736 307022 282788 307028
rect 282932 305658 282960 337146
rect 283024 328545 283052 337214
rect 283116 333282 283144 340068
rect 283208 337006 283236 340068
rect 283196 337000 283248 337006
rect 283196 336942 283248 336948
rect 283288 336728 283340 336734
rect 283288 336670 283340 336676
rect 283116 333254 283236 333282
rect 283208 331158 283236 333254
rect 283196 331152 283248 331158
rect 283196 331094 283248 331100
rect 283010 328536 283066 328545
rect 283010 328471 283066 328480
rect 283300 328030 283328 336670
rect 283392 333334 283420 340068
rect 283484 337210 283512 340068
rect 283576 337958 283604 340068
rect 283564 337952 283616 337958
rect 283564 337894 283616 337900
rect 283564 337680 283616 337686
rect 283564 337622 283616 337628
rect 283472 337204 283524 337210
rect 283472 337146 283524 337152
rect 283472 337068 283524 337074
rect 283472 337010 283524 337016
rect 283380 333328 283432 333334
rect 283380 333270 283432 333276
rect 283378 328400 283434 328409
rect 283378 328335 283434 328344
rect 283288 328024 283340 328030
rect 283288 327966 283340 327972
rect 283392 318850 283420 328335
rect 283484 319598 283512 337010
rect 283472 319592 283524 319598
rect 283472 319534 283524 319540
rect 283012 318844 283064 318850
rect 283012 318786 283064 318792
rect 283380 318844 283432 318850
rect 283380 318786 283432 318792
rect 283024 309058 283052 318786
rect 283012 309052 283064 309058
rect 283012 308994 283064 309000
rect 282920 305652 282972 305658
rect 282920 305594 282972 305600
rect 282644 291848 282696 291854
rect 282644 291790 282696 291796
rect 282092 276684 282144 276690
rect 282092 276626 282144 276632
rect 283576 6934 283604 337622
rect 283760 337074 283788 340068
rect 283748 337068 283800 337074
rect 283748 337010 283800 337016
rect 283852 335594 283880 340068
rect 283944 335730 283972 340068
rect 284128 337090 284156 340068
rect 284220 337278 284248 340068
rect 284326 340054 284432 340082
rect 284208 337272 284260 337278
rect 284208 337214 284260 337220
rect 284300 337272 284352 337278
rect 284300 337214 284352 337220
rect 284312 337090 284340 337214
rect 284024 337068 284076 337074
rect 284128 337062 284340 337090
rect 284024 337010 284076 337016
rect 284036 336122 284064 337010
rect 284116 337000 284168 337006
rect 284116 336942 284168 336948
rect 284024 336116 284076 336122
rect 284024 336058 284076 336064
rect 283944 335702 284064 335730
rect 283852 335566 283972 335594
rect 283840 331152 283892 331158
rect 283840 331094 283892 331100
rect 283656 328568 283708 328574
rect 283656 328510 283708 328516
rect 283668 323626 283696 328510
rect 283668 323598 283788 323626
rect 283760 317422 283788 323598
rect 283748 317416 283800 317422
rect 283748 317358 283800 317364
rect 283852 316742 283880 331094
rect 283840 316736 283892 316742
rect 283840 316678 283892 316684
rect 283944 304298 283972 335566
rect 284036 333266 284064 335702
rect 284024 333260 284076 333266
rect 284024 333202 284076 333208
rect 283932 304292 283984 304298
rect 283932 304234 283984 304240
rect 283748 299600 283800 299606
rect 283748 299542 283800 299548
rect 283760 298110 283788 299542
rect 283748 298104 283800 298110
rect 283748 298046 283800 298052
rect 283840 288448 283892 288454
rect 283840 288390 283892 288396
rect 283852 280106 283880 288390
rect 283760 280078 283880 280106
rect 283760 272542 283788 280078
rect 284128 273970 284156 336942
rect 284300 336796 284352 336802
rect 284300 336738 284352 336744
rect 284312 315314 284340 336738
rect 284404 333282 284432 340054
rect 284496 337006 284524 340068
rect 284484 337000 284536 337006
rect 284484 336942 284536 336948
rect 284588 336802 284616 340068
rect 284576 336796 284628 336802
rect 284576 336738 284628 336744
rect 284680 333282 284708 340068
rect 284864 338026 284892 340068
rect 284852 338020 284904 338026
rect 284852 337962 284904 337968
rect 284956 335782 284984 340068
rect 284944 335776 284996 335782
rect 284944 335718 284996 335724
rect 285048 335594 285076 340068
rect 284404 333254 284524 333282
rect 284392 328908 284444 328914
rect 284392 328850 284444 328856
rect 284300 315308 284352 315314
rect 284300 315250 284352 315256
rect 284404 301510 284432 328850
rect 284392 301504 284444 301510
rect 284392 301446 284444 301452
rect 284392 289808 284444 289814
rect 284392 289750 284444 289756
rect 284404 279206 284432 289750
rect 284392 279200 284444 279206
rect 284392 279142 284444 279148
rect 284116 273964 284168 273970
rect 284116 273906 284168 273912
rect 283748 272536 283800 272542
rect 283748 272478 283800 272484
rect 284496 271182 284524 333254
rect 284588 333254 284708 333282
rect 284772 335566 285076 335594
rect 284588 328438 284616 333254
rect 284576 328432 284628 328438
rect 284576 328374 284628 328380
rect 284576 318844 284628 318850
rect 284576 318786 284628 318792
rect 284588 313970 284616 318786
rect 284588 313942 284708 313970
rect 284680 309126 284708 313942
rect 284668 309120 284720 309126
rect 284668 309062 284720 309068
rect 284668 302184 284720 302190
rect 284668 302126 284720 302132
rect 284680 289814 284708 302126
rect 284668 289808 284720 289814
rect 284668 289750 284720 289756
rect 284484 271176 284536 271182
rect 284484 271118 284536 271124
rect 284772 268394 284800 335566
rect 284944 333260 284996 333266
rect 284944 333202 284996 333208
rect 284852 324284 284904 324290
rect 284852 324226 284904 324232
rect 284760 268388 284812 268394
rect 284760 268330 284812 268336
rect 284864 267034 284892 324226
rect 284956 290494 284984 333202
rect 285232 331838 285260 340068
rect 285220 331832 285272 331838
rect 285220 331774 285272 331780
rect 285034 321736 285090 321745
rect 285034 321671 285090 321680
rect 285048 321473 285076 321671
rect 285034 321464 285090 321473
rect 285034 321399 285090 321408
rect 285324 300150 285352 340068
rect 285416 324290 285444 340068
rect 285496 337000 285548 337006
rect 285496 336942 285548 336948
rect 285508 334694 285536 336942
rect 285496 334688 285548 334694
rect 285496 334630 285548 334636
rect 285600 330614 285628 340068
rect 285692 336938 285720 340068
rect 285798 340054 285904 340082
rect 285680 336932 285732 336938
rect 285680 336874 285732 336880
rect 285876 332926 285904 340054
rect 285968 337958 285996 340068
rect 285956 337952 286008 337958
rect 285956 337894 286008 337900
rect 286060 337210 286088 340068
rect 286048 337204 286100 337210
rect 286048 337146 286100 337152
rect 285956 336864 286008 336870
rect 285956 336806 286008 336812
rect 285864 332920 285916 332926
rect 285864 332862 285916 332868
rect 285588 330608 285640 330614
rect 285588 330550 285640 330556
rect 285404 324284 285456 324290
rect 285404 324226 285456 324232
rect 285680 323604 285732 323610
rect 285680 323546 285732 323552
rect 285312 300144 285364 300150
rect 285312 300086 285364 300092
rect 284944 290488 284996 290494
rect 284944 290430 284996 290436
rect 284944 279200 284996 279206
rect 284944 279142 284996 279148
rect 284956 269822 284984 279142
rect 284944 269816 284996 269822
rect 284944 269758 284996 269764
rect 284852 267028 284904 267034
rect 284852 266970 284904 266976
rect 283564 6928 283616 6934
rect 283564 6870 283616 6876
rect 283656 5024 283708 5030
rect 283656 4966 283708 4972
rect 281540 604 281592 610
rect 281540 546 281592 552
rect 282460 604 282512 610
rect 282460 546 282512 552
rect 282472 480 282500 546
rect 283668 480 283696 4966
rect 284760 4956 284812 4962
rect 284760 4898 284812 4904
rect 284772 480 284800 4898
rect 285692 610 285720 323546
rect 285968 297430 285996 336806
rect 286048 336796 286100 336802
rect 286048 336738 286100 336744
rect 285956 297424 286008 297430
rect 285956 297366 286008 297372
rect 286060 289134 286088 336738
rect 286048 289128 286100 289134
rect 286048 289070 286100 289076
rect 286152 262886 286180 340068
rect 286336 337686 286364 340068
rect 286324 337680 286376 337686
rect 286324 337622 286376 337628
rect 286232 337000 286284 337006
rect 286232 336942 286284 336948
rect 286140 262880 286192 262886
rect 286140 262822 286192 262828
rect 286244 261526 286272 336942
rect 286324 336932 286376 336938
rect 286324 336874 286376 336880
rect 286336 320890 286364 336874
rect 286428 336870 286456 340068
rect 286416 336864 286468 336870
rect 286416 336806 286468 336812
rect 286520 336802 286548 340068
rect 286600 337680 286652 337686
rect 286600 337622 286652 337628
rect 286508 336796 286560 336802
rect 286508 336738 286560 336744
rect 286612 333266 286640 337622
rect 286704 336802 286732 340068
rect 286692 336796 286744 336802
rect 286692 336738 286744 336744
rect 286600 333260 286652 333266
rect 286600 333202 286652 333208
rect 286796 333010 286824 340068
rect 286888 337006 286916 340068
rect 286968 337204 287020 337210
rect 286968 337146 287020 337152
rect 286876 337000 286928 337006
rect 286876 336942 286928 336948
rect 286876 336796 286928 336802
rect 286876 336738 286928 336744
rect 286612 332982 286824 333010
rect 286324 320884 286376 320890
rect 286324 320826 286376 320832
rect 286612 312594 286640 332982
rect 286784 332920 286836 332926
rect 286784 332862 286836 332868
rect 286692 326392 286744 326398
rect 286692 326334 286744 326340
rect 286704 313954 286732 326334
rect 286692 313948 286744 313954
rect 286692 313890 286744 313896
rect 286600 312588 286652 312594
rect 286600 312530 286652 312536
rect 286796 265674 286824 332862
rect 286888 329118 286916 336738
rect 286876 329112 286928 329118
rect 286876 329054 286928 329060
rect 286980 326398 287008 337146
rect 287072 336054 287100 340068
rect 287060 336048 287112 336054
rect 287060 335990 287112 335996
rect 286968 326392 287020 326398
rect 286968 326334 287020 326340
rect 287164 322250 287192 340068
rect 287152 322244 287204 322250
rect 287152 322186 287204 322192
rect 286784 265668 286836 265674
rect 286784 265610 286836 265616
rect 286232 261520 286284 261526
rect 286232 261462 286284 261468
rect 287256 260166 287284 340068
rect 287440 337686 287468 340068
rect 287428 337680 287480 337686
rect 287428 337622 287480 337628
rect 287428 337204 287480 337210
rect 287428 337146 287480 337152
rect 287440 335594 287468 337146
rect 287532 336870 287560 340068
rect 287520 336864 287572 336870
rect 287520 336806 287572 336812
rect 287624 335714 287652 340068
rect 287704 336796 287756 336802
rect 287704 336738 287756 336744
rect 287612 335708 287664 335714
rect 287612 335650 287664 335656
rect 287440 335566 287652 335594
rect 287428 333192 287480 333198
rect 287428 333134 287480 333140
rect 287440 326330 287468 333134
rect 287428 326324 287480 326330
rect 287428 326266 287480 326272
rect 287520 321632 287572 321638
rect 287520 321574 287572 321580
rect 287244 260160 287296 260166
rect 287244 260102 287296 260108
rect 287532 257378 287560 321574
rect 287520 257372 287572 257378
rect 287520 257314 287572 257320
rect 287624 22778 287652 335566
rect 287716 321638 287744 336738
rect 287808 331906 287836 340068
rect 287796 331900 287848 331906
rect 287796 331842 287848 331848
rect 287704 321632 287756 321638
rect 287704 321574 287756 321580
rect 287900 309806 287928 340068
rect 287992 336802 288020 340068
rect 288072 336864 288124 336870
rect 288072 336806 288124 336812
rect 287980 336796 288032 336802
rect 287980 336738 288032 336744
rect 288084 335594 288112 336806
rect 287992 335566 288112 335594
rect 287992 319462 288020 335566
rect 288176 333198 288204 340068
rect 288164 333192 288216 333198
rect 288164 333134 288216 333140
rect 288268 333010 288296 340068
rect 288360 337210 288388 340068
rect 288348 337204 288400 337210
rect 288348 337146 288400 337152
rect 288544 337006 288572 340068
rect 288532 337000 288584 337006
rect 288532 336942 288584 336948
rect 288636 336938 288664 340068
rect 288742 340054 288848 340082
rect 288624 336932 288676 336938
rect 288624 336874 288676 336880
rect 288084 332982 288296 333010
rect 287980 319456 288032 319462
rect 287980 319398 288032 319404
rect 287888 309800 287940 309806
rect 287888 309742 287940 309748
rect 288084 296002 288112 332982
rect 288820 332058 288848 340054
rect 288912 336870 288940 340068
rect 288900 336864 288952 336870
rect 288900 336806 288952 336812
rect 289004 332194 289032 340068
rect 289096 336802 289124 340068
rect 289084 336796 289136 336802
rect 289084 336738 289136 336744
rect 289280 334626 289308 340068
rect 289268 334620 289320 334626
rect 289268 334562 289320 334568
rect 289004 332166 289308 332194
rect 288820 332030 289032 332058
rect 288440 330540 288492 330546
rect 288440 330482 288492 330488
rect 288164 327140 288216 327146
rect 288164 327082 288216 327088
rect 288176 317422 288204 327082
rect 288164 317416 288216 317422
rect 288164 317358 288216 317364
rect 288348 310752 288400 310758
rect 288346 310720 288348 310729
rect 288400 310720 288402 310729
rect 288346 310655 288402 310664
rect 288164 307828 288216 307834
rect 288164 307770 288216 307776
rect 288176 298110 288204 307770
rect 288164 298104 288216 298110
rect 288164 298046 288216 298052
rect 288072 295996 288124 296002
rect 288072 295938 288124 295944
rect 288164 288448 288216 288454
rect 288164 288390 288216 288396
rect 288176 284968 288204 288390
rect 288176 284940 288296 284968
rect 288268 278769 288296 284940
rect 288070 278760 288126 278769
rect 288070 278695 288126 278704
rect 288254 278760 288310 278769
rect 288254 278695 288310 278704
rect 288084 269142 288112 278695
rect 288072 269136 288124 269142
rect 288072 269078 288124 269084
rect 288164 269136 288216 269142
rect 288164 269078 288216 269084
rect 288176 258738 288204 269078
rect 288164 258732 288216 258738
rect 288164 258674 288216 258680
rect 287612 22772 287664 22778
rect 287612 22714 287664 22720
rect 288348 6928 288400 6934
rect 288348 6870 288400 6876
rect 287152 4888 287204 4894
rect 287152 4830 287204 4836
rect 285680 604 285732 610
rect 285680 546 285732 552
rect 285956 604 286008 610
rect 285956 546 286008 552
rect 285968 480 285996 546
rect 287164 480 287192 4830
rect 288360 480 288388 6870
rect 288452 610 288480 330482
rect 288900 326392 288952 326398
rect 288900 326334 288952 326340
rect 288912 313970 288940 326334
rect 289004 326210 289032 332030
rect 289176 331968 289228 331974
rect 289176 331910 289228 331916
rect 289188 326398 289216 331910
rect 289176 326392 289228 326398
rect 289176 326334 289228 326340
rect 289004 326182 289216 326210
rect 289188 316690 289216 326182
rect 289280 318102 289308 332166
rect 289268 318096 289320 318102
rect 289268 318038 289320 318044
rect 289188 316662 289308 316690
rect 288912 313942 289216 313970
rect 288992 311840 289044 311846
rect 288992 311782 289044 311788
rect 289004 293162 289032 311782
rect 289188 309126 289216 313942
rect 289280 311846 289308 316662
rect 289268 311840 289320 311846
rect 289268 311782 289320 311788
rect 289176 309120 289228 309126
rect 289176 309062 289228 309068
rect 289268 309120 289320 309126
rect 289268 309062 289320 309068
rect 289280 308258 289308 309062
rect 289372 308446 289400 340068
rect 289478 340054 289584 340082
rect 289452 336796 289504 336802
rect 289452 336738 289504 336744
rect 289360 308440 289412 308446
rect 289360 308382 289412 308388
rect 289280 308230 289400 308258
rect 289372 293282 289400 308230
rect 289464 296070 289492 336738
rect 289452 296064 289504 296070
rect 289452 296006 289504 296012
rect 289556 294710 289584 340054
rect 289648 330546 289676 340068
rect 289740 331974 289768 340068
rect 289832 336802 289860 340068
rect 290004 338088 290056 338094
rect 290004 338030 290056 338036
rect 289912 337340 289964 337346
rect 289912 337282 289964 337288
rect 289820 336796 289872 336802
rect 289820 336738 289872 336744
rect 289924 334762 289952 337282
rect 290016 336190 290044 338030
rect 290832 337680 290884 337686
rect 290832 337622 290884 337628
rect 290464 337068 290516 337074
rect 290464 337010 290516 337016
rect 290004 336184 290056 336190
rect 290004 336126 290056 336132
rect 289912 334756 289964 334762
rect 289912 334698 289964 334704
rect 289728 331968 289780 331974
rect 289728 331910 289780 331916
rect 289636 330540 289688 330546
rect 289636 330482 289688 330488
rect 289636 321768 289688 321774
rect 289636 321710 289688 321716
rect 289648 321473 289676 321710
rect 289634 321464 289690 321473
rect 289634 321399 289690 321408
rect 289544 294704 289596 294710
rect 289544 294646 289596 294652
rect 289360 293276 289412 293282
rect 289360 293218 289412 293224
rect 289004 293134 289400 293162
rect 289372 287706 289400 293134
rect 289360 287700 289412 287706
rect 289360 287642 289412 287648
rect 289728 76084 289780 76090
rect 289728 76026 289780 76032
rect 289740 75993 289768 76026
rect 289726 75984 289782 75993
rect 289726 75919 289782 75928
rect 290476 15910 290504 337010
rect 290740 337000 290792 337006
rect 290740 336942 290792 336948
rect 290556 336932 290608 336938
rect 290556 336874 290608 336880
rect 290568 294642 290596 336874
rect 290648 336864 290700 336870
rect 290648 336806 290700 336812
rect 290660 323610 290688 336806
rect 290752 324970 290780 336942
rect 290844 327758 290872 337622
rect 291844 337136 291896 337142
rect 291844 337078 291896 337084
rect 291108 336796 291160 336802
rect 291108 336738 291160 336744
rect 290832 327752 290884 327758
rect 290832 327694 290884 327700
rect 290740 324964 290792 324970
rect 290740 324906 290792 324912
rect 290648 323604 290700 323610
rect 290648 323546 290700 323552
rect 290556 294636 290608 294642
rect 290556 294578 290608 294584
rect 291120 256018 291148 336738
rect 291108 256012 291160 256018
rect 291108 255954 291160 255960
rect 290464 15904 290516 15910
rect 290464 15846 290516 15852
rect 291856 13122 291884 337078
rect 291948 111790 291976 401066
rect 297456 400920 297508 400926
rect 297456 400862 297508 400868
rect 294604 400852 294656 400858
rect 294604 400794 294656 400800
rect 293960 336660 294012 336666
rect 293960 336602 294012 336608
rect 292580 333736 292632 333742
rect 292580 333678 292632 333684
rect 291936 111784 291988 111790
rect 291936 111726 291988 111732
rect 291844 13116 291896 13122
rect 291844 13058 291896 13064
rect 291936 9308 291988 9314
rect 291936 9250 291988 9256
rect 290740 4820 290792 4826
rect 290740 4762 290792 4768
rect 288440 604 288492 610
rect 288440 546 288492 552
rect 289544 604 289596 610
rect 289544 546 289596 552
rect 289556 480 289584 546
rect 290752 480 290780 4762
rect 291948 480 291976 9250
rect 292592 610 292620 333678
rect 293972 626 294000 336602
rect 294616 64870 294644 400794
rect 294696 338020 294748 338026
rect 294696 337962 294748 337968
rect 294604 64864 294656 64870
rect 294604 64806 294656 64812
rect 294708 19990 294736 337962
rect 297364 337952 297416 337958
rect 297364 337894 297416 337900
rect 296720 336592 296772 336598
rect 296720 336534 296772 336540
rect 296626 310856 296682 310865
rect 296626 310791 296682 310800
rect 296640 310758 296668 310791
rect 296628 310752 296680 310758
rect 296628 310694 296680 310700
rect 294696 19984 294748 19990
rect 294696 19926 294748 19932
rect 295524 9240 295576 9246
rect 295524 9182 295576 9188
rect 292580 604 292632 610
rect 292580 546 292632 552
rect 293132 604 293184 610
rect 293972 598 294368 626
rect 293132 546 293184 552
rect 293144 480 293172 546
rect 294340 480 294368 598
rect 295536 480 295564 9182
rect 296732 4214 296760 336534
rect 296812 332376 296864 332382
rect 296812 332318 296864 332324
rect 296720 4208 296772 4214
rect 296720 4150 296772 4156
rect 296824 1442 296852 332318
rect 297376 18630 297404 337894
rect 297468 158710 297496 400862
rect 301596 400784 301648 400790
rect 301596 400726 301648 400732
rect 298836 399968 298888 399974
rect 298836 399910 298888 399916
rect 298744 337884 298796 337890
rect 298744 337826 298796 337832
rect 298008 321768 298060 321774
rect 298006 321736 298008 321745
rect 298060 321736 298062 321745
rect 298006 321671 298062 321680
rect 297456 158704 297508 158710
rect 297456 158646 297508 158652
rect 297364 18624 297416 18630
rect 297364 18566 297416 18572
rect 298756 14482 298784 337826
rect 298848 205630 298876 399910
rect 301504 337816 301556 337822
rect 301504 337758 301556 337764
rect 300860 335096 300912 335102
rect 300860 335038 300912 335044
rect 299480 328092 299532 328098
rect 299480 328034 299532 328040
rect 298836 205624 298888 205630
rect 298836 205566 298888 205572
rect 298744 14476 298796 14482
rect 298744 14418 298796 14424
rect 299112 9172 299164 9178
rect 299112 9114 299164 9120
rect 297916 4208 297968 4214
rect 297916 4150 297968 4156
rect 296732 1414 296852 1442
rect 296732 480 296760 1414
rect 297928 480 297956 4150
rect 299124 480 299152 9114
rect 299492 610 299520 328034
rect 299570 310856 299626 310865
rect 299570 310791 299572 310800
rect 299624 310791 299626 310800
rect 299572 310762 299624 310768
rect 300872 610 300900 335038
rect 301516 11762 301544 337758
rect 301608 252550 301636 400726
rect 308404 400512 308456 400518
rect 308404 400454 308456 400460
rect 304264 400444 304316 400450
rect 304264 400386 304316 400392
rect 302976 399900 303028 399906
rect 302976 399842 303028 399848
rect 302884 337748 302936 337754
rect 302884 337690 302936 337696
rect 301596 252544 301648 252550
rect 301596 252486 301648 252492
rect 302146 227896 302202 227905
rect 302146 227831 302148 227840
rect 302200 227831 302202 227840
rect 302148 227802 302200 227808
rect 302146 76120 302202 76129
rect 302146 76055 302148 76064
rect 302200 76055 302202 76064
rect 302148 76026 302200 76032
rect 302146 29200 302202 29209
rect 302146 29135 302148 29144
rect 302200 29135 302202 29144
rect 302148 29106 302200 29112
rect 301504 11756 301556 11762
rect 301504 11698 301556 11704
rect 302896 8974 302924 337690
rect 302988 299470 303016 399842
rect 303620 329520 303672 329526
rect 303620 329462 303672 329468
rect 302976 299464 303028 299470
rect 302976 299406 303028 299412
rect 302608 8968 302660 8974
rect 302608 8910 302660 8916
rect 302884 8968 302936 8974
rect 302884 8910 302936 8916
rect 299480 604 299532 610
rect 299480 546 299532 552
rect 300308 604 300360 610
rect 300308 546 300360 552
rect 300860 604 300912 610
rect 300860 546 300912 552
rect 301412 604 301464 610
rect 301412 546 301464 552
rect 300320 480 300348 546
rect 301424 480 301452 546
rect 302620 480 302648 8910
rect 303632 610 303660 329462
rect 304276 41410 304304 400386
rect 305644 399696 305696 399702
rect 305644 399638 305696 399644
rect 305000 336524 305052 336530
rect 305000 336466 305052 336472
rect 304354 310856 304410 310865
rect 304354 310791 304356 310800
rect 304408 310791 304410 310800
rect 304356 310762 304408 310768
rect 304264 41404 304316 41410
rect 304264 41346 304316 41352
rect 303620 604 303672 610
rect 303620 546 303672 552
rect 303804 604 303856 610
rect 303804 546 303856 552
rect 303816 480 303844 546
rect 305012 480 305040 336466
rect 305656 88330 305684 399638
rect 307760 333668 307812 333674
rect 307760 333610 307812 333616
rect 306380 322516 306432 322522
rect 306380 322458 306432 322464
rect 305644 88324 305696 88330
rect 305644 88266 305696 88272
rect 306196 9104 306248 9110
rect 306196 9046 306248 9052
rect 306208 480 306236 9046
rect 306392 3482 306420 322458
rect 307772 3482 307800 333610
rect 308416 182170 308444 400454
rect 393964 398200 394016 398206
rect 393964 398142 394016 398148
rect 312542 340096 312598 340105
rect 312542 340031 312598 340040
rect 309782 338736 309838 338745
rect 309782 338671 309838 338680
rect 309046 322144 309102 322153
rect 309046 322079 309102 322088
rect 309060 321881 309088 322079
rect 309046 321872 309102 321881
rect 309046 321807 309102 321816
rect 309048 227860 309100 227866
rect 309048 227802 309100 227808
rect 309060 227769 309088 227802
rect 309046 227760 309102 227769
rect 309046 227695 309102 227704
rect 308404 182164 308456 182170
rect 308404 182106 308456 182112
rect 309796 124166 309824 338671
rect 311900 335028 311952 335034
rect 311900 334970 311952 334976
rect 310520 310004 310572 310010
rect 310520 309946 310572 309952
rect 309784 124160 309836 124166
rect 309784 124102 309836 124108
rect 309048 76084 309100 76090
rect 309048 76026 309100 76032
rect 309060 75993 309088 76026
rect 309046 75984 309102 75993
rect 309046 75919 309102 75928
rect 308956 29164 309008 29170
rect 308956 29106 309008 29112
rect 308968 29050 308996 29106
rect 309046 29064 309102 29073
rect 308968 29022 309046 29050
rect 309046 28999 309102 29008
rect 309784 9036 309836 9042
rect 309784 8978 309836 8984
rect 306392 3454 307432 3482
rect 307772 3454 308628 3482
rect 307404 480 307432 3454
rect 308600 480 308628 3454
rect 309796 480 309824 8978
rect 310532 3482 310560 309946
rect 311912 3482 311940 334970
rect 312556 218006 312584 340031
rect 315302 338872 315358 338881
rect 315302 338807 315358 338816
rect 314660 336456 314712 336462
rect 314660 336398 314712 336404
rect 313280 332308 313332 332314
rect 313280 332250 313332 332256
rect 312544 218000 312596 218006
rect 312544 217942 312596 217948
rect 313292 3482 313320 332250
rect 314568 7608 314620 7614
rect 314568 7550 314620 7556
rect 310532 3454 311020 3482
rect 311912 3454 312216 3482
rect 313292 3454 313412 3482
rect 310992 480 311020 3454
rect 312188 480 312216 3454
rect 313384 480 313412 3454
rect 314580 480 314608 7550
rect 314672 3482 314700 336398
rect 315316 264926 315344 338807
rect 320824 337680 320876 337686
rect 320824 337622 320876 337628
rect 316684 337612 316736 337618
rect 316684 337554 316736 337560
rect 316040 334960 316092 334966
rect 316040 334902 316092 334908
rect 315304 264920 315356 264926
rect 315304 264862 315356 264868
rect 316052 3618 316080 334902
rect 316696 4826 316724 337554
rect 319444 337544 319496 337550
rect 319444 337486 319496 337492
rect 318800 333600 318852 333606
rect 318800 333542 318852 333548
rect 317420 319728 317472 319734
rect 317420 319670 317472 319676
rect 316684 4820 316736 4826
rect 316684 4762 316736 4768
rect 316052 3590 317000 3618
rect 314672 3454 315804 3482
rect 315776 480 315804 3454
rect 316972 480 317000 3590
rect 317432 3482 317460 319670
rect 318812 3482 318840 333542
rect 319456 7614 319484 337486
rect 320180 330948 320232 330954
rect 320180 330890 320232 330896
rect 319444 7608 319496 7614
rect 319444 7550 319496 7556
rect 320192 3482 320220 330890
rect 320732 310820 320784 310826
rect 320732 310762 320784 310768
rect 320744 310729 320772 310762
rect 320730 310720 320786 310729
rect 320730 310655 320786 310664
rect 320836 21418 320864 337622
rect 346400 337476 346452 337482
rect 346400 337418 346452 337424
rect 327080 336388 327132 336394
rect 327080 336330 327132 336336
rect 322940 326732 322992 326738
rect 322940 326674 322992 326680
rect 321650 321872 321706 321881
rect 321650 321807 321706 321816
rect 321466 321736 321522 321745
rect 321664 321722 321692 321807
rect 321522 321694 321692 321722
rect 321466 321671 321522 321680
rect 321560 318300 321612 318306
rect 321560 318242 321612 318248
rect 321468 227928 321520 227934
rect 321466 227896 321468 227905
rect 321520 227896 321522 227905
rect 321466 227831 321522 227840
rect 321468 76152 321520 76158
rect 321466 76120 321468 76129
rect 321520 76120 321522 76129
rect 321466 76055 321522 76064
rect 321468 29232 321520 29238
rect 321466 29200 321468 29209
rect 321520 29200 321522 29209
rect 321466 29135 321522 29144
rect 320824 21412 320876 21418
rect 320824 21354 320876 21360
rect 321572 3482 321600 318242
rect 321652 29232 321704 29238
rect 321650 29200 321652 29209
rect 321704 29200 321706 29209
rect 321650 29135 321706 29144
rect 322848 5568 322900 5574
rect 322848 5510 322900 5516
rect 317432 3454 318104 3482
rect 318812 3454 319300 3482
rect 320192 3454 320496 3482
rect 321572 3454 321692 3482
rect 318076 480 318104 3454
rect 319272 480 319300 3454
rect 320468 480 320496 3454
rect 321664 480 321692 3454
rect 322860 480 322888 5510
rect 322952 3482 322980 326674
rect 324320 293344 324372 293350
rect 324320 293286 324372 293292
rect 323032 227928 323084 227934
rect 323030 227896 323032 227905
rect 323084 227896 323086 227905
rect 323030 227831 323086 227840
rect 323032 76152 323084 76158
rect 323030 76120 323032 76129
rect 323084 76120 323086 76129
rect 323030 76055 323086 76064
rect 324332 3482 324360 293286
rect 326436 5636 326488 5642
rect 326436 5578 326488 5584
rect 322952 3454 324084 3482
rect 324332 3454 325280 3482
rect 324056 480 324084 3454
rect 325252 480 325280 3454
rect 326448 480 326476 5578
rect 327092 3482 327120 336330
rect 333980 334892 334032 334898
rect 333980 334834 334032 334840
rect 331220 332240 331272 332246
rect 331220 332182 331272 332188
rect 328460 330880 328512 330886
rect 328460 330822 328512 330828
rect 328366 310856 328422 310865
rect 328366 310791 328368 310800
rect 328420 310791 328422 310800
rect 328368 310762 328420 310768
rect 328472 3482 328500 330822
rect 330024 5704 330076 5710
rect 330024 5646 330076 5652
rect 327092 3454 327672 3482
rect 328472 3454 328868 3482
rect 327644 480 327672 3454
rect 328840 480 328868 3454
rect 330036 480 330064 5646
rect 331232 480 331260 332182
rect 331312 325236 331364 325242
rect 331312 325178 331364 325184
rect 331324 3482 331352 325178
rect 333612 5772 333664 5778
rect 333612 5714 333664 5720
rect 331324 3454 332456 3482
rect 332428 480 332456 3454
rect 333624 480 333652 5714
rect 333992 3482 334020 334834
rect 342260 333532 342312 333538
rect 342260 333474 342312 333480
rect 338120 329452 338172 329458
rect 338120 329394 338172 329400
rect 335360 322448 335412 322454
rect 335360 322390 335412 322396
rect 335372 3482 335400 322390
rect 337108 5840 337160 5846
rect 337108 5782 337160 5788
rect 333992 3454 334756 3482
rect 335372 3454 335952 3482
rect 334728 480 334756 3454
rect 335924 480 335952 3454
rect 337120 480 337148 5782
rect 338132 3482 338160 329394
rect 340970 321872 341026 321881
rect 340970 321807 341026 321816
rect 340786 321736 340842 321745
rect 340984 321722 341012 321807
rect 340842 321694 341012 321722
rect 340786 321671 340842 321680
rect 340788 310752 340840 310758
rect 340786 310720 340788 310729
rect 340840 310720 340842 310729
rect 340786 310655 340842 310664
rect 339500 308576 339552 308582
rect 339500 308518 339552 308524
rect 338132 3454 338344 3482
rect 338316 480 338344 3454
rect 339512 480 339540 308518
rect 340880 10056 340932 10062
rect 340880 9998 340932 10004
rect 340696 5908 340748 5914
rect 340696 5850 340748 5856
rect 340708 480 340736 5850
rect 340892 3482 340920 9998
rect 342272 3482 342300 333474
rect 345020 10124 345072 10130
rect 345020 10066 345072 10072
rect 344284 5976 344336 5982
rect 344284 5918 344336 5924
rect 340892 3454 341932 3482
rect 342272 3454 343128 3482
rect 341904 480 341932 3454
rect 343100 480 343128 3454
rect 344296 480 344324 5918
rect 345032 3482 345060 10066
rect 346412 3482 346440 337418
rect 353300 336320 353352 336326
rect 353300 336262 353352 336268
rect 349160 323876 349212 323882
rect 349160 323818 349212 323824
rect 347686 310856 347742 310865
rect 347686 310791 347742 310800
rect 347700 310758 347728 310791
rect 347688 310752 347740 310758
rect 347688 310694 347740 310700
rect 347780 10192 347832 10198
rect 347780 10134 347832 10140
rect 347792 4214 347820 10134
rect 347872 6044 347924 6050
rect 347872 5986 347924 5992
rect 347780 4208 347832 4214
rect 347780 4150 347832 4156
rect 345032 3454 345520 3482
rect 346412 3454 346716 3482
rect 345492 480 345520 3454
rect 346688 480 346716 3454
rect 347884 480 347912 5986
rect 349068 4208 349120 4214
rect 349068 4150 349120 4156
rect 349080 480 349108 4150
rect 349172 3482 349200 323818
rect 351920 10260 351972 10266
rect 351920 10202 351972 10208
rect 351368 6112 351420 6118
rect 351368 6054 351420 6060
rect 349172 3454 350304 3482
rect 350276 480 350304 3454
rect 351380 480 351408 6054
rect 351932 3482 351960 10202
rect 351932 3454 352604 3482
rect 352576 480 352604 3454
rect 353312 1306 353340 336262
rect 356060 332172 356112 332178
rect 356060 332114 356112 332120
rect 354956 6860 355008 6866
rect 354956 6802 355008 6808
rect 353312 1278 353800 1306
rect 353772 480 353800 1278
rect 354968 480 354996 6802
rect 356072 4214 356100 332114
rect 382280 330812 382332 330818
rect 382280 330754 382332 330760
rect 367100 329384 367152 329390
rect 367100 329326 367152 329332
rect 360200 326664 360252 326670
rect 360200 326606 360252 326612
rect 359648 310820 359700 310826
rect 359648 310762 359700 310768
rect 359660 310729 359688 310762
rect 359646 310720 359702 310729
rect 359646 310655 359702 310664
rect 356152 11008 356204 11014
rect 356152 10950 356204 10956
rect 356060 4208 356112 4214
rect 356060 4150 356112 4156
rect 356164 480 356192 10950
rect 358820 10940 358872 10946
rect 358820 10882 358872 10888
rect 358544 6792 358596 6798
rect 358544 6734 358596 6740
rect 357348 4208 357400 4214
rect 357348 4150 357400 4156
rect 357360 480 357388 4150
rect 358556 480 358584 6734
rect 358832 3482 358860 10882
rect 360212 3482 360240 326606
rect 362222 322144 362278 322153
rect 362222 322079 362278 322088
rect 362236 321881 362264 322079
rect 362222 321872 362278 321881
rect 362222 321807 362278 321816
rect 364340 316940 364392 316946
rect 364340 316882 364392 316888
rect 362960 10872 363012 10878
rect 362960 10814 363012 10820
rect 362132 6724 362184 6730
rect 362132 6666 362184 6672
rect 358832 3454 359780 3482
rect 360212 3454 360976 3482
rect 359752 480 359780 3454
rect 360948 480 360976 3454
rect 362144 480 362172 6666
rect 362972 3482 363000 10814
rect 364352 3482 364380 316882
rect 367006 310856 367062 310865
rect 367006 310791 367008 310800
rect 367060 310791 367062 310800
rect 367008 310762 367060 310768
rect 365720 10804 365772 10810
rect 365720 10746 365772 10752
rect 365732 4214 365760 10746
rect 365812 6656 365864 6662
rect 365812 6598 365864 6604
rect 365720 4208 365772 4214
rect 365720 4150 365772 4156
rect 362972 3454 363368 3482
rect 364352 3454 364564 3482
rect 363340 480 363368 3454
rect 364536 480 364564 3454
rect 365824 3346 365852 6598
rect 366916 4208 366968 4214
rect 366916 4150 366968 4156
rect 365732 3318 365852 3346
rect 365732 480 365760 3318
rect 366928 480 366956 4150
rect 367112 3482 367140 329326
rect 379428 321768 379480 321774
rect 379426 321736 379428 321745
rect 379480 321736 379482 321745
rect 379426 321671 379482 321680
rect 371240 319660 371292 319666
rect 371240 319602 371292 319608
rect 369860 10736 369912 10742
rect 369860 10678 369912 10684
rect 369216 6588 369268 6594
rect 369216 6530 369268 6536
rect 367112 3454 368060 3482
rect 368032 480 368060 3454
rect 369228 480 369256 6530
rect 369872 3482 369900 10678
rect 371252 3482 371280 319602
rect 374000 315512 374052 315518
rect 374000 315454 374052 315460
rect 372804 6520 372856 6526
rect 372804 6462 372856 6468
rect 369872 3454 370452 3482
rect 371252 3454 371648 3482
rect 370424 480 370452 3454
rect 371620 480 371648 3454
rect 372816 480 372844 6462
rect 374012 4214 374040 315454
rect 379428 310752 379480 310758
rect 379426 310720 379428 310729
rect 379480 310720 379482 310729
rect 379426 310655 379482 310664
rect 378140 309936 378192 309942
rect 378140 309878 378192 309884
rect 374092 10668 374144 10674
rect 374092 10610 374144 10616
rect 374000 4208 374052 4214
rect 374000 4150 374052 4156
rect 374104 1442 374132 10610
rect 376760 10600 376812 10606
rect 376760 10542 376812 10548
rect 376392 6452 376444 6458
rect 376392 6394 376444 6400
rect 375196 4208 375248 4214
rect 375196 4150 375248 4156
rect 374012 1414 374132 1442
rect 374012 480 374040 1414
rect 375208 480 375236 4150
rect 376404 480 376432 6394
rect 376772 3482 376800 10542
rect 378152 3482 378180 309878
rect 380900 10532 380952 10538
rect 380900 10474 380952 10480
rect 379980 6384 380032 6390
rect 379980 6326 380032 6332
rect 376772 3454 377628 3482
rect 378152 3454 378824 3482
rect 377600 480 377628 3454
rect 378796 480 378824 3454
rect 379992 480 380020 6326
rect 380912 3482 380940 10474
rect 382292 3482 382320 330754
rect 393320 329316 393372 329322
rect 393320 329258 393372 329264
rect 385040 322380 385092 322386
rect 385040 322322 385092 322328
rect 383660 10464 383712 10470
rect 383660 10406 383712 10412
rect 383568 6316 383620 6322
rect 383568 6258 383620 6264
rect 380912 3454 381216 3482
rect 382292 3454 382412 3482
rect 381188 480 381216 3454
rect 382384 480 382412 3454
rect 383580 480 383608 6258
rect 383672 3482 383700 10406
rect 385052 3482 385080 322322
rect 386326 321872 386382 321881
rect 386326 321807 386382 321816
rect 386340 321774 386368 321807
rect 386328 321768 386380 321774
rect 386328 321710 386380 321716
rect 389180 314152 389232 314158
rect 389180 314094 389232 314100
rect 386326 310856 386382 310865
rect 386326 310791 386382 310800
rect 386340 310758 386368 310791
rect 386328 310752 386380 310758
rect 386328 310694 386380 310700
rect 387800 10396 387852 10402
rect 387800 10338 387852 10344
rect 387064 6248 387116 6254
rect 387064 6190 387116 6196
rect 383672 3454 384712 3482
rect 385052 3454 385908 3482
rect 384684 480 384712 3454
rect 385880 480 385908 3454
rect 387076 480 387104 6190
rect 387812 3482 387840 10338
rect 389192 3482 389220 314094
rect 390560 10328 390612 10334
rect 390560 10270 390612 10276
rect 387812 3454 388300 3482
rect 389192 3454 389496 3482
rect 388272 480 388300 3454
rect 389468 480 389496 3454
rect 390572 2854 390600 10270
rect 390652 6180 390704 6186
rect 390652 6122 390704 6128
rect 390560 2848 390612 2854
rect 390560 2790 390612 2796
rect 390664 480 390692 6122
rect 393332 3482 393360 329258
rect 393976 276010 394004 398142
rect 440240 336252 440292 336258
rect 440240 336194 440292 336200
rect 422300 334824 422352 334830
rect 422300 334766 422352 334772
rect 404360 333464 404412 333470
rect 404360 333406 404412 333412
rect 397460 332104 397512 332110
rect 397460 332046 397512 332052
rect 394700 325168 394752 325174
rect 394700 325110 394752 325116
rect 393964 276004 394016 276010
rect 393964 275946 394016 275952
rect 394712 3482 394740 325110
rect 397472 3482 397500 332046
rect 400312 328024 400364 328030
rect 400312 327966 400364 327972
rect 398840 323808 398892 323814
rect 398840 323750 398892 323756
rect 398748 310752 398800 310758
rect 398746 310720 398748 310729
rect 398800 310720 398802 310729
rect 398746 310655 398802 310664
rect 398852 3482 398880 323750
rect 400324 3482 400352 327966
rect 400862 322144 400918 322153
rect 400862 322079 400918 322088
rect 400876 321881 400904 322079
rect 400862 321872 400918 321881
rect 400862 321807 400918 321816
rect 401600 311228 401652 311234
rect 401600 311170 401652 311176
rect 401612 3482 401640 311170
rect 404372 3482 404400 333406
rect 411260 330744 411312 330750
rect 411260 330686 411312 330692
rect 408500 326596 408552 326602
rect 408500 326538 408552 326544
rect 405740 316872 405792 316878
rect 405740 316814 405792 316820
rect 405646 310856 405702 310865
rect 405646 310791 405702 310800
rect 405660 310758 405688 310791
rect 405648 310752 405700 310758
rect 405648 310694 405700 310700
rect 405752 3482 405780 316814
rect 393332 3454 394280 3482
rect 394712 3454 395476 3482
rect 397472 3454 397868 3482
rect 398852 3454 399064 3482
rect 400324 3454 401364 3482
rect 401612 3454 402560 3482
rect 404372 3454 404952 3482
rect 405752 3454 406148 3482
rect 391848 2848 391900 2854
rect 391848 2790 391900 2796
rect 393044 2848 393096 2854
rect 393044 2790 393096 2796
rect 391860 480 391888 2790
rect 393056 480 393084 2790
rect 394252 480 394280 3454
rect 395448 480 395476 3454
rect 396632 2916 396684 2922
rect 396632 2858 396684 2864
rect 396644 480 396672 2858
rect 397840 480 397868 3454
rect 399036 480 399064 3454
rect 400220 2984 400272 2990
rect 400220 2926 400272 2932
rect 400232 480 400260 2926
rect 401336 480 401364 3454
rect 402532 480 402560 3454
rect 403716 3052 403768 3058
rect 403716 2994 403768 3000
rect 403728 480 403756 2994
rect 404924 480 404952 3454
rect 406120 480 406148 3454
rect 407304 3120 407356 3126
rect 407304 3062 407356 3068
rect 407316 480 407344 3062
rect 408512 480 408540 326538
rect 408592 315444 408644 315450
rect 408592 315386 408644 315392
rect 408604 3482 408632 315386
rect 411272 3482 411300 330686
rect 415400 329248 415452 329254
rect 415400 329190 415452 329196
rect 412640 307216 412692 307222
rect 412640 307158 412692 307164
rect 412652 3482 412680 307158
rect 415306 227896 415362 227905
rect 415306 227831 415362 227840
rect 415320 227769 415348 227831
rect 415306 227760 415362 227769
rect 415306 227695 415362 227704
rect 415306 76120 415362 76129
rect 415306 76055 415362 76064
rect 415320 75993 415348 76055
rect 415306 75984 415362 75993
rect 415306 75919 415362 75928
rect 415122 29200 415178 29209
rect 415122 29135 415178 29144
rect 415136 29050 415164 29135
rect 415306 29064 415362 29073
rect 415136 29022 415306 29050
rect 415306 28999 415362 29008
rect 415412 3482 415440 329190
rect 418250 321872 418306 321881
rect 418250 321807 418306 321816
rect 418066 321736 418122 321745
rect 418264 321722 418292 321807
rect 418122 321694 418292 321722
rect 418066 321671 418122 321680
rect 418160 321088 418212 321094
rect 418160 321030 418212 321036
rect 418068 310752 418120 310758
rect 418066 310720 418068 310729
rect 418120 310720 418122 310729
rect 418066 310655 418122 310664
rect 416872 305720 416924 305726
rect 416872 305662 416924 305668
rect 408604 3454 409736 3482
rect 411272 3454 412128 3482
rect 412652 3454 413324 3482
rect 415412 3454 415716 3482
rect 409708 480 409736 3454
rect 410892 3188 410944 3194
rect 410892 3130 410944 3136
rect 410904 480 410932 3130
rect 412100 480 412128 3454
rect 413296 480 413324 3454
rect 414480 3256 414532 3262
rect 414480 3198 414532 3204
rect 414492 480 414520 3198
rect 415688 480 415716 3454
rect 416884 480 416912 305662
rect 418172 3482 418200 321030
rect 419540 291916 419592 291922
rect 419540 291858 419592 291864
rect 419552 3482 419580 291858
rect 422312 3482 422340 334766
rect 433340 332036 433392 332042
rect 433340 331978 433392 331984
rect 425152 327956 425204 327962
rect 425152 327898 425204 327904
rect 423680 314084 423732 314090
rect 423680 314026 423732 314032
rect 423692 3482 423720 314026
rect 424966 310856 425022 310865
rect 424966 310791 425022 310800
rect 424980 310758 425008 310791
rect 424968 310752 425020 310758
rect 424968 310694 425020 310700
rect 425060 4140 425112 4146
rect 425060 4082 425112 4088
rect 418172 3454 419212 3482
rect 419552 3454 420408 3482
rect 422312 3454 422800 3482
rect 423692 3454 423996 3482
rect 417976 3324 418028 3330
rect 417976 3266 418028 3272
rect 417988 480 418016 3266
rect 419184 480 419212 3454
rect 420380 480 420408 3454
rect 421564 3392 421616 3398
rect 421564 3334 421616 3340
rect 421576 480 421604 3334
rect 422772 480 422800 3454
rect 423968 480 423996 3454
rect 425072 2802 425100 4082
rect 425164 2922 425192 327898
rect 429200 325100 429252 325106
rect 429200 325042 429252 325048
rect 426440 304360 426492 304366
rect 426440 304302 426492 304308
rect 426452 3482 426480 304302
rect 428740 4072 428792 4078
rect 428740 4014 428792 4020
rect 426452 3454 427584 3482
rect 425152 2916 425204 2922
rect 425152 2858 425204 2864
rect 426348 2916 426400 2922
rect 426348 2858 426400 2864
rect 425072 2774 425192 2802
rect 425164 480 425192 2774
rect 426360 480 426388 2858
rect 427556 480 427584 3454
rect 428752 480 428780 4014
rect 429212 3482 429240 325042
rect 430580 290556 430632 290562
rect 430580 290498 430632 290504
rect 430592 3482 430620 290498
rect 432328 4004 432380 4010
rect 432328 3946 432380 3952
rect 429212 3454 429976 3482
rect 430592 3454 431172 3482
rect 429948 480 429976 3454
rect 431144 480 431172 3454
rect 432340 480 432368 3946
rect 433352 3482 433380 331978
rect 433432 326528 433484 326534
rect 433432 326470 433484 326476
rect 433444 3874 433472 326470
rect 436100 323740 436152 323746
rect 436100 323682 436152 323688
rect 435824 3936 435876 3942
rect 435824 3878 435876 3884
rect 433432 3868 433484 3874
rect 433432 3810 433484 3816
rect 434628 3868 434680 3874
rect 434628 3810 434680 3816
rect 433352 3454 433564 3482
rect 433536 480 433564 3454
rect 434640 480 434668 3810
rect 435836 480 435864 3878
rect 436112 3482 436140 323682
rect 437570 321872 437626 321881
rect 437570 321807 437626 321816
rect 437386 321736 437442 321745
rect 437584 321722 437612 321807
rect 437442 321694 437612 321722
rect 437386 321671 437442 321680
rect 437480 312724 437532 312730
rect 437480 312666 437532 312672
rect 437388 310752 437440 310758
rect 437386 310720 437388 310729
rect 437440 310720 437442 310729
rect 437386 310655 437442 310664
rect 437386 227896 437442 227905
rect 437386 227831 437388 227840
rect 437440 227831 437442 227840
rect 437388 227802 437440 227808
rect 437386 76120 437442 76129
rect 437386 76055 437388 76064
rect 437440 76055 437442 76064
rect 437388 76026 437440 76032
rect 437386 29200 437442 29209
rect 437386 29135 437388 29144
rect 437440 29135 437442 29144
rect 437388 29106 437440 29112
rect 437492 3482 437520 312666
rect 439412 4004 439464 4010
rect 439412 3946 439464 3952
rect 436112 3454 437060 3482
rect 437492 3454 438256 3482
rect 437032 480 437060 3454
rect 438228 480 438256 3454
rect 439424 480 439452 3946
rect 440252 3482 440280 336194
rect 483020 336184 483072 336190
rect 483020 336126 483072 336132
rect 465080 333396 465132 333402
rect 465080 333338 465132 333344
rect 451280 330676 451332 330682
rect 451280 330618 451332 330624
rect 443092 326460 443144 326466
rect 443092 326402 443144 326408
rect 441620 311160 441672 311166
rect 441620 311102 441672 311108
rect 441632 3482 441660 311102
rect 443000 3800 443052 3806
rect 443000 3742 443052 3748
rect 440252 3454 440648 3482
rect 441632 3454 441844 3482
rect 440620 480 440648 3454
rect 441816 480 441844 3454
rect 443012 480 443040 3742
rect 443104 3482 443132 326402
rect 447140 319592 447192 319598
rect 447140 319534 447192 319540
rect 444286 310856 444342 310865
rect 444286 310791 444342 310800
rect 444300 310758 444328 310791
rect 444288 310752 444340 310758
rect 444288 310694 444340 310700
rect 444380 303000 444432 303006
rect 444380 302942 444432 302948
rect 444288 227860 444340 227866
rect 444288 227802 444340 227808
rect 444300 227769 444328 227802
rect 444286 227760 444342 227769
rect 444286 227695 444342 227704
rect 444288 76084 444340 76090
rect 444288 76026 444340 76032
rect 444300 75993 444328 76026
rect 444286 75984 444342 75993
rect 444286 75919 444342 75928
rect 444196 29164 444248 29170
rect 444196 29106 444248 29112
rect 444208 29050 444236 29106
rect 444286 29064 444342 29073
rect 444208 29022 444286 29050
rect 444286 28999 444342 29008
rect 444392 3482 444420 302942
rect 446588 3732 446640 3738
rect 446588 3674 446640 3680
rect 443104 3454 444236 3482
rect 444392 3454 445432 3482
rect 444208 480 444236 3454
rect 445404 480 445432 3454
rect 446600 480 446628 3674
rect 447152 3482 447180 319534
rect 448520 301572 448572 301578
rect 448520 301514 448572 301520
rect 448532 3482 448560 301514
rect 450176 3664 450228 3670
rect 450176 3606 450228 3612
rect 447152 3454 447824 3482
rect 448532 3454 449020 3482
rect 447796 480 447824 3454
rect 448992 480 449020 3454
rect 450188 480 450216 3606
rect 451292 480 451320 330618
rect 462320 327888 462372 327894
rect 462320 327830 462372 327836
rect 458180 322312 458232 322318
rect 458180 322254 458232 322260
rect 456890 321872 456946 321881
rect 456890 321807 456946 321816
rect 456706 321736 456762 321745
rect 456904 321722 456932 321807
rect 456762 321694 456932 321722
rect 456706 321671 456762 321680
rect 454040 318232 454092 318238
rect 454040 318174 454092 318180
rect 451372 289196 451424 289202
rect 451372 289138 451424 289144
rect 451384 3482 451412 289138
rect 453672 3596 453724 3602
rect 453672 3538 453724 3544
rect 451384 3454 452516 3482
rect 452488 480 452516 3454
rect 453684 480 453712 3538
rect 454052 3482 454080 318174
rect 456708 310752 456760 310758
rect 456706 310720 456708 310729
rect 456760 310720 456762 310729
rect 456706 310655 456762 310664
rect 455420 300212 455472 300218
rect 455420 300154 455472 300160
rect 455432 3482 455460 300154
rect 456706 227896 456762 227905
rect 456890 227896 456946 227905
rect 456762 227854 456890 227882
rect 456706 227831 456762 227840
rect 456890 227831 456946 227840
rect 456706 76120 456762 76129
rect 456890 76120 456946 76129
rect 456762 76078 456890 76106
rect 456706 76055 456762 76064
rect 456890 76055 456946 76064
rect 456706 29200 456762 29209
rect 456890 29200 456946 29209
rect 456762 29158 456890 29186
rect 456706 29135 456762 29144
rect 456890 29135 456946 29144
rect 457260 3528 457312 3534
rect 454052 3454 454908 3482
rect 455432 3454 456104 3482
rect 457260 3470 457312 3476
rect 458192 3482 458220 322254
rect 460940 316804 460992 316810
rect 460940 316746 460992 316752
rect 459652 287768 459704 287774
rect 459652 287710 459704 287716
rect 454880 480 454908 3454
rect 456076 480 456104 3454
rect 457272 480 457300 3470
rect 458192 3454 458496 3482
rect 458468 480 458496 3454
rect 459664 480 459692 287710
rect 460952 3482 460980 316746
rect 462332 3482 462360 327830
rect 463606 310856 463662 310865
rect 463606 310791 463662 310800
rect 463620 310758 463648 310791
rect 463608 310752 463660 310758
rect 463608 310694 463660 310700
rect 464434 4040 464490 4049
rect 464434 3975 464490 3984
rect 460848 3460 460900 3466
rect 460952 3454 462084 3482
rect 462332 3454 463280 3482
rect 460848 3402 460900 3408
rect 460860 480 460888 3402
rect 462056 480 462084 3454
rect 463252 480 463280 3454
rect 464448 480 464476 3975
rect 465092 3482 465120 333338
rect 467840 329180 467892 329186
rect 467840 329122 467892 329128
rect 466460 321020 466512 321026
rect 466460 320962 466512 320968
rect 466472 3482 466500 320962
rect 467852 3534 467880 329122
rect 471980 325032 472032 325038
rect 471980 324974 472032 324980
rect 469220 298784 469272 298790
rect 469220 298726 469272 298732
rect 467930 3904 467986 3913
rect 467930 3839 467986 3848
rect 467840 3528 467892 3534
rect 465092 3454 465672 3482
rect 466472 3454 466868 3482
rect 467840 3470 467892 3476
rect 465644 480 465672 3454
rect 466840 480 466868 3454
rect 467944 480 467972 3839
rect 469128 3528 469180 3534
rect 469128 3470 469180 3476
rect 469232 3482 469260 298726
rect 471244 256012 471296 256018
rect 471244 255954 471296 255960
rect 469140 480 469168 3470
rect 469232 3454 470364 3482
rect 471256 3466 471284 255954
rect 471518 3768 471574 3777
rect 471518 3703 471574 3712
rect 470336 480 470364 3454
rect 471244 3460 471296 3466
rect 471244 3402 471296 3408
rect 471532 480 471560 3703
rect 471992 3346 472020 324974
rect 476210 321872 476266 321881
rect 476210 321807 476266 321816
rect 476026 321736 476082 321745
rect 476224 321722 476252 321807
rect 476082 321694 476252 321722
rect 476026 321671 476082 321680
rect 476120 320952 476172 320958
rect 476120 320894 476172 320900
rect 475568 310820 475620 310826
rect 475568 310762 475620 310768
rect 475580 310729 475608 310762
rect 475566 310720 475622 310729
rect 475566 310655 475622 310664
rect 473360 307148 473412 307154
rect 473360 307090 473412 307096
rect 473372 3346 473400 307090
rect 475384 294704 475436 294710
rect 475384 294646 475436 294652
rect 475106 3632 475162 3641
rect 475106 3567 475162 3576
rect 471992 3318 472756 3346
rect 473372 3318 473952 3346
rect 472728 480 472756 3318
rect 473924 480 473952 3318
rect 475120 480 475148 3567
rect 475396 3534 475424 294646
rect 476026 227896 476082 227905
rect 476026 227831 476028 227840
rect 476080 227831 476082 227840
rect 476028 227802 476080 227808
rect 475384 3528 475436 3534
rect 475384 3470 475436 3476
rect 476132 3346 476160 320894
rect 478880 315376 478932 315382
rect 478880 315318 478932 315324
rect 477500 286340 477552 286346
rect 477500 286282 477552 286288
rect 476132 3318 476344 3346
rect 476316 480 476344 3318
rect 477512 480 477540 286282
rect 478694 3496 478750 3505
rect 478694 3431 478750 3440
rect 478708 480 478736 3431
rect 478892 3346 478920 315318
rect 482926 310856 482982 310865
rect 482926 310791 482928 310800
rect 482980 310791 482982 310800
rect 482928 310762 482980 310768
rect 482284 296064 482336 296070
rect 482284 296006 482336 296012
rect 480260 284980 480312 284986
rect 480260 284922 480312 284928
rect 480272 3482 480300 284922
rect 482296 3602 482324 296006
rect 482928 227860 482980 227866
rect 482928 227802 482980 227808
rect 482940 227769 482968 227802
rect 482926 227760 482982 227769
rect 482926 227695 482982 227704
rect 482926 76120 482982 76129
rect 482926 76055 482982 76064
rect 482940 75993 482968 76055
rect 482926 75984 482982 75993
rect 482926 75919 482982 75928
rect 482284 3596 482336 3602
rect 482284 3538 482336 3544
rect 483032 3482 483060 336126
rect 484400 314016 484452 314022
rect 484400 313958 484452 313964
rect 484412 3482 484440 313958
rect 485056 171086 485084 401911
rect 489184 401872 489236 401878
rect 489184 401814 489236 401820
rect 489196 358766 489224 401814
rect 496084 400376 496136 400382
rect 496084 400318 496136 400324
rect 489184 358760 489236 358766
rect 489184 358702 489236 358708
rect 489184 337408 489236 337414
rect 489184 337350 489236 337356
rect 487160 319524 487212 319530
rect 487160 319466 487212 319472
rect 485780 283620 485832 283626
rect 485780 283562 485832 283568
rect 485044 171080 485096 171086
rect 485044 171022 485096 171028
rect 480272 3454 481128 3482
rect 483032 3454 483520 3482
rect 484412 3454 484624 3482
rect 478892 3318 479932 3346
rect 479904 480 479932 3318
rect 481100 480 481128 3454
rect 482282 3360 482338 3369
rect 482282 3295 482338 3304
rect 482296 480 482324 3295
rect 483492 480 483520 3454
rect 484596 480 484624 3454
rect 485792 480 485820 283562
rect 486976 4820 487028 4826
rect 486976 4762 487028 4768
rect 486988 480 487016 4762
rect 487172 3482 487200 319466
rect 488540 282192 488592 282198
rect 488540 282134 488592 282140
rect 488552 3618 488580 282134
rect 489196 4826 489224 337350
rect 495346 321872 495402 321881
rect 495530 321872 495586 321881
rect 495402 321830 495530 321858
rect 495346 321807 495402 321816
rect 495530 321807 495586 321816
rect 491300 312656 491352 312662
rect 491300 312598 491352 312604
rect 491206 29200 491262 29209
rect 491206 29135 491262 29144
rect 491220 28801 491248 29135
rect 491206 28792 491262 28801
rect 491206 28727 491262 28736
rect 490564 7608 490616 7614
rect 490564 7550 490616 7556
rect 489184 4820 489236 4826
rect 489184 4762 489236 4768
rect 488552 3590 489408 3618
rect 487172 3454 488212 3482
rect 488184 480 488212 3454
rect 489380 480 489408 3590
rect 490576 480 490604 7550
rect 491312 626 491340 312598
rect 495348 310752 495400 310758
rect 495346 310720 495348 310729
rect 495400 310720 495402 310729
rect 495346 310655 495402 310664
rect 494060 309868 494112 309874
rect 494060 309810 494112 309816
rect 492680 280832 492732 280838
rect 492680 280774 492732 280780
rect 491312 598 491800 626
rect 492692 610 492720 280774
rect 494072 3398 494100 309810
rect 496096 135250 496124 400318
rect 579804 393304 579856 393310
rect 579804 393246 579856 393252
rect 579816 393009 579844 393246
rect 579802 393000 579858 393009
rect 579802 392935 579858 392944
rect 580172 369844 580224 369850
rect 580172 369786 580224 369792
rect 580184 369617 580212 369786
rect 580170 369608 580226 369617
rect 580170 369543 580226 369552
rect 580080 358760 580132 358766
rect 580080 358702 580132 358708
rect 580092 357921 580120 358702
rect 580078 357912 580134 357921
rect 580078 357847 580134 357856
rect 579804 346384 579856 346390
rect 579804 346326 579856 346332
rect 579816 346089 579844 346326
rect 579802 346080 579858 346089
rect 579802 346015 579858 346024
rect 521660 336116 521712 336122
rect 521660 336058 521712 336064
rect 500960 334756 501012 334762
rect 500960 334698 501012 334704
rect 498200 308508 498252 308514
rect 498200 308450 498252 308456
rect 496084 135244 496136 135250
rect 496084 135186 496136 135192
rect 495440 134564 495492 134570
rect 495440 134506 495492 134512
rect 494152 8968 494204 8974
rect 494152 8910 494204 8916
rect 494060 3392 494112 3398
rect 494060 3334 494112 3340
rect 491772 480 491800 598
rect 492680 604 492732 610
rect 492680 546 492732 552
rect 492956 604 493008 610
rect 492956 546 493008 552
rect 492968 480 492996 546
rect 494164 480 494192 8910
rect 495348 3392 495400 3398
rect 495348 3334 495400 3340
rect 495360 480 495388 3334
rect 495452 610 495480 134506
rect 497462 29472 497518 29481
rect 497462 29407 497518 29416
rect 497476 29073 497504 29407
rect 497462 29064 497518 29073
rect 497462 28999 497518 29008
rect 497740 4820 497792 4826
rect 497740 4762 497792 4768
rect 495440 604 495492 610
rect 495440 546 495492 552
rect 496544 604 496596 610
rect 496544 546 496596 552
rect 496556 480 496584 546
rect 497752 480 497780 4762
rect 498212 610 498240 308450
rect 499580 279472 499632 279478
rect 499580 279414 499632 279420
rect 499592 3482 499620 279414
rect 500972 3482 501000 334698
rect 518900 333328 518952 333334
rect 518900 333270 518952 333276
rect 502340 327820 502392 327826
rect 502340 327762 502392 327768
rect 502246 310856 502302 310865
rect 502246 310791 502302 310800
rect 502260 310758 502288 310791
rect 502248 310752 502300 310758
rect 502248 310694 502300 310700
rect 502248 76084 502300 76090
rect 502248 76026 502300 76032
rect 502260 75857 502288 76026
rect 502246 75848 502302 75857
rect 502246 75783 502302 75792
rect 502352 3482 502380 327762
rect 509240 323672 509292 323678
rect 509240 323614 509292 323620
rect 505100 318164 505152 318170
rect 505100 318106 505152 318112
rect 502432 297492 502484 297498
rect 502432 297434 502484 297440
rect 502444 3670 502472 297434
rect 503720 11756 503772 11762
rect 503720 11698 503772 11704
rect 502432 3664 502484 3670
rect 502432 3606 502484 3612
rect 503628 3664 503680 3670
rect 503628 3606 503680 3612
rect 499592 3454 500172 3482
rect 500972 3454 501276 3482
rect 502352 3454 502472 3482
rect 498200 604 498252 610
rect 498200 546 498252 552
rect 498936 604 498988 610
rect 498936 546 498988 552
rect 498948 480 498976 546
rect 500144 480 500172 3454
rect 501248 480 501276 3454
rect 502444 480 502472 3454
rect 503640 480 503668 3606
rect 503732 3482 503760 11698
rect 505112 3482 505140 318106
rect 506480 291848 506532 291854
rect 506480 291790 506532 291796
rect 506492 3482 506520 291790
rect 507860 13116 507912 13122
rect 507860 13058 507912 13064
rect 507872 3482 507900 13058
rect 509252 3482 509280 323614
rect 514666 321872 514722 321881
rect 514850 321872 514906 321881
rect 514722 321830 514850 321858
rect 514666 321807 514722 321816
rect 514850 321807 514906 321816
rect 516140 316736 516192 316742
rect 516140 316678 516192 316684
rect 514668 310752 514720 310758
rect 514666 310720 514668 310729
rect 514720 310720 514722 310729
rect 514666 310655 514722 310664
rect 512000 307080 512052 307086
rect 512000 307022 512052 307028
rect 510620 278044 510672 278050
rect 510620 277986 510672 277992
rect 510526 76256 510582 76265
rect 510526 76191 510582 76200
rect 510540 76090 510568 76191
rect 510528 76084 510580 76090
rect 510528 76026 510580 76032
rect 510632 3482 510660 277986
rect 503732 3454 504864 3482
rect 505112 3454 506060 3482
rect 506492 3454 507256 3482
rect 507872 3454 508452 3482
rect 509252 3454 509648 3482
rect 510632 3454 510844 3482
rect 504836 480 504864 3454
rect 506032 480 506060 3454
rect 507228 480 507256 3454
rect 508424 480 508452 3454
rect 509620 480 509648 3454
rect 510816 480 510844 3454
rect 512012 3398 512040 307022
rect 513380 276684 513432 276690
rect 513380 276626 513432 276632
rect 512092 14476 512144 14482
rect 512092 14418 512144 14424
rect 512000 3392 512052 3398
rect 512000 3334 512052 3340
rect 512104 1442 512132 14418
rect 513392 3482 513420 276626
rect 514666 29200 514722 29209
rect 514666 29135 514668 29144
rect 514720 29135 514722 29144
rect 514668 29106 514720 29112
rect 514760 15904 514812 15910
rect 514760 15846 514812 15852
rect 514772 3482 514800 15846
rect 516152 3482 516180 316678
rect 517520 273964 517572 273970
rect 517520 273906 517572 273912
rect 517532 3482 517560 273906
rect 518912 3482 518940 333270
rect 521566 310856 521622 310865
rect 521566 310791 521622 310800
rect 521580 310758 521608 310791
rect 521568 310752 521620 310758
rect 521568 310694 521620 310700
rect 520280 305652 520332 305658
rect 520280 305594 520332 305600
rect 513392 3454 514432 3482
rect 514772 3454 515628 3482
rect 516152 3454 516824 3482
rect 517532 3454 517928 3482
rect 518912 3454 519124 3482
rect 513196 3392 513248 3398
rect 513196 3334 513248 3340
rect 512012 1414 512132 1442
rect 512012 480 512040 1414
rect 513208 480 513236 3334
rect 514404 480 514432 3454
rect 515600 480 515628 3454
rect 516796 480 516824 3454
rect 517900 480 517928 3454
rect 519096 480 519124 3454
rect 520292 480 520320 305594
rect 520372 272536 520424 272542
rect 520372 272478 520424 272484
rect 520384 3482 520412 272478
rect 521566 76528 521622 76537
rect 521566 76463 521622 76472
rect 521580 75993 521608 76463
rect 521566 75984 521622 75993
rect 521566 75919 521622 75928
rect 521476 29164 521528 29170
rect 521476 29106 521528 29112
rect 521488 29050 521516 29106
rect 521566 29064 521622 29073
rect 521488 29022 521566 29050
rect 521566 28999 521622 29008
rect 521672 3482 521700 336058
rect 554780 336048 554832 336054
rect 554780 335990 554832 335996
rect 528560 334688 528612 334694
rect 528560 334630 528612 334636
rect 523040 304292 523092 304298
rect 523040 304234 523092 304240
rect 523052 3482 523080 304234
rect 527180 302932 527232 302938
rect 527180 302874 527232 302880
rect 524420 290488 524472 290494
rect 524420 290430 524472 290436
rect 524432 3482 524460 290430
rect 525800 18624 525852 18630
rect 525800 18566 525852 18572
rect 525812 3482 525840 18566
rect 527192 3482 527220 302874
rect 520384 3454 521516 3482
rect 521672 3454 522712 3482
rect 523052 3454 523908 3482
rect 524432 3454 525104 3482
rect 525812 3454 526300 3482
rect 527192 3454 527496 3482
rect 521488 480 521516 3454
rect 522684 480 522712 3454
rect 523880 480 523908 3454
rect 525076 480 525104 3454
rect 526272 480 526300 3454
rect 527468 480 527496 3454
rect 528572 3398 528600 334630
rect 546500 333260 546552 333266
rect 546500 333202 546552 333208
rect 536840 331968 536892 331974
rect 536840 331910 536892 331916
rect 533986 321872 534042 321881
rect 534170 321872 534226 321881
rect 534042 321830 534170 321858
rect 533986 321807 534042 321816
rect 534170 321807 534226 321816
rect 529940 315308 529992 315314
rect 529940 315250 529992 315256
rect 528652 271176 528704 271182
rect 528652 271118 528704 271124
rect 528560 3392 528612 3398
rect 528560 3334 528612 3340
rect 528664 480 528692 271118
rect 529952 3482 529980 315250
rect 533988 310752 534040 310758
rect 533986 310720 533988 310729
rect 534040 310720 534042 310729
rect 533986 310655 534042 310664
rect 534080 301504 534132 301510
rect 534080 301446 534132 301452
rect 531320 269816 531372 269822
rect 531320 269758 531372 269764
rect 531332 3482 531360 269758
rect 533986 227896 534042 227905
rect 533986 227831 533988 227840
rect 534040 227831 534042 227840
rect 533988 227802 534040 227808
rect 533986 76120 534042 76129
rect 533986 76055 533988 76064
rect 534040 76055 534042 76064
rect 533988 76026 534040 76032
rect 533986 29200 534042 29209
rect 533986 29135 533988 29144
rect 534040 29135 534042 29144
rect 533988 29106 534040 29112
rect 532700 19984 532752 19990
rect 532700 19926 532752 19932
rect 532712 3482 532740 19926
rect 534092 3482 534120 301446
rect 535460 268388 535512 268394
rect 535460 268330 535512 268336
rect 535472 3482 535500 268330
rect 536852 3482 536880 331910
rect 539600 330608 539652 330614
rect 539600 330550 539652 330556
rect 536932 300144 536984 300150
rect 536932 300086 536984 300092
rect 536944 3670 536972 300086
rect 538220 267028 538272 267034
rect 538220 266970 538272 266976
rect 536932 3664 536984 3670
rect 536932 3606 536984 3612
rect 538128 3664 538180 3670
rect 538128 3606 538180 3612
rect 529952 3454 531084 3482
rect 531332 3454 532280 3482
rect 532712 3454 533476 3482
rect 534092 3454 534580 3482
rect 535472 3454 535776 3482
rect 536852 3454 536972 3482
rect 529848 3392 529900 3398
rect 529848 3334 529900 3340
rect 529860 480 529888 3334
rect 531056 480 531084 3454
rect 532252 480 532280 3454
rect 533448 480 533476 3454
rect 534552 480 534580 3454
rect 535748 480 535776 3454
rect 536944 480 536972 3454
rect 538140 480 538168 3606
rect 538232 3482 538260 266970
rect 539612 3482 539640 330550
rect 540980 320884 541032 320890
rect 540980 320826 541032 320832
rect 540886 310856 540942 310865
rect 540886 310791 540942 310800
rect 540900 310758 540928 310791
rect 540888 310752 540940 310758
rect 540888 310694 540940 310700
rect 540888 227860 540940 227866
rect 540888 227802 540940 227808
rect 540900 227769 540928 227802
rect 540886 227760 540942 227769
rect 540886 227695 540942 227704
rect 540888 76084 540940 76090
rect 540888 76026 540940 76032
rect 540900 75993 540928 76026
rect 540886 75984 540942 75993
rect 540886 75919 540942 75928
rect 540796 29164 540848 29170
rect 540796 29106 540848 29112
rect 540808 29050 540836 29106
rect 540886 29064 540942 29073
rect 540808 29022 540886 29050
rect 540886 28999 540942 29008
rect 540992 3482 541020 320826
rect 545120 313948 545172 313954
rect 545120 313890 545172 313896
rect 541070 310856 541126 310865
rect 541070 310791 541072 310800
rect 541124 310791 541126 310800
rect 543832 310820 543884 310826
rect 541072 310762 541124 310768
rect 543832 310762 543884 310768
rect 543844 310593 543872 310762
rect 543830 310584 543886 310593
rect 543830 310519 543886 310528
rect 542360 265668 542412 265674
rect 542360 265610 542412 265616
rect 542372 3482 542400 265610
rect 543740 21412 543792 21418
rect 543740 21354 543792 21360
rect 543752 3482 543780 21354
rect 545132 3482 545160 313890
rect 546512 3670 546540 333202
rect 550640 329112 550692 329118
rect 550640 329054 550692 329060
rect 547880 297424 547932 297430
rect 547880 297366 547932 297372
rect 546592 262880 546644 262886
rect 546592 262822 546644 262828
rect 546500 3664 546552 3670
rect 546500 3606 546552 3612
rect 546604 3482 546632 262822
rect 547696 3664 547748 3670
rect 547696 3606 547748 3612
rect 538232 3454 539364 3482
rect 539612 3454 540560 3482
rect 540992 3454 541756 3482
rect 542372 3454 542952 3482
rect 543752 3454 544148 3482
rect 545132 3454 545344 3482
rect 539336 480 539364 3454
rect 540532 480 540560 3454
rect 541728 480 541756 3454
rect 542924 480 542952 3454
rect 544120 480 544148 3454
rect 545316 480 545344 3454
rect 546512 3454 546632 3482
rect 546512 480 546540 3454
rect 547708 480 547736 3606
rect 547892 3482 547920 297366
rect 549260 289128 549312 289134
rect 549260 289070 549312 289076
rect 549272 3482 549300 289070
rect 550652 3482 550680 329054
rect 552020 312588 552072 312594
rect 552020 312530 552072 312536
rect 552032 3482 552060 312530
rect 553400 261520 553452 261526
rect 553400 261462 553452 261468
rect 553306 227896 553362 227905
rect 553306 227831 553308 227840
rect 553360 227831 553362 227840
rect 553308 227802 553360 227808
rect 553306 76120 553362 76129
rect 553306 76055 553308 76064
rect 553360 76055 553362 76064
rect 553308 76026 553360 76032
rect 553306 29200 553362 29209
rect 553306 29135 553308 29144
rect 553360 29135 553362 29144
rect 553308 29106 553360 29112
rect 553412 3482 553440 261462
rect 547892 3454 548932 3482
rect 549272 3454 550128 3482
rect 550652 3454 551232 3482
rect 552032 3454 552428 3482
rect 553412 3454 553624 3482
rect 548904 480 548932 3454
rect 550100 480 550128 3454
rect 551204 480 551232 3454
rect 552400 480 552428 3454
rect 553596 480 553624 3454
rect 554792 480 554820 335990
rect 574744 334620 574796 334626
rect 574744 334562 574796 334568
rect 560944 331900 560996 331906
rect 560944 331842 560996 331848
rect 557540 327752 557592 327758
rect 557540 327694 557592 327700
rect 554872 322244 554924 322250
rect 554872 322186 554924 322192
rect 554884 3482 554912 322186
rect 556804 319456 556856 319462
rect 556804 319398 556856 319404
rect 555422 310584 555478 310593
rect 555422 310519 555478 310528
rect 555436 310321 555464 310519
rect 555422 310312 555478 310321
rect 555422 310247 555478 310256
rect 556160 260160 556212 260166
rect 556160 260102 556212 260108
rect 556172 3618 556200 260102
rect 556816 4146 556844 319398
rect 556804 4140 556856 4146
rect 556804 4082 556856 4088
rect 556172 3590 557212 3618
rect 554884 3454 556016 3482
rect 555988 480 556016 3454
rect 557184 480 557212 3590
rect 557552 3482 557580 327694
rect 560300 258732 560352 258738
rect 560300 258674 560352 258680
rect 560208 227860 560260 227866
rect 560208 227802 560260 227808
rect 560220 227769 560248 227802
rect 560206 227760 560262 227769
rect 560206 227695 560262 227704
rect 560208 76084 560260 76090
rect 560208 76026 560260 76032
rect 560220 75993 560248 76026
rect 560206 75984 560262 75993
rect 560206 75919 560262 75928
rect 560116 29164 560168 29170
rect 560116 29106 560168 29112
rect 560128 29050 560156 29106
rect 560206 29064 560262 29073
rect 560128 29022 560206 29050
rect 560206 28999 560262 29008
rect 559564 4140 559616 4146
rect 559564 4082 559616 4088
rect 557552 3454 558408 3482
rect 558380 480 558408 3454
rect 559576 480 559604 4082
rect 560312 3482 560340 258674
rect 560312 3454 560800 3482
rect 560772 480 560800 3454
rect 560956 3398 560984 331842
rect 573364 330540 573416 330546
rect 573364 330482 573416 330488
rect 564440 326392 564492 326398
rect 564440 326334 564492 326340
rect 562874 321736 562930 321745
rect 563150 321736 563206 321745
rect 562930 321694 563150 321722
rect 562874 321671 562930 321680
rect 563150 321671 563206 321680
rect 563060 309800 563112 309806
rect 563060 309742 563112 309748
rect 563072 3482 563100 309742
rect 563152 257372 563204 257378
rect 563152 257314 563204 257320
rect 563164 3670 563192 257314
rect 563152 3664 563204 3670
rect 563152 3606 563204 3612
rect 564348 3664 564400 3670
rect 564348 3606 564400 3612
rect 563072 3454 563192 3482
rect 560944 3392 560996 3398
rect 560944 3334 560996 3340
rect 561956 3392 562008 3398
rect 561956 3334 562008 3340
rect 561968 480 561996 3334
rect 563164 480 563192 3454
rect 564360 480 564388 3606
rect 564452 3346 564480 326334
rect 568580 324964 568632 324970
rect 568580 324906 568632 324912
rect 567844 318096 567896 318102
rect 567844 318038 567896 318044
rect 565084 295996 565136 296002
rect 565084 295938 565136 295944
rect 565096 3670 565124 295938
rect 567200 22772 567252 22778
rect 567200 22714 567252 22720
rect 565084 3664 565136 3670
rect 565084 3606 565136 3612
rect 566740 3664 566792 3670
rect 566740 3606 566792 3612
rect 564452 3318 565584 3346
rect 565556 480 565584 3318
rect 566752 480 566780 3606
rect 567212 3346 567240 22714
rect 567856 3806 567884 318038
rect 567844 3800 567896 3806
rect 567844 3742 567896 3748
rect 568592 3346 568620 324906
rect 571340 323604 571392 323610
rect 571340 323546 571392 323552
rect 569960 294636 570012 294642
rect 569960 294578 570012 294584
rect 569972 3346 570000 294578
rect 571352 3602 571380 323546
rect 572626 321872 572682 321881
rect 572626 321807 572682 321816
rect 572640 321722 572668 321807
rect 572718 321736 572774 321745
rect 572640 321694 572718 321722
rect 572718 321671 572774 321680
rect 571432 287700 571484 287706
rect 571432 287642 571484 287648
rect 571340 3596 571392 3602
rect 571340 3538 571392 3544
rect 567212 3318 567884 3346
rect 568592 3318 569080 3346
rect 569972 3318 570276 3346
rect 567856 480 567884 3318
rect 569052 480 569080 3318
rect 570248 480 570276 3318
rect 571444 480 571472 287642
rect 572626 227896 572682 227905
rect 572626 227831 572628 227840
rect 572680 227831 572682 227840
rect 572628 227802 572680 227808
rect 572626 76120 572682 76129
rect 572626 76055 572628 76064
rect 572680 76055 572682 76064
rect 572628 76026 572680 76032
rect 572626 29200 572682 29209
rect 572626 29135 572628 29144
rect 572680 29135 572682 29144
rect 572628 29106 572680 29112
rect 573376 3738 573404 330482
rect 573456 293276 573508 293282
rect 573456 293218 573508 293224
rect 573364 3732 573416 3738
rect 573364 3674 573416 3680
rect 573468 3670 573496 293218
rect 573824 3800 573876 3806
rect 573824 3742 573876 3748
rect 573456 3664 573508 3670
rect 573456 3606 573508 3612
rect 572628 3596 572680 3602
rect 572628 3538 572680 3544
rect 572640 480 572668 3538
rect 573836 480 573864 3742
rect 574756 3058 574784 334562
rect 574836 308440 574888 308446
rect 574836 308382 574888 308388
rect 574848 3330 574876 308382
rect 579804 299464 579856 299470
rect 579804 299406 579856 299412
rect 579816 299169 579844 299406
rect 579802 299160 579858 299169
rect 579802 299095 579858 299104
rect 580172 276004 580224 276010
rect 580172 275946 580224 275952
rect 580184 275777 580212 275946
rect 580170 275768 580226 275777
rect 580170 275703 580226 275712
rect 580172 264920 580224 264926
rect 580172 264862 580224 264868
rect 580184 263945 580212 264862
rect 580170 263936 580226 263945
rect 580170 263871 580226 263880
rect 579804 252544 579856 252550
rect 579804 252486 579856 252492
rect 579816 252249 579844 252486
rect 579802 252240 579858 252249
rect 579802 252175 579858 252184
rect 579528 227860 579580 227866
rect 579528 227802 579580 227808
rect 579540 227769 579568 227802
rect 579526 227760 579582 227769
rect 579526 227695 579582 227704
rect 580172 218000 580224 218006
rect 580172 217942 580224 217948
rect 580184 217025 580212 217942
rect 580170 217016 580226 217025
rect 580170 216951 580226 216960
rect 579804 205624 579856 205630
rect 579804 205566 579856 205572
rect 579816 205329 579844 205566
rect 579802 205320 579858 205329
rect 579802 205255 579858 205264
rect 580172 182164 580224 182170
rect 580172 182106 580224 182112
rect 580184 181937 580212 182106
rect 580170 181928 580226 181937
rect 580170 181863 580226 181872
rect 580172 171080 580224 171086
rect 580172 171022 580224 171028
rect 580184 170105 580212 171022
rect 580170 170096 580226 170105
rect 580170 170031 580226 170040
rect 579804 158704 579856 158710
rect 579804 158646 579856 158652
rect 579816 158409 579844 158646
rect 579802 158400 579858 158409
rect 579802 158335 579858 158344
rect 580172 135244 580224 135250
rect 580172 135186 580224 135192
rect 580184 134881 580212 135186
rect 580170 134872 580226 134881
rect 580170 134807 580226 134816
rect 580172 124160 580224 124166
rect 580172 124102 580224 124108
rect 580184 123185 580212 124102
rect 580170 123176 580226 123185
rect 580170 123111 580226 123120
rect 579804 111784 579856 111790
rect 579804 111726 579856 111732
rect 579816 111489 579844 111726
rect 579802 111480 579858 111489
rect 579802 111415 579858 111424
rect 580172 88324 580224 88330
rect 580172 88266 580224 88272
rect 580184 87961 580212 88266
rect 580170 87952 580226 87961
rect 580170 87887 580226 87896
rect 579528 76084 579580 76090
rect 579528 76026 579580 76032
rect 579540 75993 579568 76026
rect 579526 75984 579582 75993
rect 579526 75919 579582 75928
rect 579804 64864 579856 64870
rect 579804 64806 579856 64812
rect 579816 64569 579844 64806
rect 579802 64560 579858 64569
rect 579802 64495 579858 64504
rect 580172 41404 580224 41410
rect 580172 41346 580224 41352
rect 580184 41041 580212 41346
rect 580170 41032 580226 41041
rect 580170 40967 580226 40976
rect 579436 29164 579488 29170
rect 579436 29106 579488 29112
rect 579448 29050 579476 29106
rect 579526 29064 579582 29073
rect 579448 29022 579526 29050
rect 579526 28999 579582 29008
rect 579804 17944 579856 17950
rect 579804 17886 579856 17892
rect 579816 17649 579844 17886
rect 579802 17640 579858 17649
rect 579802 17575 579858 17584
rect 579804 3732 579856 3738
rect 579804 3674 579856 3680
rect 578608 3392 578660 3398
rect 578608 3334 578660 3340
rect 574836 3324 574888 3330
rect 574836 3266 574888 3272
rect 577412 3324 577464 3330
rect 577412 3266 577464 3272
rect 575020 3256 575072 3262
rect 575020 3198 575072 3204
rect 574744 3052 574796 3058
rect 574744 2994 574796 3000
rect 575032 480 575060 3198
rect 576216 3052 576268 3058
rect 576216 2994 576268 3000
rect 576228 480 576256 2994
rect 577424 480 577452 3266
rect 578620 480 578648 3334
rect 579816 480 579844 3674
rect 581000 3664 581052 3670
rect 581000 3606 581052 3612
rect 581012 480 581040 3606
rect 582196 3460 582248 3466
rect 582196 3402 582248 3408
rect 582208 480 582236 3402
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8822 -960 8934 480
rect 10018 -960 10130 480
rect 11214 -960 11326 480
rect 12410 -960 12522 480
rect 13606 -960 13718 480
rect 14802 -960 14914 480
rect 15998 -960 16110 480
rect 17194 -960 17306 480
rect 18298 -960 18410 480
rect 19494 -960 19606 480
rect 20690 -960 20802 480
rect 21886 -960 21998 480
rect 23082 -960 23194 480
rect 24278 -960 24390 480
rect 25474 -960 25586 480
rect 26670 -960 26782 480
rect 27866 -960 27978 480
rect 29062 -960 29174 480
rect 30258 -960 30370 480
rect 31454 -960 31566 480
rect 32650 -960 32762 480
rect 33846 -960 33958 480
rect 34950 -960 35062 480
rect 36146 -960 36258 480
rect 37342 -960 37454 480
rect 38538 -960 38650 480
rect 39734 -960 39846 480
rect 40930 -960 41042 480
rect 42126 -960 42238 480
rect 43322 -960 43434 480
rect 44518 -960 44630 480
rect 45714 -960 45826 480
rect 46910 -960 47022 480
rect 48106 -960 48218 480
rect 49302 -960 49414 480
rect 50498 -960 50610 480
rect 51602 -960 51714 480
rect 52798 -960 52910 480
rect 53994 -960 54106 480
rect 55190 -960 55302 480
rect 56386 -960 56498 480
rect 57582 -960 57694 480
rect 58778 -960 58890 480
rect 59974 -960 60086 480
rect 61170 -960 61282 480
rect 62366 -960 62478 480
rect 63562 -960 63674 480
rect 64758 -960 64870 480
rect 65954 -960 66066 480
rect 67150 -960 67262 480
rect 68254 -960 68366 480
rect 69450 -960 69562 480
rect 70646 -960 70758 480
rect 71842 -960 71954 480
rect 73038 -960 73150 480
rect 74234 -960 74346 480
rect 75430 -960 75542 480
rect 76626 -960 76738 480
rect 77822 -960 77934 480
rect 79018 -960 79130 480
rect 80214 -960 80326 480
rect 81410 -960 81522 480
rect 82606 -960 82718 480
rect 83802 -960 83914 480
rect 84906 -960 85018 480
rect 86102 -960 86214 480
rect 87298 -960 87410 480
rect 88494 -960 88606 480
rect 89690 -960 89802 480
rect 90886 -960 90998 480
rect 92082 -960 92194 480
rect 93278 -960 93390 480
rect 94474 -960 94586 480
rect 95670 -960 95782 480
rect 96866 -960 96978 480
rect 98062 -960 98174 480
rect 99258 -960 99370 480
rect 100454 -960 100566 480
rect 101558 -960 101670 480
rect 102754 -960 102866 480
rect 103950 -960 104062 480
rect 105146 -960 105258 480
rect 106342 -960 106454 480
rect 107538 -960 107650 480
rect 108734 -960 108846 480
rect 109930 -960 110042 480
rect 111126 -960 111238 480
rect 112322 -960 112434 480
rect 113518 -960 113630 480
rect 114714 -960 114826 480
rect 115910 -960 116022 480
rect 117106 -960 117218 480
rect 118210 -960 118322 480
rect 119406 -960 119518 480
rect 120602 -960 120714 480
rect 121798 -960 121910 480
rect 122994 -960 123106 480
rect 124190 -960 124302 480
rect 125386 -960 125498 480
rect 126582 -960 126694 480
rect 127778 -960 127890 480
rect 128974 -960 129086 480
rect 130170 -960 130282 480
rect 131366 -960 131478 480
rect 132562 -960 132674 480
rect 133758 -960 133870 480
rect 134862 -960 134974 480
rect 136058 -960 136170 480
rect 137254 -960 137366 480
rect 138450 -960 138562 480
rect 139646 -960 139758 480
rect 140842 -960 140954 480
rect 142038 -960 142150 480
rect 143234 -960 143346 480
rect 144430 -960 144542 480
rect 145626 -960 145738 480
rect 146822 -960 146934 480
rect 148018 -960 148130 480
rect 149214 -960 149326 480
rect 150410 -960 150522 480
rect 151514 -960 151626 480
rect 152710 -960 152822 480
rect 153906 -960 154018 480
rect 155102 -960 155214 480
rect 156298 -960 156410 480
rect 157494 -960 157606 480
rect 158690 -960 158802 480
rect 159886 -960 159998 480
rect 161082 -960 161194 480
rect 162278 -960 162390 480
rect 163474 -960 163586 480
rect 164670 -960 164782 480
rect 165866 -960 165978 480
rect 167062 -960 167174 480
rect 168166 -960 168278 480
rect 169362 -960 169474 480
rect 170558 -960 170670 480
rect 171754 -960 171866 480
rect 172950 -960 173062 480
rect 174146 -960 174258 480
rect 175342 -960 175454 480
rect 176538 -960 176650 480
rect 177734 -960 177846 480
rect 178930 -960 179042 480
rect 180126 -960 180238 480
rect 181322 -960 181434 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184818 -960 184930 480
rect 186014 -960 186126 480
rect 187210 -960 187322 480
rect 188406 -960 188518 480
rect 189602 -960 189714 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197974 -960 198086 480
rect 199170 -960 199282 480
rect 200366 -960 200478 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206254 -960 206366 480
rect 207450 -960 207562 480
rect 208646 -960 208758 480
rect 209842 -960 209954 480
rect 211038 -960 211150 480
rect 212234 -960 212346 480
rect 213430 -960 213542 480
rect 214626 -960 214738 480
rect 215822 -960 215934 480
rect 217018 -960 217130 480
rect 218122 -960 218234 480
rect 219318 -960 219430 480
rect 220514 -960 220626 480
rect 221710 -960 221822 480
rect 222906 -960 223018 480
rect 224102 -960 224214 480
rect 225298 -960 225410 480
rect 226494 -960 226606 480
rect 227690 -960 227802 480
rect 228886 -960 228998 480
rect 230082 -960 230194 480
rect 231278 -960 231390 480
rect 232474 -960 232586 480
rect 233670 -960 233782 480
rect 234774 -960 234886 480
rect 235970 -960 236082 480
rect 237166 -960 237278 480
rect 238362 -960 238474 480
rect 239558 -960 239670 480
rect 240754 -960 240866 480
rect 241950 -960 242062 480
rect 243146 -960 243258 480
rect 244342 -960 244454 480
rect 245538 -960 245650 480
rect 246734 -960 246846 480
rect 247930 -960 248042 480
rect 249126 -960 249238 480
rect 250322 -960 250434 480
rect 251426 -960 251538 480
rect 252622 -960 252734 480
rect 253818 -960 253930 480
rect 255014 -960 255126 480
rect 256210 -960 256322 480
rect 257406 -960 257518 480
rect 258602 -960 258714 480
rect 259798 -960 259910 480
rect 260994 -960 261106 480
rect 262190 -960 262302 480
rect 263386 -960 263498 480
rect 264582 -960 264694 480
rect 265778 -960 265890 480
rect 266974 -960 267086 480
rect 268078 -960 268190 480
rect 269274 -960 269386 480
rect 270470 -960 270582 480
rect 271666 -960 271778 480
rect 272862 -960 272974 480
rect 274058 -960 274170 480
rect 275254 -960 275366 480
rect 276450 -960 276562 480
rect 277646 -960 277758 480
rect 278842 -960 278954 480
rect 280038 -960 280150 480
rect 281234 -960 281346 480
rect 282430 -960 282542 480
rect 283626 -960 283738 480
rect 284730 -960 284842 480
rect 285926 -960 286038 480
rect 287122 -960 287234 480
rect 288318 -960 288430 480
rect 289514 -960 289626 480
rect 290710 -960 290822 480
rect 291906 -960 292018 480
rect 293102 -960 293214 480
rect 294298 -960 294410 480
rect 295494 -960 295606 480
rect 296690 -960 296802 480
rect 297886 -960 297998 480
rect 299082 -960 299194 480
rect 300278 -960 300390 480
rect 301382 -960 301494 480
rect 302578 -960 302690 480
rect 303774 -960 303886 480
rect 304970 -960 305082 480
rect 306166 -960 306278 480
rect 307362 -960 307474 480
rect 308558 -960 308670 480
rect 309754 -960 309866 480
rect 310950 -960 311062 480
rect 312146 -960 312258 480
rect 313342 -960 313454 480
rect 314538 -960 314650 480
rect 315734 -960 315846 480
rect 316930 -960 317042 480
rect 318034 -960 318146 480
rect 319230 -960 319342 480
rect 320426 -960 320538 480
rect 321622 -960 321734 480
rect 322818 -960 322930 480
rect 324014 -960 324126 480
rect 325210 -960 325322 480
rect 326406 -960 326518 480
rect 327602 -960 327714 480
rect 328798 -960 328910 480
rect 329994 -960 330106 480
rect 331190 -960 331302 480
rect 332386 -960 332498 480
rect 333582 -960 333694 480
rect 334686 -960 334798 480
rect 335882 -960 335994 480
rect 337078 -960 337190 480
rect 338274 -960 338386 480
rect 339470 -960 339582 480
rect 340666 -960 340778 480
rect 341862 -960 341974 480
rect 343058 -960 343170 480
rect 344254 -960 344366 480
rect 345450 -960 345562 480
rect 346646 -960 346758 480
rect 347842 -960 347954 480
rect 349038 -960 349150 480
rect 350234 -960 350346 480
rect 351338 -960 351450 480
rect 352534 -960 352646 480
rect 353730 -960 353842 480
rect 354926 -960 355038 480
rect 356122 -960 356234 480
rect 357318 -960 357430 480
rect 358514 -960 358626 480
rect 359710 -960 359822 480
rect 360906 -960 361018 480
rect 362102 -960 362214 480
rect 363298 -960 363410 480
rect 364494 -960 364606 480
rect 365690 -960 365802 480
rect 366886 -960 366998 480
rect 367990 -960 368102 480
rect 369186 -960 369298 480
rect 370382 -960 370494 480
rect 371578 -960 371690 480
rect 372774 -960 372886 480
rect 373970 -960 374082 480
rect 375166 -960 375278 480
rect 376362 -960 376474 480
rect 377558 -960 377670 480
rect 378754 -960 378866 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384642 -960 384754 480
rect 385838 -960 385950 480
rect 387034 -960 387146 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395406 -960 395518 480
rect 396602 -960 396714 480
rect 397798 -960 397910 480
rect 398994 -960 399106 480
rect 400190 -960 400302 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403686 -960 403798 480
rect 404882 -960 404994 480
rect 406078 -960 406190 480
rect 407274 -960 407386 480
rect 408470 -960 408582 480
rect 409666 -960 409778 480
rect 410862 -960 410974 480
rect 412058 -960 412170 480
rect 413254 -960 413366 480
rect 414450 -960 414562 480
rect 415646 -960 415758 480
rect 416842 -960 416954 480
rect 417946 -960 418058 480
rect 419142 -960 419254 480
rect 420338 -960 420450 480
rect 421534 -960 421646 480
rect 422730 -960 422842 480
rect 423926 -960 424038 480
rect 425122 -960 425234 480
rect 426318 -960 426430 480
rect 427514 -960 427626 480
rect 428710 -960 428822 480
rect 429906 -960 430018 480
rect 431102 -960 431214 480
rect 432298 -960 432410 480
rect 433494 -960 433606 480
rect 434598 -960 434710 480
rect 435794 -960 435906 480
rect 436990 -960 437102 480
rect 438186 -960 438298 480
rect 439382 -960 439494 480
rect 440578 -960 440690 480
rect 441774 -960 441886 480
rect 442970 -960 443082 480
rect 444166 -960 444278 480
rect 445362 -960 445474 480
rect 446558 -960 446670 480
rect 447754 -960 447866 480
rect 448950 -960 449062 480
rect 450146 -960 450258 480
rect 451250 -960 451362 480
rect 452446 -960 452558 480
rect 453642 -960 453754 480
rect 454838 -960 454950 480
rect 456034 -960 456146 480
rect 457230 -960 457342 480
rect 458426 -960 458538 480
rect 459622 -960 459734 480
rect 460818 -960 460930 480
rect 462014 -960 462126 480
rect 463210 -960 463322 480
rect 464406 -960 464518 480
rect 465602 -960 465714 480
rect 466798 -960 466910 480
rect 467902 -960 468014 480
rect 469098 -960 469210 480
rect 470294 -960 470406 480
rect 471490 -960 471602 480
rect 472686 -960 472798 480
rect 473882 -960 473994 480
rect 475078 -960 475190 480
rect 476274 -960 476386 480
rect 477470 -960 477582 480
rect 478666 -960 478778 480
rect 479862 -960 479974 480
rect 481058 -960 481170 480
rect 482254 -960 482366 480
rect 483450 -960 483562 480
rect 484554 -960 484666 480
rect 485750 -960 485862 480
rect 486946 -960 487058 480
rect 488142 -960 488254 480
rect 489338 -960 489450 480
rect 490534 -960 490646 480
rect 491730 -960 491842 480
rect 492926 -960 493038 480
rect 494122 -960 494234 480
rect 495318 -960 495430 480
rect 496514 -960 496626 480
rect 497710 -960 497822 480
rect 498906 -960 499018 480
rect 500102 -960 500214 480
rect 501206 -960 501318 480
rect 502402 -960 502514 480
rect 503598 -960 503710 480
rect 504794 -960 504906 480
rect 505990 -960 506102 480
rect 507186 -960 507298 480
rect 508382 -960 508494 480
rect 509578 -960 509690 480
rect 510774 -960 510886 480
rect 511970 -960 512082 480
rect 513166 -960 513278 480
rect 514362 -960 514474 480
rect 515558 -960 515670 480
rect 516754 -960 516866 480
rect 517858 -960 517970 480
rect 519054 -960 519166 480
rect 520250 -960 520362 480
rect 521446 -960 521558 480
rect 522642 -960 522754 480
rect 523838 -960 523950 480
rect 525034 -960 525146 480
rect 526230 -960 526342 480
rect 527426 -960 527538 480
rect 528622 -960 528734 480
rect 529818 -960 529930 480
rect 531014 -960 531126 480
rect 532210 -960 532322 480
rect 533406 -960 533518 480
rect 534510 -960 534622 480
rect 535706 -960 535818 480
rect 536902 -960 537014 480
rect 538098 -960 538210 480
rect 539294 -960 539406 480
rect 540490 -960 540602 480
rect 541686 -960 541798 480
rect 542882 -960 542994 480
rect 544078 -960 544190 480
rect 545274 -960 545386 480
rect 546470 -960 546582 480
rect 547666 -960 547778 480
rect 548862 -960 548974 480
rect 550058 -960 550170 480
rect 551162 -960 551274 480
rect 552358 -960 552470 480
rect 553554 -960 553666 480
rect 554750 -960 554862 480
rect 555946 -960 556058 480
rect 557142 -960 557254 480
rect 558338 -960 558450 480
rect 559534 -960 559646 480
rect 560730 -960 560842 480
rect 561926 -960 562038 480
rect 563122 -960 563234 480
rect 564318 -960 564430 480
rect 565514 -960 565626 480
rect 566710 -960 566822 480
rect 567814 -960 567926 480
rect 569010 -960 569122 480
rect 570206 -960 570318 480
rect 571402 -960 571514 480
rect 572598 -960 572710 480
rect 573794 -960 573906 480
rect 574990 -960 575102 480
rect 576186 -960 576298 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 682216 3478 682272
rect 3330 653520 3386 653576
rect 3054 595992 3110 596048
rect 2962 553016 3018 553072
rect 3146 538600 3202 538656
rect 3330 495508 3386 495544
rect 3330 495488 3332 495508
rect 3332 495488 3384 495508
rect 3384 495488 3386 495508
rect 3146 481072 3202 481128
rect 3238 452376 3294 452432
rect 2962 437960 3018 438016
rect 3330 423700 3386 423736
rect 3330 423680 3332 423700
rect 3332 423680 3384 423700
rect 3384 423680 3386 423700
rect 3514 667936 3570 667992
rect 3606 624824 3662 624880
rect 3698 610408 3754 610464
rect 3882 567296 3938 567352
rect 4066 509904 4122 509960
rect 154210 482976 154266 483032
rect 154486 482976 154542 483032
rect 154118 415384 154174 415440
rect 154302 415384 154358 415440
rect 154302 415248 154358 415304
rect 154486 415248 154542 415304
rect 218886 695680 218942 695736
rect 219254 695544 219310 695600
rect 218978 540912 219034 540968
rect 219162 540912 219218 540968
rect 218978 531256 219034 531312
rect 219162 531256 219218 531312
rect 218794 521600 218850 521656
rect 218978 521600 219034 521656
rect 218978 473320 219034 473376
rect 219254 473320 219310 473376
rect 218978 425040 219034 425096
rect 219346 425040 219402 425096
rect 235814 401920 235870 401976
rect 3146 394984 3202 395040
rect 2962 366152 3018 366208
rect 3422 380568 3478 380624
rect 3422 337456 3478 337512
rect 3422 335960 3478 336016
rect 3330 323040 3386 323096
rect 3330 308760 3386 308816
rect 3146 251232 3202 251288
rect 3146 222536 3202 222592
rect 3238 179424 3294 179480
rect 2962 122032 3018 122088
rect 3238 78920 3294 78976
rect 3054 50088 3110 50144
rect 3514 294344 3570 294400
rect 3514 265648 3570 265704
rect 3974 280064 4030 280120
rect 3790 236952 3846 237008
rect 3514 208120 3570 208176
rect 3514 194520 3570 194576
rect 3514 193840 3570 193896
rect 3514 165008 3570 165064
rect 3514 151680 3570 151736
rect 3514 150728 3570 150784
rect 3514 136312 3570 136368
rect 3514 108976 3570 109032
rect 3514 107616 3570 107672
rect 3514 93200 3570 93256
rect 3514 35844 3516 35864
rect 3516 35844 3568 35864
rect 3568 35844 3570 35864
rect 3514 35808 3570 35844
rect 3422 21392 3478 21448
rect 3422 7112 3478 7168
rect 6458 3304 6514 3360
rect 14830 3440 14886 3496
rect 16026 3576 16082 3632
rect 25502 3848 25558 3904
rect 24306 3712 24362 3768
rect 32678 3984 32734 4040
rect 240322 399472 240378 399528
rect 580170 697992 580226 698048
rect 580170 686296 580226 686352
rect 580170 674600 580226 674656
rect 580170 651072 580226 651128
rect 580170 639376 580226 639432
rect 580170 627680 580226 627736
rect 580170 604152 580226 604208
rect 580170 592456 580226 592512
rect 580170 580760 580226 580816
rect 299570 560496 299626 560552
rect 299570 560360 299626 560416
rect 580170 557232 580226 557288
rect 299294 549208 299350 549264
rect 299478 549208 299534 549264
rect 580170 545536 580226 545592
rect 580170 533840 580226 533896
rect 299662 521600 299718 521656
rect 299846 521600 299902 521656
rect 580170 510312 580226 510368
rect 299478 502288 299534 502344
rect 299754 502324 299756 502344
rect 299756 502324 299808 502344
rect 299808 502324 299810 502344
rect 299754 502288 299810 502324
rect 580170 498616 580226 498672
rect 299478 492632 299534 492688
rect 299662 492652 299718 492688
rect 299662 492632 299664 492652
rect 299664 492632 299716 492652
rect 299716 492632 299718 492652
rect 580170 486784 580226 486840
rect 580170 463392 580226 463448
rect 580170 451696 580226 451752
rect 580170 439864 580226 439920
rect 580170 416472 580226 416528
rect 580170 404776 580226 404832
rect 485042 401920 485098 401976
rect 289634 401784 289690 401840
rect 231582 399336 231638 399392
rect 232962 399336 233018 399392
rect 234066 399336 234122 399392
rect 237194 399336 237250 399392
rect 237838 399336 237894 399392
rect 239402 399336 239458 399392
rect 240966 399336 241022 399392
rect 283010 399336 283066 399392
rect 284482 399336 284538 399392
rect 286138 399336 286194 399392
rect 287794 399336 287850 399392
rect 229558 241440 229614 241496
rect 229834 241440 229890 241496
rect 229558 222128 229614 222184
rect 229834 222128 229890 222184
rect 229558 202816 229614 202872
rect 229834 202816 229890 202872
rect 229558 183504 229614 183560
rect 229834 183504 229890 183560
rect 229650 154536 229706 154592
rect 229834 154536 229890 154592
rect 229466 135224 229522 135280
rect 229650 135224 229706 135280
rect 229466 115912 229522 115968
rect 229650 115912 229706 115968
rect 229466 96600 229522 96656
rect 229650 96600 229706 96656
rect 229650 67496 229706 67552
rect 229650 57976 229706 58032
rect 229098 3168 229154 3224
rect 231122 3576 231178 3632
rect 232962 3848 233018 3904
rect 232778 3712 232834 3768
rect 230662 3440 230718 3496
rect 230938 3440 230994 3496
rect 233238 3476 233240 3496
rect 233240 3476 233292 3496
rect 233292 3476 233294 3496
rect 230570 3304 230626 3360
rect 233238 3440 233294 3476
rect 234434 3984 234490 4040
rect 233790 3204 233792 3224
rect 233792 3204 233844 3224
rect 233844 3204 233846 3224
rect 233790 3168 233846 3204
rect 237654 278704 237710 278760
rect 237654 264288 237710 264344
rect 237470 219408 237526 219464
rect 237654 219408 237710 219464
rect 237562 153312 237618 153368
rect 237562 153196 237618 153232
rect 237562 153176 237564 153196
rect 237564 153176 237616 153196
rect 237616 153176 237618 153196
rect 237562 124344 237618 124400
rect 237654 124208 237710 124264
rect 238298 238856 238354 238912
rect 238114 238720 238170 238776
rect 238666 124208 238722 124264
rect 238850 219408 238906 219464
rect 238942 153196 238998 153232
rect 238942 153176 238944 153196
rect 238944 153176 238996 153196
rect 238996 153176 238998 153196
rect 238942 124208 238998 124264
rect 239126 219408 239182 219464
rect 239126 153176 239182 153232
rect 240874 237360 240930 237416
rect 240874 219408 240930 219464
rect 240874 27512 240930 27568
rect 241058 237360 241114 237416
rect 241058 219408 241114 219464
rect 241150 191800 241206 191856
rect 241334 191800 241390 191856
rect 241150 172488 241206 172544
rect 241334 172488 241390 172544
rect 241150 125704 241206 125760
rect 241058 125568 241114 125624
rect 241058 27512 241114 27568
rect 244186 228112 244242 228168
rect 244370 227976 244426 228032
rect 244278 75928 244334 75984
rect 244462 75928 244518 75984
rect 248418 227976 248474 228032
rect 248418 227568 248474 227624
rect 248878 106120 248934 106176
rect 248970 105848 249026 105904
rect 252006 335688 252062 335744
rect 251638 335416 251694 335472
rect 251362 258032 251418 258088
rect 251362 257896 251418 257952
rect 251546 202816 251602 202872
rect 251730 202816 251786 202872
rect 254122 335416 254178 335472
rect 253846 296656 253902 296712
rect 254030 296656 254086 296712
rect 253938 201456 253994 201512
rect 254122 201456 254178 201512
rect 253938 144880 253994 144936
rect 254122 144880 254178 144936
rect 254582 335416 254638 335472
rect 256422 325624 256478 325680
rect 256606 325624 256662 325680
rect 256422 316004 256424 316024
rect 256424 316004 256476 316024
rect 256476 316004 256478 316024
rect 256422 315968 256478 316004
rect 256606 316004 256608 316024
rect 256608 316004 256660 316024
rect 256660 316004 256662 316024
rect 256606 315968 256662 316004
rect 256422 132368 256478 132424
rect 256606 132368 256662 132424
rect 258538 84088 258594 84144
rect 258722 83952 258778 84008
rect 259458 227996 259514 228032
rect 259458 227976 259460 227996
rect 259460 227976 259512 227996
rect 259512 227976 259514 227996
rect 259734 220768 259790 220824
rect 259734 211112 259790 211168
rect 259734 191800 259790 191856
rect 260102 220768 260158 220824
rect 260286 220768 260342 220824
rect 259918 211112 259974 211168
rect 259918 191800 259974 191856
rect 259918 183504 259974 183560
rect 260194 211112 260250 211168
rect 260102 183504 260158 183560
rect 260194 145016 260250 145072
rect 260102 144900 260158 144936
rect 260102 144880 260104 144900
rect 260104 144880 260156 144900
rect 260156 144880 260158 144900
rect 260102 134000 260158 134056
rect 260286 133884 260342 133920
rect 260286 133864 260288 133884
rect 260288 133864 260340 133884
rect 260340 133864 260342 133884
rect 260102 17992 260158 18048
rect 260378 17992 260434 18048
rect 260562 220768 260618 220824
rect 260562 211112 260618 211168
rect 267646 310936 267702 310992
rect 267646 310528 267702 310584
rect 269026 325660 269028 325680
rect 269028 325660 269080 325680
rect 269080 325660 269082 325680
rect 269026 325624 269082 325660
rect 269210 325488 269266 325544
rect 270866 337456 270922 337512
rect 270682 337048 270738 337104
rect 270774 336742 270830 336798
rect 270406 227840 270462 227896
rect 270774 269048 270830 269104
rect 270958 269084 270960 269104
rect 270960 269084 271012 269104
rect 271012 269084 271014 269104
rect 270958 269048 271014 269084
rect 270774 249736 270830 249792
rect 270958 249736 271014 249792
rect 270774 162832 270830 162888
rect 270774 162560 270830 162616
rect 270774 153176 270830 153232
rect 270958 153176 271014 153232
rect 272154 173848 272210 173904
rect 272154 164192 272210 164248
rect 272154 74432 272210 74488
rect 272154 64912 272210 64968
rect 272338 173848 272394 173904
rect 272338 164192 272394 164248
rect 272338 74432 272394 74488
rect 272430 64912 272486 64968
rect 275190 337728 275246 337784
rect 275282 314744 275338 314800
rect 275374 229064 275430 229120
rect 275558 229064 275614 229120
rect 275834 325760 275890 325816
rect 278686 337456 278742 337512
rect 279238 337728 279294 337784
rect 278042 306312 278098 306368
rect 278318 306312 278374 306368
rect 277950 295296 278006 295352
rect 278042 277344 278098 277400
rect 278226 295296 278282 295352
rect 278318 277208 278374 277264
rect 277858 238720 277914 238776
rect 278042 238740 278098 238776
rect 278042 238720 278044 238740
rect 278044 238720 278096 238740
rect 278096 238720 278098 238740
rect 277766 229064 277822 229120
rect 277950 229064 278006 229120
rect 278042 202816 278098 202872
rect 278226 202816 278282 202872
rect 277766 180784 277822 180840
rect 277950 180784 278006 180840
rect 278134 96600 278190 96656
rect 278318 96600 278374 96656
rect 277582 3984 277638 4040
rect 277858 3848 277914 3904
rect 278226 3712 278282 3768
rect 280250 76084 280306 76120
rect 280250 76064 280252 76084
rect 280252 76064 280304 76084
rect 280304 76064 280306 76084
rect 279882 3576 279938 3632
rect 279974 3440 280030 3496
rect 279790 3304 279846 3360
rect 283010 328480 283066 328536
rect 283378 328344 283434 328400
rect 285034 321680 285090 321736
rect 285034 321408 285090 321464
rect 288346 310700 288348 310720
rect 288348 310700 288400 310720
rect 288400 310700 288402 310720
rect 288346 310664 288402 310700
rect 288070 278704 288126 278760
rect 288254 278704 288310 278760
rect 289634 321408 289690 321464
rect 289726 75928 289782 75984
rect 296626 310800 296682 310856
rect 298006 321716 298008 321736
rect 298008 321716 298060 321736
rect 298060 321716 298062 321736
rect 298006 321680 298062 321716
rect 299570 310820 299626 310856
rect 299570 310800 299572 310820
rect 299572 310800 299624 310820
rect 299624 310800 299626 310820
rect 302146 227860 302202 227896
rect 302146 227840 302148 227860
rect 302148 227840 302200 227860
rect 302200 227840 302202 227860
rect 302146 76084 302202 76120
rect 302146 76064 302148 76084
rect 302148 76064 302200 76084
rect 302200 76064 302202 76084
rect 302146 29164 302202 29200
rect 302146 29144 302148 29164
rect 302148 29144 302200 29164
rect 302200 29144 302202 29164
rect 304354 310820 304410 310856
rect 304354 310800 304356 310820
rect 304356 310800 304408 310820
rect 304408 310800 304410 310820
rect 312542 340040 312598 340096
rect 309782 338680 309838 338736
rect 309046 322088 309102 322144
rect 309046 321816 309102 321872
rect 309046 227704 309102 227760
rect 309046 75928 309102 75984
rect 309046 29008 309102 29064
rect 315302 338816 315358 338872
rect 320730 310664 320786 310720
rect 321650 321816 321706 321872
rect 321466 321680 321522 321736
rect 321466 227876 321468 227896
rect 321468 227876 321520 227896
rect 321520 227876 321522 227896
rect 321466 227840 321522 227876
rect 321466 76100 321468 76120
rect 321468 76100 321520 76120
rect 321520 76100 321522 76120
rect 321466 76064 321522 76100
rect 321466 29180 321468 29200
rect 321468 29180 321520 29200
rect 321520 29180 321522 29200
rect 321466 29144 321522 29180
rect 321650 29180 321652 29200
rect 321652 29180 321704 29200
rect 321704 29180 321706 29200
rect 321650 29144 321706 29180
rect 323030 227876 323032 227896
rect 323032 227876 323084 227896
rect 323084 227876 323086 227896
rect 323030 227840 323086 227876
rect 323030 76100 323032 76120
rect 323032 76100 323084 76120
rect 323084 76100 323086 76120
rect 323030 76064 323086 76100
rect 328366 310820 328422 310856
rect 328366 310800 328368 310820
rect 328368 310800 328420 310820
rect 328420 310800 328422 310820
rect 340970 321816 341026 321872
rect 340786 321680 340842 321736
rect 340786 310700 340788 310720
rect 340788 310700 340840 310720
rect 340840 310700 340842 310720
rect 340786 310664 340842 310700
rect 347686 310800 347742 310856
rect 359646 310664 359702 310720
rect 362222 322088 362278 322144
rect 362222 321816 362278 321872
rect 367006 310820 367062 310856
rect 367006 310800 367008 310820
rect 367008 310800 367060 310820
rect 367060 310800 367062 310820
rect 379426 321716 379428 321736
rect 379428 321716 379480 321736
rect 379480 321716 379482 321736
rect 379426 321680 379482 321716
rect 379426 310700 379428 310720
rect 379428 310700 379480 310720
rect 379480 310700 379482 310720
rect 379426 310664 379482 310700
rect 386326 321816 386382 321872
rect 386326 310800 386382 310856
rect 398746 310700 398748 310720
rect 398748 310700 398800 310720
rect 398800 310700 398802 310720
rect 398746 310664 398802 310700
rect 400862 322088 400918 322144
rect 400862 321816 400918 321872
rect 405646 310800 405702 310856
rect 415306 227840 415362 227896
rect 415306 227704 415362 227760
rect 415306 76064 415362 76120
rect 415306 75928 415362 75984
rect 415122 29144 415178 29200
rect 415306 29008 415362 29064
rect 418250 321816 418306 321872
rect 418066 321680 418122 321736
rect 418066 310700 418068 310720
rect 418068 310700 418120 310720
rect 418120 310700 418122 310720
rect 418066 310664 418122 310700
rect 424966 310800 425022 310856
rect 437570 321816 437626 321872
rect 437386 321680 437442 321736
rect 437386 310700 437388 310720
rect 437388 310700 437440 310720
rect 437440 310700 437442 310720
rect 437386 310664 437442 310700
rect 437386 227860 437442 227896
rect 437386 227840 437388 227860
rect 437388 227840 437440 227860
rect 437440 227840 437442 227860
rect 437386 76084 437442 76120
rect 437386 76064 437388 76084
rect 437388 76064 437440 76084
rect 437440 76064 437442 76084
rect 437386 29164 437442 29200
rect 437386 29144 437388 29164
rect 437388 29144 437440 29164
rect 437440 29144 437442 29164
rect 444286 310800 444342 310856
rect 444286 227704 444342 227760
rect 444286 75928 444342 75984
rect 444286 29008 444342 29064
rect 456890 321816 456946 321872
rect 456706 321680 456762 321736
rect 456706 310700 456708 310720
rect 456708 310700 456760 310720
rect 456760 310700 456762 310720
rect 456706 310664 456762 310700
rect 456706 227840 456762 227896
rect 456890 227840 456946 227896
rect 456706 76064 456762 76120
rect 456890 76064 456946 76120
rect 456706 29144 456762 29200
rect 456890 29144 456946 29200
rect 463606 310800 463662 310856
rect 464434 3984 464490 4040
rect 467930 3848 467986 3904
rect 471518 3712 471574 3768
rect 476210 321816 476266 321872
rect 476026 321680 476082 321736
rect 475566 310664 475622 310720
rect 475106 3576 475162 3632
rect 476026 227860 476082 227896
rect 476026 227840 476028 227860
rect 476028 227840 476080 227860
rect 476080 227840 476082 227860
rect 478694 3440 478750 3496
rect 482926 310820 482982 310856
rect 482926 310800 482928 310820
rect 482928 310800 482980 310820
rect 482980 310800 482982 310820
rect 482926 227704 482982 227760
rect 482926 76064 482982 76120
rect 482926 75928 482982 75984
rect 482282 3304 482338 3360
rect 495346 321816 495402 321872
rect 495530 321816 495586 321872
rect 491206 29144 491262 29200
rect 491206 28736 491262 28792
rect 495346 310700 495348 310720
rect 495348 310700 495400 310720
rect 495400 310700 495402 310720
rect 495346 310664 495402 310700
rect 579802 392944 579858 393000
rect 580170 369552 580226 369608
rect 580078 357856 580134 357912
rect 579802 346024 579858 346080
rect 497462 29416 497518 29472
rect 497462 29008 497518 29064
rect 502246 310800 502302 310856
rect 502246 75792 502302 75848
rect 514666 321816 514722 321872
rect 514850 321816 514906 321872
rect 514666 310700 514668 310720
rect 514668 310700 514720 310720
rect 514720 310700 514722 310720
rect 514666 310664 514722 310700
rect 510526 76200 510582 76256
rect 514666 29164 514722 29200
rect 514666 29144 514668 29164
rect 514668 29144 514720 29164
rect 514720 29144 514722 29164
rect 521566 310800 521622 310856
rect 521566 76472 521622 76528
rect 521566 75928 521622 75984
rect 521566 29008 521622 29064
rect 533986 321816 534042 321872
rect 534170 321816 534226 321872
rect 533986 310700 533988 310720
rect 533988 310700 534040 310720
rect 534040 310700 534042 310720
rect 533986 310664 534042 310700
rect 533986 227860 534042 227896
rect 533986 227840 533988 227860
rect 533988 227840 534040 227860
rect 534040 227840 534042 227860
rect 533986 76084 534042 76120
rect 533986 76064 533988 76084
rect 533988 76064 534040 76084
rect 534040 76064 534042 76084
rect 533986 29164 534042 29200
rect 533986 29144 533988 29164
rect 533988 29144 534040 29164
rect 534040 29144 534042 29164
rect 540886 310800 540942 310856
rect 540886 227704 540942 227760
rect 540886 75928 540942 75984
rect 540886 29008 540942 29064
rect 541070 310820 541126 310856
rect 541070 310800 541072 310820
rect 541072 310800 541124 310820
rect 541124 310800 541126 310820
rect 543830 310528 543886 310584
rect 553306 227860 553362 227896
rect 553306 227840 553308 227860
rect 553308 227840 553360 227860
rect 553360 227840 553362 227860
rect 553306 76084 553362 76120
rect 553306 76064 553308 76084
rect 553308 76064 553360 76084
rect 553360 76064 553362 76084
rect 553306 29164 553362 29200
rect 553306 29144 553308 29164
rect 553308 29144 553360 29164
rect 553360 29144 553362 29164
rect 555422 310528 555478 310584
rect 555422 310256 555478 310312
rect 560206 227704 560262 227760
rect 560206 75928 560262 75984
rect 560206 29008 560262 29064
rect 562874 321680 562930 321736
rect 563150 321680 563206 321736
rect 572626 321816 572682 321872
rect 572718 321680 572774 321736
rect 572626 227860 572682 227896
rect 572626 227840 572628 227860
rect 572628 227840 572680 227860
rect 572680 227840 572682 227860
rect 572626 76084 572682 76120
rect 572626 76064 572628 76084
rect 572628 76064 572680 76084
rect 572680 76064 572682 76084
rect 572626 29164 572682 29200
rect 572626 29144 572628 29164
rect 572628 29144 572680 29164
rect 572680 29144 572682 29164
rect 579802 299104 579858 299160
rect 580170 275712 580226 275768
rect 580170 263880 580226 263936
rect 579802 252184 579858 252240
rect 579526 227704 579582 227760
rect 580170 216960 580226 217016
rect 579802 205264 579858 205320
rect 580170 181872 580226 181928
rect 580170 170040 580226 170096
rect 579802 158344 579858 158400
rect 580170 134816 580226 134872
rect 580170 123120 580226 123176
rect 579802 111424 579858 111480
rect 580170 87896 580226 87952
rect 579526 75928 579582 75984
rect 579802 64504 579858 64560
rect 580170 40976 580226 41032
rect 579526 29008 579582 29064
rect 579802 17584 579858 17640
<< metal3 >>
rect 580165 698050 580231 698053
rect 583520 698050 584960 698140
rect 580165 698048 584960 698050
rect 580165 697992 580170 698048
rect 580226 697992 584960 698048
rect 580165 697990 584960 697992
rect 580165 697987 580231 697990
rect 583520 697900 584960 697990
rect -960 696540 480 696780
rect 218881 695738 218947 695741
rect 218881 695736 219450 695738
rect 218881 695680 218886 695736
rect 218942 695680 219450 695736
rect 218881 695678 219450 695680
rect 218881 695675 218947 695678
rect 219249 695602 219315 695605
rect 219390 695602 219450 695678
rect 219249 695600 219450 695602
rect 219249 695544 219254 695600
rect 219310 695544 219450 695600
rect 219249 695542 219450 695544
rect 219249 695539 219315 695542
rect 580165 686354 580231 686357
rect 583520 686354 584960 686444
rect 580165 686352 584960 686354
rect 580165 686296 580170 686352
rect 580226 686296 584960 686352
rect 580165 686294 584960 686296
rect 580165 686291 580231 686294
rect 583520 686204 584960 686294
rect -960 682274 480 682364
rect 3417 682274 3483 682277
rect -960 682272 3483 682274
rect -960 682216 3422 682272
rect 3478 682216 3483 682272
rect -960 682214 3483 682216
rect -960 682124 480 682214
rect 3417 682211 3483 682214
rect 580165 674658 580231 674661
rect 583520 674658 584960 674748
rect 580165 674656 584960 674658
rect 580165 674600 580170 674656
rect 580226 674600 584960 674656
rect 580165 674598 584960 674600
rect 580165 674595 580231 674598
rect 583520 674508 584960 674598
rect -960 667994 480 668084
rect 3509 667994 3575 667997
rect -960 667992 3575 667994
rect -960 667936 3514 667992
rect 3570 667936 3575 667992
rect -960 667934 3575 667936
rect -960 667844 480 667934
rect 3509 667931 3575 667934
rect 583520 662676 584960 662916
rect -960 653578 480 653668
rect 3325 653578 3391 653581
rect -960 653576 3391 653578
rect -960 653520 3330 653576
rect 3386 653520 3391 653576
rect -960 653518 3391 653520
rect -960 653428 480 653518
rect 3325 653515 3391 653518
rect 580165 651130 580231 651133
rect 583520 651130 584960 651220
rect 580165 651128 584960 651130
rect 580165 651072 580170 651128
rect 580226 651072 584960 651128
rect 580165 651070 584960 651072
rect 580165 651067 580231 651070
rect 583520 650980 584960 651070
rect 580165 639434 580231 639437
rect 583520 639434 584960 639524
rect 580165 639432 584960 639434
rect 580165 639376 580170 639432
rect 580226 639376 584960 639432
rect 580165 639374 584960 639376
rect 580165 639371 580231 639374
rect 583520 639284 584960 639374
rect -960 639012 480 639252
rect 580165 627738 580231 627741
rect 583520 627738 584960 627828
rect 580165 627736 584960 627738
rect 580165 627680 580170 627736
rect 580226 627680 584960 627736
rect 580165 627678 584960 627680
rect 580165 627675 580231 627678
rect 583520 627588 584960 627678
rect -960 624882 480 624972
rect 3601 624882 3667 624885
rect -960 624880 3667 624882
rect -960 624824 3606 624880
rect 3662 624824 3667 624880
rect -960 624822 3667 624824
rect -960 624732 480 624822
rect 3601 624819 3667 624822
rect 583520 615756 584960 615996
rect -960 610466 480 610556
rect 3693 610466 3759 610469
rect -960 610464 3759 610466
rect -960 610408 3698 610464
rect 3754 610408 3759 610464
rect -960 610406 3759 610408
rect -960 610316 480 610406
rect 3693 610403 3759 610406
rect 580165 604210 580231 604213
rect 583520 604210 584960 604300
rect 580165 604208 584960 604210
rect 580165 604152 580170 604208
rect 580226 604152 584960 604208
rect 580165 604150 584960 604152
rect 580165 604147 580231 604150
rect 583520 604060 584960 604150
rect -960 596050 480 596140
rect 3049 596050 3115 596053
rect -960 596048 3115 596050
rect -960 595992 3054 596048
rect 3110 595992 3115 596048
rect -960 595990 3115 595992
rect -960 595900 480 595990
rect 3049 595987 3115 595990
rect 580165 592514 580231 592517
rect 583520 592514 584960 592604
rect 580165 592512 584960 592514
rect 580165 592456 580170 592512
rect 580226 592456 584960 592512
rect 580165 592454 584960 592456
rect 580165 592451 580231 592454
rect 583520 592364 584960 592454
rect -960 581620 480 581860
rect 580165 580818 580231 580821
rect 583520 580818 584960 580908
rect 580165 580816 584960 580818
rect 580165 580760 580170 580816
rect 580226 580760 584960 580816
rect 580165 580758 584960 580760
rect 580165 580755 580231 580758
rect 583520 580668 584960 580758
rect 583520 568836 584960 569076
rect -960 567354 480 567444
rect 3877 567354 3943 567357
rect -960 567352 3943 567354
rect -960 567296 3882 567352
rect 3938 567296 3943 567352
rect -960 567294 3943 567296
rect -960 567204 480 567294
rect 3877 567291 3943 567294
rect 299565 560554 299631 560557
rect 299430 560552 299631 560554
rect 299430 560496 299570 560552
rect 299626 560496 299631 560552
rect 299430 560494 299631 560496
rect 299430 560418 299490 560494
rect 299565 560491 299631 560494
rect 299565 560418 299631 560421
rect 299430 560416 299631 560418
rect 299430 560360 299570 560416
rect 299626 560360 299631 560416
rect 299430 560358 299631 560360
rect 299565 560355 299631 560358
rect 580165 557290 580231 557293
rect 583520 557290 584960 557380
rect 580165 557288 584960 557290
rect 580165 557232 580170 557288
rect 580226 557232 584960 557288
rect 580165 557230 584960 557232
rect 580165 557227 580231 557230
rect 583520 557140 584960 557230
rect -960 553074 480 553164
rect 2957 553074 3023 553077
rect -960 553072 3023 553074
rect -960 553016 2962 553072
rect 3018 553016 3023 553072
rect -960 553014 3023 553016
rect -960 552924 480 553014
rect 2957 553011 3023 553014
rect 299289 549266 299355 549269
rect 299473 549266 299539 549269
rect 299289 549264 299539 549266
rect 299289 549208 299294 549264
rect 299350 549208 299478 549264
rect 299534 549208 299539 549264
rect 299289 549206 299539 549208
rect 299289 549203 299355 549206
rect 299473 549203 299539 549206
rect 580165 545594 580231 545597
rect 583520 545594 584960 545684
rect 580165 545592 584960 545594
rect 580165 545536 580170 545592
rect 580226 545536 584960 545592
rect 580165 545534 584960 545536
rect 580165 545531 580231 545534
rect 583520 545444 584960 545534
rect 218973 540970 219039 540973
rect 219157 540970 219223 540973
rect 218973 540968 219223 540970
rect 218973 540912 218978 540968
rect 219034 540912 219162 540968
rect 219218 540912 219223 540968
rect 218973 540910 219223 540912
rect 218973 540907 219039 540910
rect 219157 540907 219223 540910
rect -960 538658 480 538748
rect 3141 538658 3207 538661
rect -960 538656 3207 538658
rect -960 538600 3146 538656
rect 3202 538600 3207 538656
rect -960 538598 3207 538600
rect -960 538508 480 538598
rect 3141 538595 3207 538598
rect 580165 533898 580231 533901
rect 583520 533898 584960 533988
rect 580165 533896 584960 533898
rect 580165 533840 580170 533896
rect 580226 533840 584960 533896
rect 580165 533838 584960 533840
rect 580165 533835 580231 533838
rect 583520 533748 584960 533838
rect 218973 531314 219039 531317
rect 219157 531314 219223 531317
rect 218973 531312 219223 531314
rect 218973 531256 218978 531312
rect 219034 531256 219162 531312
rect 219218 531256 219223 531312
rect 218973 531254 219223 531256
rect 218973 531251 219039 531254
rect 219157 531251 219223 531254
rect -960 524092 480 524332
rect 583520 521916 584960 522156
rect 218789 521658 218855 521661
rect 218973 521658 219039 521661
rect 218789 521656 219039 521658
rect 218789 521600 218794 521656
rect 218850 521600 218978 521656
rect 219034 521600 219039 521656
rect 218789 521598 219039 521600
rect 218789 521595 218855 521598
rect 218973 521595 219039 521598
rect 299657 521658 299723 521661
rect 299841 521658 299907 521661
rect 299657 521656 299907 521658
rect 299657 521600 299662 521656
rect 299718 521600 299846 521656
rect 299902 521600 299907 521656
rect 299657 521598 299907 521600
rect 299657 521595 299723 521598
rect 299841 521595 299907 521598
rect 580165 510370 580231 510373
rect 583520 510370 584960 510460
rect 580165 510368 584960 510370
rect 580165 510312 580170 510368
rect 580226 510312 584960 510368
rect 580165 510310 584960 510312
rect 580165 510307 580231 510310
rect 583520 510220 584960 510310
rect -960 509962 480 510052
rect 4061 509962 4127 509965
rect -960 509960 4127 509962
rect -960 509904 4066 509960
rect 4122 509904 4127 509960
rect -960 509902 4127 509904
rect -960 509812 480 509902
rect 4061 509899 4127 509902
rect 299473 502346 299539 502349
rect 299749 502346 299815 502349
rect 299473 502344 299815 502346
rect 299473 502288 299478 502344
rect 299534 502288 299754 502344
rect 299810 502288 299815 502344
rect 299473 502286 299815 502288
rect 299473 502283 299539 502286
rect 299749 502283 299815 502286
rect 580165 498674 580231 498677
rect 583520 498674 584960 498764
rect 580165 498672 584960 498674
rect 580165 498616 580170 498672
rect 580226 498616 584960 498672
rect 580165 498614 584960 498616
rect 580165 498611 580231 498614
rect 583520 498524 584960 498614
rect -960 495546 480 495636
rect 3325 495546 3391 495549
rect -960 495544 3391 495546
rect -960 495488 3330 495544
rect 3386 495488 3391 495544
rect -960 495486 3391 495488
rect -960 495396 480 495486
rect 3325 495483 3391 495486
rect 299473 492690 299539 492693
rect 299657 492690 299723 492693
rect 299473 492688 299723 492690
rect 299473 492632 299478 492688
rect 299534 492632 299662 492688
rect 299718 492632 299723 492688
rect 299473 492630 299723 492632
rect 299473 492627 299539 492630
rect 299657 492627 299723 492630
rect 580165 486842 580231 486845
rect 583520 486842 584960 486932
rect 580165 486840 584960 486842
rect 580165 486784 580170 486840
rect 580226 486784 584960 486840
rect 580165 486782 584960 486784
rect 580165 486779 580231 486782
rect 583520 486692 584960 486782
rect 154205 483034 154271 483037
rect 154481 483034 154547 483037
rect 154205 483032 154547 483034
rect 154205 482976 154210 483032
rect 154266 482976 154486 483032
rect 154542 482976 154547 483032
rect 154205 482974 154547 482976
rect 154205 482971 154271 482974
rect 154481 482971 154547 482974
rect -960 481130 480 481220
rect 3141 481130 3207 481133
rect -960 481128 3207 481130
rect -960 481072 3146 481128
rect 3202 481072 3207 481128
rect -960 481070 3207 481072
rect -960 480980 480 481070
rect 3141 481067 3207 481070
rect 583520 474996 584960 475236
rect 218973 473378 219039 473381
rect 219249 473378 219315 473381
rect 218973 473376 219315 473378
rect 218973 473320 218978 473376
rect 219034 473320 219254 473376
rect 219310 473320 219315 473376
rect 218973 473318 219315 473320
rect 218973 473315 219039 473318
rect 219249 473315 219315 473318
rect -960 466700 480 466940
rect 580165 463450 580231 463453
rect 583520 463450 584960 463540
rect 580165 463448 584960 463450
rect 580165 463392 580170 463448
rect 580226 463392 584960 463448
rect 580165 463390 584960 463392
rect 580165 463387 580231 463390
rect 583520 463300 584960 463390
rect -960 452434 480 452524
rect 3233 452434 3299 452437
rect -960 452432 3299 452434
rect -960 452376 3238 452432
rect 3294 452376 3299 452432
rect -960 452374 3299 452376
rect -960 452284 480 452374
rect 3233 452371 3299 452374
rect 580165 451754 580231 451757
rect 583520 451754 584960 451844
rect 580165 451752 584960 451754
rect 580165 451696 580170 451752
rect 580226 451696 584960 451752
rect 580165 451694 584960 451696
rect 580165 451691 580231 451694
rect 583520 451604 584960 451694
rect 580165 439922 580231 439925
rect 583520 439922 584960 440012
rect 580165 439920 584960 439922
rect 580165 439864 580170 439920
rect 580226 439864 584960 439920
rect 580165 439862 584960 439864
rect 580165 439859 580231 439862
rect 583520 439772 584960 439862
rect -960 438018 480 438108
rect 2957 438018 3023 438021
rect -960 438016 3023 438018
rect -960 437960 2962 438016
rect 3018 437960 3023 438016
rect -960 437958 3023 437960
rect -960 437868 480 437958
rect 2957 437955 3023 437958
rect 583520 428076 584960 428316
rect 218973 425098 219039 425101
rect 219341 425098 219407 425101
rect 218973 425096 219407 425098
rect 218973 425040 218978 425096
rect 219034 425040 219346 425096
rect 219402 425040 219407 425096
rect 218973 425038 219407 425040
rect 218973 425035 219039 425038
rect 219341 425035 219407 425038
rect -960 423738 480 423828
rect 3325 423738 3391 423741
rect -960 423736 3391 423738
rect -960 423680 3330 423736
rect 3386 423680 3391 423736
rect -960 423678 3391 423680
rect -960 423588 480 423678
rect 3325 423675 3391 423678
rect 580165 416530 580231 416533
rect 583520 416530 584960 416620
rect 580165 416528 584960 416530
rect 580165 416472 580170 416528
rect 580226 416472 584960 416528
rect 580165 416470 584960 416472
rect 580165 416467 580231 416470
rect 583520 416380 584960 416470
rect 154113 415442 154179 415445
rect 154297 415442 154363 415445
rect 154113 415440 154363 415442
rect 154113 415384 154118 415440
rect 154174 415384 154302 415440
rect 154358 415384 154363 415440
rect 154113 415382 154363 415384
rect 154113 415379 154179 415382
rect 154297 415379 154363 415382
rect 154297 415306 154363 415309
rect 154481 415306 154547 415309
rect 154297 415304 154547 415306
rect 154297 415248 154302 415304
rect 154358 415248 154486 415304
rect 154542 415248 154547 415304
rect 154297 415246 154547 415248
rect 154297 415243 154363 415246
rect 154481 415243 154547 415246
rect -960 409172 480 409412
rect 580165 404834 580231 404837
rect 583520 404834 584960 404924
rect 580165 404832 584960 404834
rect 580165 404776 580170 404832
rect 580226 404776 584960 404832
rect 580165 404774 584960 404776
rect 580165 404771 580231 404774
rect 583520 404684 584960 404774
rect 235809 401978 235875 401981
rect 485037 401978 485103 401981
rect 235809 401976 485103 401978
rect 235809 401920 235814 401976
rect 235870 401920 485042 401976
rect 485098 401920 485103 401976
rect 235809 401918 485103 401920
rect 235809 401915 235875 401918
rect 485037 401915 485103 401918
rect 262806 401780 262812 401844
rect 262876 401842 262882 401844
rect 289629 401842 289695 401845
rect 262876 401840 289695 401842
rect 262876 401784 289634 401840
rect 289690 401784 289695 401840
rect 262876 401782 289695 401784
rect 262876 401780 262882 401782
rect 289629 401779 289695 401782
rect 240317 399530 240383 399533
rect 243486 399530 243492 399532
rect 240317 399528 243492 399530
rect 240317 399472 240322 399528
rect 240378 399472 243492 399528
rect 240317 399470 243492 399472
rect 240317 399467 240383 399470
rect 243486 399468 243492 399470
rect 243556 399468 243562 399532
rect 231577 399394 231643 399397
rect 232957 399396 233023 399397
rect 231710 399394 231716 399396
rect 231577 399392 231716 399394
rect 231577 399336 231582 399392
rect 231638 399336 231716 399392
rect 231577 399334 231716 399336
rect 231577 399331 231643 399334
rect 231710 399332 231716 399334
rect 231780 399332 231786 399396
rect 232957 399392 233004 399396
rect 233068 399394 233074 399396
rect 232957 399336 232962 399392
rect 232957 399332 233004 399336
rect 233068 399334 233114 399394
rect 233068 399332 233074 399334
rect 233918 399332 233924 399396
rect 233988 399394 233994 399396
rect 234061 399394 234127 399397
rect 233988 399392 234127 399394
rect 233988 399336 234066 399392
rect 234122 399336 234127 399392
rect 233988 399334 234127 399336
rect 233988 399332 233994 399334
rect 232957 399331 233023 399332
rect 234061 399331 234127 399334
rect 237189 399396 237255 399397
rect 237189 399392 237236 399396
rect 237300 399394 237306 399396
rect 237833 399394 237899 399397
rect 238150 399394 238156 399396
rect 237189 399336 237194 399392
rect 237189 399332 237236 399336
rect 237300 399334 237346 399394
rect 237833 399392 238156 399394
rect 237833 399336 237838 399392
rect 237894 399336 238156 399392
rect 237833 399334 238156 399336
rect 237300 399332 237306 399334
rect 237189 399331 237255 399332
rect 237833 399331 237899 399334
rect 238150 399332 238156 399334
rect 238220 399332 238226 399396
rect 239397 399394 239463 399397
rect 239990 399394 239996 399396
rect 239397 399392 239996 399394
rect 239397 399336 239402 399392
rect 239458 399336 239996 399392
rect 239397 399334 239996 399336
rect 239397 399331 239463 399334
rect 239990 399332 239996 399334
rect 240060 399332 240066 399396
rect 240961 399394 241027 399397
rect 241278 399394 241284 399396
rect 240961 399392 241284 399394
rect 240961 399336 240966 399392
rect 241022 399336 241284 399392
rect 240961 399334 241284 399336
rect 240961 399331 241027 399334
rect 241278 399332 241284 399334
rect 241348 399332 241354 399396
rect 282862 399332 282868 399396
rect 282932 399394 282938 399396
rect 283005 399394 283071 399397
rect 282932 399392 283071 399394
rect 282932 399336 283010 399392
rect 283066 399336 283071 399392
rect 282932 399334 283071 399336
rect 282932 399332 282938 399334
rect 283005 399331 283071 399334
rect 284334 399332 284340 399396
rect 284404 399394 284410 399396
rect 284477 399394 284543 399397
rect 284404 399392 284543 399394
rect 284404 399336 284482 399392
rect 284538 399336 284543 399392
rect 284404 399334 284543 399336
rect 284404 399332 284410 399334
rect 284477 399331 284543 399334
rect 285622 399332 285628 399396
rect 285692 399394 285698 399396
rect 286133 399394 286199 399397
rect 285692 399392 286199 399394
rect 285692 399336 286138 399392
rect 286194 399336 286199 399392
rect 285692 399334 286199 399336
rect 285692 399332 285698 399334
rect 286133 399331 286199 399334
rect 287094 399332 287100 399396
rect 287164 399394 287170 399396
rect 287789 399394 287855 399397
rect 287164 399392 287855 399394
rect 287164 399336 287794 399392
rect 287850 399336 287855 399392
rect 287164 399334 287855 399336
rect 287164 399332 287170 399334
rect 287789 399331 287855 399334
rect -960 395042 480 395132
rect 3141 395042 3207 395045
rect -960 395040 3207 395042
rect -960 394984 3146 395040
rect 3202 394984 3207 395040
rect -960 394982 3207 394984
rect -960 394892 480 394982
rect 3141 394979 3207 394982
rect 579797 393002 579863 393005
rect 583520 393002 584960 393092
rect 579797 393000 584960 393002
rect 579797 392944 579802 393000
rect 579858 392944 584960 393000
rect 579797 392942 584960 392944
rect 579797 392939 579863 392942
rect 583520 392852 584960 392942
rect 583520 381156 584960 381396
rect -960 380626 480 380716
rect 3417 380626 3483 380629
rect -960 380624 3483 380626
rect -960 380568 3422 380624
rect 3478 380568 3483 380624
rect -960 380566 3483 380568
rect -960 380476 480 380566
rect 3417 380563 3483 380566
rect 580165 369610 580231 369613
rect 583520 369610 584960 369700
rect 580165 369608 584960 369610
rect 580165 369552 580170 369608
rect 580226 369552 584960 369608
rect 580165 369550 584960 369552
rect 580165 369547 580231 369550
rect 583520 369460 584960 369550
rect -960 366210 480 366300
rect 2957 366210 3023 366213
rect -960 366208 3023 366210
rect -960 366152 2962 366208
rect 3018 366152 3023 366208
rect -960 366150 3023 366152
rect -960 366060 480 366150
rect 2957 366147 3023 366150
rect 580073 357914 580139 357917
rect 583520 357914 584960 358004
rect 580073 357912 584960 357914
rect 580073 357856 580078 357912
rect 580134 357856 584960 357912
rect 580073 357854 584960 357856
rect 580073 357851 580139 357854
rect 583520 357764 584960 357854
rect -960 351780 480 352020
rect 579797 346082 579863 346085
rect 583520 346082 584960 346172
rect 579797 346080 584960 346082
rect 579797 346024 579802 346080
rect 579858 346024 584960 346080
rect 579797 346022 584960 346024
rect 579797 346019 579863 346022
rect 583520 345932 584960 346022
rect 238150 340036 238156 340100
rect 238220 340098 238226 340100
rect 312537 340098 312603 340101
rect 238220 340096 312603 340098
rect 238220 340040 312542 340096
rect 312598 340040 312603 340096
rect 238220 340038 312603 340040
rect 238220 340036 238226 340038
rect 312537 340035 312603 340038
rect 239990 338812 239996 338876
rect 240060 338874 240066 338876
rect 315297 338874 315363 338877
rect 240060 338872 315363 338874
rect 240060 338816 315302 338872
rect 315358 338816 315363 338872
rect 240060 338814 315363 338816
rect 240060 338812 240066 338814
rect 315297 338811 315363 338814
rect 233918 338676 233924 338740
rect 233988 338738 233994 338740
rect 309777 338738 309843 338741
rect 233988 338736 309843 338738
rect 233988 338680 309782 338736
rect 309838 338680 309843 338736
rect 233988 338678 309843 338680
rect 233988 338676 233994 338678
rect 309777 338675 309843 338678
rect 275185 337786 275251 337789
rect 279233 337786 279299 337789
rect 275185 337784 279299 337786
rect 275185 337728 275190 337784
rect 275246 337728 279238 337784
rect 279294 337728 279299 337784
rect 275185 337726 279299 337728
rect 275185 337723 275251 337726
rect 279233 337723 279299 337726
rect -960 337514 480 337604
rect 3417 337514 3483 337517
rect -960 337512 3483 337514
rect -960 337456 3422 337512
rect 3478 337456 3483 337512
rect -960 337454 3483 337456
rect -960 337364 480 337454
rect 3417 337451 3483 337454
rect 270861 337514 270927 337517
rect 278681 337514 278747 337517
rect 270861 337512 278747 337514
rect 270861 337456 270866 337512
rect 270922 337456 278686 337512
rect 278742 337456 278747 337512
rect 270861 337454 278747 337456
rect 270861 337451 270927 337454
rect 278681 337451 278747 337454
rect 270677 337106 270743 337109
rect 270677 337104 270970 337106
rect 270677 337048 270682 337104
rect 270738 337048 270970 337104
rect 270677 337046 270970 337048
rect 270677 337043 270743 337046
rect 270769 336800 270835 336803
rect 270910 336800 270970 337046
rect 270769 336798 270970 336800
rect 270769 336742 270774 336798
rect 270830 336742 270970 336798
rect 270769 336740 270970 336742
rect 270769 336737 270835 336740
rect 3417 336018 3483 336021
rect 262806 336018 262812 336020
rect 3417 336016 262812 336018
rect 3417 335960 3422 336016
rect 3478 335960 262812 336016
rect 3417 335958 262812 335960
rect 3417 335955 3483 335958
rect 262806 335956 262812 335958
rect 262876 335956 262882 336020
rect 252001 335746 252067 335749
rect 251958 335744 252067 335746
rect 251958 335688 252006 335744
rect 252062 335688 252067 335744
rect 251958 335683 252067 335688
rect 251633 335474 251699 335477
rect 251958 335474 252018 335683
rect 251633 335472 252018 335474
rect 251633 335416 251638 335472
rect 251694 335416 252018 335472
rect 251633 335414 252018 335416
rect 254117 335474 254183 335477
rect 254577 335474 254643 335477
rect 254117 335472 254643 335474
rect 254117 335416 254122 335472
rect 254178 335416 254582 335472
rect 254638 335416 254643 335472
rect 254117 335414 254643 335416
rect 251633 335411 251699 335414
rect 254117 335411 254183 335414
rect 254577 335411 254643 335414
rect 583520 334236 584960 334476
rect 283005 328538 283071 328541
rect 283005 328536 283298 328538
rect 283005 328480 283010 328536
rect 283066 328480 283298 328536
rect 283005 328478 283298 328480
rect 283005 328475 283071 328478
rect 283238 328402 283298 328478
rect 283373 328402 283439 328405
rect 283238 328400 283439 328402
rect 283238 328344 283378 328400
rect 283434 328344 283439 328400
rect 283238 328342 283439 328344
rect 283373 328339 283439 328342
rect 275829 325818 275895 325821
rect 275326 325816 275895 325818
rect 275326 325760 275834 325816
rect 275890 325760 275895 325816
rect 275326 325758 275895 325760
rect 256417 325682 256483 325685
rect 256601 325682 256667 325685
rect 256417 325680 256667 325682
rect 256417 325624 256422 325680
rect 256478 325624 256606 325680
rect 256662 325624 256667 325680
rect 256417 325622 256667 325624
rect 256417 325619 256483 325622
rect 256601 325619 256667 325622
rect 269021 325682 269087 325685
rect 275326 325684 275386 325758
rect 275829 325755 275895 325758
rect 269021 325680 269130 325682
rect 269021 325624 269026 325680
rect 269082 325624 269130 325680
rect 269021 325619 269130 325624
rect 275318 325620 275324 325684
rect 275388 325620 275394 325684
rect 269070 325546 269130 325619
rect 269205 325546 269271 325549
rect 269070 325544 269271 325546
rect 269070 325488 269210 325544
rect 269266 325488 269271 325544
rect 269070 325486 269271 325488
rect 269205 325483 269271 325486
rect -960 323098 480 323188
rect 3325 323098 3391 323101
rect -960 323096 3391 323098
rect -960 323040 3330 323096
rect 3386 323040 3391 323096
rect -960 323038 3391 323040
rect -960 322948 480 323038
rect 3325 323035 3391 323038
rect 583520 322690 584960 322780
rect 583342 322630 584960 322690
rect 299422 322084 299428 322148
rect 299492 322146 299498 322148
rect 309041 322146 309107 322149
rect 299492 322144 309107 322146
rect 299492 322088 309046 322144
rect 309102 322088 309107 322144
rect 299492 322086 309107 322088
rect 299492 322084 299498 322086
rect 309041 322083 309107 322086
rect 357382 322084 357388 322148
rect 357452 322146 357458 322148
rect 362217 322146 362283 322149
rect 357452 322144 362283 322146
rect 357452 322088 362222 322144
rect 362278 322088 362283 322144
rect 357452 322086 362283 322088
rect 357452 322084 357458 322086
rect 362217 322083 362283 322086
rect 396022 322084 396028 322148
rect 396092 322146 396098 322148
rect 400857 322146 400923 322149
rect 396092 322144 400923 322146
rect 396092 322088 400862 322144
rect 400918 322088 400923 322144
rect 396092 322086 400923 322088
rect 396092 322084 396098 322086
rect 400857 322083 400923 322086
rect 309041 321874 309107 321877
rect 321645 321874 321711 321877
rect 340965 321874 341031 321877
rect 362217 321874 362283 321877
rect 386321 321874 386387 321877
rect 400857 321874 400923 321877
rect 418245 321874 418311 321877
rect 437565 321874 437631 321877
rect 456885 321874 456951 321877
rect 476205 321874 476271 321877
rect 495341 321874 495407 321877
rect 251038 321814 280170 321874
rect 243486 321540 243492 321604
rect 243556 321602 243562 321604
rect 251038 321602 251098 321814
rect 280110 321738 280170 321814
rect 309041 321872 312002 321874
rect 309041 321816 309046 321872
rect 309102 321816 312002 321872
rect 309041 321814 312002 321816
rect 309041 321811 309107 321814
rect 285029 321738 285095 321741
rect 280110 321736 285095 321738
rect 280110 321680 285034 321736
rect 285090 321680 285095 321736
rect 280110 321678 285095 321680
rect 285029 321675 285095 321678
rect 298001 321738 298067 321741
rect 299422 321738 299428 321740
rect 298001 321736 299428 321738
rect 298001 321680 298006 321736
rect 298062 321680 299428 321736
rect 298001 321678 299428 321680
rect 298001 321675 298067 321678
rect 299422 321676 299428 321678
rect 299492 321676 299498 321740
rect 311942 321738 312002 321814
rect 321645 321872 331322 321874
rect 321645 321816 321650 321872
rect 321706 321816 331322 321872
rect 321645 321814 331322 321816
rect 321645 321811 321711 321814
rect 321461 321738 321527 321741
rect 311942 321736 321527 321738
rect 311942 321680 321466 321736
rect 321522 321680 321527 321736
rect 311942 321678 321527 321680
rect 331262 321738 331322 321814
rect 340965 321872 350642 321874
rect 340965 321816 340970 321872
rect 341026 321816 350642 321872
rect 340965 321814 350642 321816
rect 340965 321811 341031 321814
rect 340781 321738 340847 321741
rect 331262 321736 340847 321738
rect 331262 321680 340786 321736
rect 340842 321680 340847 321736
rect 331262 321678 340847 321680
rect 350582 321738 350642 321814
rect 362217 321872 369962 321874
rect 362217 321816 362222 321872
rect 362278 321816 369962 321872
rect 362217 321814 369962 321816
rect 362217 321811 362283 321814
rect 357382 321738 357388 321740
rect 350582 321678 357388 321738
rect 321461 321675 321527 321678
rect 340781 321675 340847 321678
rect 357382 321676 357388 321678
rect 357452 321676 357458 321740
rect 369902 321738 369962 321814
rect 386321 321872 389282 321874
rect 386321 321816 386326 321872
rect 386382 321816 389282 321872
rect 386321 321814 389282 321816
rect 386321 321811 386387 321814
rect 379421 321738 379487 321741
rect 369902 321736 379487 321738
rect 369902 321680 379426 321736
rect 379482 321680 379487 321736
rect 369902 321678 379487 321680
rect 389222 321738 389282 321814
rect 400857 321872 408602 321874
rect 400857 321816 400862 321872
rect 400918 321816 408602 321872
rect 400857 321814 408602 321816
rect 400857 321811 400923 321814
rect 396022 321738 396028 321740
rect 389222 321678 396028 321738
rect 379421 321675 379487 321678
rect 396022 321676 396028 321678
rect 396092 321676 396098 321740
rect 408542 321738 408602 321814
rect 418245 321872 427922 321874
rect 418245 321816 418250 321872
rect 418306 321816 427922 321872
rect 418245 321814 427922 321816
rect 418245 321811 418311 321814
rect 418061 321738 418127 321741
rect 408542 321736 418127 321738
rect 408542 321680 418066 321736
rect 418122 321680 418127 321736
rect 408542 321678 418127 321680
rect 427862 321738 427922 321814
rect 437565 321872 447242 321874
rect 437565 321816 437570 321872
rect 437626 321816 447242 321872
rect 437565 321814 447242 321816
rect 437565 321811 437631 321814
rect 437381 321738 437447 321741
rect 427862 321736 437447 321738
rect 427862 321680 437386 321736
rect 437442 321680 437447 321736
rect 427862 321678 437447 321680
rect 447182 321738 447242 321814
rect 456885 321872 466562 321874
rect 456885 321816 456890 321872
rect 456946 321816 466562 321872
rect 456885 321814 466562 321816
rect 456885 321811 456951 321814
rect 456701 321738 456767 321741
rect 447182 321736 456767 321738
rect 447182 321680 456706 321736
rect 456762 321680 456767 321736
rect 447182 321678 456767 321680
rect 466502 321738 466562 321814
rect 476205 321872 485882 321874
rect 476205 321816 476210 321872
rect 476266 321816 485882 321872
rect 476205 321814 485882 321816
rect 476205 321811 476271 321814
rect 476021 321738 476087 321741
rect 466502 321736 476087 321738
rect 466502 321680 476026 321736
rect 476082 321680 476087 321736
rect 466502 321678 476087 321680
rect 485822 321738 485882 321814
rect 495022 321872 495407 321874
rect 495022 321816 495346 321872
rect 495402 321816 495407 321872
rect 495022 321814 495407 321816
rect 495022 321738 495082 321814
rect 495341 321811 495407 321814
rect 495525 321874 495591 321877
rect 514661 321874 514727 321877
rect 495525 321872 505202 321874
rect 495525 321816 495530 321872
rect 495586 321816 505202 321872
rect 495525 321814 505202 321816
rect 495525 321811 495591 321814
rect 485822 321678 495082 321738
rect 505142 321738 505202 321814
rect 514342 321872 514727 321874
rect 514342 321816 514666 321872
rect 514722 321816 514727 321872
rect 514342 321814 514727 321816
rect 514342 321738 514402 321814
rect 514661 321811 514727 321814
rect 514845 321874 514911 321877
rect 533981 321874 534047 321877
rect 514845 321872 524522 321874
rect 514845 321816 514850 321872
rect 514906 321816 524522 321872
rect 514845 321814 524522 321816
rect 514845 321811 514911 321814
rect 505142 321678 514402 321738
rect 524462 321738 524522 321814
rect 533662 321872 534047 321874
rect 533662 321816 533986 321872
rect 534042 321816 534047 321872
rect 533662 321814 534047 321816
rect 533662 321738 533722 321814
rect 533981 321811 534047 321814
rect 534165 321874 534231 321877
rect 572621 321874 572687 321877
rect 534165 321872 553410 321874
rect 534165 321816 534170 321872
rect 534226 321816 553410 321872
rect 534165 321814 553410 321816
rect 534165 321811 534231 321814
rect 524462 321678 533722 321738
rect 553350 321738 553410 321814
rect 569910 321872 572687 321874
rect 569910 321816 572626 321872
rect 572682 321816 572687 321872
rect 569910 321814 572687 321816
rect 562869 321738 562935 321741
rect 553350 321736 562935 321738
rect 553350 321680 562874 321736
rect 562930 321680 562935 321736
rect 553350 321678 562935 321680
rect 418061 321675 418127 321678
rect 437381 321675 437447 321678
rect 456701 321675 456767 321678
rect 476021 321675 476087 321678
rect 562869 321675 562935 321678
rect 563145 321738 563211 321741
rect 569910 321738 569970 321814
rect 572621 321811 572687 321814
rect 563145 321736 569970 321738
rect 563145 321680 563150 321736
rect 563206 321680 569970 321736
rect 563145 321678 569970 321680
rect 572713 321738 572779 321741
rect 583342 321738 583402 322630
rect 583520 322540 584960 322630
rect 572713 321736 583402 321738
rect 572713 321680 572718 321736
rect 572774 321680 583402 321736
rect 572713 321678 583402 321680
rect 563145 321675 563211 321678
rect 572713 321675 572779 321678
rect 243556 321542 251098 321602
rect 243556 321540 243562 321542
rect 285029 321466 285095 321469
rect 289629 321466 289695 321469
rect 285029 321464 289695 321466
rect 285029 321408 285034 321464
rect 285090 321408 289634 321464
rect 289690 321408 289695 321464
rect 285029 321406 289695 321408
rect 285029 321403 285095 321406
rect 289629 321403 289695 321406
rect 256417 316026 256483 316029
rect 256601 316026 256667 316029
rect 256417 316024 256667 316026
rect 256417 315968 256422 316024
rect 256478 315968 256606 316024
rect 256662 315968 256667 316024
rect 256417 315966 256667 315968
rect 256417 315963 256483 315966
rect 256601 315963 256667 315966
rect 275318 314938 275324 314940
rect 275280 314876 275324 314938
rect 275388 314876 275394 314940
rect 275280 314805 275340 314876
rect 275277 314800 275343 314805
rect 275277 314744 275282 314800
rect 275338 314744 275343 314800
rect 275277 314739 275343 314744
rect 241278 310932 241284 310996
rect 241348 310994 241354 310996
rect 257838 310994 257844 310996
rect 241348 310934 257844 310994
rect 241348 310932 241354 310934
rect 257838 310932 257844 310934
rect 257908 310932 257914 310996
rect 258022 310932 258028 310996
rect 258092 310994 258098 310996
rect 267641 310994 267707 310997
rect 258092 310992 267707 310994
rect 258092 310936 267646 310992
rect 267702 310936 267707 310992
rect 258092 310934 267707 310936
rect 258092 310932 258098 310934
rect 267641 310931 267707 310934
rect 296621 310858 296687 310861
rect 299565 310858 299631 310861
rect 296621 310856 299631 310858
rect 296621 310800 296626 310856
rect 296682 310800 299570 310856
rect 299626 310800 299631 310856
rect 296621 310798 299631 310800
rect 296621 310795 296687 310798
rect 299565 310795 299631 310798
rect 304349 310858 304415 310861
rect 328361 310858 328427 310861
rect 347681 310858 347747 310861
rect 367001 310858 367067 310861
rect 386321 310858 386387 310861
rect 405641 310858 405707 310861
rect 424961 310858 425027 310861
rect 444281 310858 444347 310861
rect 463601 310858 463667 310861
rect 482921 310858 482987 310861
rect 502241 310858 502307 310861
rect 521561 310858 521627 310861
rect 540881 310858 540947 310861
rect 541065 310858 541131 310861
rect 304349 310856 312002 310858
rect 304349 310800 304354 310856
rect 304410 310800 312002 310856
rect 304349 310798 312002 310800
rect 304349 310795 304415 310798
rect 257838 310660 257844 310724
rect 257908 310722 257914 310724
rect 258022 310722 258028 310724
rect 257908 310662 258028 310722
rect 257908 310660 257914 310662
rect 258022 310660 258028 310662
rect 258092 310660 258098 310724
rect 288341 310722 288407 310725
rect 278822 310720 288407 310722
rect 278822 310664 288346 310720
rect 288402 310664 288407 310720
rect 278822 310662 288407 310664
rect 311942 310722 312002 310798
rect 328361 310856 331322 310858
rect 328361 310800 328366 310856
rect 328422 310800 331322 310856
rect 328361 310798 331322 310800
rect 328361 310795 328427 310798
rect 320725 310722 320791 310725
rect 311942 310720 320791 310722
rect 311942 310664 320730 310720
rect 320786 310664 320791 310720
rect 311942 310662 320791 310664
rect 331262 310722 331322 310798
rect 347681 310856 350642 310858
rect 347681 310800 347686 310856
rect 347742 310800 350642 310856
rect 347681 310798 350642 310800
rect 347681 310795 347747 310798
rect 340781 310722 340847 310725
rect 331262 310720 340847 310722
rect 331262 310664 340786 310720
rect 340842 310664 340847 310720
rect 331262 310662 340847 310664
rect 350582 310722 350642 310798
rect 367001 310856 369962 310858
rect 367001 310800 367006 310856
rect 367062 310800 369962 310856
rect 367001 310798 369962 310800
rect 367001 310795 367067 310798
rect 359641 310722 359707 310725
rect 350582 310720 359707 310722
rect 350582 310664 359646 310720
rect 359702 310664 359707 310720
rect 350582 310662 359707 310664
rect 369902 310722 369962 310798
rect 386321 310856 389282 310858
rect 386321 310800 386326 310856
rect 386382 310800 389282 310856
rect 386321 310798 389282 310800
rect 386321 310795 386387 310798
rect 379421 310722 379487 310725
rect 369902 310720 379487 310722
rect 369902 310664 379426 310720
rect 379482 310664 379487 310720
rect 369902 310662 379487 310664
rect 389222 310722 389282 310798
rect 405641 310856 408602 310858
rect 405641 310800 405646 310856
rect 405702 310800 408602 310856
rect 405641 310798 408602 310800
rect 405641 310795 405707 310798
rect 398741 310722 398807 310725
rect 389222 310720 398807 310722
rect 389222 310664 398746 310720
rect 398802 310664 398807 310720
rect 389222 310662 398807 310664
rect 408542 310722 408602 310798
rect 424961 310856 427922 310858
rect 424961 310800 424966 310856
rect 425022 310800 427922 310856
rect 424961 310798 427922 310800
rect 424961 310795 425027 310798
rect 418061 310722 418127 310725
rect 408542 310720 418127 310722
rect 408542 310664 418066 310720
rect 418122 310664 418127 310720
rect 408542 310662 418127 310664
rect 427862 310722 427922 310798
rect 444281 310856 447242 310858
rect 444281 310800 444286 310856
rect 444342 310800 447242 310856
rect 444281 310798 447242 310800
rect 444281 310795 444347 310798
rect 437381 310722 437447 310725
rect 427862 310720 437447 310722
rect 427862 310664 437386 310720
rect 437442 310664 437447 310720
rect 427862 310662 437447 310664
rect 447182 310722 447242 310798
rect 463601 310856 466562 310858
rect 463601 310800 463606 310856
rect 463662 310800 466562 310856
rect 463601 310798 466562 310800
rect 463601 310795 463667 310798
rect 456701 310722 456767 310725
rect 447182 310720 456767 310722
rect 447182 310664 456706 310720
rect 456762 310664 456767 310720
rect 447182 310662 456767 310664
rect 466502 310722 466562 310798
rect 482921 310856 485882 310858
rect 482921 310800 482926 310856
rect 482982 310800 485882 310856
rect 482921 310798 485882 310800
rect 482921 310795 482987 310798
rect 475561 310722 475627 310725
rect 466502 310720 475627 310722
rect 466502 310664 475566 310720
rect 475622 310664 475627 310720
rect 466502 310662 475627 310664
rect 485822 310722 485882 310798
rect 502241 310856 505202 310858
rect 502241 310800 502246 310856
rect 502302 310800 505202 310856
rect 502241 310798 505202 310800
rect 502241 310795 502307 310798
rect 495341 310722 495407 310725
rect 485822 310720 495407 310722
rect 485822 310664 495346 310720
rect 495402 310664 495407 310720
rect 485822 310662 495407 310664
rect 505142 310722 505202 310798
rect 521561 310856 524522 310858
rect 521561 310800 521566 310856
rect 521622 310800 524522 310856
rect 521561 310798 524522 310800
rect 521561 310795 521627 310798
rect 514661 310722 514727 310725
rect 505142 310720 514727 310722
rect 505142 310664 514666 310720
rect 514722 310664 514727 310720
rect 505142 310662 514727 310664
rect 524462 310722 524522 310798
rect 540881 310856 541131 310858
rect 540881 310800 540886 310856
rect 540942 310800 541070 310856
rect 541126 310800 541131 310856
rect 540881 310798 541131 310800
rect 540881 310795 540947 310798
rect 541065 310795 541131 310798
rect 560334 310796 560340 310860
rect 560404 310796 560410 310860
rect 583520 310858 584960 310948
rect 583342 310798 584960 310858
rect 533981 310722 534047 310725
rect 560342 310722 560402 310796
rect 524462 310720 534047 310722
rect 524462 310664 533986 310720
rect 534042 310664 534047 310720
rect 524462 310662 534047 310664
rect 267641 310586 267707 310589
rect 278822 310586 278882 310662
rect 288341 310659 288407 310662
rect 320725 310659 320791 310662
rect 340781 310659 340847 310662
rect 359641 310659 359707 310662
rect 379421 310659 379487 310662
rect 398741 310659 398807 310662
rect 418061 310659 418127 310662
rect 437381 310659 437447 310662
rect 456701 310659 456767 310662
rect 475561 310659 475627 310662
rect 495341 310659 495407 310662
rect 514661 310659 514727 310662
rect 533981 310659 534047 310662
rect 560158 310662 560402 310722
rect 267641 310584 278882 310586
rect 267641 310528 267646 310584
rect 267702 310528 278882 310584
rect 267641 310526 278882 310528
rect 543825 310586 543891 310589
rect 550582 310586 550588 310588
rect 543825 310584 550588 310586
rect 543825 310528 543830 310584
rect 543886 310528 550588 310584
rect 543825 310526 550588 310528
rect 267641 310523 267707 310526
rect 543825 310523 543891 310526
rect 550582 310524 550588 310526
rect 550652 310524 550658 310588
rect 555417 310586 555483 310589
rect 560158 310586 560218 310662
rect 560518 310660 560524 310724
rect 560588 310722 560594 310724
rect 583342 310722 583402 310798
rect 560588 310662 576778 310722
rect 560588 310660 560594 310662
rect 555417 310584 560218 310586
rect 555417 310528 555422 310584
rect 555478 310528 560218 310584
rect 555417 310526 560218 310528
rect 576718 310586 576778 310662
rect 576902 310662 583402 310722
rect 583520 310708 584960 310798
rect 576902 310586 576962 310662
rect 576718 310526 576962 310586
rect 555417 310523 555483 310526
rect 550582 310252 550588 310316
rect 550652 310314 550658 310316
rect 555417 310314 555483 310317
rect 550652 310312 555483 310314
rect 550652 310256 555422 310312
rect 555478 310256 555483 310312
rect 550652 310254 555483 310256
rect 550652 310252 550658 310254
rect 555417 310251 555483 310254
rect -960 308818 480 308908
rect 3325 308818 3391 308821
rect -960 308816 3391 308818
rect -960 308760 3330 308816
rect 3386 308760 3391 308816
rect -960 308758 3391 308760
rect -960 308668 480 308758
rect 3325 308755 3391 308758
rect 278037 306370 278103 306373
rect 278313 306370 278379 306373
rect 278037 306368 278379 306370
rect 278037 306312 278042 306368
rect 278098 306312 278318 306368
rect 278374 306312 278379 306368
rect 278037 306310 278379 306312
rect 278037 306307 278103 306310
rect 278313 306307 278379 306310
rect 579797 299162 579863 299165
rect 583520 299162 584960 299252
rect 579797 299160 584960 299162
rect 579797 299104 579802 299160
rect 579858 299104 584960 299160
rect 579797 299102 584960 299104
rect 579797 299099 579863 299102
rect 583520 299012 584960 299102
rect 253841 296714 253907 296717
rect 254025 296714 254091 296717
rect 253841 296712 254091 296714
rect 253841 296656 253846 296712
rect 253902 296656 254030 296712
rect 254086 296656 254091 296712
rect 253841 296654 254091 296656
rect 253841 296651 253907 296654
rect 254025 296651 254091 296654
rect 277945 295354 278011 295357
rect 278221 295354 278287 295357
rect 277945 295352 278287 295354
rect 277945 295296 277950 295352
rect 278006 295296 278226 295352
rect 278282 295296 278287 295352
rect 277945 295294 278287 295296
rect 277945 295291 278011 295294
rect 278221 295291 278287 295294
rect -960 294402 480 294492
rect 3509 294402 3575 294405
rect -960 294400 3575 294402
rect -960 294344 3514 294400
rect 3570 294344 3575 294400
rect -960 294342 3575 294344
rect -960 294252 480 294342
rect 3509 294339 3575 294342
rect 583520 287316 584960 287556
rect -960 280122 480 280212
rect 3969 280122 4035 280125
rect -960 280120 4035 280122
rect -960 280064 3974 280120
rect 4030 280064 4035 280120
rect -960 280062 4035 280064
rect -960 279972 480 280062
rect 3969 280059 4035 280062
rect 237649 278762 237715 278765
rect 237782 278762 237788 278764
rect 237649 278760 237788 278762
rect 237649 278704 237654 278760
rect 237710 278704 237788 278760
rect 237649 278702 237788 278704
rect 237649 278699 237715 278702
rect 237782 278700 237788 278702
rect 237852 278700 237858 278764
rect 288065 278762 288131 278765
rect 288249 278762 288315 278765
rect 288065 278760 288315 278762
rect 288065 278704 288070 278760
rect 288126 278704 288254 278760
rect 288310 278704 288315 278760
rect 288065 278702 288315 278704
rect 288065 278699 288131 278702
rect 288249 278699 288315 278702
rect 278037 277402 278103 277405
rect 277902 277400 278103 277402
rect 277902 277344 278042 277400
rect 278098 277344 278103 277400
rect 277902 277342 278103 277344
rect 277902 277266 277962 277342
rect 278037 277339 278103 277342
rect 278313 277266 278379 277269
rect 277902 277264 278379 277266
rect 277902 277208 278318 277264
rect 278374 277208 278379 277264
rect 277902 277206 278379 277208
rect 278313 277203 278379 277206
rect 580165 275770 580231 275773
rect 583520 275770 584960 275860
rect 580165 275768 584960 275770
rect 580165 275712 580170 275768
rect 580226 275712 584960 275768
rect 580165 275710 584960 275712
rect 580165 275707 580231 275710
rect 583520 275620 584960 275710
rect 270769 269106 270835 269109
rect 270953 269106 271019 269109
rect 270769 269104 271019 269106
rect 270769 269048 270774 269104
rect 270830 269048 270958 269104
rect 271014 269048 271019 269104
rect 270769 269046 271019 269048
rect 270769 269043 270835 269046
rect 270953 269043 271019 269046
rect -960 265706 480 265796
rect 3509 265706 3575 265709
rect -960 265704 3575 265706
rect -960 265648 3514 265704
rect 3570 265648 3575 265704
rect -960 265646 3575 265648
rect -960 265556 480 265646
rect 3509 265643 3575 265646
rect 237649 264346 237715 264349
rect 237782 264346 237788 264348
rect 237649 264344 237788 264346
rect 237649 264288 237654 264344
rect 237710 264288 237788 264344
rect 237649 264286 237788 264288
rect 237649 264283 237715 264286
rect 237782 264284 237788 264286
rect 237852 264284 237858 264348
rect 580165 263938 580231 263941
rect 583520 263938 584960 264028
rect 580165 263936 584960 263938
rect 580165 263880 580170 263936
rect 580226 263880 584960 263936
rect 580165 263878 584960 263880
rect 580165 263875 580231 263878
rect 583520 263788 584960 263878
rect 251357 258090 251423 258093
rect 251357 258088 251466 258090
rect 251357 258032 251362 258088
rect 251418 258032 251466 258088
rect 251357 258027 251466 258032
rect 251406 257957 251466 258027
rect 251357 257952 251466 257957
rect 251357 257896 251362 257952
rect 251418 257896 251466 257952
rect 251357 257894 251466 257896
rect 251357 257891 251423 257894
rect 579797 252242 579863 252245
rect 583520 252242 584960 252332
rect 579797 252240 584960 252242
rect 579797 252184 579802 252240
rect 579858 252184 584960 252240
rect 579797 252182 584960 252184
rect 579797 252179 579863 252182
rect 583520 252092 584960 252182
rect -960 251290 480 251380
rect 3141 251290 3207 251293
rect -960 251288 3207 251290
rect -960 251232 3146 251288
rect 3202 251232 3207 251288
rect -960 251230 3207 251232
rect -960 251140 480 251230
rect 3141 251227 3207 251230
rect 270769 249794 270835 249797
rect 270953 249794 271019 249797
rect 270769 249792 271019 249794
rect 270769 249736 270774 249792
rect 270830 249736 270958 249792
rect 271014 249736 271019 249792
rect 270769 249734 271019 249736
rect 270769 249731 270835 249734
rect 270953 249731 271019 249734
rect 229553 241498 229619 241501
rect 229829 241498 229895 241501
rect 229553 241496 229895 241498
rect 229553 241440 229558 241496
rect 229614 241440 229834 241496
rect 229890 241440 229895 241496
rect 229553 241438 229895 241440
rect 229553 241435 229619 241438
rect 229829 241435 229895 241438
rect 583520 240396 584960 240636
rect 238293 238914 238359 238917
rect 237974 238912 238359 238914
rect 237974 238856 238298 238912
rect 238354 238856 238359 238912
rect 237974 238854 238359 238856
rect 237974 238778 238034 238854
rect 238293 238851 238359 238854
rect 238109 238778 238175 238781
rect 237974 238776 238175 238778
rect 237974 238720 238114 238776
rect 238170 238720 238175 238776
rect 237974 238718 238175 238720
rect 238109 238715 238175 238718
rect 277853 238778 277919 238781
rect 278037 238778 278103 238781
rect 277853 238776 278103 238778
rect 277853 238720 277858 238776
rect 277914 238720 278042 238776
rect 278098 238720 278103 238776
rect 277853 238718 278103 238720
rect 277853 238715 277919 238718
rect 278037 238715 278103 238718
rect 240869 237418 240935 237421
rect 241053 237418 241119 237421
rect 240869 237416 241119 237418
rect 240869 237360 240874 237416
rect 240930 237360 241058 237416
rect 241114 237360 241119 237416
rect 240869 237358 241119 237360
rect 240869 237355 240935 237358
rect 241053 237355 241119 237358
rect -960 237010 480 237100
rect 3785 237010 3851 237013
rect -960 237008 3851 237010
rect -960 236952 3790 237008
rect 3846 236952 3851 237008
rect -960 236950 3851 236952
rect -960 236860 480 236950
rect 3785 236947 3851 236950
rect 275369 229122 275435 229125
rect 275553 229122 275619 229125
rect 275369 229120 275619 229122
rect 275369 229064 275374 229120
rect 275430 229064 275558 229120
rect 275614 229064 275619 229120
rect 275369 229062 275619 229064
rect 275369 229059 275435 229062
rect 275553 229059 275619 229062
rect 277761 229122 277827 229125
rect 277945 229122 278011 229125
rect 277761 229120 278011 229122
rect 277761 229064 277766 229120
rect 277822 229064 277950 229120
rect 278006 229064 278011 229120
rect 277761 229062 278011 229064
rect 277761 229059 277827 229062
rect 277945 229059 278011 229062
rect 583520 228850 584960 228940
rect 583342 228790 584960 228850
rect 237230 228108 237236 228172
rect 237300 228170 237306 228172
rect 244181 228170 244247 228173
rect 237300 228168 244247 228170
rect 237300 228112 244186 228168
rect 244242 228112 244247 228168
rect 237300 228110 244247 228112
rect 237300 228108 237306 228110
rect 244181 228107 244247 228110
rect 244365 228034 244431 228037
rect 248413 228034 248479 228037
rect 244365 228032 248479 228034
rect 244365 227976 244370 228032
rect 244426 227976 248418 228032
rect 248474 227976 248479 228032
rect 244365 227974 248479 227976
rect 244365 227971 244431 227974
rect 248413 227971 248479 227974
rect 257838 227972 257844 228036
rect 257908 228034 257914 228036
rect 259453 228034 259519 228037
rect 257908 228032 259519 228034
rect 257908 227976 259458 228032
rect 259514 227976 259519 228032
rect 257908 227974 259519 227976
rect 257908 227972 257914 227974
rect 259453 227971 259519 227974
rect 273302 227974 282930 228034
rect 270401 227898 270467 227901
rect 273302 227898 273362 227974
rect 270401 227896 273362 227898
rect 270401 227840 270406 227896
rect 270462 227840 273362 227896
rect 270401 227838 273362 227840
rect 270401 227835 270467 227838
rect 282870 227762 282930 227974
rect 335310 227974 344938 228034
rect 302141 227898 302207 227901
rect 321461 227898 321527 227901
rect 292622 227896 302207 227898
rect 292622 227840 302146 227896
rect 302202 227840 302207 227896
rect 292622 227838 302207 227840
rect 292622 227762 292682 227838
rect 302141 227835 302207 227838
rect 311942 227896 321527 227898
rect 311942 227840 321466 227896
rect 321522 227840 321527 227896
rect 311942 227838 321527 227840
rect 282870 227702 292682 227762
rect 309041 227762 309107 227765
rect 311942 227762 312002 227838
rect 321461 227835 321527 227838
rect 323025 227898 323091 227901
rect 323025 227896 331138 227898
rect 323025 227840 323030 227896
rect 323086 227840 331138 227896
rect 323025 227838 331138 227840
rect 323025 227835 323091 227838
rect 309041 227760 312002 227762
rect 309041 227704 309046 227760
rect 309102 227704 312002 227760
rect 309041 227702 312002 227704
rect 331078 227762 331138 227838
rect 335310 227762 335370 227974
rect 331078 227702 335370 227762
rect 344878 227762 344938 227974
rect 345062 227974 354690 228034
rect 345062 227762 345122 227974
rect 354630 227898 354690 227974
rect 364382 227974 374010 228034
rect 354630 227838 364258 227898
rect 344878 227702 345122 227762
rect 364198 227762 364258 227838
rect 364382 227762 364442 227974
rect 373950 227898 374010 227974
rect 383702 227974 405842 228034
rect 373950 227838 383578 227898
rect 364198 227702 364442 227762
rect 383518 227762 383578 227838
rect 383702 227762 383762 227974
rect 405782 227898 405842 227974
rect 495390 227974 514770 228034
rect 415301 227898 415367 227901
rect 437381 227898 437447 227901
rect 456701 227898 456767 227901
rect 405782 227896 415367 227898
rect 405782 227840 415306 227896
rect 415362 227840 415367 227896
rect 405782 227838 415367 227840
rect 415301 227835 415367 227838
rect 427862 227896 437447 227898
rect 427862 227840 437386 227896
rect 437442 227840 437447 227896
rect 427862 227838 437447 227840
rect 383518 227702 383762 227762
rect 415301 227762 415367 227765
rect 427862 227762 427922 227838
rect 437381 227835 437447 227838
rect 447182 227896 456767 227898
rect 447182 227840 456706 227896
rect 456762 227840 456767 227896
rect 447182 227838 456767 227840
rect 415301 227760 427922 227762
rect 415301 227704 415306 227760
rect 415362 227704 427922 227760
rect 415301 227702 427922 227704
rect 444281 227762 444347 227765
rect 447182 227762 447242 227838
rect 456701 227835 456767 227838
rect 456885 227898 456951 227901
rect 476021 227898 476087 227901
rect 456885 227896 466378 227898
rect 456885 227840 456890 227896
rect 456946 227840 466378 227896
rect 456885 227838 466378 227840
rect 456885 227835 456951 227838
rect 444281 227760 447242 227762
rect 444281 227704 444286 227760
rect 444342 227704 447242 227760
rect 444281 227702 447242 227704
rect 466318 227762 466378 227838
rect 466502 227896 476087 227898
rect 466502 227840 476026 227896
rect 476082 227840 476087 227896
rect 466502 227838 476087 227840
rect 466502 227762 466562 227838
rect 476021 227835 476087 227838
rect 466318 227702 466562 227762
rect 482921 227762 482987 227765
rect 495390 227762 495450 227974
rect 482921 227760 495450 227762
rect 482921 227704 482926 227760
rect 482982 227704 495450 227760
rect 482921 227702 495450 227704
rect 514710 227762 514770 227974
rect 533981 227898 534047 227901
rect 553301 227898 553367 227901
rect 572621 227898 572687 227901
rect 524462 227896 534047 227898
rect 524462 227840 533986 227896
rect 534042 227840 534047 227896
rect 524462 227838 534047 227840
rect 524462 227762 524522 227838
rect 533981 227835 534047 227838
rect 543782 227896 553367 227898
rect 543782 227840 553306 227896
rect 553362 227840 553367 227896
rect 543782 227838 553367 227840
rect 514710 227702 524522 227762
rect 540881 227762 540947 227765
rect 543782 227762 543842 227838
rect 553301 227835 553367 227838
rect 563102 227896 572687 227898
rect 563102 227840 572626 227896
rect 572682 227840 572687 227896
rect 563102 227838 572687 227840
rect 540881 227760 543842 227762
rect 540881 227704 540886 227760
rect 540942 227704 543842 227760
rect 540881 227702 543842 227704
rect 560201 227762 560267 227765
rect 563102 227762 563162 227838
rect 572621 227835 572687 227838
rect 560201 227760 563162 227762
rect 560201 227704 560206 227760
rect 560262 227704 563162 227760
rect 560201 227702 563162 227704
rect 579521 227762 579587 227765
rect 583342 227762 583402 228790
rect 583520 228700 584960 228790
rect 579521 227760 583402 227762
rect 579521 227704 579526 227760
rect 579582 227704 583402 227760
rect 579521 227702 583402 227704
rect 309041 227699 309107 227702
rect 415301 227699 415367 227702
rect 444281 227699 444347 227702
rect 482921 227699 482987 227702
rect 540881 227699 540947 227702
rect 560201 227699 560267 227702
rect 579521 227699 579587 227702
rect 248413 227626 248479 227629
rect 257838 227626 257844 227628
rect 248413 227624 257844 227626
rect 248413 227568 248418 227624
rect 248474 227568 257844 227624
rect 248413 227566 257844 227568
rect 248413 227563 248479 227566
rect 257838 227564 257844 227566
rect 257908 227564 257914 227628
rect -960 222594 480 222684
rect 3141 222594 3207 222597
rect -960 222592 3207 222594
rect -960 222536 3146 222592
rect 3202 222536 3207 222592
rect -960 222534 3207 222536
rect -960 222444 480 222534
rect 3141 222531 3207 222534
rect 229553 222186 229619 222189
rect 229829 222186 229895 222189
rect 229553 222184 229895 222186
rect 229553 222128 229558 222184
rect 229614 222128 229834 222184
rect 229890 222128 229895 222184
rect 229553 222126 229895 222128
rect 229553 222123 229619 222126
rect 229829 222123 229895 222126
rect 259729 220826 259795 220829
rect 260097 220826 260163 220829
rect 259729 220824 260163 220826
rect 259729 220768 259734 220824
rect 259790 220768 260102 220824
rect 260158 220768 260163 220824
rect 259729 220766 260163 220768
rect 259729 220763 259795 220766
rect 260097 220763 260163 220766
rect 260281 220826 260347 220829
rect 260557 220826 260623 220829
rect 260281 220824 260623 220826
rect 260281 220768 260286 220824
rect 260342 220768 260562 220824
rect 260618 220768 260623 220824
rect 260281 220766 260623 220768
rect 260281 220763 260347 220766
rect 260557 220763 260623 220766
rect 237465 219466 237531 219469
rect 237649 219466 237715 219469
rect 237465 219464 237715 219466
rect 237465 219408 237470 219464
rect 237526 219408 237654 219464
rect 237710 219408 237715 219464
rect 237465 219406 237715 219408
rect 237465 219403 237531 219406
rect 237649 219403 237715 219406
rect 238845 219466 238911 219469
rect 239121 219466 239187 219469
rect 238845 219464 239187 219466
rect 238845 219408 238850 219464
rect 238906 219408 239126 219464
rect 239182 219408 239187 219464
rect 238845 219406 239187 219408
rect 238845 219403 238911 219406
rect 239121 219403 239187 219406
rect 240869 219466 240935 219469
rect 241053 219466 241119 219469
rect 240869 219464 241119 219466
rect 240869 219408 240874 219464
rect 240930 219408 241058 219464
rect 241114 219408 241119 219464
rect 240869 219406 241119 219408
rect 240869 219403 240935 219406
rect 241053 219403 241119 219406
rect 580165 217018 580231 217021
rect 583520 217018 584960 217108
rect 580165 217016 584960 217018
rect 580165 216960 580170 217016
rect 580226 216960 584960 217016
rect 580165 216958 584960 216960
rect 580165 216955 580231 216958
rect 583520 216868 584960 216958
rect 259729 211170 259795 211173
rect 259913 211170 259979 211173
rect 259729 211168 259979 211170
rect 259729 211112 259734 211168
rect 259790 211112 259918 211168
rect 259974 211112 259979 211168
rect 259729 211110 259979 211112
rect 259729 211107 259795 211110
rect 259913 211107 259979 211110
rect 260189 211170 260255 211173
rect 260557 211170 260623 211173
rect 260189 211168 260623 211170
rect 260189 211112 260194 211168
rect 260250 211112 260562 211168
rect 260618 211112 260623 211168
rect 260189 211110 260623 211112
rect 260189 211107 260255 211110
rect 260557 211107 260623 211110
rect -960 208178 480 208268
rect 3509 208178 3575 208181
rect -960 208176 3575 208178
rect -960 208120 3514 208176
rect 3570 208120 3575 208176
rect -960 208118 3575 208120
rect -960 208028 480 208118
rect 3509 208115 3575 208118
rect 579797 205322 579863 205325
rect 583520 205322 584960 205412
rect 579797 205320 584960 205322
rect 579797 205264 579802 205320
rect 579858 205264 584960 205320
rect 579797 205262 584960 205264
rect 579797 205259 579863 205262
rect 583520 205172 584960 205262
rect 229553 202874 229619 202877
rect 229829 202874 229895 202877
rect 229553 202872 229895 202874
rect 229553 202816 229558 202872
rect 229614 202816 229834 202872
rect 229890 202816 229895 202872
rect 229553 202814 229895 202816
rect 229553 202811 229619 202814
rect 229829 202811 229895 202814
rect 251541 202874 251607 202877
rect 251725 202874 251791 202877
rect 251541 202872 251791 202874
rect 251541 202816 251546 202872
rect 251602 202816 251730 202872
rect 251786 202816 251791 202872
rect 251541 202814 251791 202816
rect 251541 202811 251607 202814
rect 251725 202811 251791 202814
rect 278037 202874 278103 202877
rect 278221 202874 278287 202877
rect 278037 202872 278287 202874
rect 278037 202816 278042 202872
rect 278098 202816 278226 202872
rect 278282 202816 278287 202872
rect 278037 202814 278287 202816
rect 278037 202811 278103 202814
rect 278221 202811 278287 202814
rect 253933 201514 253999 201517
rect 254117 201514 254183 201517
rect 253933 201512 254183 201514
rect 253933 201456 253938 201512
rect 253994 201456 254122 201512
rect 254178 201456 254183 201512
rect 253933 201454 254183 201456
rect 253933 201451 253999 201454
rect 254117 201451 254183 201454
rect 3509 194578 3575 194581
rect 282862 194578 282868 194580
rect 3509 194576 282868 194578
rect 3509 194520 3514 194576
rect 3570 194520 282868 194576
rect 3509 194518 282868 194520
rect 3509 194515 3575 194518
rect 282862 194516 282868 194518
rect 282932 194516 282938 194580
rect -960 193898 480 193988
rect 3509 193898 3575 193901
rect -960 193896 3575 193898
rect -960 193840 3514 193896
rect 3570 193840 3575 193896
rect -960 193838 3575 193840
rect -960 193748 480 193838
rect 3509 193835 3575 193838
rect 583520 193476 584960 193716
rect 241145 191858 241211 191861
rect 241329 191858 241395 191861
rect 241145 191856 241395 191858
rect 241145 191800 241150 191856
rect 241206 191800 241334 191856
rect 241390 191800 241395 191856
rect 241145 191798 241395 191800
rect 241145 191795 241211 191798
rect 241329 191795 241395 191798
rect 259729 191858 259795 191861
rect 259913 191858 259979 191861
rect 259729 191856 259979 191858
rect 259729 191800 259734 191856
rect 259790 191800 259918 191856
rect 259974 191800 259979 191856
rect 259729 191798 259979 191800
rect 259729 191795 259795 191798
rect 259913 191795 259979 191798
rect 229553 183562 229619 183565
rect 229829 183562 229895 183565
rect 229553 183560 229895 183562
rect 229553 183504 229558 183560
rect 229614 183504 229834 183560
rect 229890 183504 229895 183560
rect 229553 183502 229895 183504
rect 229553 183499 229619 183502
rect 229829 183499 229895 183502
rect 259913 183562 259979 183565
rect 260097 183562 260163 183565
rect 259913 183560 260163 183562
rect 259913 183504 259918 183560
rect 259974 183504 260102 183560
rect 260158 183504 260163 183560
rect 259913 183502 260163 183504
rect 259913 183499 259979 183502
rect 260097 183499 260163 183502
rect 580165 181930 580231 181933
rect 583520 181930 584960 182020
rect 580165 181928 584960 181930
rect 580165 181872 580170 181928
rect 580226 181872 584960 181928
rect 580165 181870 584960 181872
rect 580165 181867 580231 181870
rect 583520 181780 584960 181870
rect 277761 180842 277827 180845
rect 277945 180842 278011 180845
rect 277761 180840 278011 180842
rect 277761 180784 277766 180840
rect 277822 180784 277950 180840
rect 278006 180784 278011 180840
rect 277761 180782 278011 180784
rect 277761 180779 277827 180782
rect 277945 180779 278011 180782
rect -960 179482 480 179572
rect 3233 179482 3299 179485
rect -960 179480 3299 179482
rect -960 179424 3238 179480
rect 3294 179424 3299 179480
rect -960 179422 3299 179424
rect -960 179332 480 179422
rect 3233 179419 3299 179422
rect 272149 173906 272215 173909
rect 272333 173906 272399 173909
rect 272149 173904 272399 173906
rect 272149 173848 272154 173904
rect 272210 173848 272338 173904
rect 272394 173848 272399 173904
rect 272149 173846 272399 173848
rect 272149 173843 272215 173846
rect 272333 173843 272399 173846
rect 241145 172546 241211 172549
rect 241329 172546 241395 172549
rect 241145 172544 241395 172546
rect 241145 172488 241150 172544
rect 241206 172488 241334 172544
rect 241390 172488 241395 172544
rect 241145 172486 241395 172488
rect 241145 172483 241211 172486
rect 241329 172483 241395 172486
rect 580165 170098 580231 170101
rect 583520 170098 584960 170188
rect 580165 170096 584960 170098
rect 580165 170040 580170 170096
rect 580226 170040 584960 170096
rect 580165 170038 584960 170040
rect 580165 170035 580231 170038
rect 583520 169948 584960 170038
rect -960 165066 480 165156
rect 3509 165066 3575 165069
rect -960 165064 3575 165066
rect -960 165008 3514 165064
rect 3570 165008 3575 165064
rect -960 165006 3575 165008
rect -960 164916 480 165006
rect 3509 165003 3575 165006
rect 272149 164250 272215 164253
rect 272333 164250 272399 164253
rect 272149 164248 272399 164250
rect 272149 164192 272154 164248
rect 272210 164192 272338 164248
rect 272394 164192 272399 164248
rect 272149 164190 272399 164192
rect 272149 164187 272215 164190
rect 272333 164187 272399 164190
rect 270769 162890 270835 162893
rect 270769 162888 270970 162890
rect 270769 162832 270774 162888
rect 270830 162832 270970 162888
rect 270769 162830 270970 162832
rect 270769 162827 270835 162830
rect 270769 162618 270835 162621
rect 270910 162618 270970 162830
rect 270769 162616 270970 162618
rect 270769 162560 270774 162616
rect 270830 162560 270970 162616
rect 270769 162558 270970 162560
rect 270769 162555 270835 162558
rect 579797 158402 579863 158405
rect 583520 158402 584960 158492
rect 579797 158400 584960 158402
rect 579797 158344 579802 158400
rect 579858 158344 584960 158400
rect 579797 158342 584960 158344
rect 579797 158339 579863 158342
rect 583520 158252 584960 158342
rect 229645 154594 229711 154597
rect 229829 154594 229895 154597
rect 229645 154592 229895 154594
rect 229645 154536 229650 154592
rect 229706 154536 229834 154592
rect 229890 154536 229895 154592
rect 229645 154534 229895 154536
rect 229645 154531 229711 154534
rect 229829 154531 229895 154534
rect 237557 153370 237623 153373
rect 237557 153368 237666 153370
rect 237557 153312 237562 153368
rect 237618 153312 237666 153368
rect 237557 153307 237666 153312
rect 237606 153237 237666 153307
rect 237557 153232 237666 153237
rect 237557 153176 237562 153232
rect 237618 153176 237666 153232
rect 237557 153174 237666 153176
rect 238937 153234 239003 153237
rect 239121 153234 239187 153237
rect 238937 153232 239187 153234
rect 238937 153176 238942 153232
rect 238998 153176 239126 153232
rect 239182 153176 239187 153232
rect 238937 153174 239187 153176
rect 237557 153171 237623 153174
rect 238937 153171 239003 153174
rect 239121 153171 239187 153174
rect 270769 153234 270835 153237
rect 270953 153234 271019 153237
rect 270769 153232 271019 153234
rect 270769 153176 270774 153232
rect 270830 153176 270958 153232
rect 271014 153176 271019 153232
rect 270769 153174 271019 153176
rect 270769 153171 270835 153174
rect 270953 153171 271019 153174
rect 3509 151738 3575 151741
rect 284334 151738 284340 151740
rect 3509 151736 284340 151738
rect 3509 151680 3514 151736
rect 3570 151680 284340 151736
rect 3509 151678 284340 151680
rect 3509 151675 3575 151678
rect 284334 151676 284340 151678
rect 284404 151676 284410 151740
rect -960 150786 480 150876
rect 3509 150786 3575 150789
rect -960 150784 3575 150786
rect -960 150728 3514 150784
rect 3570 150728 3575 150784
rect -960 150726 3575 150728
rect -960 150636 480 150726
rect 3509 150723 3575 150726
rect 583520 146556 584960 146796
rect 260189 145074 260255 145077
rect 260054 145072 260255 145074
rect 260054 145016 260194 145072
rect 260250 145016 260255 145072
rect 260054 145014 260255 145016
rect 260054 144941 260114 145014
rect 260189 145011 260255 145014
rect 253933 144938 253999 144941
rect 254117 144938 254183 144941
rect 253933 144936 254183 144938
rect 253933 144880 253938 144936
rect 253994 144880 254122 144936
rect 254178 144880 254183 144936
rect 253933 144878 254183 144880
rect 260054 144936 260163 144941
rect 260054 144880 260102 144936
rect 260158 144880 260163 144936
rect 260054 144878 260163 144880
rect 253933 144875 253999 144878
rect 254117 144875 254183 144878
rect 260097 144875 260163 144878
rect -960 136370 480 136460
rect 3509 136370 3575 136373
rect -960 136368 3575 136370
rect -960 136312 3514 136368
rect 3570 136312 3575 136368
rect -960 136310 3575 136312
rect -960 136220 480 136310
rect 3509 136307 3575 136310
rect 229461 135282 229527 135285
rect 229645 135282 229711 135285
rect 229461 135280 229711 135282
rect 229461 135224 229466 135280
rect 229522 135224 229650 135280
rect 229706 135224 229711 135280
rect 229461 135222 229711 135224
rect 229461 135219 229527 135222
rect 229645 135219 229711 135222
rect 580165 134874 580231 134877
rect 583520 134874 584960 134964
rect 580165 134872 584960 134874
rect 580165 134816 580170 134872
rect 580226 134816 584960 134872
rect 580165 134814 584960 134816
rect 580165 134811 580231 134814
rect 583520 134724 584960 134814
rect 260097 134058 260163 134061
rect 260097 134056 260298 134058
rect 260097 134000 260102 134056
rect 260158 134000 260298 134056
rect 260097 133998 260298 134000
rect 260097 133995 260163 133998
rect 260238 133925 260298 133998
rect 260238 133920 260347 133925
rect 260238 133864 260286 133920
rect 260342 133864 260347 133920
rect 260238 133862 260347 133864
rect 260281 133859 260347 133862
rect 256417 132426 256483 132429
rect 256601 132426 256667 132429
rect 256417 132424 256667 132426
rect 256417 132368 256422 132424
rect 256478 132368 256606 132424
rect 256662 132368 256667 132424
rect 256417 132366 256667 132368
rect 256417 132363 256483 132366
rect 256601 132363 256667 132366
rect 241145 125762 241211 125765
rect 241102 125760 241211 125762
rect 241102 125704 241150 125760
rect 241206 125704 241211 125760
rect 241102 125699 241211 125704
rect 241102 125629 241162 125699
rect 241053 125624 241162 125629
rect 241053 125568 241058 125624
rect 241114 125568 241162 125624
rect 241053 125566 241162 125568
rect 241053 125563 241119 125566
rect 237557 124402 237623 124405
rect 237557 124400 237666 124402
rect 237557 124344 237562 124400
rect 237618 124344 237666 124400
rect 237557 124339 237666 124344
rect 237606 124269 237666 124339
rect 237606 124264 237715 124269
rect 237606 124208 237654 124264
rect 237710 124208 237715 124264
rect 237606 124206 237715 124208
rect 237649 124203 237715 124206
rect 238661 124266 238727 124269
rect 238937 124266 239003 124269
rect 238661 124264 239003 124266
rect 238661 124208 238666 124264
rect 238722 124208 238942 124264
rect 238998 124208 239003 124264
rect 238661 124206 239003 124208
rect 238661 124203 238727 124206
rect 238937 124203 239003 124206
rect 580165 123178 580231 123181
rect 583520 123178 584960 123268
rect 580165 123176 584960 123178
rect 580165 123120 580170 123176
rect 580226 123120 584960 123176
rect 580165 123118 584960 123120
rect 580165 123115 580231 123118
rect 583520 123028 584960 123118
rect -960 122090 480 122180
rect 2957 122090 3023 122093
rect -960 122088 3023 122090
rect -960 122032 2962 122088
rect 3018 122032 3023 122088
rect -960 122030 3023 122032
rect -960 121940 480 122030
rect 2957 122027 3023 122030
rect 229461 115970 229527 115973
rect 229645 115970 229711 115973
rect 229461 115968 229711 115970
rect 229461 115912 229466 115968
rect 229522 115912 229650 115968
rect 229706 115912 229711 115968
rect 229461 115910 229711 115912
rect 229461 115907 229527 115910
rect 229645 115907 229711 115910
rect 579797 111482 579863 111485
rect 583520 111482 584960 111572
rect 579797 111480 584960 111482
rect 579797 111424 579802 111480
rect 579858 111424 584960 111480
rect 579797 111422 584960 111424
rect 579797 111419 579863 111422
rect 583520 111332 584960 111422
rect 3509 109034 3575 109037
rect 285622 109034 285628 109036
rect 3509 109032 285628 109034
rect 3509 108976 3514 109032
rect 3570 108976 285628 109032
rect 3509 108974 285628 108976
rect 3509 108971 3575 108974
rect 285622 108972 285628 108974
rect 285692 108972 285698 109036
rect -960 107674 480 107764
rect 3509 107674 3575 107677
rect -960 107672 3575 107674
rect -960 107616 3514 107672
rect 3570 107616 3575 107672
rect -960 107614 3575 107616
rect -960 107524 480 107614
rect 3509 107611 3575 107614
rect 248873 106178 248939 106181
rect 248873 106176 249074 106178
rect 248873 106120 248878 106176
rect 248934 106120 249074 106176
rect 248873 106118 249074 106120
rect 248873 106115 248939 106118
rect 249014 105909 249074 106118
rect 248965 105904 249074 105909
rect 248965 105848 248970 105904
rect 249026 105848 249074 105904
rect 248965 105846 249074 105848
rect 248965 105843 249031 105846
rect 583520 99636 584960 99876
rect 229461 96658 229527 96661
rect 229645 96658 229711 96661
rect 229461 96656 229711 96658
rect 229461 96600 229466 96656
rect 229522 96600 229650 96656
rect 229706 96600 229711 96656
rect 229461 96598 229711 96600
rect 229461 96595 229527 96598
rect 229645 96595 229711 96598
rect 278129 96658 278195 96661
rect 278313 96658 278379 96661
rect 278129 96656 278379 96658
rect 278129 96600 278134 96656
rect 278190 96600 278318 96656
rect 278374 96600 278379 96656
rect 278129 96598 278379 96600
rect 278129 96595 278195 96598
rect 278313 96595 278379 96598
rect -960 93258 480 93348
rect 3509 93258 3575 93261
rect -960 93256 3575 93258
rect -960 93200 3514 93256
rect 3570 93200 3575 93256
rect -960 93198 3575 93200
rect -960 93108 480 93198
rect 3509 93195 3575 93198
rect 580165 87954 580231 87957
rect 583520 87954 584960 88044
rect 580165 87952 584960 87954
rect 580165 87896 580170 87952
rect 580226 87896 584960 87952
rect 580165 87894 584960 87896
rect 580165 87891 580231 87894
rect 583520 87804 584960 87894
rect 258533 84146 258599 84149
rect 258398 84144 258599 84146
rect 258398 84088 258538 84144
rect 258594 84088 258599 84144
rect 258398 84086 258599 84088
rect 258398 84010 258458 84086
rect 258533 84083 258599 84086
rect 258717 84010 258783 84013
rect 258398 84008 258783 84010
rect 258398 83952 258722 84008
rect 258778 83952 258783 84008
rect 258398 83950 258783 83952
rect 258717 83947 258783 83950
rect -960 78978 480 79068
rect 3233 78978 3299 78981
rect -960 78976 3299 78978
rect -960 78920 3238 78976
rect 3294 78920 3299 78976
rect -960 78918 3299 78920
rect -960 78828 480 78918
rect 3233 78915 3299 78918
rect 521561 76530 521627 76533
rect 511950 76528 521627 76530
rect 511950 76472 521566 76528
rect 521622 76472 521627 76528
rect 511950 76470 521627 76472
rect 232998 76196 233004 76260
rect 233068 76258 233074 76260
rect 241462 76258 241468 76260
rect 233068 76198 241468 76258
rect 233068 76196 233074 76198
rect 241462 76196 241468 76198
rect 241532 76196 241538 76260
rect 510521 76258 510587 76261
rect 511950 76258 512010 76470
rect 521561 76467 521627 76470
rect 583520 76258 584960 76348
rect 335310 76198 344938 76258
rect 260966 76060 260972 76124
rect 261036 76122 261042 76124
rect 280245 76122 280311 76125
rect 302141 76122 302207 76125
rect 321461 76122 321527 76125
rect 261036 76120 280311 76122
rect 261036 76064 280250 76120
rect 280306 76064 280311 76120
rect 261036 76062 280311 76064
rect 261036 76060 261042 76062
rect 280245 76059 280311 76062
rect 292622 76120 302207 76122
rect 292622 76064 302146 76120
rect 302202 76064 302207 76120
rect 292622 76062 302207 76064
rect 241462 75924 241468 75988
rect 241532 75986 241538 75988
rect 244273 75986 244339 75989
rect 241532 75984 244339 75986
rect 241532 75928 244278 75984
rect 244334 75928 244339 75984
rect 241532 75926 244339 75928
rect 241532 75924 241538 75926
rect 244273 75923 244339 75926
rect 244457 75986 244523 75989
rect 260782 75986 260788 75988
rect 244457 75984 260788 75986
rect 244457 75928 244462 75984
rect 244518 75928 260788 75984
rect 244457 75926 260788 75928
rect 244457 75923 244523 75926
rect 260782 75924 260788 75926
rect 260852 75924 260858 75988
rect 289721 75986 289787 75989
rect 292622 75986 292682 76062
rect 302141 76059 302207 76062
rect 311942 76120 321527 76122
rect 311942 76064 321466 76120
rect 321522 76064 321527 76120
rect 311942 76062 321527 76064
rect 289721 75984 292682 75986
rect 289721 75928 289726 75984
rect 289782 75928 292682 75984
rect 289721 75926 292682 75928
rect 309041 75986 309107 75989
rect 311942 75986 312002 76062
rect 321461 76059 321527 76062
rect 323025 76122 323091 76125
rect 323025 76120 331138 76122
rect 323025 76064 323030 76120
rect 323086 76064 331138 76120
rect 323025 76062 331138 76064
rect 323025 76059 323091 76062
rect 309041 75984 312002 75986
rect 309041 75928 309046 75984
rect 309102 75928 312002 75984
rect 309041 75926 312002 75928
rect 331078 75986 331138 76062
rect 335310 75986 335370 76198
rect 331078 75926 335370 75986
rect 344878 75986 344938 76198
rect 345062 76198 354690 76258
rect 345062 75986 345122 76198
rect 354630 76122 354690 76198
rect 364382 76198 374010 76258
rect 354630 76062 364258 76122
rect 344878 75926 345122 75986
rect 364198 75986 364258 76062
rect 364382 75986 364442 76198
rect 373950 76122 374010 76198
rect 383702 76198 405842 76258
rect 373950 76062 383578 76122
rect 364198 75926 364442 75986
rect 383518 75986 383578 76062
rect 383702 75986 383762 76198
rect 405782 76122 405842 76198
rect 510521 76256 512010 76258
rect 510521 76200 510526 76256
rect 510582 76200 512010 76256
rect 510521 76198 512010 76200
rect 583342 76198 584960 76258
rect 510521 76195 510587 76198
rect 415301 76122 415367 76125
rect 437381 76122 437447 76125
rect 456701 76122 456767 76125
rect 405782 76120 415367 76122
rect 405782 76064 415306 76120
rect 415362 76064 415367 76120
rect 405782 76062 415367 76064
rect 415301 76059 415367 76062
rect 427862 76120 437447 76122
rect 427862 76064 437386 76120
rect 437442 76064 437447 76120
rect 427862 76062 437447 76064
rect 383518 75926 383762 75986
rect 415301 75986 415367 75989
rect 427862 75986 427922 76062
rect 437381 76059 437447 76062
rect 447182 76120 456767 76122
rect 447182 76064 456706 76120
rect 456762 76064 456767 76120
rect 447182 76062 456767 76064
rect 415301 75984 427922 75986
rect 415301 75928 415306 75984
rect 415362 75928 427922 75984
rect 415301 75926 427922 75928
rect 444281 75986 444347 75989
rect 447182 75986 447242 76062
rect 456701 76059 456767 76062
rect 456885 76122 456951 76125
rect 482921 76122 482987 76125
rect 492622 76122 492628 76124
rect 456885 76120 466378 76122
rect 456885 76064 456890 76120
rect 456946 76064 466378 76120
rect 456885 76062 466378 76064
rect 456885 76059 456951 76062
rect 444281 75984 447242 75986
rect 444281 75928 444286 75984
rect 444342 75928 447242 75984
rect 444281 75926 447242 75928
rect 466318 75986 466378 76062
rect 466502 76120 482987 76122
rect 466502 76064 482926 76120
rect 482982 76064 482987 76120
rect 466502 76062 482987 76064
rect 466502 75986 466562 76062
rect 482921 76059 482987 76062
rect 483062 76062 492628 76122
rect 466318 75926 466562 75986
rect 482921 75986 482987 75989
rect 483062 75986 483122 76062
rect 492622 76060 492628 76062
rect 492692 76060 492698 76124
rect 533981 76122 534047 76125
rect 553301 76122 553367 76125
rect 572621 76122 572687 76125
rect 524462 76120 534047 76122
rect 524462 76064 533986 76120
rect 534042 76064 534047 76120
rect 524462 76062 534047 76064
rect 482921 75984 483122 75986
rect 482921 75928 482926 75984
rect 482982 75928 483122 75984
rect 482921 75926 483122 75928
rect 521561 75986 521627 75989
rect 524462 75986 524522 76062
rect 533981 76059 534047 76062
rect 543782 76120 553367 76122
rect 543782 76064 553306 76120
rect 553362 76064 553367 76120
rect 543782 76062 553367 76064
rect 521561 75984 524522 75986
rect 521561 75928 521566 75984
rect 521622 75928 524522 75984
rect 521561 75926 524522 75928
rect 540881 75986 540947 75989
rect 543782 75986 543842 76062
rect 553301 76059 553367 76062
rect 563102 76120 572687 76122
rect 563102 76064 572626 76120
rect 572682 76064 572687 76120
rect 563102 76062 572687 76064
rect 540881 75984 543842 75986
rect 540881 75928 540886 75984
rect 540942 75928 543842 75984
rect 540881 75926 543842 75928
rect 560201 75986 560267 75989
rect 563102 75986 563162 76062
rect 572621 76059 572687 76062
rect 560201 75984 563162 75986
rect 560201 75928 560206 75984
rect 560262 75928 563162 75984
rect 560201 75926 563162 75928
rect 579521 75986 579587 75989
rect 583342 75986 583402 76198
rect 583520 76108 584960 76198
rect 579521 75984 583402 75986
rect 579521 75928 579526 75984
rect 579582 75928 583402 75984
rect 579521 75926 583402 75928
rect 289721 75923 289787 75926
rect 309041 75923 309107 75926
rect 415301 75923 415367 75926
rect 444281 75923 444347 75926
rect 482921 75923 482987 75926
rect 521561 75923 521627 75926
rect 540881 75923 540947 75926
rect 560201 75923 560267 75926
rect 579521 75923 579587 75926
rect 492622 75788 492628 75852
rect 492692 75850 492698 75852
rect 502241 75850 502307 75853
rect 492692 75848 502307 75850
rect 492692 75792 502246 75848
rect 502302 75792 502307 75848
rect 492692 75790 502307 75792
rect 492692 75788 492698 75790
rect 502241 75787 502307 75790
rect 272149 74490 272215 74493
rect 272333 74490 272399 74493
rect 272149 74488 272399 74490
rect 272149 74432 272154 74488
rect 272210 74432 272338 74488
rect 272394 74432 272399 74488
rect 272149 74430 272399 74432
rect 272149 74427 272215 74430
rect 272333 74427 272399 74430
rect 229502 67492 229508 67556
rect 229572 67554 229578 67556
rect 229645 67554 229711 67557
rect 229572 67552 229711 67554
rect 229572 67496 229650 67552
rect 229706 67496 229711 67552
rect 229572 67494 229711 67496
rect 229572 67492 229578 67494
rect 229645 67491 229711 67494
rect 272149 64970 272215 64973
rect 272425 64970 272491 64973
rect 272149 64968 272491 64970
rect 272149 64912 272154 64968
rect 272210 64912 272430 64968
rect 272486 64912 272491 64968
rect 272149 64910 272491 64912
rect 272149 64907 272215 64910
rect 272425 64907 272491 64910
rect 287094 64834 287100 64836
rect 614 64774 287100 64834
rect -960 64562 480 64652
rect 614 64562 674 64774
rect 287094 64772 287100 64774
rect 287164 64772 287170 64836
rect -960 64502 674 64562
rect 579797 64562 579863 64565
rect 583520 64562 584960 64652
rect 579797 64560 584960 64562
rect 579797 64504 579802 64560
rect 579858 64504 584960 64560
rect 579797 64502 584960 64504
rect -960 64412 480 64502
rect 579797 64499 579863 64502
rect 583520 64412 584960 64502
rect 229645 58036 229711 58037
rect 229645 58032 229692 58036
rect 229756 58034 229762 58036
rect 229645 57976 229650 58032
rect 229645 57972 229692 57976
rect 229756 57974 229802 58034
rect 229756 57972 229762 57974
rect 229645 57971 229711 57972
rect 583520 52716 584960 52956
rect -960 50146 480 50236
rect 3049 50146 3115 50149
rect -960 50144 3115 50146
rect -960 50088 3054 50144
rect 3110 50088 3115 50144
rect -960 50086 3115 50088
rect -960 49996 480 50086
rect 3049 50083 3115 50086
rect 580165 41034 580231 41037
rect 583520 41034 584960 41124
rect 580165 41032 584960 41034
rect 580165 40976 580170 41032
rect 580226 40976 584960 41032
rect 580165 40974 584960 40976
rect 580165 40971 580231 40974
rect 583520 40884 584960 40974
rect -960 35866 480 35956
rect 3509 35866 3575 35869
rect -960 35864 3575 35866
rect -960 35808 3514 35864
rect 3570 35808 3575 35864
rect -960 35806 3575 35808
rect -960 35716 480 35806
rect 3509 35803 3575 35806
rect 497457 29474 497523 29477
rect 492630 29472 497523 29474
rect 492630 29416 497462 29472
rect 497518 29416 497523 29472
rect 492630 29414 497523 29416
rect 269062 29276 269068 29340
rect 269132 29338 269138 29340
rect 269132 29278 282930 29338
rect 269132 29276 269138 29278
rect 231710 29140 231716 29204
rect 231780 29202 231786 29204
rect 249742 29202 249748 29204
rect 231780 29142 249748 29202
rect 231780 29140 231786 29142
rect 249742 29140 249748 29142
rect 249812 29140 249818 29204
rect 249926 29004 249932 29068
rect 249996 29066 250002 29068
rect 269062 29066 269068 29068
rect 249996 29006 269068 29066
rect 249996 29004 250002 29006
rect 269062 29004 269068 29006
rect 269132 29004 269138 29068
rect 282870 29066 282930 29278
rect 335310 29278 344938 29338
rect 302141 29202 302207 29205
rect 321461 29202 321527 29205
rect 292622 29200 302207 29202
rect 292622 29144 302146 29200
rect 302202 29144 302207 29200
rect 292622 29142 302207 29144
rect 292622 29066 292682 29142
rect 302141 29139 302207 29142
rect 311942 29200 321527 29202
rect 311942 29144 321466 29200
rect 321522 29144 321527 29200
rect 311942 29142 321527 29144
rect 282870 29006 292682 29066
rect 309041 29066 309107 29069
rect 311942 29066 312002 29142
rect 321461 29139 321527 29142
rect 321645 29202 321711 29205
rect 321645 29200 331138 29202
rect 321645 29144 321650 29200
rect 321706 29144 331138 29200
rect 321645 29142 331138 29144
rect 321645 29139 321711 29142
rect 309041 29064 312002 29066
rect 309041 29008 309046 29064
rect 309102 29008 312002 29064
rect 309041 29006 312002 29008
rect 331078 29066 331138 29142
rect 335310 29066 335370 29278
rect 331078 29006 335370 29066
rect 344878 29066 344938 29278
rect 345062 29278 354690 29338
rect 345062 29066 345122 29278
rect 354630 29202 354690 29278
rect 364382 29278 374010 29338
rect 354630 29142 364258 29202
rect 344878 29006 345122 29066
rect 364198 29066 364258 29142
rect 364382 29066 364442 29278
rect 373950 29202 374010 29278
rect 383702 29278 405842 29338
rect 373950 29142 383578 29202
rect 364198 29006 364442 29066
rect 383518 29066 383578 29142
rect 383702 29066 383762 29278
rect 405782 29202 405842 29278
rect 415117 29202 415183 29205
rect 437381 29202 437447 29205
rect 456701 29202 456767 29205
rect 405782 29200 415183 29202
rect 405782 29144 415122 29200
rect 415178 29144 415183 29200
rect 405782 29142 415183 29144
rect 415117 29139 415183 29142
rect 427862 29200 437447 29202
rect 427862 29144 437386 29200
rect 437442 29144 437447 29200
rect 427862 29142 437447 29144
rect 383518 29006 383762 29066
rect 415301 29066 415367 29069
rect 427862 29066 427922 29142
rect 437381 29139 437447 29142
rect 447182 29200 456767 29202
rect 447182 29144 456706 29200
rect 456762 29144 456767 29200
rect 447182 29142 456767 29144
rect 415301 29064 427922 29066
rect 415301 29008 415306 29064
rect 415362 29008 427922 29064
rect 415301 29006 427922 29008
rect 444281 29066 444347 29069
rect 447182 29066 447242 29142
rect 456701 29139 456767 29142
rect 456885 29202 456951 29205
rect 491201 29202 491267 29205
rect 492630 29202 492690 29414
rect 497457 29411 497523 29414
rect 583520 29338 584960 29428
rect 583342 29278 584960 29338
rect 514661 29202 514727 29205
rect 533981 29202 534047 29205
rect 553301 29202 553367 29205
rect 572621 29202 572687 29205
rect 456885 29200 466378 29202
rect 456885 29144 456890 29200
rect 456946 29144 466378 29200
rect 456885 29142 466378 29144
rect 456885 29139 456951 29142
rect 444281 29064 447242 29066
rect 444281 29008 444286 29064
rect 444342 29008 447242 29064
rect 444281 29006 447242 29008
rect 466318 29066 466378 29142
rect 466502 29142 478154 29202
rect 466502 29066 466562 29142
rect 466318 29006 466562 29066
rect 478094 29066 478154 29142
rect 491201 29200 492690 29202
rect 491201 29144 491206 29200
rect 491262 29144 492690 29200
rect 491201 29142 492690 29144
rect 505142 29200 514727 29202
rect 505142 29144 514666 29200
rect 514722 29144 514727 29200
rect 505142 29142 514727 29144
rect 491201 29139 491267 29142
rect 481582 29066 481588 29068
rect 478094 29006 481588 29066
rect 309041 29003 309107 29006
rect 415301 29003 415367 29006
rect 444281 29003 444347 29006
rect 481582 29004 481588 29006
rect 481652 29004 481658 29068
rect 497457 29066 497523 29069
rect 505142 29066 505202 29142
rect 514661 29139 514727 29142
rect 524462 29200 534047 29202
rect 524462 29144 533986 29200
rect 534042 29144 534047 29200
rect 524462 29142 534047 29144
rect 497457 29064 505202 29066
rect 497457 29008 497462 29064
rect 497518 29008 505202 29064
rect 497457 29006 505202 29008
rect 521561 29066 521627 29069
rect 524462 29066 524522 29142
rect 533981 29139 534047 29142
rect 543782 29200 553367 29202
rect 543782 29144 553306 29200
rect 553362 29144 553367 29200
rect 543782 29142 553367 29144
rect 521561 29064 524522 29066
rect 521561 29008 521566 29064
rect 521622 29008 524522 29064
rect 521561 29006 524522 29008
rect 540881 29066 540947 29069
rect 543782 29066 543842 29142
rect 553301 29139 553367 29142
rect 563102 29200 572687 29202
rect 563102 29144 572626 29200
rect 572682 29144 572687 29200
rect 563102 29142 572687 29144
rect 540881 29064 543842 29066
rect 540881 29008 540886 29064
rect 540942 29008 543842 29064
rect 540881 29006 543842 29008
rect 560201 29066 560267 29069
rect 563102 29066 563162 29142
rect 572621 29139 572687 29142
rect 560201 29064 563162 29066
rect 560201 29008 560206 29064
rect 560262 29008 563162 29064
rect 560201 29006 563162 29008
rect 579521 29066 579587 29069
rect 583342 29066 583402 29278
rect 583520 29188 584960 29278
rect 579521 29064 583402 29066
rect 579521 29008 579526 29064
rect 579582 29008 583402 29064
rect 579521 29006 583402 29008
rect 497457 29003 497523 29006
rect 521561 29003 521627 29006
rect 540881 29003 540947 29006
rect 560201 29003 560267 29006
rect 579521 29003 579587 29006
rect 481582 28732 481588 28796
rect 481652 28794 481658 28796
rect 491201 28794 491267 28797
rect 481652 28792 491267 28794
rect 481652 28736 491206 28792
rect 491262 28736 491267 28792
rect 481652 28734 491267 28736
rect 481652 28732 481658 28734
rect 491201 28731 491267 28734
rect 240869 27570 240935 27573
rect 241053 27570 241119 27573
rect 240869 27568 241119 27570
rect 240869 27512 240874 27568
rect 240930 27512 241058 27568
rect 241114 27512 241119 27568
rect 240869 27510 241119 27512
rect 240869 27507 240935 27510
rect 241053 27507 241119 27510
rect -960 21450 480 21540
rect 3417 21450 3483 21453
rect -960 21448 3483 21450
rect -960 21392 3422 21448
rect 3478 21392 3483 21448
rect -960 21390 3483 21392
rect -960 21300 480 21390
rect 3417 21387 3483 21390
rect 260097 18050 260163 18053
rect 260373 18050 260439 18053
rect 260097 18048 260439 18050
rect 260097 17992 260102 18048
rect 260158 17992 260378 18048
rect 260434 17992 260439 18048
rect 260097 17990 260439 17992
rect 260097 17987 260163 17990
rect 260373 17987 260439 17990
rect 579797 17642 579863 17645
rect 583520 17642 584960 17732
rect 579797 17640 584960 17642
rect 579797 17584 579802 17640
rect 579858 17584 584960 17640
rect 579797 17582 584960 17584
rect 579797 17579 579863 17582
rect 583520 17492 584960 17582
rect -960 7170 480 7260
rect 3417 7170 3483 7173
rect -960 7168 3483 7170
rect -960 7112 3422 7168
rect 3478 7112 3483 7168
rect -960 7110 3483 7112
rect -960 7020 480 7110
rect 3417 7107 3483 7110
rect 583520 5796 584960 6036
rect 32673 4042 32739 4045
rect 234429 4042 234495 4045
rect 32673 4040 234495 4042
rect 32673 3984 32678 4040
rect 32734 3984 234434 4040
rect 234490 3984 234495 4040
rect 32673 3982 234495 3984
rect 32673 3979 32739 3982
rect 234429 3979 234495 3982
rect 277577 4042 277643 4045
rect 464429 4042 464495 4045
rect 277577 4040 464495 4042
rect 277577 3984 277582 4040
rect 277638 3984 464434 4040
rect 464490 3984 464495 4040
rect 277577 3982 464495 3984
rect 277577 3979 277643 3982
rect 464429 3979 464495 3982
rect 25497 3906 25563 3909
rect 232957 3906 233023 3909
rect 25497 3904 233023 3906
rect 25497 3848 25502 3904
rect 25558 3848 232962 3904
rect 233018 3848 233023 3904
rect 25497 3846 233023 3848
rect 25497 3843 25563 3846
rect 232957 3843 233023 3846
rect 277853 3906 277919 3909
rect 467925 3906 467991 3909
rect 277853 3904 467991 3906
rect 277853 3848 277858 3904
rect 277914 3848 467930 3904
rect 467986 3848 467991 3904
rect 277853 3846 467991 3848
rect 277853 3843 277919 3846
rect 467925 3843 467991 3846
rect 24301 3770 24367 3773
rect 232773 3770 232839 3773
rect 24301 3768 232839 3770
rect 24301 3712 24306 3768
rect 24362 3712 232778 3768
rect 232834 3712 232839 3768
rect 24301 3710 232839 3712
rect 24301 3707 24367 3710
rect 232773 3707 232839 3710
rect 278221 3770 278287 3773
rect 471513 3770 471579 3773
rect 278221 3768 471579 3770
rect 278221 3712 278226 3768
rect 278282 3712 471518 3768
rect 471574 3712 471579 3768
rect 278221 3710 471579 3712
rect 278221 3707 278287 3710
rect 471513 3707 471579 3710
rect 16021 3634 16087 3637
rect 231117 3634 231183 3637
rect 16021 3632 231183 3634
rect 16021 3576 16026 3632
rect 16082 3576 231122 3632
rect 231178 3576 231183 3632
rect 16021 3574 231183 3576
rect 16021 3571 16087 3574
rect 231117 3571 231183 3574
rect 279877 3634 279943 3637
rect 475101 3634 475167 3637
rect 279877 3632 475167 3634
rect 279877 3576 279882 3632
rect 279938 3576 475106 3632
rect 475162 3576 475167 3632
rect 279877 3574 475167 3576
rect 279877 3571 279943 3574
rect 475101 3571 475167 3574
rect 14825 3498 14891 3501
rect 230657 3498 230723 3501
rect 14825 3496 230723 3498
rect 14825 3440 14830 3496
rect 14886 3440 230662 3496
rect 230718 3440 230723 3496
rect 14825 3438 230723 3440
rect 14825 3435 14891 3438
rect 230657 3435 230723 3438
rect 230933 3498 230999 3501
rect 233233 3498 233299 3501
rect 230933 3496 233299 3498
rect 230933 3440 230938 3496
rect 230994 3440 233238 3496
rect 233294 3440 233299 3496
rect 230933 3438 233299 3440
rect 230933 3435 230999 3438
rect 233233 3435 233299 3438
rect 279969 3498 280035 3501
rect 478689 3498 478755 3501
rect 279969 3496 478755 3498
rect 279969 3440 279974 3496
rect 280030 3440 478694 3496
rect 478750 3440 478755 3496
rect 279969 3438 478755 3440
rect 279969 3435 280035 3438
rect 478689 3435 478755 3438
rect 6453 3362 6519 3365
rect 230565 3362 230631 3365
rect 6453 3360 230631 3362
rect 6453 3304 6458 3360
rect 6514 3304 230570 3360
rect 230626 3304 230631 3360
rect 6453 3302 230631 3304
rect 6453 3299 6519 3302
rect 230565 3299 230631 3302
rect 279785 3362 279851 3365
rect 482277 3362 482343 3365
rect 279785 3360 482343 3362
rect 279785 3304 279790 3360
rect 279846 3304 482282 3360
rect 482338 3304 482343 3360
rect 279785 3302 482343 3304
rect 279785 3299 279851 3302
rect 482277 3299 482343 3302
rect 229093 3226 229159 3229
rect 233785 3226 233851 3229
rect 229093 3224 233851 3226
rect 229093 3168 229098 3224
rect 229154 3168 233790 3224
rect 233846 3168 233851 3224
rect 229093 3166 233851 3168
rect 229093 3163 229159 3166
rect 233785 3163 233851 3166
<< via3 >>
rect 262812 401780 262876 401844
rect 243492 399468 243556 399532
rect 231716 399332 231780 399396
rect 233004 399392 233068 399396
rect 233004 399336 233018 399392
rect 233018 399336 233068 399392
rect 233004 399332 233068 399336
rect 233924 399332 233988 399396
rect 237236 399392 237300 399396
rect 237236 399336 237250 399392
rect 237250 399336 237300 399392
rect 237236 399332 237300 399336
rect 238156 399332 238220 399396
rect 239996 399332 240060 399396
rect 241284 399332 241348 399396
rect 282868 399332 282932 399396
rect 284340 399332 284404 399396
rect 285628 399332 285692 399396
rect 287100 399332 287164 399396
rect 238156 340036 238220 340100
rect 239996 338812 240060 338876
rect 233924 338676 233988 338740
rect 262812 335956 262876 336020
rect 275324 325620 275388 325684
rect 299428 322084 299492 322148
rect 357388 322084 357452 322148
rect 396028 322084 396092 322148
rect 243492 321540 243556 321604
rect 299428 321676 299492 321740
rect 357388 321676 357452 321740
rect 396028 321676 396092 321740
rect 275324 314876 275388 314940
rect 241284 310932 241348 310996
rect 257844 310932 257908 310996
rect 258028 310932 258092 310996
rect 257844 310660 257908 310724
rect 258028 310660 258092 310724
rect 560340 310796 560404 310860
rect 550588 310524 550652 310588
rect 560524 310660 560588 310724
rect 550588 310252 550652 310316
rect 237788 278700 237852 278764
rect 237788 264284 237852 264348
rect 237236 228108 237300 228172
rect 257844 227972 257908 228036
rect 257844 227564 257908 227628
rect 282868 194516 282932 194580
rect 284340 151676 284404 151740
rect 285628 108972 285692 109036
rect 233004 76196 233068 76260
rect 241468 76196 241532 76260
rect 260972 76060 261036 76124
rect 241468 75924 241532 75988
rect 260788 75924 260852 75988
rect 492628 76060 492692 76124
rect 492628 75788 492692 75852
rect 229508 67492 229572 67556
rect 287100 64772 287164 64836
rect 229692 58032 229756 58036
rect 229692 57976 229706 58032
rect 229706 57976 229756 58032
rect 229692 57972 229756 57976
rect 269068 29276 269132 29340
rect 231716 29140 231780 29204
rect 249748 29140 249812 29204
rect 249932 29004 249996 29068
rect 269068 29004 269132 29068
rect 481588 29004 481652 29068
rect 481588 28732 481652 28796
<< metal4 >>
rect -8436 711278 -7836 711300
rect -8436 711042 -8254 711278
rect -8018 711042 -7836 711278
rect -8436 710958 -7836 711042
rect -8436 710722 -8254 710958
rect -8018 710722 -7836 710958
rect -8436 679254 -7836 710722
rect -8436 679018 -8254 679254
rect -8018 679018 -7836 679254
rect -8436 678934 -7836 679018
rect -8436 678698 -8254 678934
rect -8018 678698 -7836 678934
rect -8436 643254 -7836 678698
rect -8436 643018 -8254 643254
rect -8018 643018 -7836 643254
rect -8436 642934 -7836 643018
rect -8436 642698 -8254 642934
rect -8018 642698 -7836 642934
rect -8436 607254 -7836 642698
rect -8436 607018 -8254 607254
rect -8018 607018 -7836 607254
rect -8436 606934 -7836 607018
rect -8436 606698 -8254 606934
rect -8018 606698 -7836 606934
rect -8436 571254 -7836 606698
rect -8436 571018 -8254 571254
rect -8018 571018 -7836 571254
rect -8436 570934 -7836 571018
rect -8436 570698 -8254 570934
rect -8018 570698 -7836 570934
rect -8436 535254 -7836 570698
rect -8436 535018 -8254 535254
rect -8018 535018 -7836 535254
rect -8436 534934 -7836 535018
rect -8436 534698 -8254 534934
rect -8018 534698 -7836 534934
rect -8436 499254 -7836 534698
rect -8436 499018 -8254 499254
rect -8018 499018 -7836 499254
rect -8436 498934 -7836 499018
rect -8436 498698 -8254 498934
rect -8018 498698 -7836 498934
rect -8436 463254 -7836 498698
rect -8436 463018 -8254 463254
rect -8018 463018 -7836 463254
rect -8436 462934 -7836 463018
rect -8436 462698 -8254 462934
rect -8018 462698 -7836 462934
rect -8436 427254 -7836 462698
rect -8436 427018 -8254 427254
rect -8018 427018 -7836 427254
rect -8436 426934 -7836 427018
rect -8436 426698 -8254 426934
rect -8018 426698 -7836 426934
rect -8436 391254 -7836 426698
rect -8436 391018 -8254 391254
rect -8018 391018 -7836 391254
rect -8436 390934 -7836 391018
rect -8436 390698 -8254 390934
rect -8018 390698 -7836 390934
rect -8436 355254 -7836 390698
rect -8436 355018 -8254 355254
rect -8018 355018 -7836 355254
rect -8436 354934 -7836 355018
rect -8436 354698 -8254 354934
rect -8018 354698 -7836 354934
rect -8436 319254 -7836 354698
rect -8436 319018 -8254 319254
rect -8018 319018 -7836 319254
rect -8436 318934 -7836 319018
rect -8436 318698 -8254 318934
rect -8018 318698 -7836 318934
rect -8436 283254 -7836 318698
rect -8436 283018 -8254 283254
rect -8018 283018 -7836 283254
rect -8436 282934 -7836 283018
rect -8436 282698 -8254 282934
rect -8018 282698 -7836 282934
rect -8436 247254 -7836 282698
rect -8436 247018 -8254 247254
rect -8018 247018 -7836 247254
rect -8436 246934 -7836 247018
rect -8436 246698 -8254 246934
rect -8018 246698 -7836 246934
rect -8436 211254 -7836 246698
rect -8436 211018 -8254 211254
rect -8018 211018 -7836 211254
rect -8436 210934 -7836 211018
rect -8436 210698 -8254 210934
rect -8018 210698 -7836 210934
rect -8436 175254 -7836 210698
rect -8436 175018 -8254 175254
rect -8018 175018 -7836 175254
rect -8436 174934 -7836 175018
rect -8436 174698 -8254 174934
rect -8018 174698 -7836 174934
rect -8436 139254 -7836 174698
rect -8436 139018 -8254 139254
rect -8018 139018 -7836 139254
rect -8436 138934 -7836 139018
rect -8436 138698 -8254 138934
rect -8018 138698 -7836 138934
rect -8436 103254 -7836 138698
rect -8436 103018 -8254 103254
rect -8018 103018 -7836 103254
rect -8436 102934 -7836 103018
rect -8436 102698 -8254 102934
rect -8018 102698 -7836 102934
rect -8436 67254 -7836 102698
rect -8436 67018 -8254 67254
rect -8018 67018 -7836 67254
rect -8436 66934 -7836 67018
rect -8436 66698 -8254 66934
rect -8018 66698 -7836 66934
rect -8436 31254 -7836 66698
rect -8436 31018 -8254 31254
rect -8018 31018 -7836 31254
rect -8436 30934 -7836 31018
rect -8436 30698 -8254 30934
rect -8018 30698 -7836 30934
rect -8436 -6786 -7836 30698
rect -7516 710358 -6916 710380
rect -7516 710122 -7334 710358
rect -7098 710122 -6916 710358
rect -7516 710038 -6916 710122
rect -7516 709802 -7334 710038
rect -7098 709802 -6916 710038
rect -7516 697254 -6916 709802
rect 11604 710358 12204 711300
rect 11604 710122 11786 710358
rect 12022 710122 12204 710358
rect 11604 710038 12204 710122
rect 11604 709802 11786 710038
rect 12022 709802 12204 710038
rect -7516 697018 -7334 697254
rect -7098 697018 -6916 697254
rect -7516 696934 -6916 697018
rect -7516 696698 -7334 696934
rect -7098 696698 -6916 696934
rect -7516 661254 -6916 696698
rect -7516 661018 -7334 661254
rect -7098 661018 -6916 661254
rect -7516 660934 -6916 661018
rect -7516 660698 -7334 660934
rect -7098 660698 -6916 660934
rect -7516 625254 -6916 660698
rect -7516 625018 -7334 625254
rect -7098 625018 -6916 625254
rect -7516 624934 -6916 625018
rect -7516 624698 -7334 624934
rect -7098 624698 -6916 624934
rect -7516 589254 -6916 624698
rect -7516 589018 -7334 589254
rect -7098 589018 -6916 589254
rect -7516 588934 -6916 589018
rect -7516 588698 -7334 588934
rect -7098 588698 -6916 588934
rect -7516 553254 -6916 588698
rect -7516 553018 -7334 553254
rect -7098 553018 -6916 553254
rect -7516 552934 -6916 553018
rect -7516 552698 -7334 552934
rect -7098 552698 -6916 552934
rect -7516 517254 -6916 552698
rect -7516 517018 -7334 517254
rect -7098 517018 -6916 517254
rect -7516 516934 -6916 517018
rect -7516 516698 -7334 516934
rect -7098 516698 -6916 516934
rect -7516 481254 -6916 516698
rect -7516 481018 -7334 481254
rect -7098 481018 -6916 481254
rect -7516 480934 -6916 481018
rect -7516 480698 -7334 480934
rect -7098 480698 -6916 480934
rect -7516 445254 -6916 480698
rect -7516 445018 -7334 445254
rect -7098 445018 -6916 445254
rect -7516 444934 -6916 445018
rect -7516 444698 -7334 444934
rect -7098 444698 -6916 444934
rect -7516 409254 -6916 444698
rect -7516 409018 -7334 409254
rect -7098 409018 -6916 409254
rect -7516 408934 -6916 409018
rect -7516 408698 -7334 408934
rect -7098 408698 -6916 408934
rect -7516 373254 -6916 408698
rect -7516 373018 -7334 373254
rect -7098 373018 -6916 373254
rect -7516 372934 -6916 373018
rect -7516 372698 -7334 372934
rect -7098 372698 -6916 372934
rect -7516 337254 -6916 372698
rect -7516 337018 -7334 337254
rect -7098 337018 -6916 337254
rect -7516 336934 -6916 337018
rect -7516 336698 -7334 336934
rect -7098 336698 -6916 336934
rect -7516 301254 -6916 336698
rect -7516 301018 -7334 301254
rect -7098 301018 -6916 301254
rect -7516 300934 -6916 301018
rect -7516 300698 -7334 300934
rect -7098 300698 -6916 300934
rect -7516 265254 -6916 300698
rect -7516 265018 -7334 265254
rect -7098 265018 -6916 265254
rect -7516 264934 -6916 265018
rect -7516 264698 -7334 264934
rect -7098 264698 -6916 264934
rect -7516 229254 -6916 264698
rect -7516 229018 -7334 229254
rect -7098 229018 -6916 229254
rect -7516 228934 -6916 229018
rect -7516 228698 -7334 228934
rect -7098 228698 -6916 228934
rect -7516 193254 -6916 228698
rect -7516 193018 -7334 193254
rect -7098 193018 -6916 193254
rect -7516 192934 -6916 193018
rect -7516 192698 -7334 192934
rect -7098 192698 -6916 192934
rect -7516 157254 -6916 192698
rect -7516 157018 -7334 157254
rect -7098 157018 -6916 157254
rect -7516 156934 -6916 157018
rect -7516 156698 -7334 156934
rect -7098 156698 -6916 156934
rect -7516 121254 -6916 156698
rect -7516 121018 -7334 121254
rect -7098 121018 -6916 121254
rect -7516 120934 -6916 121018
rect -7516 120698 -7334 120934
rect -7098 120698 -6916 120934
rect -7516 85254 -6916 120698
rect -7516 85018 -7334 85254
rect -7098 85018 -6916 85254
rect -7516 84934 -6916 85018
rect -7516 84698 -7334 84934
rect -7098 84698 -6916 84934
rect -7516 49254 -6916 84698
rect -7516 49018 -7334 49254
rect -7098 49018 -6916 49254
rect -7516 48934 -6916 49018
rect -7516 48698 -7334 48934
rect -7098 48698 -6916 48934
rect -7516 13254 -6916 48698
rect -7516 13018 -7334 13254
rect -7098 13018 -6916 13254
rect -7516 12934 -6916 13018
rect -7516 12698 -7334 12934
rect -7098 12698 -6916 12934
rect -7516 -5866 -6916 12698
rect -6596 709438 -5996 709460
rect -6596 709202 -6414 709438
rect -6178 709202 -5996 709438
rect -6596 709118 -5996 709202
rect -6596 708882 -6414 709118
rect -6178 708882 -5996 709118
rect -6596 675654 -5996 708882
rect -6596 675418 -6414 675654
rect -6178 675418 -5996 675654
rect -6596 675334 -5996 675418
rect -6596 675098 -6414 675334
rect -6178 675098 -5996 675334
rect -6596 639654 -5996 675098
rect -6596 639418 -6414 639654
rect -6178 639418 -5996 639654
rect -6596 639334 -5996 639418
rect -6596 639098 -6414 639334
rect -6178 639098 -5996 639334
rect -6596 603654 -5996 639098
rect -6596 603418 -6414 603654
rect -6178 603418 -5996 603654
rect -6596 603334 -5996 603418
rect -6596 603098 -6414 603334
rect -6178 603098 -5996 603334
rect -6596 567654 -5996 603098
rect -6596 567418 -6414 567654
rect -6178 567418 -5996 567654
rect -6596 567334 -5996 567418
rect -6596 567098 -6414 567334
rect -6178 567098 -5996 567334
rect -6596 531654 -5996 567098
rect -6596 531418 -6414 531654
rect -6178 531418 -5996 531654
rect -6596 531334 -5996 531418
rect -6596 531098 -6414 531334
rect -6178 531098 -5996 531334
rect -6596 495654 -5996 531098
rect -6596 495418 -6414 495654
rect -6178 495418 -5996 495654
rect -6596 495334 -5996 495418
rect -6596 495098 -6414 495334
rect -6178 495098 -5996 495334
rect -6596 459654 -5996 495098
rect -6596 459418 -6414 459654
rect -6178 459418 -5996 459654
rect -6596 459334 -5996 459418
rect -6596 459098 -6414 459334
rect -6178 459098 -5996 459334
rect -6596 423654 -5996 459098
rect -6596 423418 -6414 423654
rect -6178 423418 -5996 423654
rect -6596 423334 -5996 423418
rect -6596 423098 -6414 423334
rect -6178 423098 -5996 423334
rect -6596 387654 -5996 423098
rect -6596 387418 -6414 387654
rect -6178 387418 -5996 387654
rect -6596 387334 -5996 387418
rect -6596 387098 -6414 387334
rect -6178 387098 -5996 387334
rect -6596 351654 -5996 387098
rect -6596 351418 -6414 351654
rect -6178 351418 -5996 351654
rect -6596 351334 -5996 351418
rect -6596 351098 -6414 351334
rect -6178 351098 -5996 351334
rect -6596 315654 -5996 351098
rect -6596 315418 -6414 315654
rect -6178 315418 -5996 315654
rect -6596 315334 -5996 315418
rect -6596 315098 -6414 315334
rect -6178 315098 -5996 315334
rect -6596 279654 -5996 315098
rect -6596 279418 -6414 279654
rect -6178 279418 -5996 279654
rect -6596 279334 -5996 279418
rect -6596 279098 -6414 279334
rect -6178 279098 -5996 279334
rect -6596 243654 -5996 279098
rect -6596 243418 -6414 243654
rect -6178 243418 -5996 243654
rect -6596 243334 -5996 243418
rect -6596 243098 -6414 243334
rect -6178 243098 -5996 243334
rect -6596 207654 -5996 243098
rect -6596 207418 -6414 207654
rect -6178 207418 -5996 207654
rect -6596 207334 -5996 207418
rect -6596 207098 -6414 207334
rect -6178 207098 -5996 207334
rect -6596 171654 -5996 207098
rect -6596 171418 -6414 171654
rect -6178 171418 -5996 171654
rect -6596 171334 -5996 171418
rect -6596 171098 -6414 171334
rect -6178 171098 -5996 171334
rect -6596 135654 -5996 171098
rect -6596 135418 -6414 135654
rect -6178 135418 -5996 135654
rect -6596 135334 -5996 135418
rect -6596 135098 -6414 135334
rect -6178 135098 -5996 135334
rect -6596 99654 -5996 135098
rect -6596 99418 -6414 99654
rect -6178 99418 -5996 99654
rect -6596 99334 -5996 99418
rect -6596 99098 -6414 99334
rect -6178 99098 -5996 99334
rect -6596 63654 -5996 99098
rect -6596 63418 -6414 63654
rect -6178 63418 -5996 63654
rect -6596 63334 -5996 63418
rect -6596 63098 -6414 63334
rect -6178 63098 -5996 63334
rect -6596 27654 -5996 63098
rect -6596 27418 -6414 27654
rect -6178 27418 -5996 27654
rect -6596 27334 -5996 27418
rect -6596 27098 -6414 27334
rect -6178 27098 -5996 27334
rect -6596 -4946 -5996 27098
rect -5676 708518 -5076 708540
rect -5676 708282 -5494 708518
rect -5258 708282 -5076 708518
rect -5676 708198 -5076 708282
rect -5676 707962 -5494 708198
rect -5258 707962 -5076 708198
rect -5676 693654 -5076 707962
rect 8004 708518 8604 709460
rect 8004 708282 8186 708518
rect 8422 708282 8604 708518
rect 8004 708198 8604 708282
rect 8004 707962 8186 708198
rect 8422 707962 8604 708198
rect -5676 693418 -5494 693654
rect -5258 693418 -5076 693654
rect -5676 693334 -5076 693418
rect -5676 693098 -5494 693334
rect -5258 693098 -5076 693334
rect -5676 657654 -5076 693098
rect -5676 657418 -5494 657654
rect -5258 657418 -5076 657654
rect -5676 657334 -5076 657418
rect -5676 657098 -5494 657334
rect -5258 657098 -5076 657334
rect -5676 621654 -5076 657098
rect -5676 621418 -5494 621654
rect -5258 621418 -5076 621654
rect -5676 621334 -5076 621418
rect -5676 621098 -5494 621334
rect -5258 621098 -5076 621334
rect -5676 585654 -5076 621098
rect -5676 585418 -5494 585654
rect -5258 585418 -5076 585654
rect -5676 585334 -5076 585418
rect -5676 585098 -5494 585334
rect -5258 585098 -5076 585334
rect -5676 549654 -5076 585098
rect -5676 549418 -5494 549654
rect -5258 549418 -5076 549654
rect -5676 549334 -5076 549418
rect -5676 549098 -5494 549334
rect -5258 549098 -5076 549334
rect -5676 513654 -5076 549098
rect -5676 513418 -5494 513654
rect -5258 513418 -5076 513654
rect -5676 513334 -5076 513418
rect -5676 513098 -5494 513334
rect -5258 513098 -5076 513334
rect -5676 477654 -5076 513098
rect -5676 477418 -5494 477654
rect -5258 477418 -5076 477654
rect -5676 477334 -5076 477418
rect -5676 477098 -5494 477334
rect -5258 477098 -5076 477334
rect -5676 441654 -5076 477098
rect -5676 441418 -5494 441654
rect -5258 441418 -5076 441654
rect -5676 441334 -5076 441418
rect -5676 441098 -5494 441334
rect -5258 441098 -5076 441334
rect -5676 405654 -5076 441098
rect -5676 405418 -5494 405654
rect -5258 405418 -5076 405654
rect -5676 405334 -5076 405418
rect -5676 405098 -5494 405334
rect -5258 405098 -5076 405334
rect -5676 369654 -5076 405098
rect -5676 369418 -5494 369654
rect -5258 369418 -5076 369654
rect -5676 369334 -5076 369418
rect -5676 369098 -5494 369334
rect -5258 369098 -5076 369334
rect -5676 333654 -5076 369098
rect -5676 333418 -5494 333654
rect -5258 333418 -5076 333654
rect -5676 333334 -5076 333418
rect -5676 333098 -5494 333334
rect -5258 333098 -5076 333334
rect -5676 297654 -5076 333098
rect -5676 297418 -5494 297654
rect -5258 297418 -5076 297654
rect -5676 297334 -5076 297418
rect -5676 297098 -5494 297334
rect -5258 297098 -5076 297334
rect -5676 261654 -5076 297098
rect -5676 261418 -5494 261654
rect -5258 261418 -5076 261654
rect -5676 261334 -5076 261418
rect -5676 261098 -5494 261334
rect -5258 261098 -5076 261334
rect -5676 225654 -5076 261098
rect -5676 225418 -5494 225654
rect -5258 225418 -5076 225654
rect -5676 225334 -5076 225418
rect -5676 225098 -5494 225334
rect -5258 225098 -5076 225334
rect -5676 189654 -5076 225098
rect -5676 189418 -5494 189654
rect -5258 189418 -5076 189654
rect -5676 189334 -5076 189418
rect -5676 189098 -5494 189334
rect -5258 189098 -5076 189334
rect -5676 153654 -5076 189098
rect -5676 153418 -5494 153654
rect -5258 153418 -5076 153654
rect -5676 153334 -5076 153418
rect -5676 153098 -5494 153334
rect -5258 153098 -5076 153334
rect -5676 117654 -5076 153098
rect -5676 117418 -5494 117654
rect -5258 117418 -5076 117654
rect -5676 117334 -5076 117418
rect -5676 117098 -5494 117334
rect -5258 117098 -5076 117334
rect -5676 81654 -5076 117098
rect -5676 81418 -5494 81654
rect -5258 81418 -5076 81654
rect -5676 81334 -5076 81418
rect -5676 81098 -5494 81334
rect -5258 81098 -5076 81334
rect -5676 45654 -5076 81098
rect -5676 45418 -5494 45654
rect -5258 45418 -5076 45654
rect -5676 45334 -5076 45418
rect -5676 45098 -5494 45334
rect -5258 45098 -5076 45334
rect -5676 9654 -5076 45098
rect -5676 9418 -5494 9654
rect -5258 9418 -5076 9654
rect -5676 9334 -5076 9418
rect -5676 9098 -5494 9334
rect -5258 9098 -5076 9334
rect -5676 -4026 -5076 9098
rect -4756 707598 -4156 707620
rect -4756 707362 -4574 707598
rect -4338 707362 -4156 707598
rect -4756 707278 -4156 707362
rect -4756 707042 -4574 707278
rect -4338 707042 -4156 707278
rect -4756 672054 -4156 707042
rect -4756 671818 -4574 672054
rect -4338 671818 -4156 672054
rect -4756 671734 -4156 671818
rect -4756 671498 -4574 671734
rect -4338 671498 -4156 671734
rect -4756 636054 -4156 671498
rect -4756 635818 -4574 636054
rect -4338 635818 -4156 636054
rect -4756 635734 -4156 635818
rect -4756 635498 -4574 635734
rect -4338 635498 -4156 635734
rect -4756 600054 -4156 635498
rect -4756 599818 -4574 600054
rect -4338 599818 -4156 600054
rect -4756 599734 -4156 599818
rect -4756 599498 -4574 599734
rect -4338 599498 -4156 599734
rect -4756 564054 -4156 599498
rect -4756 563818 -4574 564054
rect -4338 563818 -4156 564054
rect -4756 563734 -4156 563818
rect -4756 563498 -4574 563734
rect -4338 563498 -4156 563734
rect -4756 528054 -4156 563498
rect -4756 527818 -4574 528054
rect -4338 527818 -4156 528054
rect -4756 527734 -4156 527818
rect -4756 527498 -4574 527734
rect -4338 527498 -4156 527734
rect -4756 492054 -4156 527498
rect -4756 491818 -4574 492054
rect -4338 491818 -4156 492054
rect -4756 491734 -4156 491818
rect -4756 491498 -4574 491734
rect -4338 491498 -4156 491734
rect -4756 456054 -4156 491498
rect -4756 455818 -4574 456054
rect -4338 455818 -4156 456054
rect -4756 455734 -4156 455818
rect -4756 455498 -4574 455734
rect -4338 455498 -4156 455734
rect -4756 420054 -4156 455498
rect -4756 419818 -4574 420054
rect -4338 419818 -4156 420054
rect -4756 419734 -4156 419818
rect -4756 419498 -4574 419734
rect -4338 419498 -4156 419734
rect -4756 384054 -4156 419498
rect -4756 383818 -4574 384054
rect -4338 383818 -4156 384054
rect -4756 383734 -4156 383818
rect -4756 383498 -4574 383734
rect -4338 383498 -4156 383734
rect -4756 348054 -4156 383498
rect -4756 347818 -4574 348054
rect -4338 347818 -4156 348054
rect -4756 347734 -4156 347818
rect -4756 347498 -4574 347734
rect -4338 347498 -4156 347734
rect -4756 312054 -4156 347498
rect -4756 311818 -4574 312054
rect -4338 311818 -4156 312054
rect -4756 311734 -4156 311818
rect -4756 311498 -4574 311734
rect -4338 311498 -4156 311734
rect -4756 276054 -4156 311498
rect -4756 275818 -4574 276054
rect -4338 275818 -4156 276054
rect -4756 275734 -4156 275818
rect -4756 275498 -4574 275734
rect -4338 275498 -4156 275734
rect -4756 240054 -4156 275498
rect -4756 239818 -4574 240054
rect -4338 239818 -4156 240054
rect -4756 239734 -4156 239818
rect -4756 239498 -4574 239734
rect -4338 239498 -4156 239734
rect -4756 204054 -4156 239498
rect -4756 203818 -4574 204054
rect -4338 203818 -4156 204054
rect -4756 203734 -4156 203818
rect -4756 203498 -4574 203734
rect -4338 203498 -4156 203734
rect -4756 168054 -4156 203498
rect -4756 167818 -4574 168054
rect -4338 167818 -4156 168054
rect -4756 167734 -4156 167818
rect -4756 167498 -4574 167734
rect -4338 167498 -4156 167734
rect -4756 132054 -4156 167498
rect -4756 131818 -4574 132054
rect -4338 131818 -4156 132054
rect -4756 131734 -4156 131818
rect -4756 131498 -4574 131734
rect -4338 131498 -4156 131734
rect -4756 96054 -4156 131498
rect -4756 95818 -4574 96054
rect -4338 95818 -4156 96054
rect -4756 95734 -4156 95818
rect -4756 95498 -4574 95734
rect -4338 95498 -4156 95734
rect -4756 60054 -4156 95498
rect -4756 59818 -4574 60054
rect -4338 59818 -4156 60054
rect -4756 59734 -4156 59818
rect -4756 59498 -4574 59734
rect -4338 59498 -4156 59734
rect -4756 24054 -4156 59498
rect -4756 23818 -4574 24054
rect -4338 23818 -4156 24054
rect -4756 23734 -4156 23818
rect -4756 23498 -4574 23734
rect -4338 23498 -4156 23734
rect -4756 -3106 -4156 23498
rect -3836 706678 -3236 706700
rect -3836 706442 -3654 706678
rect -3418 706442 -3236 706678
rect -3836 706358 -3236 706442
rect -3836 706122 -3654 706358
rect -3418 706122 -3236 706358
rect -3836 690054 -3236 706122
rect 4404 706678 5004 707620
rect 4404 706442 4586 706678
rect 4822 706442 5004 706678
rect 4404 706358 5004 706442
rect 4404 706122 4586 706358
rect 4822 706122 5004 706358
rect -3836 689818 -3654 690054
rect -3418 689818 -3236 690054
rect -3836 689734 -3236 689818
rect -3836 689498 -3654 689734
rect -3418 689498 -3236 689734
rect -3836 654054 -3236 689498
rect -3836 653818 -3654 654054
rect -3418 653818 -3236 654054
rect -3836 653734 -3236 653818
rect -3836 653498 -3654 653734
rect -3418 653498 -3236 653734
rect -3836 618054 -3236 653498
rect -3836 617818 -3654 618054
rect -3418 617818 -3236 618054
rect -3836 617734 -3236 617818
rect -3836 617498 -3654 617734
rect -3418 617498 -3236 617734
rect -3836 582054 -3236 617498
rect -3836 581818 -3654 582054
rect -3418 581818 -3236 582054
rect -3836 581734 -3236 581818
rect -3836 581498 -3654 581734
rect -3418 581498 -3236 581734
rect -3836 546054 -3236 581498
rect -3836 545818 -3654 546054
rect -3418 545818 -3236 546054
rect -3836 545734 -3236 545818
rect -3836 545498 -3654 545734
rect -3418 545498 -3236 545734
rect -3836 510054 -3236 545498
rect -3836 509818 -3654 510054
rect -3418 509818 -3236 510054
rect -3836 509734 -3236 509818
rect -3836 509498 -3654 509734
rect -3418 509498 -3236 509734
rect -3836 474054 -3236 509498
rect -3836 473818 -3654 474054
rect -3418 473818 -3236 474054
rect -3836 473734 -3236 473818
rect -3836 473498 -3654 473734
rect -3418 473498 -3236 473734
rect -3836 438054 -3236 473498
rect -3836 437818 -3654 438054
rect -3418 437818 -3236 438054
rect -3836 437734 -3236 437818
rect -3836 437498 -3654 437734
rect -3418 437498 -3236 437734
rect -3836 402054 -3236 437498
rect -3836 401818 -3654 402054
rect -3418 401818 -3236 402054
rect -3836 401734 -3236 401818
rect -3836 401498 -3654 401734
rect -3418 401498 -3236 401734
rect -3836 366054 -3236 401498
rect -3836 365818 -3654 366054
rect -3418 365818 -3236 366054
rect -3836 365734 -3236 365818
rect -3836 365498 -3654 365734
rect -3418 365498 -3236 365734
rect -3836 330054 -3236 365498
rect -3836 329818 -3654 330054
rect -3418 329818 -3236 330054
rect -3836 329734 -3236 329818
rect -3836 329498 -3654 329734
rect -3418 329498 -3236 329734
rect -3836 294054 -3236 329498
rect -3836 293818 -3654 294054
rect -3418 293818 -3236 294054
rect -3836 293734 -3236 293818
rect -3836 293498 -3654 293734
rect -3418 293498 -3236 293734
rect -3836 258054 -3236 293498
rect -3836 257818 -3654 258054
rect -3418 257818 -3236 258054
rect -3836 257734 -3236 257818
rect -3836 257498 -3654 257734
rect -3418 257498 -3236 257734
rect -3836 222054 -3236 257498
rect -3836 221818 -3654 222054
rect -3418 221818 -3236 222054
rect -3836 221734 -3236 221818
rect -3836 221498 -3654 221734
rect -3418 221498 -3236 221734
rect -3836 186054 -3236 221498
rect -3836 185818 -3654 186054
rect -3418 185818 -3236 186054
rect -3836 185734 -3236 185818
rect -3836 185498 -3654 185734
rect -3418 185498 -3236 185734
rect -3836 150054 -3236 185498
rect -3836 149818 -3654 150054
rect -3418 149818 -3236 150054
rect -3836 149734 -3236 149818
rect -3836 149498 -3654 149734
rect -3418 149498 -3236 149734
rect -3836 114054 -3236 149498
rect -3836 113818 -3654 114054
rect -3418 113818 -3236 114054
rect -3836 113734 -3236 113818
rect -3836 113498 -3654 113734
rect -3418 113498 -3236 113734
rect -3836 78054 -3236 113498
rect -3836 77818 -3654 78054
rect -3418 77818 -3236 78054
rect -3836 77734 -3236 77818
rect -3836 77498 -3654 77734
rect -3418 77498 -3236 77734
rect -3836 42054 -3236 77498
rect -3836 41818 -3654 42054
rect -3418 41818 -3236 42054
rect -3836 41734 -3236 41818
rect -3836 41498 -3654 41734
rect -3418 41498 -3236 41734
rect -3836 6054 -3236 41498
rect -3836 5818 -3654 6054
rect -3418 5818 -3236 6054
rect -3836 5734 -3236 5818
rect -3836 5498 -3654 5734
rect -3418 5498 -3236 5734
rect -3836 -2186 -3236 5498
rect -2916 705758 -2316 705780
rect -2916 705522 -2734 705758
rect -2498 705522 -2316 705758
rect -2916 705438 -2316 705522
rect -2916 705202 -2734 705438
rect -2498 705202 -2316 705438
rect -2916 668454 -2316 705202
rect -2916 668218 -2734 668454
rect -2498 668218 -2316 668454
rect -2916 668134 -2316 668218
rect -2916 667898 -2734 668134
rect -2498 667898 -2316 668134
rect -2916 632454 -2316 667898
rect -2916 632218 -2734 632454
rect -2498 632218 -2316 632454
rect -2916 632134 -2316 632218
rect -2916 631898 -2734 632134
rect -2498 631898 -2316 632134
rect -2916 596454 -2316 631898
rect -2916 596218 -2734 596454
rect -2498 596218 -2316 596454
rect -2916 596134 -2316 596218
rect -2916 595898 -2734 596134
rect -2498 595898 -2316 596134
rect -2916 560454 -2316 595898
rect -2916 560218 -2734 560454
rect -2498 560218 -2316 560454
rect -2916 560134 -2316 560218
rect -2916 559898 -2734 560134
rect -2498 559898 -2316 560134
rect -2916 524454 -2316 559898
rect -2916 524218 -2734 524454
rect -2498 524218 -2316 524454
rect -2916 524134 -2316 524218
rect -2916 523898 -2734 524134
rect -2498 523898 -2316 524134
rect -2916 488454 -2316 523898
rect -2916 488218 -2734 488454
rect -2498 488218 -2316 488454
rect -2916 488134 -2316 488218
rect -2916 487898 -2734 488134
rect -2498 487898 -2316 488134
rect -2916 452454 -2316 487898
rect -2916 452218 -2734 452454
rect -2498 452218 -2316 452454
rect -2916 452134 -2316 452218
rect -2916 451898 -2734 452134
rect -2498 451898 -2316 452134
rect -2916 416454 -2316 451898
rect -2916 416218 -2734 416454
rect -2498 416218 -2316 416454
rect -2916 416134 -2316 416218
rect -2916 415898 -2734 416134
rect -2498 415898 -2316 416134
rect -2916 380454 -2316 415898
rect -2916 380218 -2734 380454
rect -2498 380218 -2316 380454
rect -2916 380134 -2316 380218
rect -2916 379898 -2734 380134
rect -2498 379898 -2316 380134
rect -2916 344454 -2316 379898
rect -2916 344218 -2734 344454
rect -2498 344218 -2316 344454
rect -2916 344134 -2316 344218
rect -2916 343898 -2734 344134
rect -2498 343898 -2316 344134
rect -2916 308454 -2316 343898
rect -2916 308218 -2734 308454
rect -2498 308218 -2316 308454
rect -2916 308134 -2316 308218
rect -2916 307898 -2734 308134
rect -2498 307898 -2316 308134
rect -2916 272454 -2316 307898
rect -2916 272218 -2734 272454
rect -2498 272218 -2316 272454
rect -2916 272134 -2316 272218
rect -2916 271898 -2734 272134
rect -2498 271898 -2316 272134
rect -2916 236454 -2316 271898
rect -2916 236218 -2734 236454
rect -2498 236218 -2316 236454
rect -2916 236134 -2316 236218
rect -2916 235898 -2734 236134
rect -2498 235898 -2316 236134
rect -2916 200454 -2316 235898
rect -2916 200218 -2734 200454
rect -2498 200218 -2316 200454
rect -2916 200134 -2316 200218
rect -2916 199898 -2734 200134
rect -2498 199898 -2316 200134
rect -2916 164454 -2316 199898
rect -2916 164218 -2734 164454
rect -2498 164218 -2316 164454
rect -2916 164134 -2316 164218
rect -2916 163898 -2734 164134
rect -2498 163898 -2316 164134
rect -2916 128454 -2316 163898
rect -2916 128218 -2734 128454
rect -2498 128218 -2316 128454
rect -2916 128134 -2316 128218
rect -2916 127898 -2734 128134
rect -2498 127898 -2316 128134
rect -2916 92454 -2316 127898
rect -2916 92218 -2734 92454
rect -2498 92218 -2316 92454
rect -2916 92134 -2316 92218
rect -2916 91898 -2734 92134
rect -2498 91898 -2316 92134
rect -2916 56454 -2316 91898
rect -2916 56218 -2734 56454
rect -2498 56218 -2316 56454
rect -2916 56134 -2316 56218
rect -2916 55898 -2734 56134
rect -2498 55898 -2316 56134
rect -2916 20454 -2316 55898
rect -2916 20218 -2734 20454
rect -2498 20218 -2316 20454
rect -2916 20134 -2316 20218
rect -2916 19898 -2734 20134
rect -2498 19898 -2316 20134
rect -2916 -1266 -2316 19898
rect -1996 704838 -1396 704860
rect -1996 704602 -1814 704838
rect -1578 704602 -1396 704838
rect -1996 704518 -1396 704602
rect -1996 704282 -1814 704518
rect -1578 704282 -1396 704518
rect -1996 686454 -1396 704282
rect -1996 686218 -1814 686454
rect -1578 686218 -1396 686454
rect -1996 686134 -1396 686218
rect -1996 685898 -1814 686134
rect -1578 685898 -1396 686134
rect -1996 650454 -1396 685898
rect -1996 650218 -1814 650454
rect -1578 650218 -1396 650454
rect -1996 650134 -1396 650218
rect -1996 649898 -1814 650134
rect -1578 649898 -1396 650134
rect -1996 614454 -1396 649898
rect -1996 614218 -1814 614454
rect -1578 614218 -1396 614454
rect -1996 614134 -1396 614218
rect -1996 613898 -1814 614134
rect -1578 613898 -1396 614134
rect -1996 578454 -1396 613898
rect -1996 578218 -1814 578454
rect -1578 578218 -1396 578454
rect -1996 578134 -1396 578218
rect -1996 577898 -1814 578134
rect -1578 577898 -1396 578134
rect -1996 542454 -1396 577898
rect -1996 542218 -1814 542454
rect -1578 542218 -1396 542454
rect -1996 542134 -1396 542218
rect -1996 541898 -1814 542134
rect -1578 541898 -1396 542134
rect -1996 506454 -1396 541898
rect -1996 506218 -1814 506454
rect -1578 506218 -1396 506454
rect -1996 506134 -1396 506218
rect -1996 505898 -1814 506134
rect -1578 505898 -1396 506134
rect -1996 470454 -1396 505898
rect -1996 470218 -1814 470454
rect -1578 470218 -1396 470454
rect -1996 470134 -1396 470218
rect -1996 469898 -1814 470134
rect -1578 469898 -1396 470134
rect -1996 434454 -1396 469898
rect -1996 434218 -1814 434454
rect -1578 434218 -1396 434454
rect -1996 434134 -1396 434218
rect -1996 433898 -1814 434134
rect -1578 433898 -1396 434134
rect -1996 398454 -1396 433898
rect -1996 398218 -1814 398454
rect -1578 398218 -1396 398454
rect -1996 398134 -1396 398218
rect -1996 397898 -1814 398134
rect -1578 397898 -1396 398134
rect -1996 362454 -1396 397898
rect -1996 362218 -1814 362454
rect -1578 362218 -1396 362454
rect -1996 362134 -1396 362218
rect -1996 361898 -1814 362134
rect -1578 361898 -1396 362134
rect -1996 326454 -1396 361898
rect -1996 326218 -1814 326454
rect -1578 326218 -1396 326454
rect -1996 326134 -1396 326218
rect -1996 325898 -1814 326134
rect -1578 325898 -1396 326134
rect -1996 290454 -1396 325898
rect -1996 290218 -1814 290454
rect -1578 290218 -1396 290454
rect -1996 290134 -1396 290218
rect -1996 289898 -1814 290134
rect -1578 289898 -1396 290134
rect -1996 254454 -1396 289898
rect -1996 254218 -1814 254454
rect -1578 254218 -1396 254454
rect -1996 254134 -1396 254218
rect -1996 253898 -1814 254134
rect -1578 253898 -1396 254134
rect -1996 218454 -1396 253898
rect -1996 218218 -1814 218454
rect -1578 218218 -1396 218454
rect -1996 218134 -1396 218218
rect -1996 217898 -1814 218134
rect -1578 217898 -1396 218134
rect -1996 182454 -1396 217898
rect -1996 182218 -1814 182454
rect -1578 182218 -1396 182454
rect -1996 182134 -1396 182218
rect -1996 181898 -1814 182134
rect -1578 181898 -1396 182134
rect -1996 146454 -1396 181898
rect -1996 146218 -1814 146454
rect -1578 146218 -1396 146454
rect -1996 146134 -1396 146218
rect -1996 145898 -1814 146134
rect -1578 145898 -1396 146134
rect -1996 110454 -1396 145898
rect -1996 110218 -1814 110454
rect -1578 110218 -1396 110454
rect -1996 110134 -1396 110218
rect -1996 109898 -1814 110134
rect -1578 109898 -1396 110134
rect -1996 74454 -1396 109898
rect -1996 74218 -1814 74454
rect -1578 74218 -1396 74454
rect -1996 74134 -1396 74218
rect -1996 73898 -1814 74134
rect -1578 73898 -1396 74134
rect -1996 38454 -1396 73898
rect -1996 38218 -1814 38454
rect -1578 38218 -1396 38454
rect -1996 38134 -1396 38218
rect -1996 37898 -1814 38134
rect -1578 37898 -1396 38134
rect -1996 2454 -1396 37898
rect -1996 2218 -1814 2454
rect -1578 2218 -1396 2454
rect -1996 2134 -1396 2218
rect -1996 1898 -1814 2134
rect -1578 1898 -1396 2134
rect -1996 -346 -1396 1898
rect -1996 -582 -1814 -346
rect -1578 -582 -1396 -346
rect -1996 -666 -1396 -582
rect -1996 -902 -1814 -666
rect -1578 -902 -1396 -666
rect -1996 -924 -1396 -902
rect 804 704838 1404 705780
rect 804 704602 986 704838
rect 1222 704602 1404 704838
rect 804 704518 1404 704602
rect 804 704282 986 704518
rect 1222 704282 1404 704518
rect 804 686454 1404 704282
rect 804 686218 986 686454
rect 1222 686218 1404 686454
rect 804 686134 1404 686218
rect 804 685898 986 686134
rect 1222 685898 1404 686134
rect 804 650454 1404 685898
rect 804 650218 986 650454
rect 1222 650218 1404 650454
rect 804 650134 1404 650218
rect 804 649898 986 650134
rect 1222 649898 1404 650134
rect 804 614454 1404 649898
rect 804 614218 986 614454
rect 1222 614218 1404 614454
rect 804 614134 1404 614218
rect 804 613898 986 614134
rect 1222 613898 1404 614134
rect 804 578454 1404 613898
rect 804 578218 986 578454
rect 1222 578218 1404 578454
rect 804 578134 1404 578218
rect 804 577898 986 578134
rect 1222 577898 1404 578134
rect 804 542454 1404 577898
rect 804 542218 986 542454
rect 1222 542218 1404 542454
rect 804 542134 1404 542218
rect 804 541898 986 542134
rect 1222 541898 1404 542134
rect 804 506454 1404 541898
rect 804 506218 986 506454
rect 1222 506218 1404 506454
rect 804 506134 1404 506218
rect 804 505898 986 506134
rect 1222 505898 1404 506134
rect 804 470454 1404 505898
rect 804 470218 986 470454
rect 1222 470218 1404 470454
rect 804 470134 1404 470218
rect 804 469898 986 470134
rect 1222 469898 1404 470134
rect 804 434454 1404 469898
rect 804 434218 986 434454
rect 1222 434218 1404 434454
rect 804 434134 1404 434218
rect 804 433898 986 434134
rect 1222 433898 1404 434134
rect 804 398454 1404 433898
rect 804 398218 986 398454
rect 1222 398218 1404 398454
rect 804 398134 1404 398218
rect 804 397898 986 398134
rect 1222 397898 1404 398134
rect 804 362454 1404 397898
rect 804 362218 986 362454
rect 1222 362218 1404 362454
rect 804 362134 1404 362218
rect 804 361898 986 362134
rect 1222 361898 1404 362134
rect 804 326454 1404 361898
rect 804 326218 986 326454
rect 1222 326218 1404 326454
rect 804 326134 1404 326218
rect 804 325898 986 326134
rect 1222 325898 1404 326134
rect 804 290454 1404 325898
rect 804 290218 986 290454
rect 1222 290218 1404 290454
rect 804 290134 1404 290218
rect 804 289898 986 290134
rect 1222 289898 1404 290134
rect 804 254454 1404 289898
rect 804 254218 986 254454
rect 1222 254218 1404 254454
rect 804 254134 1404 254218
rect 804 253898 986 254134
rect 1222 253898 1404 254134
rect 804 218454 1404 253898
rect 804 218218 986 218454
rect 1222 218218 1404 218454
rect 804 218134 1404 218218
rect 804 217898 986 218134
rect 1222 217898 1404 218134
rect 804 182454 1404 217898
rect 804 182218 986 182454
rect 1222 182218 1404 182454
rect 804 182134 1404 182218
rect 804 181898 986 182134
rect 1222 181898 1404 182134
rect 804 146454 1404 181898
rect 804 146218 986 146454
rect 1222 146218 1404 146454
rect 804 146134 1404 146218
rect 804 145898 986 146134
rect 1222 145898 1404 146134
rect 804 110454 1404 145898
rect 804 110218 986 110454
rect 1222 110218 1404 110454
rect 804 110134 1404 110218
rect 804 109898 986 110134
rect 1222 109898 1404 110134
rect 804 74454 1404 109898
rect 804 74218 986 74454
rect 1222 74218 1404 74454
rect 804 74134 1404 74218
rect 804 73898 986 74134
rect 1222 73898 1404 74134
rect 804 38454 1404 73898
rect 804 38218 986 38454
rect 1222 38218 1404 38454
rect 804 38134 1404 38218
rect 804 37898 986 38134
rect 1222 37898 1404 38134
rect 804 2454 1404 37898
rect 804 2218 986 2454
rect 1222 2218 1404 2454
rect 804 2134 1404 2218
rect 804 1898 986 2134
rect 1222 1898 1404 2134
rect 804 -346 1404 1898
rect 804 -582 986 -346
rect 1222 -582 1404 -346
rect 804 -666 1404 -582
rect 804 -902 986 -666
rect 1222 -902 1404 -666
rect -2916 -1502 -2734 -1266
rect -2498 -1502 -2316 -1266
rect -2916 -1586 -2316 -1502
rect -2916 -1822 -2734 -1586
rect -2498 -1822 -2316 -1586
rect -2916 -1844 -2316 -1822
rect 804 -1844 1404 -902
rect 4404 690054 5004 706122
rect 4404 689818 4586 690054
rect 4822 689818 5004 690054
rect 4404 689734 5004 689818
rect 4404 689498 4586 689734
rect 4822 689498 5004 689734
rect 4404 654054 5004 689498
rect 4404 653818 4586 654054
rect 4822 653818 5004 654054
rect 4404 653734 5004 653818
rect 4404 653498 4586 653734
rect 4822 653498 5004 653734
rect 4404 618054 5004 653498
rect 4404 617818 4586 618054
rect 4822 617818 5004 618054
rect 4404 617734 5004 617818
rect 4404 617498 4586 617734
rect 4822 617498 5004 617734
rect 4404 582054 5004 617498
rect 4404 581818 4586 582054
rect 4822 581818 5004 582054
rect 4404 581734 5004 581818
rect 4404 581498 4586 581734
rect 4822 581498 5004 581734
rect 4404 546054 5004 581498
rect 4404 545818 4586 546054
rect 4822 545818 5004 546054
rect 4404 545734 5004 545818
rect 4404 545498 4586 545734
rect 4822 545498 5004 545734
rect 4404 510054 5004 545498
rect 4404 509818 4586 510054
rect 4822 509818 5004 510054
rect 4404 509734 5004 509818
rect 4404 509498 4586 509734
rect 4822 509498 5004 509734
rect 4404 474054 5004 509498
rect 4404 473818 4586 474054
rect 4822 473818 5004 474054
rect 4404 473734 5004 473818
rect 4404 473498 4586 473734
rect 4822 473498 5004 473734
rect 4404 438054 5004 473498
rect 4404 437818 4586 438054
rect 4822 437818 5004 438054
rect 4404 437734 5004 437818
rect 4404 437498 4586 437734
rect 4822 437498 5004 437734
rect 4404 402054 5004 437498
rect 4404 401818 4586 402054
rect 4822 401818 5004 402054
rect 4404 401734 5004 401818
rect 4404 401498 4586 401734
rect 4822 401498 5004 401734
rect 4404 366054 5004 401498
rect 4404 365818 4586 366054
rect 4822 365818 5004 366054
rect 4404 365734 5004 365818
rect 4404 365498 4586 365734
rect 4822 365498 5004 365734
rect 4404 330054 5004 365498
rect 4404 329818 4586 330054
rect 4822 329818 5004 330054
rect 4404 329734 5004 329818
rect 4404 329498 4586 329734
rect 4822 329498 5004 329734
rect 4404 294054 5004 329498
rect 4404 293818 4586 294054
rect 4822 293818 5004 294054
rect 4404 293734 5004 293818
rect 4404 293498 4586 293734
rect 4822 293498 5004 293734
rect 4404 258054 5004 293498
rect 4404 257818 4586 258054
rect 4822 257818 5004 258054
rect 4404 257734 5004 257818
rect 4404 257498 4586 257734
rect 4822 257498 5004 257734
rect 4404 222054 5004 257498
rect 4404 221818 4586 222054
rect 4822 221818 5004 222054
rect 4404 221734 5004 221818
rect 4404 221498 4586 221734
rect 4822 221498 5004 221734
rect 4404 186054 5004 221498
rect 4404 185818 4586 186054
rect 4822 185818 5004 186054
rect 4404 185734 5004 185818
rect 4404 185498 4586 185734
rect 4822 185498 5004 185734
rect 4404 150054 5004 185498
rect 4404 149818 4586 150054
rect 4822 149818 5004 150054
rect 4404 149734 5004 149818
rect 4404 149498 4586 149734
rect 4822 149498 5004 149734
rect 4404 114054 5004 149498
rect 4404 113818 4586 114054
rect 4822 113818 5004 114054
rect 4404 113734 5004 113818
rect 4404 113498 4586 113734
rect 4822 113498 5004 113734
rect 4404 78054 5004 113498
rect 4404 77818 4586 78054
rect 4822 77818 5004 78054
rect 4404 77734 5004 77818
rect 4404 77498 4586 77734
rect 4822 77498 5004 77734
rect 4404 42054 5004 77498
rect 4404 41818 4586 42054
rect 4822 41818 5004 42054
rect 4404 41734 5004 41818
rect 4404 41498 4586 41734
rect 4822 41498 5004 41734
rect 4404 6054 5004 41498
rect 4404 5818 4586 6054
rect 4822 5818 5004 6054
rect 4404 5734 5004 5818
rect 4404 5498 4586 5734
rect 4822 5498 5004 5734
rect -3836 -2422 -3654 -2186
rect -3418 -2422 -3236 -2186
rect -3836 -2506 -3236 -2422
rect -3836 -2742 -3654 -2506
rect -3418 -2742 -3236 -2506
rect -3836 -2764 -3236 -2742
rect 4404 -2186 5004 5498
rect 4404 -2422 4586 -2186
rect 4822 -2422 5004 -2186
rect 4404 -2506 5004 -2422
rect 4404 -2742 4586 -2506
rect 4822 -2742 5004 -2506
rect -4756 -3342 -4574 -3106
rect -4338 -3342 -4156 -3106
rect -4756 -3426 -4156 -3342
rect -4756 -3662 -4574 -3426
rect -4338 -3662 -4156 -3426
rect -4756 -3684 -4156 -3662
rect 4404 -3684 5004 -2742
rect 8004 693654 8604 707962
rect 8004 693418 8186 693654
rect 8422 693418 8604 693654
rect 8004 693334 8604 693418
rect 8004 693098 8186 693334
rect 8422 693098 8604 693334
rect 8004 657654 8604 693098
rect 8004 657418 8186 657654
rect 8422 657418 8604 657654
rect 8004 657334 8604 657418
rect 8004 657098 8186 657334
rect 8422 657098 8604 657334
rect 8004 621654 8604 657098
rect 8004 621418 8186 621654
rect 8422 621418 8604 621654
rect 8004 621334 8604 621418
rect 8004 621098 8186 621334
rect 8422 621098 8604 621334
rect 8004 585654 8604 621098
rect 8004 585418 8186 585654
rect 8422 585418 8604 585654
rect 8004 585334 8604 585418
rect 8004 585098 8186 585334
rect 8422 585098 8604 585334
rect 8004 549654 8604 585098
rect 8004 549418 8186 549654
rect 8422 549418 8604 549654
rect 8004 549334 8604 549418
rect 8004 549098 8186 549334
rect 8422 549098 8604 549334
rect 8004 513654 8604 549098
rect 8004 513418 8186 513654
rect 8422 513418 8604 513654
rect 8004 513334 8604 513418
rect 8004 513098 8186 513334
rect 8422 513098 8604 513334
rect 8004 477654 8604 513098
rect 8004 477418 8186 477654
rect 8422 477418 8604 477654
rect 8004 477334 8604 477418
rect 8004 477098 8186 477334
rect 8422 477098 8604 477334
rect 8004 441654 8604 477098
rect 8004 441418 8186 441654
rect 8422 441418 8604 441654
rect 8004 441334 8604 441418
rect 8004 441098 8186 441334
rect 8422 441098 8604 441334
rect 8004 405654 8604 441098
rect 8004 405418 8186 405654
rect 8422 405418 8604 405654
rect 8004 405334 8604 405418
rect 8004 405098 8186 405334
rect 8422 405098 8604 405334
rect 8004 369654 8604 405098
rect 8004 369418 8186 369654
rect 8422 369418 8604 369654
rect 8004 369334 8604 369418
rect 8004 369098 8186 369334
rect 8422 369098 8604 369334
rect 8004 333654 8604 369098
rect 8004 333418 8186 333654
rect 8422 333418 8604 333654
rect 8004 333334 8604 333418
rect 8004 333098 8186 333334
rect 8422 333098 8604 333334
rect 8004 297654 8604 333098
rect 8004 297418 8186 297654
rect 8422 297418 8604 297654
rect 8004 297334 8604 297418
rect 8004 297098 8186 297334
rect 8422 297098 8604 297334
rect 8004 261654 8604 297098
rect 8004 261418 8186 261654
rect 8422 261418 8604 261654
rect 8004 261334 8604 261418
rect 8004 261098 8186 261334
rect 8422 261098 8604 261334
rect 8004 225654 8604 261098
rect 8004 225418 8186 225654
rect 8422 225418 8604 225654
rect 8004 225334 8604 225418
rect 8004 225098 8186 225334
rect 8422 225098 8604 225334
rect 8004 189654 8604 225098
rect 8004 189418 8186 189654
rect 8422 189418 8604 189654
rect 8004 189334 8604 189418
rect 8004 189098 8186 189334
rect 8422 189098 8604 189334
rect 8004 153654 8604 189098
rect 8004 153418 8186 153654
rect 8422 153418 8604 153654
rect 8004 153334 8604 153418
rect 8004 153098 8186 153334
rect 8422 153098 8604 153334
rect 8004 117654 8604 153098
rect 8004 117418 8186 117654
rect 8422 117418 8604 117654
rect 8004 117334 8604 117418
rect 8004 117098 8186 117334
rect 8422 117098 8604 117334
rect 8004 81654 8604 117098
rect 8004 81418 8186 81654
rect 8422 81418 8604 81654
rect 8004 81334 8604 81418
rect 8004 81098 8186 81334
rect 8422 81098 8604 81334
rect 8004 45654 8604 81098
rect 8004 45418 8186 45654
rect 8422 45418 8604 45654
rect 8004 45334 8604 45418
rect 8004 45098 8186 45334
rect 8422 45098 8604 45334
rect 8004 9654 8604 45098
rect 8004 9418 8186 9654
rect 8422 9418 8604 9654
rect 8004 9334 8604 9418
rect 8004 9098 8186 9334
rect 8422 9098 8604 9334
rect -5676 -4262 -5494 -4026
rect -5258 -4262 -5076 -4026
rect -5676 -4346 -5076 -4262
rect -5676 -4582 -5494 -4346
rect -5258 -4582 -5076 -4346
rect -5676 -4604 -5076 -4582
rect 8004 -4026 8604 9098
rect 8004 -4262 8186 -4026
rect 8422 -4262 8604 -4026
rect 8004 -4346 8604 -4262
rect 8004 -4582 8186 -4346
rect 8422 -4582 8604 -4346
rect -6596 -5182 -6414 -4946
rect -6178 -5182 -5996 -4946
rect -6596 -5266 -5996 -5182
rect -6596 -5502 -6414 -5266
rect -6178 -5502 -5996 -5266
rect -6596 -5524 -5996 -5502
rect 8004 -5524 8604 -4582
rect 11604 697254 12204 709802
rect 29604 711278 30204 711300
rect 29604 711042 29786 711278
rect 30022 711042 30204 711278
rect 29604 710958 30204 711042
rect 29604 710722 29786 710958
rect 30022 710722 30204 710958
rect 26004 709438 26604 709460
rect 26004 709202 26186 709438
rect 26422 709202 26604 709438
rect 26004 709118 26604 709202
rect 26004 708882 26186 709118
rect 26422 708882 26604 709118
rect 22404 707598 23004 707620
rect 22404 707362 22586 707598
rect 22822 707362 23004 707598
rect 22404 707278 23004 707362
rect 22404 707042 22586 707278
rect 22822 707042 23004 707278
rect 11604 697018 11786 697254
rect 12022 697018 12204 697254
rect 11604 696934 12204 697018
rect 11604 696698 11786 696934
rect 12022 696698 12204 696934
rect 11604 661254 12204 696698
rect 11604 661018 11786 661254
rect 12022 661018 12204 661254
rect 11604 660934 12204 661018
rect 11604 660698 11786 660934
rect 12022 660698 12204 660934
rect 11604 625254 12204 660698
rect 11604 625018 11786 625254
rect 12022 625018 12204 625254
rect 11604 624934 12204 625018
rect 11604 624698 11786 624934
rect 12022 624698 12204 624934
rect 11604 589254 12204 624698
rect 11604 589018 11786 589254
rect 12022 589018 12204 589254
rect 11604 588934 12204 589018
rect 11604 588698 11786 588934
rect 12022 588698 12204 588934
rect 11604 553254 12204 588698
rect 11604 553018 11786 553254
rect 12022 553018 12204 553254
rect 11604 552934 12204 553018
rect 11604 552698 11786 552934
rect 12022 552698 12204 552934
rect 11604 517254 12204 552698
rect 11604 517018 11786 517254
rect 12022 517018 12204 517254
rect 11604 516934 12204 517018
rect 11604 516698 11786 516934
rect 12022 516698 12204 516934
rect 11604 481254 12204 516698
rect 11604 481018 11786 481254
rect 12022 481018 12204 481254
rect 11604 480934 12204 481018
rect 11604 480698 11786 480934
rect 12022 480698 12204 480934
rect 11604 445254 12204 480698
rect 11604 445018 11786 445254
rect 12022 445018 12204 445254
rect 11604 444934 12204 445018
rect 11604 444698 11786 444934
rect 12022 444698 12204 444934
rect 11604 409254 12204 444698
rect 11604 409018 11786 409254
rect 12022 409018 12204 409254
rect 11604 408934 12204 409018
rect 11604 408698 11786 408934
rect 12022 408698 12204 408934
rect 11604 373254 12204 408698
rect 11604 373018 11786 373254
rect 12022 373018 12204 373254
rect 11604 372934 12204 373018
rect 11604 372698 11786 372934
rect 12022 372698 12204 372934
rect 11604 337254 12204 372698
rect 11604 337018 11786 337254
rect 12022 337018 12204 337254
rect 11604 336934 12204 337018
rect 11604 336698 11786 336934
rect 12022 336698 12204 336934
rect 11604 301254 12204 336698
rect 11604 301018 11786 301254
rect 12022 301018 12204 301254
rect 11604 300934 12204 301018
rect 11604 300698 11786 300934
rect 12022 300698 12204 300934
rect 11604 265254 12204 300698
rect 11604 265018 11786 265254
rect 12022 265018 12204 265254
rect 11604 264934 12204 265018
rect 11604 264698 11786 264934
rect 12022 264698 12204 264934
rect 11604 229254 12204 264698
rect 11604 229018 11786 229254
rect 12022 229018 12204 229254
rect 11604 228934 12204 229018
rect 11604 228698 11786 228934
rect 12022 228698 12204 228934
rect 11604 193254 12204 228698
rect 11604 193018 11786 193254
rect 12022 193018 12204 193254
rect 11604 192934 12204 193018
rect 11604 192698 11786 192934
rect 12022 192698 12204 192934
rect 11604 157254 12204 192698
rect 11604 157018 11786 157254
rect 12022 157018 12204 157254
rect 11604 156934 12204 157018
rect 11604 156698 11786 156934
rect 12022 156698 12204 156934
rect 11604 121254 12204 156698
rect 11604 121018 11786 121254
rect 12022 121018 12204 121254
rect 11604 120934 12204 121018
rect 11604 120698 11786 120934
rect 12022 120698 12204 120934
rect 11604 85254 12204 120698
rect 11604 85018 11786 85254
rect 12022 85018 12204 85254
rect 11604 84934 12204 85018
rect 11604 84698 11786 84934
rect 12022 84698 12204 84934
rect 11604 49254 12204 84698
rect 11604 49018 11786 49254
rect 12022 49018 12204 49254
rect 11604 48934 12204 49018
rect 11604 48698 11786 48934
rect 12022 48698 12204 48934
rect 11604 13254 12204 48698
rect 11604 13018 11786 13254
rect 12022 13018 12204 13254
rect 11604 12934 12204 13018
rect 11604 12698 11786 12934
rect 12022 12698 12204 12934
rect -7516 -6102 -7334 -5866
rect -7098 -6102 -6916 -5866
rect -7516 -6186 -6916 -6102
rect -7516 -6422 -7334 -6186
rect -7098 -6422 -6916 -6186
rect -7516 -6444 -6916 -6422
rect 11604 -5866 12204 12698
rect 18804 705758 19404 705780
rect 18804 705522 18986 705758
rect 19222 705522 19404 705758
rect 18804 705438 19404 705522
rect 18804 705202 18986 705438
rect 19222 705202 19404 705438
rect 18804 668454 19404 705202
rect 18804 668218 18986 668454
rect 19222 668218 19404 668454
rect 18804 668134 19404 668218
rect 18804 667898 18986 668134
rect 19222 667898 19404 668134
rect 18804 632454 19404 667898
rect 18804 632218 18986 632454
rect 19222 632218 19404 632454
rect 18804 632134 19404 632218
rect 18804 631898 18986 632134
rect 19222 631898 19404 632134
rect 18804 596454 19404 631898
rect 18804 596218 18986 596454
rect 19222 596218 19404 596454
rect 18804 596134 19404 596218
rect 18804 595898 18986 596134
rect 19222 595898 19404 596134
rect 18804 560454 19404 595898
rect 18804 560218 18986 560454
rect 19222 560218 19404 560454
rect 18804 560134 19404 560218
rect 18804 559898 18986 560134
rect 19222 559898 19404 560134
rect 18804 524454 19404 559898
rect 18804 524218 18986 524454
rect 19222 524218 19404 524454
rect 18804 524134 19404 524218
rect 18804 523898 18986 524134
rect 19222 523898 19404 524134
rect 18804 488454 19404 523898
rect 18804 488218 18986 488454
rect 19222 488218 19404 488454
rect 18804 488134 19404 488218
rect 18804 487898 18986 488134
rect 19222 487898 19404 488134
rect 18804 452454 19404 487898
rect 18804 452218 18986 452454
rect 19222 452218 19404 452454
rect 18804 452134 19404 452218
rect 18804 451898 18986 452134
rect 19222 451898 19404 452134
rect 18804 416454 19404 451898
rect 18804 416218 18986 416454
rect 19222 416218 19404 416454
rect 18804 416134 19404 416218
rect 18804 415898 18986 416134
rect 19222 415898 19404 416134
rect 18804 380454 19404 415898
rect 18804 380218 18986 380454
rect 19222 380218 19404 380454
rect 18804 380134 19404 380218
rect 18804 379898 18986 380134
rect 19222 379898 19404 380134
rect 18804 344454 19404 379898
rect 18804 344218 18986 344454
rect 19222 344218 19404 344454
rect 18804 344134 19404 344218
rect 18804 343898 18986 344134
rect 19222 343898 19404 344134
rect 18804 308454 19404 343898
rect 18804 308218 18986 308454
rect 19222 308218 19404 308454
rect 18804 308134 19404 308218
rect 18804 307898 18986 308134
rect 19222 307898 19404 308134
rect 18804 272454 19404 307898
rect 18804 272218 18986 272454
rect 19222 272218 19404 272454
rect 18804 272134 19404 272218
rect 18804 271898 18986 272134
rect 19222 271898 19404 272134
rect 18804 236454 19404 271898
rect 18804 236218 18986 236454
rect 19222 236218 19404 236454
rect 18804 236134 19404 236218
rect 18804 235898 18986 236134
rect 19222 235898 19404 236134
rect 18804 200454 19404 235898
rect 18804 200218 18986 200454
rect 19222 200218 19404 200454
rect 18804 200134 19404 200218
rect 18804 199898 18986 200134
rect 19222 199898 19404 200134
rect 18804 164454 19404 199898
rect 18804 164218 18986 164454
rect 19222 164218 19404 164454
rect 18804 164134 19404 164218
rect 18804 163898 18986 164134
rect 19222 163898 19404 164134
rect 18804 128454 19404 163898
rect 18804 128218 18986 128454
rect 19222 128218 19404 128454
rect 18804 128134 19404 128218
rect 18804 127898 18986 128134
rect 19222 127898 19404 128134
rect 18804 92454 19404 127898
rect 18804 92218 18986 92454
rect 19222 92218 19404 92454
rect 18804 92134 19404 92218
rect 18804 91898 18986 92134
rect 19222 91898 19404 92134
rect 18804 56454 19404 91898
rect 18804 56218 18986 56454
rect 19222 56218 19404 56454
rect 18804 56134 19404 56218
rect 18804 55898 18986 56134
rect 19222 55898 19404 56134
rect 18804 20454 19404 55898
rect 18804 20218 18986 20454
rect 19222 20218 19404 20454
rect 18804 20134 19404 20218
rect 18804 19898 18986 20134
rect 19222 19898 19404 20134
rect 18804 -1266 19404 19898
rect 18804 -1502 18986 -1266
rect 19222 -1502 19404 -1266
rect 18804 -1586 19404 -1502
rect 18804 -1822 18986 -1586
rect 19222 -1822 19404 -1586
rect 18804 -1844 19404 -1822
rect 22404 672054 23004 707042
rect 22404 671818 22586 672054
rect 22822 671818 23004 672054
rect 22404 671734 23004 671818
rect 22404 671498 22586 671734
rect 22822 671498 23004 671734
rect 22404 636054 23004 671498
rect 22404 635818 22586 636054
rect 22822 635818 23004 636054
rect 22404 635734 23004 635818
rect 22404 635498 22586 635734
rect 22822 635498 23004 635734
rect 22404 600054 23004 635498
rect 22404 599818 22586 600054
rect 22822 599818 23004 600054
rect 22404 599734 23004 599818
rect 22404 599498 22586 599734
rect 22822 599498 23004 599734
rect 22404 564054 23004 599498
rect 22404 563818 22586 564054
rect 22822 563818 23004 564054
rect 22404 563734 23004 563818
rect 22404 563498 22586 563734
rect 22822 563498 23004 563734
rect 22404 528054 23004 563498
rect 22404 527818 22586 528054
rect 22822 527818 23004 528054
rect 22404 527734 23004 527818
rect 22404 527498 22586 527734
rect 22822 527498 23004 527734
rect 22404 492054 23004 527498
rect 22404 491818 22586 492054
rect 22822 491818 23004 492054
rect 22404 491734 23004 491818
rect 22404 491498 22586 491734
rect 22822 491498 23004 491734
rect 22404 456054 23004 491498
rect 22404 455818 22586 456054
rect 22822 455818 23004 456054
rect 22404 455734 23004 455818
rect 22404 455498 22586 455734
rect 22822 455498 23004 455734
rect 22404 420054 23004 455498
rect 22404 419818 22586 420054
rect 22822 419818 23004 420054
rect 22404 419734 23004 419818
rect 22404 419498 22586 419734
rect 22822 419498 23004 419734
rect 22404 384054 23004 419498
rect 22404 383818 22586 384054
rect 22822 383818 23004 384054
rect 22404 383734 23004 383818
rect 22404 383498 22586 383734
rect 22822 383498 23004 383734
rect 22404 348054 23004 383498
rect 22404 347818 22586 348054
rect 22822 347818 23004 348054
rect 22404 347734 23004 347818
rect 22404 347498 22586 347734
rect 22822 347498 23004 347734
rect 22404 312054 23004 347498
rect 22404 311818 22586 312054
rect 22822 311818 23004 312054
rect 22404 311734 23004 311818
rect 22404 311498 22586 311734
rect 22822 311498 23004 311734
rect 22404 276054 23004 311498
rect 22404 275818 22586 276054
rect 22822 275818 23004 276054
rect 22404 275734 23004 275818
rect 22404 275498 22586 275734
rect 22822 275498 23004 275734
rect 22404 240054 23004 275498
rect 22404 239818 22586 240054
rect 22822 239818 23004 240054
rect 22404 239734 23004 239818
rect 22404 239498 22586 239734
rect 22822 239498 23004 239734
rect 22404 204054 23004 239498
rect 22404 203818 22586 204054
rect 22822 203818 23004 204054
rect 22404 203734 23004 203818
rect 22404 203498 22586 203734
rect 22822 203498 23004 203734
rect 22404 168054 23004 203498
rect 22404 167818 22586 168054
rect 22822 167818 23004 168054
rect 22404 167734 23004 167818
rect 22404 167498 22586 167734
rect 22822 167498 23004 167734
rect 22404 132054 23004 167498
rect 22404 131818 22586 132054
rect 22822 131818 23004 132054
rect 22404 131734 23004 131818
rect 22404 131498 22586 131734
rect 22822 131498 23004 131734
rect 22404 96054 23004 131498
rect 22404 95818 22586 96054
rect 22822 95818 23004 96054
rect 22404 95734 23004 95818
rect 22404 95498 22586 95734
rect 22822 95498 23004 95734
rect 22404 60054 23004 95498
rect 22404 59818 22586 60054
rect 22822 59818 23004 60054
rect 22404 59734 23004 59818
rect 22404 59498 22586 59734
rect 22822 59498 23004 59734
rect 22404 24054 23004 59498
rect 22404 23818 22586 24054
rect 22822 23818 23004 24054
rect 22404 23734 23004 23818
rect 22404 23498 22586 23734
rect 22822 23498 23004 23734
rect 22404 -3106 23004 23498
rect 22404 -3342 22586 -3106
rect 22822 -3342 23004 -3106
rect 22404 -3426 23004 -3342
rect 22404 -3662 22586 -3426
rect 22822 -3662 23004 -3426
rect 22404 -3684 23004 -3662
rect 26004 675654 26604 708882
rect 26004 675418 26186 675654
rect 26422 675418 26604 675654
rect 26004 675334 26604 675418
rect 26004 675098 26186 675334
rect 26422 675098 26604 675334
rect 26004 639654 26604 675098
rect 26004 639418 26186 639654
rect 26422 639418 26604 639654
rect 26004 639334 26604 639418
rect 26004 639098 26186 639334
rect 26422 639098 26604 639334
rect 26004 603654 26604 639098
rect 26004 603418 26186 603654
rect 26422 603418 26604 603654
rect 26004 603334 26604 603418
rect 26004 603098 26186 603334
rect 26422 603098 26604 603334
rect 26004 567654 26604 603098
rect 26004 567418 26186 567654
rect 26422 567418 26604 567654
rect 26004 567334 26604 567418
rect 26004 567098 26186 567334
rect 26422 567098 26604 567334
rect 26004 531654 26604 567098
rect 26004 531418 26186 531654
rect 26422 531418 26604 531654
rect 26004 531334 26604 531418
rect 26004 531098 26186 531334
rect 26422 531098 26604 531334
rect 26004 495654 26604 531098
rect 26004 495418 26186 495654
rect 26422 495418 26604 495654
rect 26004 495334 26604 495418
rect 26004 495098 26186 495334
rect 26422 495098 26604 495334
rect 26004 459654 26604 495098
rect 26004 459418 26186 459654
rect 26422 459418 26604 459654
rect 26004 459334 26604 459418
rect 26004 459098 26186 459334
rect 26422 459098 26604 459334
rect 26004 423654 26604 459098
rect 26004 423418 26186 423654
rect 26422 423418 26604 423654
rect 26004 423334 26604 423418
rect 26004 423098 26186 423334
rect 26422 423098 26604 423334
rect 26004 387654 26604 423098
rect 26004 387418 26186 387654
rect 26422 387418 26604 387654
rect 26004 387334 26604 387418
rect 26004 387098 26186 387334
rect 26422 387098 26604 387334
rect 26004 351654 26604 387098
rect 26004 351418 26186 351654
rect 26422 351418 26604 351654
rect 26004 351334 26604 351418
rect 26004 351098 26186 351334
rect 26422 351098 26604 351334
rect 26004 315654 26604 351098
rect 26004 315418 26186 315654
rect 26422 315418 26604 315654
rect 26004 315334 26604 315418
rect 26004 315098 26186 315334
rect 26422 315098 26604 315334
rect 26004 279654 26604 315098
rect 26004 279418 26186 279654
rect 26422 279418 26604 279654
rect 26004 279334 26604 279418
rect 26004 279098 26186 279334
rect 26422 279098 26604 279334
rect 26004 243654 26604 279098
rect 26004 243418 26186 243654
rect 26422 243418 26604 243654
rect 26004 243334 26604 243418
rect 26004 243098 26186 243334
rect 26422 243098 26604 243334
rect 26004 207654 26604 243098
rect 26004 207418 26186 207654
rect 26422 207418 26604 207654
rect 26004 207334 26604 207418
rect 26004 207098 26186 207334
rect 26422 207098 26604 207334
rect 26004 171654 26604 207098
rect 26004 171418 26186 171654
rect 26422 171418 26604 171654
rect 26004 171334 26604 171418
rect 26004 171098 26186 171334
rect 26422 171098 26604 171334
rect 26004 135654 26604 171098
rect 26004 135418 26186 135654
rect 26422 135418 26604 135654
rect 26004 135334 26604 135418
rect 26004 135098 26186 135334
rect 26422 135098 26604 135334
rect 26004 99654 26604 135098
rect 26004 99418 26186 99654
rect 26422 99418 26604 99654
rect 26004 99334 26604 99418
rect 26004 99098 26186 99334
rect 26422 99098 26604 99334
rect 26004 63654 26604 99098
rect 26004 63418 26186 63654
rect 26422 63418 26604 63654
rect 26004 63334 26604 63418
rect 26004 63098 26186 63334
rect 26422 63098 26604 63334
rect 26004 27654 26604 63098
rect 26004 27418 26186 27654
rect 26422 27418 26604 27654
rect 26004 27334 26604 27418
rect 26004 27098 26186 27334
rect 26422 27098 26604 27334
rect 26004 -4946 26604 27098
rect 26004 -5182 26186 -4946
rect 26422 -5182 26604 -4946
rect 26004 -5266 26604 -5182
rect 26004 -5502 26186 -5266
rect 26422 -5502 26604 -5266
rect 26004 -5524 26604 -5502
rect 29604 679254 30204 710722
rect 47604 710358 48204 711300
rect 47604 710122 47786 710358
rect 48022 710122 48204 710358
rect 47604 710038 48204 710122
rect 47604 709802 47786 710038
rect 48022 709802 48204 710038
rect 44004 708518 44604 709460
rect 44004 708282 44186 708518
rect 44422 708282 44604 708518
rect 44004 708198 44604 708282
rect 44004 707962 44186 708198
rect 44422 707962 44604 708198
rect 40404 706678 41004 707620
rect 40404 706442 40586 706678
rect 40822 706442 41004 706678
rect 40404 706358 41004 706442
rect 40404 706122 40586 706358
rect 40822 706122 41004 706358
rect 29604 679018 29786 679254
rect 30022 679018 30204 679254
rect 29604 678934 30204 679018
rect 29604 678698 29786 678934
rect 30022 678698 30204 678934
rect 29604 643254 30204 678698
rect 29604 643018 29786 643254
rect 30022 643018 30204 643254
rect 29604 642934 30204 643018
rect 29604 642698 29786 642934
rect 30022 642698 30204 642934
rect 29604 607254 30204 642698
rect 29604 607018 29786 607254
rect 30022 607018 30204 607254
rect 29604 606934 30204 607018
rect 29604 606698 29786 606934
rect 30022 606698 30204 606934
rect 29604 571254 30204 606698
rect 29604 571018 29786 571254
rect 30022 571018 30204 571254
rect 29604 570934 30204 571018
rect 29604 570698 29786 570934
rect 30022 570698 30204 570934
rect 29604 535254 30204 570698
rect 29604 535018 29786 535254
rect 30022 535018 30204 535254
rect 29604 534934 30204 535018
rect 29604 534698 29786 534934
rect 30022 534698 30204 534934
rect 29604 499254 30204 534698
rect 29604 499018 29786 499254
rect 30022 499018 30204 499254
rect 29604 498934 30204 499018
rect 29604 498698 29786 498934
rect 30022 498698 30204 498934
rect 29604 463254 30204 498698
rect 29604 463018 29786 463254
rect 30022 463018 30204 463254
rect 29604 462934 30204 463018
rect 29604 462698 29786 462934
rect 30022 462698 30204 462934
rect 29604 427254 30204 462698
rect 29604 427018 29786 427254
rect 30022 427018 30204 427254
rect 29604 426934 30204 427018
rect 29604 426698 29786 426934
rect 30022 426698 30204 426934
rect 29604 391254 30204 426698
rect 29604 391018 29786 391254
rect 30022 391018 30204 391254
rect 29604 390934 30204 391018
rect 29604 390698 29786 390934
rect 30022 390698 30204 390934
rect 29604 355254 30204 390698
rect 29604 355018 29786 355254
rect 30022 355018 30204 355254
rect 29604 354934 30204 355018
rect 29604 354698 29786 354934
rect 30022 354698 30204 354934
rect 29604 319254 30204 354698
rect 29604 319018 29786 319254
rect 30022 319018 30204 319254
rect 29604 318934 30204 319018
rect 29604 318698 29786 318934
rect 30022 318698 30204 318934
rect 29604 283254 30204 318698
rect 29604 283018 29786 283254
rect 30022 283018 30204 283254
rect 29604 282934 30204 283018
rect 29604 282698 29786 282934
rect 30022 282698 30204 282934
rect 29604 247254 30204 282698
rect 29604 247018 29786 247254
rect 30022 247018 30204 247254
rect 29604 246934 30204 247018
rect 29604 246698 29786 246934
rect 30022 246698 30204 246934
rect 29604 211254 30204 246698
rect 29604 211018 29786 211254
rect 30022 211018 30204 211254
rect 29604 210934 30204 211018
rect 29604 210698 29786 210934
rect 30022 210698 30204 210934
rect 29604 175254 30204 210698
rect 29604 175018 29786 175254
rect 30022 175018 30204 175254
rect 29604 174934 30204 175018
rect 29604 174698 29786 174934
rect 30022 174698 30204 174934
rect 29604 139254 30204 174698
rect 29604 139018 29786 139254
rect 30022 139018 30204 139254
rect 29604 138934 30204 139018
rect 29604 138698 29786 138934
rect 30022 138698 30204 138934
rect 29604 103254 30204 138698
rect 29604 103018 29786 103254
rect 30022 103018 30204 103254
rect 29604 102934 30204 103018
rect 29604 102698 29786 102934
rect 30022 102698 30204 102934
rect 29604 67254 30204 102698
rect 29604 67018 29786 67254
rect 30022 67018 30204 67254
rect 29604 66934 30204 67018
rect 29604 66698 29786 66934
rect 30022 66698 30204 66934
rect 29604 31254 30204 66698
rect 29604 31018 29786 31254
rect 30022 31018 30204 31254
rect 29604 30934 30204 31018
rect 29604 30698 29786 30934
rect 30022 30698 30204 30934
rect 11604 -6102 11786 -5866
rect 12022 -6102 12204 -5866
rect 11604 -6186 12204 -6102
rect 11604 -6422 11786 -6186
rect 12022 -6422 12204 -6186
rect -8436 -7022 -8254 -6786
rect -8018 -7022 -7836 -6786
rect -8436 -7106 -7836 -7022
rect -8436 -7342 -8254 -7106
rect -8018 -7342 -7836 -7106
rect -8436 -7364 -7836 -7342
rect 11604 -7364 12204 -6422
rect 29604 -6786 30204 30698
rect 36804 704838 37404 705780
rect 36804 704602 36986 704838
rect 37222 704602 37404 704838
rect 36804 704518 37404 704602
rect 36804 704282 36986 704518
rect 37222 704282 37404 704518
rect 36804 686454 37404 704282
rect 36804 686218 36986 686454
rect 37222 686218 37404 686454
rect 36804 686134 37404 686218
rect 36804 685898 36986 686134
rect 37222 685898 37404 686134
rect 36804 650454 37404 685898
rect 36804 650218 36986 650454
rect 37222 650218 37404 650454
rect 36804 650134 37404 650218
rect 36804 649898 36986 650134
rect 37222 649898 37404 650134
rect 36804 614454 37404 649898
rect 36804 614218 36986 614454
rect 37222 614218 37404 614454
rect 36804 614134 37404 614218
rect 36804 613898 36986 614134
rect 37222 613898 37404 614134
rect 36804 578454 37404 613898
rect 36804 578218 36986 578454
rect 37222 578218 37404 578454
rect 36804 578134 37404 578218
rect 36804 577898 36986 578134
rect 37222 577898 37404 578134
rect 36804 542454 37404 577898
rect 36804 542218 36986 542454
rect 37222 542218 37404 542454
rect 36804 542134 37404 542218
rect 36804 541898 36986 542134
rect 37222 541898 37404 542134
rect 36804 506454 37404 541898
rect 36804 506218 36986 506454
rect 37222 506218 37404 506454
rect 36804 506134 37404 506218
rect 36804 505898 36986 506134
rect 37222 505898 37404 506134
rect 36804 470454 37404 505898
rect 36804 470218 36986 470454
rect 37222 470218 37404 470454
rect 36804 470134 37404 470218
rect 36804 469898 36986 470134
rect 37222 469898 37404 470134
rect 36804 434454 37404 469898
rect 36804 434218 36986 434454
rect 37222 434218 37404 434454
rect 36804 434134 37404 434218
rect 36804 433898 36986 434134
rect 37222 433898 37404 434134
rect 36804 398454 37404 433898
rect 36804 398218 36986 398454
rect 37222 398218 37404 398454
rect 36804 398134 37404 398218
rect 36804 397898 36986 398134
rect 37222 397898 37404 398134
rect 36804 362454 37404 397898
rect 36804 362218 36986 362454
rect 37222 362218 37404 362454
rect 36804 362134 37404 362218
rect 36804 361898 36986 362134
rect 37222 361898 37404 362134
rect 36804 326454 37404 361898
rect 36804 326218 36986 326454
rect 37222 326218 37404 326454
rect 36804 326134 37404 326218
rect 36804 325898 36986 326134
rect 37222 325898 37404 326134
rect 36804 290454 37404 325898
rect 36804 290218 36986 290454
rect 37222 290218 37404 290454
rect 36804 290134 37404 290218
rect 36804 289898 36986 290134
rect 37222 289898 37404 290134
rect 36804 254454 37404 289898
rect 36804 254218 36986 254454
rect 37222 254218 37404 254454
rect 36804 254134 37404 254218
rect 36804 253898 36986 254134
rect 37222 253898 37404 254134
rect 36804 218454 37404 253898
rect 36804 218218 36986 218454
rect 37222 218218 37404 218454
rect 36804 218134 37404 218218
rect 36804 217898 36986 218134
rect 37222 217898 37404 218134
rect 36804 182454 37404 217898
rect 36804 182218 36986 182454
rect 37222 182218 37404 182454
rect 36804 182134 37404 182218
rect 36804 181898 36986 182134
rect 37222 181898 37404 182134
rect 36804 146454 37404 181898
rect 36804 146218 36986 146454
rect 37222 146218 37404 146454
rect 36804 146134 37404 146218
rect 36804 145898 36986 146134
rect 37222 145898 37404 146134
rect 36804 110454 37404 145898
rect 36804 110218 36986 110454
rect 37222 110218 37404 110454
rect 36804 110134 37404 110218
rect 36804 109898 36986 110134
rect 37222 109898 37404 110134
rect 36804 74454 37404 109898
rect 36804 74218 36986 74454
rect 37222 74218 37404 74454
rect 36804 74134 37404 74218
rect 36804 73898 36986 74134
rect 37222 73898 37404 74134
rect 36804 38454 37404 73898
rect 36804 38218 36986 38454
rect 37222 38218 37404 38454
rect 36804 38134 37404 38218
rect 36804 37898 36986 38134
rect 37222 37898 37404 38134
rect 36804 2454 37404 37898
rect 36804 2218 36986 2454
rect 37222 2218 37404 2454
rect 36804 2134 37404 2218
rect 36804 1898 36986 2134
rect 37222 1898 37404 2134
rect 36804 -346 37404 1898
rect 36804 -582 36986 -346
rect 37222 -582 37404 -346
rect 36804 -666 37404 -582
rect 36804 -902 36986 -666
rect 37222 -902 37404 -666
rect 36804 -1844 37404 -902
rect 40404 690054 41004 706122
rect 40404 689818 40586 690054
rect 40822 689818 41004 690054
rect 40404 689734 41004 689818
rect 40404 689498 40586 689734
rect 40822 689498 41004 689734
rect 40404 654054 41004 689498
rect 40404 653818 40586 654054
rect 40822 653818 41004 654054
rect 40404 653734 41004 653818
rect 40404 653498 40586 653734
rect 40822 653498 41004 653734
rect 40404 618054 41004 653498
rect 40404 617818 40586 618054
rect 40822 617818 41004 618054
rect 40404 617734 41004 617818
rect 40404 617498 40586 617734
rect 40822 617498 41004 617734
rect 40404 582054 41004 617498
rect 40404 581818 40586 582054
rect 40822 581818 41004 582054
rect 40404 581734 41004 581818
rect 40404 581498 40586 581734
rect 40822 581498 41004 581734
rect 40404 546054 41004 581498
rect 40404 545818 40586 546054
rect 40822 545818 41004 546054
rect 40404 545734 41004 545818
rect 40404 545498 40586 545734
rect 40822 545498 41004 545734
rect 40404 510054 41004 545498
rect 40404 509818 40586 510054
rect 40822 509818 41004 510054
rect 40404 509734 41004 509818
rect 40404 509498 40586 509734
rect 40822 509498 41004 509734
rect 40404 474054 41004 509498
rect 40404 473818 40586 474054
rect 40822 473818 41004 474054
rect 40404 473734 41004 473818
rect 40404 473498 40586 473734
rect 40822 473498 41004 473734
rect 40404 438054 41004 473498
rect 40404 437818 40586 438054
rect 40822 437818 41004 438054
rect 40404 437734 41004 437818
rect 40404 437498 40586 437734
rect 40822 437498 41004 437734
rect 40404 402054 41004 437498
rect 40404 401818 40586 402054
rect 40822 401818 41004 402054
rect 40404 401734 41004 401818
rect 40404 401498 40586 401734
rect 40822 401498 41004 401734
rect 40404 366054 41004 401498
rect 40404 365818 40586 366054
rect 40822 365818 41004 366054
rect 40404 365734 41004 365818
rect 40404 365498 40586 365734
rect 40822 365498 41004 365734
rect 40404 330054 41004 365498
rect 40404 329818 40586 330054
rect 40822 329818 41004 330054
rect 40404 329734 41004 329818
rect 40404 329498 40586 329734
rect 40822 329498 41004 329734
rect 40404 294054 41004 329498
rect 40404 293818 40586 294054
rect 40822 293818 41004 294054
rect 40404 293734 41004 293818
rect 40404 293498 40586 293734
rect 40822 293498 41004 293734
rect 40404 258054 41004 293498
rect 40404 257818 40586 258054
rect 40822 257818 41004 258054
rect 40404 257734 41004 257818
rect 40404 257498 40586 257734
rect 40822 257498 41004 257734
rect 40404 222054 41004 257498
rect 40404 221818 40586 222054
rect 40822 221818 41004 222054
rect 40404 221734 41004 221818
rect 40404 221498 40586 221734
rect 40822 221498 41004 221734
rect 40404 186054 41004 221498
rect 40404 185818 40586 186054
rect 40822 185818 41004 186054
rect 40404 185734 41004 185818
rect 40404 185498 40586 185734
rect 40822 185498 41004 185734
rect 40404 150054 41004 185498
rect 40404 149818 40586 150054
rect 40822 149818 41004 150054
rect 40404 149734 41004 149818
rect 40404 149498 40586 149734
rect 40822 149498 41004 149734
rect 40404 114054 41004 149498
rect 40404 113818 40586 114054
rect 40822 113818 41004 114054
rect 40404 113734 41004 113818
rect 40404 113498 40586 113734
rect 40822 113498 41004 113734
rect 40404 78054 41004 113498
rect 40404 77818 40586 78054
rect 40822 77818 41004 78054
rect 40404 77734 41004 77818
rect 40404 77498 40586 77734
rect 40822 77498 41004 77734
rect 40404 42054 41004 77498
rect 40404 41818 40586 42054
rect 40822 41818 41004 42054
rect 40404 41734 41004 41818
rect 40404 41498 40586 41734
rect 40822 41498 41004 41734
rect 40404 6054 41004 41498
rect 40404 5818 40586 6054
rect 40822 5818 41004 6054
rect 40404 5734 41004 5818
rect 40404 5498 40586 5734
rect 40822 5498 41004 5734
rect 40404 -2186 41004 5498
rect 40404 -2422 40586 -2186
rect 40822 -2422 41004 -2186
rect 40404 -2506 41004 -2422
rect 40404 -2742 40586 -2506
rect 40822 -2742 41004 -2506
rect 40404 -3684 41004 -2742
rect 44004 693654 44604 707962
rect 44004 693418 44186 693654
rect 44422 693418 44604 693654
rect 44004 693334 44604 693418
rect 44004 693098 44186 693334
rect 44422 693098 44604 693334
rect 44004 657654 44604 693098
rect 44004 657418 44186 657654
rect 44422 657418 44604 657654
rect 44004 657334 44604 657418
rect 44004 657098 44186 657334
rect 44422 657098 44604 657334
rect 44004 621654 44604 657098
rect 44004 621418 44186 621654
rect 44422 621418 44604 621654
rect 44004 621334 44604 621418
rect 44004 621098 44186 621334
rect 44422 621098 44604 621334
rect 44004 585654 44604 621098
rect 44004 585418 44186 585654
rect 44422 585418 44604 585654
rect 44004 585334 44604 585418
rect 44004 585098 44186 585334
rect 44422 585098 44604 585334
rect 44004 549654 44604 585098
rect 44004 549418 44186 549654
rect 44422 549418 44604 549654
rect 44004 549334 44604 549418
rect 44004 549098 44186 549334
rect 44422 549098 44604 549334
rect 44004 513654 44604 549098
rect 44004 513418 44186 513654
rect 44422 513418 44604 513654
rect 44004 513334 44604 513418
rect 44004 513098 44186 513334
rect 44422 513098 44604 513334
rect 44004 477654 44604 513098
rect 44004 477418 44186 477654
rect 44422 477418 44604 477654
rect 44004 477334 44604 477418
rect 44004 477098 44186 477334
rect 44422 477098 44604 477334
rect 44004 441654 44604 477098
rect 44004 441418 44186 441654
rect 44422 441418 44604 441654
rect 44004 441334 44604 441418
rect 44004 441098 44186 441334
rect 44422 441098 44604 441334
rect 44004 405654 44604 441098
rect 44004 405418 44186 405654
rect 44422 405418 44604 405654
rect 44004 405334 44604 405418
rect 44004 405098 44186 405334
rect 44422 405098 44604 405334
rect 44004 369654 44604 405098
rect 44004 369418 44186 369654
rect 44422 369418 44604 369654
rect 44004 369334 44604 369418
rect 44004 369098 44186 369334
rect 44422 369098 44604 369334
rect 44004 333654 44604 369098
rect 44004 333418 44186 333654
rect 44422 333418 44604 333654
rect 44004 333334 44604 333418
rect 44004 333098 44186 333334
rect 44422 333098 44604 333334
rect 44004 297654 44604 333098
rect 44004 297418 44186 297654
rect 44422 297418 44604 297654
rect 44004 297334 44604 297418
rect 44004 297098 44186 297334
rect 44422 297098 44604 297334
rect 44004 261654 44604 297098
rect 44004 261418 44186 261654
rect 44422 261418 44604 261654
rect 44004 261334 44604 261418
rect 44004 261098 44186 261334
rect 44422 261098 44604 261334
rect 44004 225654 44604 261098
rect 44004 225418 44186 225654
rect 44422 225418 44604 225654
rect 44004 225334 44604 225418
rect 44004 225098 44186 225334
rect 44422 225098 44604 225334
rect 44004 189654 44604 225098
rect 44004 189418 44186 189654
rect 44422 189418 44604 189654
rect 44004 189334 44604 189418
rect 44004 189098 44186 189334
rect 44422 189098 44604 189334
rect 44004 153654 44604 189098
rect 44004 153418 44186 153654
rect 44422 153418 44604 153654
rect 44004 153334 44604 153418
rect 44004 153098 44186 153334
rect 44422 153098 44604 153334
rect 44004 117654 44604 153098
rect 44004 117418 44186 117654
rect 44422 117418 44604 117654
rect 44004 117334 44604 117418
rect 44004 117098 44186 117334
rect 44422 117098 44604 117334
rect 44004 81654 44604 117098
rect 44004 81418 44186 81654
rect 44422 81418 44604 81654
rect 44004 81334 44604 81418
rect 44004 81098 44186 81334
rect 44422 81098 44604 81334
rect 44004 45654 44604 81098
rect 44004 45418 44186 45654
rect 44422 45418 44604 45654
rect 44004 45334 44604 45418
rect 44004 45098 44186 45334
rect 44422 45098 44604 45334
rect 44004 9654 44604 45098
rect 44004 9418 44186 9654
rect 44422 9418 44604 9654
rect 44004 9334 44604 9418
rect 44004 9098 44186 9334
rect 44422 9098 44604 9334
rect 44004 -4026 44604 9098
rect 44004 -4262 44186 -4026
rect 44422 -4262 44604 -4026
rect 44004 -4346 44604 -4262
rect 44004 -4582 44186 -4346
rect 44422 -4582 44604 -4346
rect 44004 -5524 44604 -4582
rect 47604 697254 48204 709802
rect 65604 711278 66204 711300
rect 65604 711042 65786 711278
rect 66022 711042 66204 711278
rect 65604 710958 66204 711042
rect 65604 710722 65786 710958
rect 66022 710722 66204 710958
rect 62004 709438 62604 709460
rect 62004 709202 62186 709438
rect 62422 709202 62604 709438
rect 62004 709118 62604 709202
rect 62004 708882 62186 709118
rect 62422 708882 62604 709118
rect 58404 707598 59004 707620
rect 58404 707362 58586 707598
rect 58822 707362 59004 707598
rect 58404 707278 59004 707362
rect 58404 707042 58586 707278
rect 58822 707042 59004 707278
rect 47604 697018 47786 697254
rect 48022 697018 48204 697254
rect 47604 696934 48204 697018
rect 47604 696698 47786 696934
rect 48022 696698 48204 696934
rect 47604 661254 48204 696698
rect 47604 661018 47786 661254
rect 48022 661018 48204 661254
rect 47604 660934 48204 661018
rect 47604 660698 47786 660934
rect 48022 660698 48204 660934
rect 47604 625254 48204 660698
rect 47604 625018 47786 625254
rect 48022 625018 48204 625254
rect 47604 624934 48204 625018
rect 47604 624698 47786 624934
rect 48022 624698 48204 624934
rect 47604 589254 48204 624698
rect 47604 589018 47786 589254
rect 48022 589018 48204 589254
rect 47604 588934 48204 589018
rect 47604 588698 47786 588934
rect 48022 588698 48204 588934
rect 47604 553254 48204 588698
rect 47604 553018 47786 553254
rect 48022 553018 48204 553254
rect 47604 552934 48204 553018
rect 47604 552698 47786 552934
rect 48022 552698 48204 552934
rect 47604 517254 48204 552698
rect 47604 517018 47786 517254
rect 48022 517018 48204 517254
rect 47604 516934 48204 517018
rect 47604 516698 47786 516934
rect 48022 516698 48204 516934
rect 47604 481254 48204 516698
rect 47604 481018 47786 481254
rect 48022 481018 48204 481254
rect 47604 480934 48204 481018
rect 47604 480698 47786 480934
rect 48022 480698 48204 480934
rect 47604 445254 48204 480698
rect 47604 445018 47786 445254
rect 48022 445018 48204 445254
rect 47604 444934 48204 445018
rect 47604 444698 47786 444934
rect 48022 444698 48204 444934
rect 47604 409254 48204 444698
rect 47604 409018 47786 409254
rect 48022 409018 48204 409254
rect 47604 408934 48204 409018
rect 47604 408698 47786 408934
rect 48022 408698 48204 408934
rect 47604 373254 48204 408698
rect 47604 373018 47786 373254
rect 48022 373018 48204 373254
rect 47604 372934 48204 373018
rect 47604 372698 47786 372934
rect 48022 372698 48204 372934
rect 47604 337254 48204 372698
rect 47604 337018 47786 337254
rect 48022 337018 48204 337254
rect 47604 336934 48204 337018
rect 47604 336698 47786 336934
rect 48022 336698 48204 336934
rect 47604 301254 48204 336698
rect 47604 301018 47786 301254
rect 48022 301018 48204 301254
rect 47604 300934 48204 301018
rect 47604 300698 47786 300934
rect 48022 300698 48204 300934
rect 47604 265254 48204 300698
rect 47604 265018 47786 265254
rect 48022 265018 48204 265254
rect 47604 264934 48204 265018
rect 47604 264698 47786 264934
rect 48022 264698 48204 264934
rect 47604 229254 48204 264698
rect 47604 229018 47786 229254
rect 48022 229018 48204 229254
rect 47604 228934 48204 229018
rect 47604 228698 47786 228934
rect 48022 228698 48204 228934
rect 47604 193254 48204 228698
rect 47604 193018 47786 193254
rect 48022 193018 48204 193254
rect 47604 192934 48204 193018
rect 47604 192698 47786 192934
rect 48022 192698 48204 192934
rect 47604 157254 48204 192698
rect 47604 157018 47786 157254
rect 48022 157018 48204 157254
rect 47604 156934 48204 157018
rect 47604 156698 47786 156934
rect 48022 156698 48204 156934
rect 47604 121254 48204 156698
rect 47604 121018 47786 121254
rect 48022 121018 48204 121254
rect 47604 120934 48204 121018
rect 47604 120698 47786 120934
rect 48022 120698 48204 120934
rect 47604 85254 48204 120698
rect 47604 85018 47786 85254
rect 48022 85018 48204 85254
rect 47604 84934 48204 85018
rect 47604 84698 47786 84934
rect 48022 84698 48204 84934
rect 47604 49254 48204 84698
rect 47604 49018 47786 49254
rect 48022 49018 48204 49254
rect 47604 48934 48204 49018
rect 47604 48698 47786 48934
rect 48022 48698 48204 48934
rect 47604 13254 48204 48698
rect 47604 13018 47786 13254
rect 48022 13018 48204 13254
rect 47604 12934 48204 13018
rect 47604 12698 47786 12934
rect 48022 12698 48204 12934
rect 29604 -7022 29786 -6786
rect 30022 -7022 30204 -6786
rect 29604 -7106 30204 -7022
rect 29604 -7342 29786 -7106
rect 30022 -7342 30204 -7106
rect 29604 -7364 30204 -7342
rect 47604 -5866 48204 12698
rect 54804 705758 55404 705780
rect 54804 705522 54986 705758
rect 55222 705522 55404 705758
rect 54804 705438 55404 705522
rect 54804 705202 54986 705438
rect 55222 705202 55404 705438
rect 54804 668454 55404 705202
rect 54804 668218 54986 668454
rect 55222 668218 55404 668454
rect 54804 668134 55404 668218
rect 54804 667898 54986 668134
rect 55222 667898 55404 668134
rect 54804 632454 55404 667898
rect 54804 632218 54986 632454
rect 55222 632218 55404 632454
rect 54804 632134 55404 632218
rect 54804 631898 54986 632134
rect 55222 631898 55404 632134
rect 54804 596454 55404 631898
rect 54804 596218 54986 596454
rect 55222 596218 55404 596454
rect 54804 596134 55404 596218
rect 54804 595898 54986 596134
rect 55222 595898 55404 596134
rect 54804 560454 55404 595898
rect 54804 560218 54986 560454
rect 55222 560218 55404 560454
rect 54804 560134 55404 560218
rect 54804 559898 54986 560134
rect 55222 559898 55404 560134
rect 54804 524454 55404 559898
rect 54804 524218 54986 524454
rect 55222 524218 55404 524454
rect 54804 524134 55404 524218
rect 54804 523898 54986 524134
rect 55222 523898 55404 524134
rect 54804 488454 55404 523898
rect 54804 488218 54986 488454
rect 55222 488218 55404 488454
rect 54804 488134 55404 488218
rect 54804 487898 54986 488134
rect 55222 487898 55404 488134
rect 54804 452454 55404 487898
rect 54804 452218 54986 452454
rect 55222 452218 55404 452454
rect 54804 452134 55404 452218
rect 54804 451898 54986 452134
rect 55222 451898 55404 452134
rect 54804 416454 55404 451898
rect 54804 416218 54986 416454
rect 55222 416218 55404 416454
rect 54804 416134 55404 416218
rect 54804 415898 54986 416134
rect 55222 415898 55404 416134
rect 54804 380454 55404 415898
rect 54804 380218 54986 380454
rect 55222 380218 55404 380454
rect 54804 380134 55404 380218
rect 54804 379898 54986 380134
rect 55222 379898 55404 380134
rect 54804 344454 55404 379898
rect 54804 344218 54986 344454
rect 55222 344218 55404 344454
rect 54804 344134 55404 344218
rect 54804 343898 54986 344134
rect 55222 343898 55404 344134
rect 54804 308454 55404 343898
rect 54804 308218 54986 308454
rect 55222 308218 55404 308454
rect 54804 308134 55404 308218
rect 54804 307898 54986 308134
rect 55222 307898 55404 308134
rect 54804 272454 55404 307898
rect 54804 272218 54986 272454
rect 55222 272218 55404 272454
rect 54804 272134 55404 272218
rect 54804 271898 54986 272134
rect 55222 271898 55404 272134
rect 54804 236454 55404 271898
rect 54804 236218 54986 236454
rect 55222 236218 55404 236454
rect 54804 236134 55404 236218
rect 54804 235898 54986 236134
rect 55222 235898 55404 236134
rect 54804 200454 55404 235898
rect 54804 200218 54986 200454
rect 55222 200218 55404 200454
rect 54804 200134 55404 200218
rect 54804 199898 54986 200134
rect 55222 199898 55404 200134
rect 54804 164454 55404 199898
rect 54804 164218 54986 164454
rect 55222 164218 55404 164454
rect 54804 164134 55404 164218
rect 54804 163898 54986 164134
rect 55222 163898 55404 164134
rect 54804 128454 55404 163898
rect 54804 128218 54986 128454
rect 55222 128218 55404 128454
rect 54804 128134 55404 128218
rect 54804 127898 54986 128134
rect 55222 127898 55404 128134
rect 54804 92454 55404 127898
rect 54804 92218 54986 92454
rect 55222 92218 55404 92454
rect 54804 92134 55404 92218
rect 54804 91898 54986 92134
rect 55222 91898 55404 92134
rect 54804 56454 55404 91898
rect 54804 56218 54986 56454
rect 55222 56218 55404 56454
rect 54804 56134 55404 56218
rect 54804 55898 54986 56134
rect 55222 55898 55404 56134
rect 54804 20454 55404 55898
rect 54804 20218 54986 20454
rect 55222 20218 55404 20454
rect 54804 20134 55404 20218
rect 54804 19898 54986 20134
rect 55222 19898 55404 20134
rect 54804 -1266 55404 19898
rect 54804 -1502 54986 -1266
rect 55222 -1502 55404 -1266
rect 54804 -1586 55404 -1502
rect 54804 -1822 54986 -1586
rect 55222 -1822 55404 -1586
rect 54804 -1844 55404 -1822
rect 58404 672054 59004 707042
rect 58404 671818 58586 672054
rect 58822 671818 59004 672054
rect 58404 671734 59004 671818
rect 58404 671498 58586 671734
rect 58822 671498 59004 671734
rect 58404 636054 59004 671498
rect 58404 635818 58586 636054
rect 58822 635818 59004 636054
rect 58404 635734 59004 635818
rect 58404 635498 58586 635734
rect 58822 635498 59004 635734
rect 58404 600054 59004 635498
rect 58404 599818 58586 600054
rect 58822 599818 59004 600054
rect 58404 599734 59004 599818
rect 58404 599498 58586 599734
rect 58822 599498 59004 599734
rect 58404 564054 59004 599498
rect 58404 563818 58586 564054
rect 58822 563818 59004 564054
rect 58404 563734 59004 563818
rect 58404 563498 58586 563734
rect 58822 563498 59004 563734
rect 58404 528054 59004 563498
rect 58404 527818 58586 528054
rect 58822 527818 59004 528054
rect 58404 527734 59004 527818
rect 58404 527498 58586 527734
rect 58822 527498 59004 527734
rect 58404 492054 59004 527498
rect 58404 491818 58586 492054
rect 58822 491818 59004 492054
rect 58404 491734 59004 491818
rect 58404 491498 58586 491734
rect 58822 491498 59004 491734
rect 58404 456054 59004 491498
rect 58404 455818 58586 456054
rect 58822 455818 59004 456054
rect 58404 455734 59004 455818
rect 58404 455498 58586 455734
rect 58822 455498 59004 455734
rect 58404 420054 59004 455498
rect 58404 419818 58586 420054
rect 58822 419818 59004 420054
rect 58404 419734 59004 419818
rect 58404 419498 58586 419734
rect 58822 419498 59004 419734
rect 58404 384054 59004 419498
rect 58404 383818 58586 384054
rect 58822 383818 59004 384054
rect 58404 383734 59004 383818
rect 58404 383498 58586 383734
rect 58822 383498 59004 383734
rect 58404 348054 59004 383498
rect 58404 347818 58586 348054
rect 58822 347818 59004 348054
rect 58404 347734 59004 347818
rect 58404 347498 58586 347734
rect 58822 347498 59004 347734
rect 58404 312054 59004 347498
rect 58404 311818 58586 312054
rect 58822 311818 59004 312054
rect 58404 311734 59004 311818
rect 58404 311498 58586 311734
rect 58822 311498 59004 311734
rect 58404 276054 59004 311498
rect 58404 275818 58586 276054
rect 58822 275818 59004 276054
rect 58404 275734 59004 275818
rect 58404 275498 58586 275734
rect 58822 275498 59004 275734
rect 58404 240054 59004 275498
rect 58404 239818 58586 240054
rect 58822 239818 59004 240054
rect 58404 239734 59004 239818
rect 58404 239498 58586 239734
rect 58822 239498 59004 239734
rect 58404 204054 59004 239498
rect 58404 203818 58586 204054
rect 58822 203818 59004 204054
rect 58404 203734 59004 203818
rect 58404 203498 58586 203734
rect 58822 203498 59004 203734
rect 58404 168054 59004 203498
rect 58404 167818 58586 168054
rect 58822 167818 59004 168054
rect 58404 167734 59004 167818
rect 58404 167498 58586 167734
rect 58822 167498 59004 167734
rect 58404 132054 59004 167498
rect 58404 131818 58586 132054
rect 58822 131818 59004 132054
rect 58404 131734 59004 131818
rect 58404 131498 58586 131734
rect 58822 131498 59004 131734
rect 58404 96054 59004 131498
rect 58404 95818 58586 96054
rect 58822 95818 59004 96054
rect 58404 95734 59004 95818
rect 58404 95498 58586 95734
rect 58822 95498 59004 95734
rect 58404 60054 59004 95498
rect 58404 59818 58586 60054
rect 58822 59818 59004 60054
rect 58404 59734 59004 59818
rect 58404 59498 58586 59734
rect 58822 59498 59004 59734
rect 58404 24054 59004 59498
rect 58404 23818 58586 24054
rect 58822 23818 59004 24054
rect 58404 23734 59004 23818
rect 58404 23498 58586 23734
rect 58822 23498 59004 23734
rect 58404 -3106 59004 23498
rect 58404 -3342 58586 -3106
rect 58822 -3342 59004 -3106
rect 58404 -3426 59004 -3342
rect 58404 -3662 58586 -3426
rect 58822 -3662 59004 -3426
rect 58404 -3684 59004 -3662
rect 62004 675654 62604 708882
rect 62004 675418 62186 675654
rect 62422 675418 62604 675654
rect 62004 675334 62604 675418
rect 62004 675098 62186 675334
rect 62422 675098 62604 675334
rect 62004 639654 62604 675098
rect 62004 639418 62186 639654
rect 62422 639418 62604 639654
rect 62004 639334 62604 639418
rect 62004 639098 62186 639334
rect 62422 639098 62604 639334
rect 62004 603654 62604 639098
rect 62004 603418 62186 603654
rect 62422 603418 62604 603654
rect 62004 603334 62604 603418
rect 62004 603098 62186 603334
rect 62422 603098 62604 603334
rect 62004 567654 62604 603098
rect 62004 567418 62186 567654
rect 62422 567418 62604 567654
rect 62004 567334 62604 567418
rect 62004 567098 62186 567334
rect 62422 567098 62604 567334
rect 62004 531654 62604 567098
rect 62004 531418 62186 531654
rect 62422 531418 62604 531654
rect 62004 531334 62604 531418
rect 62004 531098 62186 531334
rect 62422 531098 62604 531334
rect 62004 495654 62604 531098
rect 62004 495418 62186 495654
rect 62422 495418 62604 495654
rect 62004 495334 62604 495418
rect 62004 495098 62186 495334
rect 62422 495098 62604 495334
rect 62004 459654 62604 495098
rect 62004 459418 62186 459654
rect 62422 459418 62604 459654
rect 62004 459334 62604 459418
rect 62004 459098 62186 459334
rect 62422 459098 62604 459334
rect 62004 423654 62604 459098
rect 62004 423418 62186 423654
rect 62422 423418 62604 423654
rect 62004 423334 62604 423418
rect 62004 423098 62186 423334
rect 62422 423098 62604 423334
rect 62004 387654 62604 423098
rect 62004 387418 62186 387654
rect 62422 387418 62604 387654
rect 62004 387334 62604 387418
rect 62004 387098 62186 387334
rect 62422 387098 62604 387334
rect 62004 351654 62604 387098
rect 62004 351418 62186 351654
rect 62422 351418 62604 351654
rect 62004 351334 62604 351418
rect 62004 351098 62186 351334
rect 62422 351098 62604 351334
rect 62004 315654 62604 351098
rect 62004 315418 62186 315654
rect 62422 315418 62604 315654
rect 62004 315334 62604 315418
rect 62004 315098 62186 315334
rect 62422 315098 62604 315334
rect 62004 279654 62604 315098
rect 62004 279418 62186 279654
rect 62422 279418 62604 279654
rect 62004 279334 62604 279418
rect 62004 279098 62186 279334
rect 62422 279098 62604 279334
rect 62004 243654 62604 279098
rect 62004 243418 62186 243654
rect 62422 243418 62604 243654
rect 62004 243334 62604 243418
rect 62004 243098 62186 243334
rect 62422 243098 62604 243334
rect 62004 207654 62604 243098
rect 62004 207418 62186 207654
rect 62422 207418 62604 207654
rect 62004 207334 62604 207418
rect 62004 207098 62186 207334
rect 62422 207098 62604 207334
rect 62004 171654 62604 207098
rect 62004 171418 62186 171654
rect 62422 171418 62604 171654
rect 62004 171334 62604 171418
rect 62004 171098 62186 171334
rect 62422 171098 62604 171334
rect 62004 135654 62604 171098
rect 62004 135418 62186 135654
rect 62422 135418 62604 135654
rect 62004 135334 62604 135418
rect 62004 135098 62186 135334
rect 62422 135098 62604 135334
rect 62004 99654 62604 135098
rect 62004 99418 62186 99654
rect 62422 99418 62604 99654
rect 62004 99334 62604 99418
rect 62004 99098 62186 99334
rect 62422 99098 62604 99334
rect 62004 63654 62604 99098
rect 62004 63418 62186 63654
rect 62422 63418 62604 63654
rect 62004 63334 62604 63418
rect 62004 63098 62186 63334
rect 62422 63098 62604 63334
rect 62004 27654 62604 63098
rect 62004 27418 62186 27654
rect 62422 27418 62604 27654
rect 62004 27334 62604 27418
rect 62004 27098 62186 27334
rect 62422 27098 62604 27334
rect 62004 -4946 62604 27098
rect 62004 -5182 62186 -4946
rect 62422 -5182 62604 -4946
rect 62004 -5266 62604 -5182
rect 62004 -5502 62186 -5266
rect 62422 -5502 62604 -5266
rect 62004 -5524 62604 -5502
rect 65604 679254 66204 710722
rect 83604 710358 84204 711300
rect 83604 710122 83786 710358
rect 84022 710122 84204 710358
rect 83604 710038 84204 710122
rect 83604 709802 83786 710038
rect 84022 709802 84204 710038
rect 80004 708518 80604 709460
rect 80004 708282 80186 708518
rect 80422 708282 80604 708518
rect 80004 708198 80604 708282
rect 80004 707962 80186 708198
rect 80422 707962 80604 708198
rect 76404 706678 77004 707620
rect 76404 706442 76586 706678
rect 76822 706442 77004 706678
rect 76404 706358 77004 706442
rect 76404 706122 76586 706358
rect 76822 706122 77004 706358
rect 65604 679018 65786 679254
rect 66022 679018 66204 679254
rect 65604 678934 66204 679018
rect 65604 678698 65786 678934
rect 66022 678698 66204 678934
rect 65604 643254 66204 678698
rect 65604 643018 65786 643254
rect 66022 643018 66204 643254
rect 65604 642934 66204 643018
rect 65604 642698 65786 642934
rect 66022 642698 66204 642934
rect 65604 607254 66204 642698
rect 65604 607018 65786 607254
rect 66022 607018 66204 607254
rect 65604 606934 66204 607018
rect 65604 606698 65786 606934
rect 66022 606698 66204 606934
rect 65604 571254 66204 606698
rect 65604 571018 65786 571254
rect 66022 571018 66204 571254
rect 65604 570934 66204 571018
rect 65604 570698 65786 570934
rect 66022 570698 66204 570934
rect 65604 535254 66204 570698
rect 65604 535018 65786 535254
rect 66022 535018 66204 535254
rect 65604 534934 66204 535018
rect 65604 534698 65786 534934
rect 66022 534698 66204 534934
rect 65604 499254 66204 534698
rect 65604 499018 65786 499254
rect 66022 499018 66204 499254
rect 65604 498934 66204 499018
rect 65604 498698 65786 498934
rect 66022 498698 66204 498934
rect 65604 463254 66204 498698
rect 65604 463018 65786 463254
rect 66022 463018 66204 463254
rect 65604 462934 66204 463018
rect 65604 462698 65786 462934
rect 66022 462698 66204 462934
rect 65604 427254 66204 462698
rect 65604 427018 65786 427254
rect 66022 427018 66204 427254
rect 65604 426934 66204 427018
rect 65604 426698 65786 426934
rect 66022 426698 66204 426934
rect 65604 391254 66204 426698
rect 65604 391018 65786 391254
rect 66022 391018 66204 391254
rect 65604 390934 66204 391018
rect 65604 390698 65786 390934
rect 66022 390698 66204 390934
rect 65604 355254 66204 390698
rect 65604 355018 65786 355254
rect 66022 355018 66204 355254
rect 65604 354934 66204 355018
rect 65604 354698 65786 354934
rect 66022 354698 66204 354934
rect 65604 319254 66204 354698
rect 65604 319018 65786 319254
rect 66022 319018 66204 319254
rect 65604 318934 66204 319018
rect 65604 318698 65786 318934
rect 66022 318698 66204 318934
rect 65604 283254 66204 318698
rect 65604 283018 65786 283254
rect 66022 283018 66204 283254
rect 65604 282934 66204 283018
rect 65604 282698 65786 282934
rect 66022 282698 66204 282934
rect 65604 247254 66204 282698
rect 65604 247018 65786 247254
rect 66022 247018 66204 247254
rect 65604 246934 66204 247018
rect 65604 246698 65786 246934
rect 66022 246698 66204 246934
rect 65604 211254 66204 246698
rect 65604 211018 65786 211254
rect 66022 211018 66204 211254
rect 65604 210934 66204 211018
rect 65604 210698 65786 210934
rect 66022 210698 66204 210934
rect 65604 175254 66204 210698
rect 65604 175018 65786 175254
rect 66022 175018 66204 175254
rect 65604 174934 66204 175018
rect 65604 174698 65786 174934
rect 66022 174698 66204 174934
rect 65604 139254 66204 174698
rect 65604 139018 65786 139254
rect 66022 139018 66204 139254
rect 65604 138934 66204 139018
rect 65604 138698 65786 138934
rect 66022 138698 66204 138934
rect 65604 103254 66204 138698
rect 65604 103018 65786 103254
rect 66022 103018 66204 103254
rect 65604 102934 66204 103018
rect 65604 102698 65786 102934
rect 66022 102698 66204 102934
rect 65604 67254 66204 102698
rect 65604 67018 65786 67254
rect 66022 67018 66204 67254
rect 65604 66934 66204 67018
rect 65604 66698 65786 66934
rect 66022 66698 66204 66934
rect 65604 31254 66204 66698
rect 65604 31018 65786 31254
rect 66022 31018 66204 31254
rect 65604 30934 66204 31018
rect 65604 30698 65786 30934
rect 66022 30698 66204 30934
rect 47604 -6102 47786 -5866
rect 48022 -6102 48204 -5866
rect 47604 -6186 48204 -6102
rect 47604 -6422 47786 -6186
rect 48022 -6422 48204 -6186
rect 47604 -7364 48204 -6422
rect 65604 -6786 66204 30698
rect 72804 704838 73404 705780
rect 72804 704602 72986 704838
rect 73222 704602 73404 704838
rect 72804 704518 73404 704602
rect 72804 704282 72986 704518
rect 73222 704282 73404 704518
rect 72804 686454 73404 704282
rect 72804 686218 72986 686454
rect 73222 686218 73404 686454
rect 72804 686134 73404 686218
rect 72804 685898 72986 686134
rect 73222 685898 73404 686134
rect 72804 650454 73404 685898
rect 72804 650218 72986 650454
rect 73222 650218 73404 650454
rect 72804 650134 73404 650218
rect 72804 649898 72986 650134
rect 73222 649898 73404 650134
rect 72804 614454 73404 649898
rect 72804 614218 72986 614454
rect 73222 614218 73404 614454
rect 72804 614134 73404 614218
rect 72804 613898 72986 614134
rect 73222 613898 73404 614134
rect 72804 578454 73404 613898
rect 72804 578218 72986 578454
rect 73222 578218 73404 578454
rect 72804 578134 73404 578218
rect 72804 577898 72986 578134
rect 73222 577898 73404 578134
rect 72804 542454 73404 577898
rect 72804 542218 72986 542454
rect 73222 542218 73404 542454
rect 72804 542134 73404 542218
rect 72804 541898 72986 542134
rect 73222 541898 73404 542134
rect 72804 506454 73404 541898
rect 72804 506218 72986 506454
rect 73222 506218 73404 506454
rect 72804 506134 73404 506218
rect 72804 505898 72986 506134
rect 73222 505898 73404 506134
rect 72804 470454 73404 505898
rect 72804 470218 72986 470454
rect 73222 470218 73404 470454
rect 72804 470134 73404 470218
rect 72804 469898 72986 470134
rect 73222 469898 73404 470134
rect 72804 434454 73404 469898
rect 72804 434218 72986 434454
rect 73222 434218 73404 434454
rect 72804 434134 73404 434218
rect 72804 433898 72986 434134
rect 73222 433898 73404 434134
rect 72804 398454 73404 433898
rect 72804 398218 72986 398454
rect 73222 398218 73404 398454
rect 72804 398134 73404 398218
rect 72804 397898 72986 398134
rect 73222 397898 73404 398134
rect 72804 362454 73404 397898
rect 72804 362218 72986 362454
rect 73222 362218 73404 362454
rect 72804 362134 73404 362218
rect 72804 361898 72986 362134
rect 73222 361898 73404 362134
rect 72804 326454 73404 361898
rect 72804 326218 72986 326454
rect 73222 326218 73404 326454
rect 72804 326134 73404 326218
rect 72804 325898 72986 326134
rect 73222 325898 73404 326134
rect 72804 290454 73404 325898
rect 72804 290218 72986 290454
rect 73222 290218 73404 290454
rect 72804 290134 73404 290218
rect 72804 289898 72986 290134
rect 73222 289898 73404 290134
rect 72804 254454 73404 289898
rect 72804 254218 72986 254454
rect 73222 254218 73404 254454
rect 72804 254134 73404 254218
rect 72804 253898 72986 254134
rect 73222 253898 73404 254134
rect 72804 218454 73404 253898
rect 72804 218218 72986 218454
rect 73222 218218 73404 218454
rect 72804 218134 73404 218218
rect 72804 217898 72986 218134
rect 73222 217898 73404 218134
rect 72804 182454 73404 217898
rect 72804 182218 72986 182454
rect 73222 182218 73404 182454
rect 72804 182134 73404 182218
rect 72804 181898 72986 182134
rect 73222 181898 73404 182134
rect 72804 146454 73404 181898
rect 72804 146218 72986 146454
rect 73222 146218 73404 146454
rect 72804 146134 73404 146218
rect 72804 145898 72986 146134
rect 73222 145898 73404 146134
rect 72804 110454 73404 145898
rect 72804 110218 72986 110454
rect 73222 110218 73404 110454
rect 72804 110134 73404 110218
rect 72804 109898 72986 110134
rect 73222 109898 73404 110134
rect 72804 74454 73404 109898
rect 72804 74218 72986 74454
rect 73222 74218 73404 74454
rect 72804 74134 73404 74218
rect 72804 73898 72986 74134
rect 73222 73898 73404 74134
rect 72804 38454 73404 73898
rect 72804 38218 72986 38454
rect 73222 38218 73404 38454
rect 72804 38134 73404 38218
rect 72804 37898 72986 38134
rect 73222 37898 73404 38134
rect 72804 2454 73404 37898
rect 72804 2218 72986 2454
rect 73222 2218 73404 2454
rect 72804 2134 73404 2218
rect 72804 1898 72986 2134
rect 73222 1898 73404 2134
rect 72804 -346 73404 1898
rect 72804 -582 72986 -346
rect 73222 -582 73404 -346
rect 72804 -666 73404 -582
rect 72804 -902 72986 -666
rect 73222 -902 73404 -666
rect 72804 -1844 73404 -902
rect 76404 690054 77004 706122
rect 76404 689818 76586 690054
rect 76822 689818 77004 690054
rect 76404 689734 77004 689818
rect 76404 689498 76586 689734
rect 76822 689498 77004 689734
rect 76404 654054 77004 689498
rect 76404 653818 76586 654054
rect 76822 653818 77004 654054
rect 76404 653734 77004 653818
rect 76404 653498 76586 653734
rect 76822 653498 77004 653734
rect 76404 618054 77004 653498
rect 76404 617818 76586 618054
rect 76822 617818 77004 618054
rect 76404 617734 77004 617818
rect 76404 617498 76586 617734
rect 76822 617498 77004 617734
rect 76404 582054 77004 617498
rect 76404 581818 76586 582054
rect 76822 581818 77004 582054
rect 76404 581734 77004 581818
rect 76404 581498 76586 581734
rect 76822 581498 77004 581734
rect 76404 546054 77004 581498
rect 76404 545818 76586 546054
rect 76822 545818 77004 546054
rect 76404 545734 77004 545818
rect 76404 545498 76586 545734
rect 76822 545498 77004 545734
rect 76404 510054 77004 545498
rect 76404 509818 76586 510054
rect 76822 509818 77004 510054
rect 76404 509734 77004 509818
rect 76404 509498 76586 509734
rect 76822 509498 77004 509734
rect 76404 474054 77004 509498
rect 76404 473818 76586 474054
rect 76822 473818 77004 474054
rect 76404 473734 77004 473818
rect 76404 473498 76586 473734
rect 76822 473498 77004 473734
rect 76404 438054 77004 473498
rect 76404 437818 76586 438054
rect 76822 437818 77004 438054
rect 76404 437734 77004 437818
rect 76404 437498 76586 437734
rect 76822 437498 77004 437734
rect 76404 402054 77004 437498
rect 76404 401818 76586 402054
rect 76822 401818 77004 402054
rect 76404 401734 77004 401818
rect 76404 401498 76586 401734
rect 76822 401498 77004 401734
rect 76404 366054 77004 401498
rect 76404 365818 76586 366054
rect 76822 365818 77004 366054
rect 76404 365734 77004 365818
rect 76404 365498 76586 365734
rect 76822 365498 77004 365734
rect 76404 330054 77004 365498
rect 76404 329818 76586 330054
rect 76822 329818 77004 330054
rect 76404 329734 77004 329818
rect 76404 329498 76586 329734
rect 76822 329498 77004 329734
rect 76404 294054 77004 329498
rect 76404 293818 76586 294054
rect 76822 293818 77004 294054
rect 76404 293734 77004 293818
rect 76404 293498 76586 293734
rect 76822 293498 77004 293734
rect 76404 258054 77004 293498
rect 76404 257818 76586 258054
rect 76822 257818 77004 258054
rect 76404 257734 77004 257818
rect 76404 257498 76586 257734
rect 76822 257498 77004 257734
rect 76404 222054 77004 257498
rect 76404 221818 76586 222054
rect 76822 221818 77004 222054
rect 76404 221734 77004 221818
rect 76404 221498 76586 221734
rect 76822 221498 77004 221734
rect 76404 186054 77004 221498
rect 76404 185818 76586 186054
rect 76822 185818 77004 186054
rect 76404 185734 77004 185818
rect 76404 185498 76586 185734
rect 76822 185498 77004 185734
rect 76404 150054 77004 185498
rect 76404 149818 76586 150054
rect 76822 149818 77004 150054
rect 76404 149734 77004 149818
rect 76404 149498 76586 149734
rect 76822 149498 77004 149734
rect 76404 114054 77004 149498
rect 76404 113818 76586 114054
rect 76822 113818 77004 114054
rect 76404 113734 77004 113818
rect 76404 113498 76586 113734
rect 76822 113498 77004 113734
rect 76404 78054 77004 113498
rect 76404 77818 76586 78054
rect 76822 77818 77004 78054
rect 76404 77734 77004 77818
rect 76404 77498 76586 77734
rect 76822 77498 77004 77734
rect 76404 42054 77004 77498
rect 76404 41818 76586 42054
rect 76822 41818 77004 42054
rect 76404 41734 77004 41818
rect 76404 41498 76586 41734
rect 76822 41498 77004 41734
rect 76404 6054 77004 41498
rect 76404 5818 76586 6054
rect 76822 5818 77004 6054
rect 76404 5734 77004 5818
rect 76404 5498 76586 5734
rect 76822 5498 77004 5734
rect 76404 -2186 77004 5498
rect 76404 -2422 76586 -2186
rect 76822 -2422 77004 -2186
rect 76404 -2506 77004 -2422
rect 76404 -2742 76586 -2506
rect 76822 -2742 77004 -2506
rect 76404 -3684 77004 -2742
rect 80004 693654 80604 707962
rect 80004 693418 80186 693654
rect 80422 693418 80604 693654
rect 80004 693334 80604 693418
rect 80004 693098 80186 693334
rect 80422 693098 80604 693334
rect 80004 657654 80604 693098
rect 80004 657418 80186 657654
rect 80422 657418 80604 657654
rect 80004 657334 80604 657418
rect 80004 657098 80186 657334
rect 80422 657098 80604 657334
rect 80004 621654 80604 657098
rect 80004 621418 80186 621654
rect 80422 621418 80604 621654
rect 80004 621334 80604 621418
rect 80004 621098 80186 621334
rect 80422 621098 80604 621334
rect 80004 585654 80604 621098
rect 80004 585418 80186 585654
rect 80422 585418 80604 585654
rect 80004 585334 80604 585418
rect 80004 585098 80186 585334
rect 80422 585098 80604 585334
rect 80004 549654 80604 585098
rect 80004 549418 80186 549654
rect 80422 549418 80604 549654
rect 80004 549334 80604 549418
rect 80004 549098 80186 549334
rect 80422 549098 80604 549334
rect 80004 513654 80604 549098
rect 80004 513418 80186 513654
rect 80422 513418 80604 513654
rect 80004 513334 80604 513418
rect 80004 513098 80186 513334
rect 80422 513098 80604 513334
rect 80004 477654 80604 513098
rect 80004 477418 80186 477654
rect 80422 477418 80604 477654
rect 80004 477334 80604 477418
rect 80004 477098 80186 477334
rect 80422 477098 80604 477334
rect 80004 441654 80604 477098
rect 80004 441418 80186 441654
rect 80422 441418 80604 441654
rect 80004 441334 80604 441418
rect 80004 441098 80186 441334
rect 80422 441098 80604 441334
rect 80004 405654 80604 441098
rect 80004 405418 80186 405654
rect 80422 405418 80604 405654
rect 80004 405334 80604 405418
rect 80004 405098 80186 405334
rect 80422 405098 80604 405334
rect 80004 369654 80604 405098
rect 80004 369418 80186 369654
rect 80422 369418 80604 369654
rect 80004 369334 80604 369418
rect 80004 369098 80186 369334
rect 80422 369098 80604 369334
rect 80004 333654 80604 369098
rect 80004 333418 80186 333654
rect 80422 333418 80604 333654
rect 80004 333334 80604 333418
rect 80004 333098 80186 333334
rect 80422 333098 80604 333334
rect 80004 297654 80604 333098
rect 80004 297418 80186 297654
rect 80422 297418 80604 297654
rect 80004 297334 80604 297418
rect 80004 297098 80186 297334
rect 80422 297098 80604 297334
rect 80004 261654 80604 297098
rect 80004 261418 80186 261654
rect 80422 261418 80604 261654
rect 80004 261334 80604 261418
rect 80004 261098 80186 261334
rect 80422 261098 80604 261334
rect 80004 225654 80604 261098
rect 80004 225418 80186 225654
rect 80422 225418 80604 225654
rect 80004 225334 80604 225418
rect 80004 225098 80186 225334
rect 80422 225098 80604 225334
rect 80004 189654 80604 225098
rect 80004 189418 80186 189654
rect 80422 189418 80604 189654
rect 80004 189334 80604 189418
rect 80004 189098 80186 189334
rect 80422 189098 80604 189334
rect 80004 153654 80604 189098
rect 80004 153418 80186 153654
rect 80422 153418 80604 153654
rect 80004 153334 80604 153418
rect 80004 153098 80186 153334
rect 80422 153098 80604 153334
rect 80004 117654 80604 153098
rect 80004 117418 80186 117654
rect 80422 117418 80604 117654
rect 80004 117334 80604 117418
rect 80004 117098 80186 117334
rect 80422 117098 80604 117334
rect 80004 81654 80604 117098
rect 80004 81418 80186 81654
rect 80422 81418 80604 81654
rect 80004 81334 80604 81418
rect 80004 81098 80186 81334
rect 80422 81098 80604 81334
rect 80004 45654 80604 81098
rect 80004 45418 80186 45654
rect 80422 45418 80604 45654
rect 80004 45334 80604 45418
rect 80004 45098 80186 45334
rect 80422 45098 80604 45334
rect 80004 9654 80604 45098
rect 80004 9418 80186 9654
rect 80422 9418 80604 9654
rect 80004 9334 80604 9418
rect 80004 9098 80186 9334
rect 80422 9098 80604 9334
rect 80004 -4026 80604 9098
rect 80004 -4262 80186 -4026
rect 80422 -4262 80604 -4026
rect 80004 -4346 80604 -4262
rect 80004 -4582 80186 -4346
rect 80422 -4582 80604 -4346
rect 80004 -5524 80604 -4582
rect 83604 697254 84204 709802
rect 101604 711278 102204 711300
rect 101604 711042 101786 711278
rect 102022 711042 102204 711278
rect 101604 710958 102204 711042
rect 101604 710722 101786 710958
rect 102022 710722 102204 710958
rect 98004 709438 98604 709460
rect 98004 709202 98186 709438
rect 98422 709202 98604 709438
rect 98004 709118 98604 709202
rect 98004 708882 98186 709118
rect 98422 708882 98604 709118
rect 94404 707598 95004 707620
rect 94404 707362 94586 707598
rect 94822 707362 95004 707598
rect 94404 707278 95004 707362
rect 94404 707042 94586 707278
rect 94822 707042 95004 707278
rect 83604 697018 83786 697254
rect 84022 697018 84204 697254
rect 83604 696934 84204 697018
rect 83604 696698 83786 696934
rect 84022 696698 84204 696934
rect 83604 661254 84204 696698
rect 83604 661018 83786 661254
rect 84022 661018 84204 661254
rect 83604 660934 84204 661018
rect 83604 660698 83786 660934
rect 84022 660698 84204 660934
rect 83604 625254 84204 660698
rect 83604 625018 83786 625254
rect 84022 625018 84204 625254
rect 83604 624934 84204 625018
rect 83604 624698 83786 624934
rect 84022 624698 84204 624934
rect 83604 589254 84204 624698
rect 83604 589018 83786 589254
rect 84022 589018 84204 589254
rect 83604 588934 84204 589018
rect 83604 588698 83786 588934
rect 84022 588698 84204 588934
rect 83604 553254 84204 588698
rect 83604 553018 83786 553254
rect 84022 553018 84204 553254
rect 83604 552934 84204 553018
rect 83604 552698 83786 552934
rect 84022 552698 84204 552934
rect 83604 517254 84204 552698
rect 83604 517018 83786 517254
rect 84022 517018 84204 517254
rect 83604 516934 84204 517018
rect 83604 516698 83786 516934
rect 84022 516698 84204 516934
rect 83604 481254 84204 516698
rect 83604 481018 83786 481254
rect 84022 481018 84204 481254
rect 83604 480934 84204 481018
rect 83604 480698 83786 480934
rect 84022 480698 84204 480934
rect 83604 445254 84204 480698
rect 83604 445018 83786 445254
rect 84022 445018 84204 445254
rect 83604 444934 84204 445018
rect 83604 444698 83786 444934
rect 84022 444698 84204 444934
rect 83604 409254 84204 444698
rect 83604 409018 83786 409254
rect 84022 409018 84204 409254
rect 83604 408934 84204 409018
rect 83604 408698 83786 408934
rect 84022 408698 84204 408934
rect 83604 373254 84204 408698
rect 83604 373018 83786 373254
rect 84022 373018 84204 373254
rect 83604 372934 84204 373018
rect 83604 372698 83786 372934
rect 84022 372698 84204 372934
rect 83604 337254 84204 372698
rect 83604 337018 83786 337254
rect 84022 337018 84204 337254
rect 83604 336934 84204 337018
rect 83604 336698 83786 336934
rect 84022 336698 84204 336934
rect 83604 301254 84204 336698
rect 83604 301018 83786 301254
rect 84022 301018 84204 301254
rect 83604 300934 84204 301018
rect 83604 300698 83786 300934
rect 84022 300698 84204 300934
rect 83604 265254 84204 300698
rect 83604 265018 83786 265254
rect 84022 265018 84204 265254
rect 83604 264934 84204 265018
rect 83604 264698 83786 264934
rect 84022 264698 84204 264934
rect 83604 229254 84204 264698
rect 83604 229018 83786 229254
rect 84022 229018 84204 229254
rect 83604 228934 84204 229018
rect 83604 228698 83786 228934
rect 84022 228698 84204 228934
rect 83604 193254 84204 228698
rect 83604 193018 83786 193254
rect 84022 193018 84204 193254
rect 83604 192934 84204 193018
rect 83604 192698 83786 192934
rect 84022 192698 84204 192934
rect 83604 157254 84204 192698
rect 83604 157018 83786 157254
rect 84022 157018 84204 157254
rect 83604 156934 84204 157018
rect 83604 156698 83786 156934
rect 84022 156698 84204 156934
rect 83604 121254 84204 156698
rect 83604 121018 83786 121254
rect 84022 121018 84204 121254
rect 83604 120934 84204 121018
rect 83604 120698 83786 120934
rect 84022 120698 84204 120934
rect 83604 85254 84204 120698
rect 83604 85018 83786 85254
rect 84022 85018 84204 85254
rect 83604 84934 84204 85018
rect 83604 84698 83786 84934
rect 84022 84698 84204 84934
rect 83604 49254 84204 84698
rect 83604 49018 83786 49254
rect 84022 49018 84204 49254
rect 83604 48934 84204 49018
rect 83604 48698 83786 48934
rect 84022 48698 84204 48934
rect 83604 13254 84204 48698
rect 83604 13018 83786 13254
rect 84022 13018 84204 13254
rect 83604 12934 84204 13018
rect 83604 12698 83786 12934
rect 84022 12698 84204 12934
rect 65604 -7022 65786 -6786
rect 66022 -7022 66204 -6786
rect 65604 -7106 66204 -7022
rect 65604 -7342 65786 -7106
rect 66022 -7342 66204 -7106
rect 65604 -7364 66204 -7342
rect 83604 -5866 84204 12698
rect 90804 705758 91404 705780
rect 90804 705522 90986 705758
rect 91222 705522 91404 705758
rect 90804 705438 91404 705522
rect 90804 705202 90986 705438
rect 91222 705202 91404 705438
rect 90804 668454 91404 705202
rect 90804 668218 90986 668454
rect 91222 668218 91404 668454
rect 90804 668134 91404 668218
rect 90804 667898 90986 668134
rect 91222 667898 91404 668134
rect 90804 632454 91404 667898
rect 90804 632218 90986 632454
rect 91222 632218 91404 632454
rect 90804 632134 91404 632218
rect 90804 631898 90986 632134
rect 91222 631898 91404 632134
rect 90804 596454 91404 631898
rect 90804 596218 90986 596454
rect 91222 596218 91404 596454
rect 90804 596134 91404 596218
rect 90804 595898 90986 596134
rect 91222 595898 91404 596134
rect 90804 560454 91404 595898
rect 90804 560218 90986 560454
rect 91222 560218 91404 560454
rect 90804 560134 91404 560218
rect 90804 559898 90986 560134
rect 91222 559898 91404 560134
rect 90804 524454 91404 559898
rect 90804 524218 90986 524454
rect 91222 524218 91404 524454
rect 90804 524134 91404 524218
rect 90804 523898 90986 524134
rect 91222 523898 91404 524134
rect 90804 488454 91404 523898
rect 90804 488218 90986 488454
rect 91222 488218 91404 488454
rect 90804 488134 91404 488218
rect 90804 487898 90986 488134
rect 91222 487898 91404 488134
rect 90804 452454 91404 487898
rect 90804 452218 90986 452454
rect 91222 452218 91404 452454
rect 90804 452134 91404 452218
rect 90804 451898 90986 452134
rect 91222 451898 91404 452134
rect 90804 416454 91404 451898
rect 90804 416218 90986 416454
rect 91222 416218 91404 416454
rect 90804 416134 91404 416218
rect 90804 415898 90986 416134
rect 91222 415898 91404 416134
rect 90804 380454 91404 415898
rect 90804 380218 90986 380454
rect 91222 380218 91404 380454
rect 90804 380134 91404 380218
rect 90804 379898 90986 380134
rect 91222 379898 91404 380134
rect 90804 344454 91404 379898
rect 90804 344218 90986 344454
rect 91222 344218 91404 344454
rect 90804 344134 91404 344218
rect 90804 343898 90986 344134
rect 91222 343898 91404 344134
rect 90804 308454 91404 343898
rect 90804 308218 90986 308454
rect 91222 308218 91404 308454
rect 90804 308134 91404 308218
rect 90804 307898 90986 308134
rect 91222 307898 91404 308134
rect 90804 272454 91404 307898
rect 90804 272218 90986 272454
rect 91222 272218 91404 272454
rect 90804 272134 91404 272218
rect 90804 271898 90986 272134
rect 91222 271898 91404 272134
rect 90804 236454 91404 271898
rect 90804 236218 90986 236454
rect 91222 236218 91404 236454
rect 90804 236134 91404 236218
rect 90804 235898 90986 236134
rect 91222 235898 91404 236134
rect 90804 200454 91404 235898
rect 90804 200218 90986 200454
rect 91222 200218 91404 200454
rect 90804 200134 91404 200218
rect 90804 199898 90986 200134
rect 91222 199898 91404 200134
rect 90804 164454 91404 199898
rect 90804 164218 90986 164454
rect 91222 164218 91404 164454
rect 90804 164134 91404 164218
rect 90804 163898 90986 164134
rect 91222 163898 91404 164134
rect 90804 128454 91404 163898
rect 90804 128218 90986 128454
rect 91222 128218 91404 128454
rect 90804 128134 91404 128218
rect 90804 127898 90986 128134
rect 91222 127898 91404 128134
rect 90804 92454 91404 127898
rect 90804 92218 90986 92454
rect 91222 92218 91404 92454
rect 90804 92134 91404 92218
rect 90804 91898 90986 92134
rect 91222 91898 91404 92134
rect 90804 56454 91404 91898
rect 90804 56218 90986 56454
rect 91222 56218 91404 56454
rect 90804 56134 91404 56218
rect 90804 55898 90986 56134
rect 91222 55898 91404 56134
rect 90804 20454 91404 55898
rect 90804 20218 90986 20454
rect 91222 20218 91404 20454
rect 90804 20134 91404 20218
rect 90804 19898 90986 20134
rect 91222 19898 91404 20134
rect 90804 -1266 91404 19898
rect 90804 -1502 90986 -1266
rect 91222 -1502 91404 -1266
rect 90804 -1586 91404 -1502
rect 90804 -1822 90986 -1586
rect 91222 -1822 91404 -1586
rect 90804 -1844 91404 -1822
rect 94404 672054 95004 707042
rect 94404 671818 94586 672054
rect 94822 671818 95004 672054
rect 94404 671734 95004 671818
rect 94404 671498 94586 671734
rect 94822 671498 95004 671734
rect 94404 636054 95004 671498
rect 94404 635818 94586 636054
rect 94822 635818 95004 636054
rect 94404 635734 95004 635818
rect 94404 635498 94586 635734
rect 94822 635498 95004 635734
rect 94404 600054 95004 635498
rect 94404 599818 94586 600054
rect 94822 599818 95004 600054
rect 94404 599734 95004 599818
rect 94404 599498 94586 599734
rect 94822 599498 95004 599734
rect 94404 564054 95004 599498
rect 94404 563818 94586 564054
rect 94822 563818 95004 564054
rect 94404 563734 95004 563818
rect 94404 563498 94586 563734
rect 94822 563498 95004 563734
rect 94404 528054 95004 563498
rect 94404 527818 94586 528054
rect 94822 527818 95004 528054
rect 94404 527734 95004 527818
rect 94404 527498 94586 527734
rect 94822 527498 95004 527734
rect 94404 492054 95004 527498
rect 94404 491818 94586 492054
rect 94822 491818 95004 492054
rect 94404 491734 95004 491818
rect 94404 491498 94586 491734
rect 94822 491498 95004 491734
rect 94404 456054 95004 491498
rect 94404 455818 94586 456054
rect 94822 455818 95004 456054
rect 94404 455734 95004 455818
rect 94404 455498 94586 455734
rect 94822 455498 95004 455734
rect 94404 420054 95004 455498
rect 94404 419818 94586 420054
rect 94822 419818 95004 420054
rect 94404 419734 95004 419818
rect 94404 419498 94586 419734
rect 94822 419498 95004 419734
rect 94404 384054 95004 419498
rect 94404 383818 94586 384054
rect 94822 383818 95004 384054
rect 94404 383734 95004 383818
rect 94404 383498 94586 383734
rect 94822 383498 95004 383734
rect 94404 348054 95004 383498
rect 94404 347818 94586 348054
rect 94822 347818 95004 348054
rect 94404 347734 95004 347818
rect 94404 347498 94586 347734
rect 94822 347498 95004 347734
rect 94404 312054 95004 347498
rect 94404 311818 94586 312054
rect 94822 311818 95004 312054
rect 94404 311734 95004 311818
rect 94404 311498 94586 311734
rect 94822 311498 95004 311734
rect 94404 276054 95004 311498
rect 94404 275818 94586 276054
rect 94822 275818 95004 276054
rect 94404 275734 95004 275818
rect 94404 275498 94586 275734
rect 94822 275498 95004 275734
rect 94404 240054 95004 275498
rect 94404 239818 94586 240054
rect 94822 239818 95004 240054
rect 94404 239734 95004 239818
rect 94404 239498 94586 239734
rect 94822 239498 95004 239734
rect 94404 204054 95004 239498
rect 94404 203818 94586 204054
rect 94822 203818 95004 204054
rect 94404 203734 95004 203818
rect 94404 203498 94586 203734
rect 94822 203498 95004 203734
rect 94404 168054 95004 203498
rect 94404 167818 94586 168054
rect 94822 167818 95004 168054
rect 94404 167734 95004 167818
rect 94404 167498 94586 167734
rect 94822 167498 95004 167734
rect 94404 132054 95004 167498
rect 94404 131818 94586 132054
rect 94822 131818 95004 132054
rect 94404 131734 95004 131818
rect 94404 131498 94586 131734
rect 94822 131498 95004 131734
rect 94404 96054 95004 131498
rect 94404 95818 94586 96054
rect 94822 95818 95004 96054
rect 94404 95734 95004 95818
rect 94404 95498 94586 95734
rect 94822 95498 95004 95734
rect 94404 60054 95004 95498
rect 94404 59818 94586 60054
rect 94822 59818 95004 60054
rect 94404 59734 95004 59818
rect 94404 59498 94586 59734
rect 94822 59498 95004 59734
rect 94404 24054 95004 59498
rect 94404 23818 94586 24054
rect 94822 23818 95004 24054
rect 94404 23734 95004 23818
rect 94404 23498 94586 23734
rect 94822 23498 95004 23734
rect 94404 -3106 95004 23498
rect 94404 -3342 94586 -3106
rect 94822 -3342 95004 -3106
rect 94404 -3426 95004 -3342
rect 94404 -3662 94586 -3426
rect 94822 -3662 95004 -3426
rect 94404 -3684 95004 -3662
rect 98004 675654 98604 708882
rect 98004 675418 98186 675654
rect 98422 675418 98604 675654
rect 98004 675334 98604 675418
rect 98004 675098 98186 675334
rect 98422 675098 98604 675334
rect 98004 639654 98604 675098
rect 98004 639418 98186 639654
rect 98422 639418 98604 639654
rect 98004 639334 98604 639418
rect 98004 639098 98186 639334
rect 98422 639098 98604 639334
rect 98004 603654 98604 639098
rect 98004 603418 98186 603654
rect 98422 603418 98604 603654
rect 98004 603334 98604 603418
rect 98004 603098 98186 603334
rect 98422 603098 98604 603334
rect 98004 567654 98604 603098
rect 98004 567418 98186 567654
rect 98422 567418 98604 567654
rect 98004 567334 98604 567418
rect 98004 567098 98186 567334
rect 98422 567098 98604 567334
rect 98004 531654 98604 567098
rect 98004 531418 98186 531654
rect 98422 531418 98604 531654
rect 98004 531334 98604 531418
rect 98004 531098 98186 531334
rect 98422 531098 98604 531334
rect 98004 495654 98604 531098
rect 98004 495418 98186 495654
rect 98422 495418 98604 495654
rect 98004 495334 98604 495418
rect 98004 495098 98186 495334
rect 98422 495098 98604 495334
rect 98004 459654 98604 495098
rect 98004 459418 98186 459654
rect 98422 459418 98604 459654
rect 98004 459334 98604 459418
rect 98004 459098 98186 459334
rect 98422 459098 98604 459334
rect 98004 423654 98604 459098
rect 98004 423418 98186 423654
rect 98422 423418 98604 423654
rect 98004 423334 98604 423418
rect 98004 423098 98186 423334
rect 98422 423098 98604 423334
rect 98004 387654 98604 423098
rect 98004 387418 98186 387654
rect 98422 387418 98604 387654
rect 98004 387334 98604 387418
rect 98004 387098 98186 387334
rect 98422 387098 98604 387334
rect 98004 351654 98604 387098
rect 98004 351418 98186 351654
rect 98422 351418 98604 351654
rect 98004 351334 98604 351418
rect 98004 351098 98186 351334
rect 98422 351098 98604 351334
rect 98004 315654 98604 351098
rect 98004 315418 98186 315654
rect 98422 315418 98604 315654
rect 98004 315334 98604 315418
rect 98004 315098 98186 315334
rect 98422 315098 98604 315334
rect 98004 279654 98604 315098
rect 98004 279418 98186 279654
rect 98422 279418 98604 279654
rect 98004 279334 98604 279418
rect 98004 279098 98186 279334
rect 98422 279098 98604 279334
rect 98004 243654 98604 279098
rect 98004 243418 98186 243654
rect 98422 243418 98604 243654
rect 98004 243334 98604 243418
rect 98004 243098 98186 243334
rect 98422 243098 98604 243334
rect 98004 207654 98604 243098
rect 98004 207418 98186 207654
rect 98422 207418 98604 207654
rect 98004 207334 98604 207418
rect 98004 207098 98186 207334
rect 98422 207098 98604 207334
rect 98004 171654 98604 207098
rect 98004 171418 98186 171654
rect 98422 171418 98604 171654
rect 98004 171334 98604 171418
rect 98004 171098 98186 171334
rect 98422 171098 98604 171334
rect 98004 135654 98604 171098
rect 98004 135418 98186 135654
rect 98422 135418 98604 135654
rect 98004 135334 98604 135418
rect 98004 135098 98186 135334
rect 98422 135098 98604 135334
rect 98004 99654 98604 135098
rect 98004 99418 98186 99654
rect 98422 99418 98604 99654
rect 98004 99334 98604 99418
rect 98004 99098 98186 99334
rect 98422 99098 98604 99334
rect 98004 63654 98604 99098
rect 98004 63418 98186 63654
rect 98422 63418 98604 63654
rect 98004 63334 98604 63418
rect 98004 63098 98186 63334
rect 98422 63098 98604 63334
rect 98004 27654 98604 63098
rect 98004 27418 98186 27654
rect 98422 27418 98604 27654
rect 98004 27334 98604 27418
rect 98004 27098 98186 27334
rect 98422 27098 98604 27334
rect 98004 -4946 98604 27098
rect 98004 -5182 98186 -4946
rect 98422 -5182 98604 -4946
rect 98004 -5266 98604 -5182
rect 98004 -5502 98186 -5266
rect 98422 -5502 98604 -5266
rect 98004 -5524 98604 -5502
rect 101604 679254 102204 710722
rect 119604 710358 120204 711300
rect 119604 710122 119786 710358
rect 120022 710122 120204 710358
rect 119604 710038 120204 710122
rect 119604 709802 119786 710038
rect 120022 709802 120204 710038
rect 116004 708518 116604 709460
rect 116004 708282 116186 708518
rect 116422 708282 116604 708518
rect 116004 708198 116604 708282
rect 116004 707962 116186 708198
rect 116422 707962 116604 708198
rect 112404 706678 113004 707620
rect 112404 706442 112586 706678
rect 112822 706442 113004 706678
rect 112404 706358 113004 706442
rect 112404 706122 112586 706358
rect 112822 706122 113004 706358
rect 101604 679018 101786 679254
rect 102022 679018 102204 679254
rect 101604 678934 102204 679018
rect 101604 678698 101786 678934
rect 102022 678698 102204 678934
rect 101604 643254 102204 678698
rect 101604 643018 101786 643254
rect 102022 643018 102204 643254
rect 101604 642934 102204 643018
rect 101604 642698 101786 642934
rect 102022 642698 102204 642934
rect 101604 607254 102204 642698
rect 101604 607018 101786 607254
rect 102022 607018 102204 607254
rect 101604 606934 102204 607018
rect 101604 606698 101786 606934
rect 102022 606698 102204 606934
rect 101604 571254 102204 606698
rect 101604 571018 101786 571254
rect 102022 571018 102204 571254
rect 101604 570934 102204 571018
rect 101604 570698 101786 570934
rect 102022 570698 102204 570934
rect 101604 535254 102204 570698
rect 101604 535018 101786 535254
rect 102022 535018 102204 535254
rect 101604 534934 102204 535018
rect 101604 534698 101786 534934
rect 102022 534698 102204 534934
rect 101604 499254 102204 534698
rect 101604 499018 101786 499254
rect 102022 499018 102204 499254
rect 101604 498934 102204 499018
rect 101604 498698 101786 498934
rect 102022 498698 102204 498934
rect 101604 463254 102204 498698
rect 101604 463018 101786 463254
rect 102022 463018 102204 463254
rect 101604 462934 102204 463018
rect 101604 462698 101786 462934
rect 102022 462698 102204 462934
rect 101604 427254 102204 462698
rect 101604 427018 101786 427254
rect 102022 427018 102204 427254
rect 101604 426934 102204 427018
rect 101604 426698 101786 426934
rect 102022 426698 102204 426934
rect 101604 391254 102204 426698
rect 101604 391018 101786 391254
rect 102022 391018 102204 391254
rect 101604 390934 102204 391018
rect 101604 390698 101786 390934
rect 102022 390698 102204 390934
rect 101604 355254 102204 390698
rect 101604 355018 101786 355254
rect 102022 355018 102204 355254
rect 101604 354934 102204 355018
rect 101604 354698 101786 354934
rect 102022 354698 102204 354934
rect 101604 319254 102204 354698
rect 101604 319018 101786 319254
rect 102022 319018 102204 319254
rect 101604 318934 102204 319018
rect 101604 318698 101786 318934
rect 102022 318698 102204 318934
rect 101604 283254 102204 318698
rect 101604 283018 101786 283254
rect 102022 283018 102204 283254
rect 101604 282934 102204 283018
rect 101604 282698 101786 282934
rect 102022 282698 102204 282934
rect 101604 247254 102204 282698
rect 101604 247018 101786 247254
rect 102022 247018 102204 247254
rect 101604 246934 102204 247018
rect 101604 246698 101786 246934
rect 102022 246698 102204 246934
rect 101604 211254 102204 246698
rect 101604 211018 101786 211254
rect 102022 211018 102204 211254
rect 101604 210934 102204 211018
rect 101604 210698 101786 210934
rect 102022 210698 102204 210934
rect 101604 175254 102204 210698
rect 101604 175018 101786 175254
rect 102022 175018 102204 175254
rect 101604 174934 102204 175018
rect 101604 174698 101786 174934
rect 102022 174698 102204 174934
rect 101604 139254 102204 174698
rect 101604 139018 101786 139254
rect 102022 139018 102204 139254
rect 101604 138934 102204 139018
rect 101604 138698 101786 138934
rect 102022 138698 102204 138934
rect 101604 103254 102204 138698
rect 101604 103018 101786 103254
rect 102022 103018 102204 103254
rect 101604 102934 102204 103018
rect 101604 102698 101786 102934
rect 102022 102698 102204 102934
rect 101604 67254 102204 102698
rect 101604 67018 101786 67254
rect 102022 67018 102204 67254
rect 101604 66934 102204 67018
rect 101604 66698 101786 66934
rect 102022 66698 102204 66934
rect 101604 31254 102204 66698
rect 101604 31018 101786 31254
rect 102022 31018 102204 31254
rect 101604 30934 102204 31018
rect 101604 30698 101786 30934
rect 102022 30698 102204 30934
rect 83604 -6102 83786 -5866
rect 84022 -6102 84204 -5866
rect 83604 -6186 84204 -6102
rect 83604 -6422 83786 -6186
rect 84022 -6422 84204 -6186
rect 83604 -7364 84204 -6422
rect 101604 -6786 102204 30698
rect 108804 704838 109404 705780
rect 108804 704602 108986 704838
rect 109222 704602 109404 704838
rect 108804 704518 109404 704602
rect 108804 704282 108986 704518
rect 109222 704282 109404 704518
rect 108804 686454 109404 704282
rect 108804 686218 108986 686454
rect 109222 686218 109404 686454
rect 108804 686134 109404 686218
rect 108804 685898 108986 686134
rect 109222 685898 109404 686134
rect 108804 650454 109404 685898
rect 108804 650218 108986 650454
rect 109222 650218 109404 650454
rect 108804 650134 109404 650218
rect 108804 649898 108986 650134
rect 109222 649898 109404 650134
rect 108804 614454 109404 649898
rect 108804 614218 108986 614454
rect 109222 614218 109404 614454
rect 108804 614134 109404 614218
rect 108804 613898 108986 614134
rect 109222 613898 109404 614134
rect 108804 578454 109404 613898
rect 108804 578218 108986 578454
rect 109222 578218 109404 578454
rect 108804 578134 109404 578218
rect 108804 577898 108986 578134
rect 109222 577898 109404 578134
rect 108804 542454 109404 577898
rect 108804 542218 108986 542454
rect 109222 542218 109404 542454
rect 108804 542134 109404 542218
rect 108804 541898 108986 542134
rect 109222 541898 109404 542134
rect 108804 506454 109404 541898
rect 108804 506218 108986 506454
rect 109222 506218 109404 506454
rect 108804 506134 109404 506218
rect 108804 505898 108986 506134
rect 109222 505898 109404 506134
rect 108804 470454 109404 505898
rect 108804 470218 108986 470454
rect 109222 470218 109404 470454
rect 108804 470134 109404 470218
rect 108804 469898 108986 470134
rect 109222 469898 109404 470134
rect 108804 434454 109404 469898
rect 108804 434218 108986 434454
rect 109222 434218 109404 434454
rect 108804 434134 109404 434218
rect 108804 433898 108986 434134
rect 109222 433898 109404 434134
rect 108804 398454 109404 433898
rect 108804 398218 108986 398454
rect 109222 398218 109404 398454
rect 108804 398134 109404 398218
rect 108804 397898 108986 398134
rect 109222 397898 109404 398134
rect 108804 362454 109404 397898
rect 108804 362218 108986 362454
rect 109222 362218 109404 362454
rect 108804 362134 109404 362218
rect 108804 361898 108986 362134
rect 109222 361898 109404 362134
rect 108804 326454 109404 361898
rect 108804 326218 108986 326454
rect 109222 326218 109404 326454
rect 108804 326134 109404 326218
rect 108804 325898 108986 326134
rect 109222 325898 109404 326134
rect 108804 290454 109404 325898
rect 108804 290218 108986 290454
rect 109222 290218 109404 290454
rect 108804 290134 109404 290218
rect 108804 289898 108986 290134
rect 109222 289898 109404 290134
rect 108804 254454 109404 289898
rect 108804 254218 108986 254454
rect 109222 254218 109404 254454
rect 108804 254134 109404 254218
rect 108804 253898 108986 254134
rect 109222 253898 109404 254134
rect 108804 218454 109404 253898
rect 108804 218218 108986 218454
rect 109222 218218 109404 218454
rect 108804 218134 109404 218218
rect 108804 217898 108986 218134
rect 109222 217898 109404 218134
rect 108804 182454 109404 217898
rect 108804 182218 108986 182454
rect 109222 182218 109404 182454
rect 108804 182134 109404 182218
rect 108804 181898 108986 182134
rect 109222 181898 109404 182134
rect 108804 146454 109404 181898
rect 108804 146218 108986 146454
rect 109222 146218 109404 146454
rect 108804 146134 109404 146218
rect 108804 145898 108986 146134
rect 109222 145898 109404 146134
rect 108804 110454 109404 145898
rect 108804 110218 108986 110454
rect 109222 110218 109404 110454
rect 108804 110134 109404 110218
rect 108804 109898 108986 110134
rect 109222 109898 109404 110134
rect 108804 74454 109404 109898
rect 108804 74218 108986 74454
rect 109222 74218 109404 74454
rect 108804 74134 109404 74218
rect 108804 73898 108986 74134
rect 109222 73898 109404 74134
rect 108804 38454 109404 73898
rect 108804 38218 108986 38454
rect 109222 38218 109404 38454
rect 108804 38134 109404 38218
rect 108804 37898 108986 38134
rect 109222 37898 109404 38134
rect 108804 2454 109404 37898
rect 108804 2218 108986 2454
rect 109222 2218 109404 2454
rect 108804 2134 109404 2218
rect 108804 1898 108986 2134
rect 109222 1898 109404 2134
rect 108804 -346 109404 1898
rect 108804 -582 108986 -346
rect 109222 -582 109404 -346
rect 108804 -666 109404 -582
rect 108804 -902 108986 -666
rect 109222 -902 109404 -666
rect 108804 -1844 109404 -902
rect 112404 690054 113004 706122
rect 112404 689818 112586 690054
rect 112822 689818 113004 690054
rect 112404 689734 113004 689818
rect 112404 689498 112586 689734
rect 112822 689498 113004 689734
rect 112404 654054 113004 689498
rect 112404 653818 112586 654054
rect 112822 653818 113004 654054
rect 112404 653734 113004 653818
rect 112404 653498 112586 653734
rect 112822 653498 113004 653734
rect 112404 618054 113004 653498
rect 112404 617818 112586 618054
rect 112822 617818 113004 618054
rect 112404 617734 113004 617818
rect 112404 617498 112586 617734
rect 112822 617498 113004 617734
rect 112404 582054 113004 617498
rect 112404 581818 112586 582054
rect 112822 581818 113004 582054
rect 112404 581734 113004 581818
rect 112404 581498 112586 581734
rect 112822 581498 113004 581734
rect 112404 546054 113004 581498
rect 112404 545818 112586 546054
rect 112822 545818 113004 546054
rect 112404 545734 113004 545818
rect 112404 545498 112586 545734
rect 112822 545498 113004 545734
rect 112404 510054 113004 545498
rect 112404 509818 112586 510054
rect 112822 509818 113004 510054
rect 112404 509734 113004 509818
rect 112404 509498 112586 509734
rect 112822 509498 113004 509734
rect 112404 474054 113004 509498
rect 112404 473818 112586 474054
rect 112822 473818 113004 474054
rect 112404 473734 113004 473818
rect 112404 473498 112586 473734
rect 112822 473498 113004 473734
rect 112404 438054 113004 473498
rect 112404 437818 112586 438054
rect 112822 437818 113004 438054
rect 112404 437734 113004 437818
rect 112404 437498 112586 437734
rect 112822 437498 113004 437734
rect 112404 402054 113004 437498
rect 112404 401818 112586 402054
rect 112822 401818 113004 402054
rect 112404 401734 113004 401818
rect 112404 401498 112586 401734
rect 112822 401498 113004 401734
rect 112404 366054 113004 401498
rect 112404 365818 112586 366054
rect 112822 365818 113004 366054
rect 112404 365734 113004 365818
rect 112404 365498 112586 365734
rect 112822 365498 113004 365734
rect 112404 330054 113004 365498
rect 112404 329818 112586 330054
rect 112822 329818 113004 330054
rect 112404 329734 113004 329818
rect 112404 329498 112586 329734
rect 112822 329498 113004 329734
rect 112404 294054 113004 329498
rect 112404 293818 112586 294054
rect 112822 293818 113004 294054
rect 112404 293734 113004 293818
rect 112404 293498 112586 293734
rect 112822 293498 113004 293734
rect 112404 258054 113004 293498
rect 112404 257818 112586 258054
rect 112822 257818 113004 258054
rect 112404 257734 113004 257818
rect 112404 257498 112586 257734
rect 112822 257498 113004 257734
rect 112404 222054 113004 257498
rect 112404 221818 112586 222054
rect 112822 221818 113004 222054
rect 112404 221734 113004 221818
rect 112404 221498 112586 221734
rect 112822 221498 113004 221734
rect 112404 186054 113004 221498
rect 112404 185818 112586 186054
rect 112822 185818 113004 186054
rect 112404 185734 113004 185818
rect 112404 185498 112586 185734
rect 112822 185498 113004 185734
rect 112404 150054 113004 185498
rect 112404 149818 112586 150054
rect 112822 149818 113004 150054
rect 112404 149734 113004 149818
rect 112404 149498 112586 149734
rect 112822 149498 113004 149734
rect 112404 114054 113004 149498
rect 112404 113818 112586 114054
rect 112822 113818 113004 114054
rect 112404 113734 113004 113818
rect 112404 113498 112586 113734
rect 112822 113498 113004 113734
rect 112404 78054 113004 113498
rect 112404 77818 112586 78054
rect 112822 77818 113004 78054
rect 112404 77734 113004 77818
rect 112404 77498 112586 77734
rect 112822 77498 113004 77734
rect 112404 42054 113004 77498
rect 112404 41818 112586 42054
rect 112822 41818 113004 42054
rect 112404 41734 113004 41818
rect 112404 41498 112586 41734
rect 112822 41498 113004 41734
rect 112404 6054 113004 41498
rect 112404 5818 112586 6054
rect 112822 5818 113004 6054
rect 112404 5734 113004 5818
rect 112404 5498 112586 5734
rect 112822 5498 113004 5734
rect 112404 -2186 113004 5498
rect 112404 -2422 112586 -2186
rect 112822 -2422 113004 -2186
rect 112404 -2506 113004 -2422
rect 112404 -2742 112586 -2506
rect 112822 -2742 113004 -2506
rect 112404 -3684 113004 -2742
rect 116004 693654 116604 707962
rect 116004 693418 116186 693654
rect 116422 693418 116604 693654
rect 116004 693334 116604 693418
rect 116004 693098 116186 693334
rect 116422 693098 116604 693334
rect 116004 657654 116604 693098
rect 116004 657418 116186 657654
rect 116422 657418 116604 657654
rect 116004 657334 116604 657418
rect 116004 657098 116186 657334
rect 116422 657098 116604 657334
rect 116004 621654 116604 657098
rect 116004 621418 116186 621654
rect 116422 621418 116604 621654
rect 116004 621334 116604 621418
rect 116004 621098 116186 621334
rect 116422 621098 116604 621334
rect 116004 585654 116604 621098
rect 116004 585418 116186 585654
rect 116422 585418 116604 585654
rect 116004 585334 116604 585418
rect 116004 585098 116186 585334
rect 116422 585098 116604 585334
rect 116004 549654 116604 585098
rect 116004 549418 116186 549654
rect 116422 549418 116604 549654
rect 116004 549334 116604 549418
rect 116004 549098 116186 549334
rect 116422 549098 116604 549334
rect 116004 513654 116604 549098
rect 116004 513418 116186 513654
rect 116422 513418 116604 513654
rect 116004 513334 116604 513418
rect 116004 513098 116186 513334
rect 116422 513098 116604 513334
rect 116004 477654 116604 513098
rect 116004 477418 116186 477654
rect 116422 477418 116604 477654
rect 116004 477334 116604 477418
rect 116004 477098 116186 477334
rect 116422 477098 116604 477334
rect 116004 441654 116604 477098
rect 116004 441418 116186 441654
rect 116422 441418 116604 441654
rect 116004 441334 116604 441418
rect 116004 441098 116186 441334
rect 116422 441098 116604 441334
rect 116004 405654 116604 441098
rect 116004 405418 116186 405654
rect 116422 405418 116604 405654
rect 116004 405334 116604 405418
rect 116004 405098 116186 405334
rect 116422 405098 116604 405334
rect 116004 369654 116604 405098
rect 116004 369418 116186 369654
rect 116422 369418 116604 369654
rect 116004 369334 116604 369418
rect 116004 369098 116186 369334
rect 116422 369098 116604 369334
rect 116004 333654 116604 369098
rect 116004 333418 116186 333654
rect 116422 333418 116604 333654
rect 116004 333334 116604 333418
rect 116004 333098 116186 333334
rect 116422 333098 116604 333334
rect 116004 297654 116604 333098
rect 116004 297418 116186 297654
rect 116422 297418 116604 297654
rect 116004 297334 116604 297418
rect 116004 297098 116186 297334
rect 116422 297098 116604 297334
rect 116004 261654 116604 297098
rect 116004 261418 116186 261654
rect 116422 261418 116604 261654
rect 116004 261334 116604 261418
rect 116004 261098 116186 261334
rect 116422 261098 116604 261334
rect 116004 225654 116604 261098
rect 116004 225418 116186 225654
rect 116422 225418 116604 225654
rect 116004 225334 116604 225418
rect 116004 225098 116186 225334
rect 116422 225098 116604 225334
rect 116004 189654 116604 225098
rect 116004 189418 116186 189654
rect 116422 189418 116604 189654
rect 116004 189334 116604 189418
rect 116004 189098 116186 189334
rect 116422 189098 116604 189334
rect 116004 153654 116604 189098
rect 116004 153418 116186 153654
rect 116422 153418 116604 153654
rect 116004 153334 116604 153418
rect 116004 153098 116186 153334
rect 116422 153098 116604 153334
rect 116004 117654 116604 153098
rect 116004 117418 116186 117654
rect 116422 117418 116604 117654
rect 116004 117334 116604 117418
rect 116004 117098 116186 117334
rect 116422 117098 116604 117334
rect 116004 81654 116604 117098
rect 116004 81418 116186 81654
rect 116422 81418 116604 81654
rect 116004 81334 116604 81418
rect 116004 81098 116186 81334
rect 116422 81098 116604 81334
rect 116004 45654 116604 81098
rect 116004 45418 116186 45654
rect 116422 45418 116604 45654
rect 116004 45334 116604 45418
rect 116004 45098 116186 45334
rect 116422 45098 116604 45334
rect 116004 9654 116604 45098
rect 116004 9418 116186 9654
rect 116422 9418 116604 9654
rect 116004 9334 116604 9418
rect 116004 9098 116186 9334
rect 116422 9098 116604 9334
rect 116004 -4026 116604 9098
rect 116004 -4262 116186 -4026
rect 116422 -4262 116604 -4026
rect 116004 -4346 116604 -4262
rect 116004 -4582 116186 -4346
rect 116422 -4582 116604 -4346
rect 116004 -5524 116604 -4582
rect 119604 697254 120204 709802
rect 137604 711278 138204 711300
rect 137604 711042 137786 711278
rect 138022 711042 138204 711278
rect 137604 710958 138204 711042
rect 137604 710722 137786 710958
rect 138022 710722 138204 710958
rect 134004 709438 134604 709460
rect 134004 709202 134186 709438
rect 134422 709202 134604 709438
rect 134004 709118 134604 709202
rect 134004 708882 134186 709118
rect 134422 708882 134604 709118
rect 130404 707598 131004 707620
rect 130404 707362 130586 707598
rect 130822 707362 131004 707598
rect 130404 707278 131004 707362
rect 130404 707042 130586 707278
rect 130822 707042 131004 707278
rect 119604 697018 119786 697254
rect 120022 697018 120204 697254
rect 119604 696934 120204 697018
rect 119604 696698 119786 696934
rect 120022 696698 120204 696934
rect 119604 661254 120204 696698
rect 119604 661018 119786 661254
rect 120022 661018 120204 661254
rect 119604 660934 120204 661018
rect 119604 660698 119786 660934
rect 120022 660698 120204 660934
rect 119604 625254 120204 660698
rect 119604 625018 119786 625254
rect 120022 625018 120204 625254
rect 119604 624934 120204 625018
rect 119604 624698 119786 624934
rect 120022 624698 120204 624934
rect 119604 589254 120204 624698
rect 119604 589018 119786 589254
rect 120022 589018 120204 589254
rect 119604 588934 120204 589018
rect 119604 588698 119786 588934
rect 120022 588698 120204 588934
rect 119604 553254 120204 588698
rect 119604 553018 119786 553254
rect 120022 553018 120204 553254
rect 119604 552934 120204 553018
rect 119604 552698 119786 552934
rect 120022 552698 120204 552934
rect 119604 517254 120204 552698
rect 119604 517018 119786 517254
rect 120022 517018 120204 517254
rect 119604 516934 120204 517018
rect 119604 516698 119786 516934
rect 120022 516698 120204 516934
rect 119604 481254 120204 516698
rect 119604 481018 119786 481254
rect 120022 481018 120204 481254
rect 119604 480934 120204 481018
rect 119604 480698 119786 480934
rect 120022 480698 120204 480934
rect 119604 445254 120204 480698
rect 119604 445018 119786 445254
rect 120022 445018 120204 445254
rect 119604 444934 120204 445018
rect 119604 444698 119786 444934
rect 120022 444698 120204 444934
rect 119604 409254 120204 444698
rect 119604 409018 119786 409254
rect 120022 409018 120204 409254
rect 119604 408934 120204 409018
rect 119604 408698 119786 408934
rect 120022 408698 120204 408934
rect 119604 373254 120204 408698
rect 119604 373018 119786 373254
rect 120022 373018 120204 373254
rect 119604 372934 120204 373018
rect 119604 372698 119786 372934
rect 120022 372698 120204 372934
rect 119604 337254 120204 372698
rect 119604 337018 119786 337254
rect 120022 337018 120204 337254
rect 119604 336934 120204 337018
rect 119604 336698 119786 336934
rect 120022 336698 120204 336934
rect 119604 301254 120204 336698
rect 119604 301018 119786 301254
rect 120022 301018 120204 301254
rect 119604 300934 120204 301018
rect 119604 300698 119786 300934
rect 120022 300698 120204 300934
rect 119604 265254 120204 300698
rect 119604 265018 119786 265254
rect 120022 265018 120204 265254
rect 119604 264934 120204 265018
rect 119604 264698 119786 264934
rect 120022 264698 120204 264934
rect 119604 229254 120204 264698
rect 119604 229018 119786 229254
rect 120022 229018 120204 229254
rect 119604 228934 120204 229018
rect 119604 228698 119786 228934
rect 120022 228698 120204 228934
rect 119604 193254 120204 228698
rect 119604 193018 119786 193254
rect 120022 193018 120204 193254
rect 119604 192934 120204 193018
rect 119604 192698 119786 192934
rect 120022 192698 120204 192934
rect 119604 157254 120204 192698
rect 119604 157018 119786 157254
rect 120022 157018 120204 157254
rect 119604 156934 120204 157018
rect 119604 156698 119786 156934
rect 120022 156698 120204 156934
rect 119604 121254 120204 156698
rect 119604 121018 119786 121254
rect 120022 121018 120204 121254
rect 119604 120934 120204 121018
rect 119604 120698 119786 120934
rect 120022 120698 120204 120934
rect 119604 85254 120204 120698
rect 119604 85018 119786 85254
rect 120022 85018 120204 85254
rect 119604 84934 120204 85018
rect 119604 84698 119786 84934
rect 120022 84698 120204 84934
rect 119604 49254 120204 84698
rect 119604 49018 119786 49254
rect 120022 49018 120204 49254
rect 119604 48934 120204 49018
rect 119604 48698 119786 48934
rect 120022 48698 120204 48934
rect 119604 13254 120204 48698
rect 119604 13018 119786 13254
rect 120022 13018 120204 13254
rect 119604 12934 120204 13018
rect 119604 12698 119786 12934
rect 120022 12698 120204 12934
rect 101604 -7022 101786 -6786
rect 102022 -7022 102204 -6786
rect 101604 -7106 102204 -7022
rect 101604 -7342 101786 -7106
rect 102022 -7342 102204 -7106
rect 101604 -7364 102204 -7342
rect 119604 -5866 120204 12698
rect 126804 705758 127404 705780
rect 126804 705522 126986 705758
rect 127222 705522 127404 705758
rect 126804 705438 127404 705522
rect 126804 705202 126986 705438
rect 127222 705202 127404 705438
rect 126804 668454 127404 705202
rect 126804 668218 126986 668454
rect 127222 668218 127404 668454
rect 126804 668134 127404 668218
rect 126804 667898 126986 668134
rect 127222 667898 127404 668134
rect 126804 632454 127404 667898
rect 126804 632218 126986 632454
rect 127222 632218 127404 632454
rect 126804 632134 127404 632218
rect 126804 631898 126986 632134
rect 127222 631898 127404 632134
rect 126804 596454 127404 631898
rect 126804 596218 126986 596454
rect 127222 596218 127404 596454
rect 126804 596134 127404 596218
rect 126804 595898 126986 596134
rect 127222 595898 127404 596134
rect 126804 560454 127404 595898
rect 126804 560218 126986 560454
rect 127222 560218 127404 560454
rect 126804 560134 127404 560218
rect 126804 559898 126986 560134
rect 127222 559898 127404 560134
rect 126804 524454 127404 559898
rect 126804 524218 126986 524454
rect 127222 524218 127404 524454
rect 126804 524134 127404 524218
rect 126804 523898 126986 524134
rect 127222 523898 127404 524134
rect 126804 488454 127404 523898
rect 126804 488218 126986 488454
rect 127222 488218 127404 488454
rect 126804 488134 127404 488218
rect 126804 487898 126986 488134
rect 127222 487898 127404 488134
rect 126804 452454 127404 487898
rect 126804 452218 126986 452454
rect 127222 452218 127404 452454
rect 126804 452134 127404 452218
rect 126804 451898 126986 452134
rect 127222 451898 127404 452134
rect 126804 416454 127404 451898
rect 126804 416218 126986 416454
rect 127222 416218 127404 416454
rect 126804 416134 127404 416218
rect 126804 415898 126986 416134
rect 127222 415898 127404 416134
rect 126804 380454 127404 415898
rect 126804 380218 126986 380454
rect 127222 380218 127404 380454
rect 126804 380134 127404 380218
rect 126804 379898 126986 380134
rect 127222 379898 127404 380134
rect 126804 344454 127404 379898
rect 126804 344218 126986 344454
rect 127222 344218 127404 344454
rect 126804 344134 127404 344218
rect 126804 343898 126986 344134
rect 127222 343898 127404 344134
rect 126804 308454 127404 343898
rect 126804 308218 126986 308454
rect 127222 308218 127404 308454
rect 126804 308134 127404 308218
rect 126804 307898 126986 308134
rect 127222 307898 127404 308134
rect 126804 272454 127404 307898
rect 126804 272218 126986 272454
rect 127222 272218 127404 272454
rect 126804 272134 127404 272218
rect 126804 271898 126986 272134
rect 127222 271898 127404 272134
rect 126804 236454 127404 271898
rect 126804 236218 126986 236454
rect 127222 236218 127404 236454
rect 126804 236134 127404 236218
rect 126804 235898 126986 236134
rect 127222 235898 127404 236134
rect 126804 200454 127404 235898
rect 126804 200218 126986 200454
rect 127222 200218 127404 200454
rect 126804 200134 127404 200218
rect 126804 199898 126986 200134
rect 127222 199898 127404 200134
rect 126804 164454 127404 199898
rect 126804 164218 126986 164454
rect 127222 164218 127404 164454
rect 126804 164134 127404 164218
rect 126804 163898 126986 164134
rect 127222 163898 127404 164134
rect 126804 128454 127404 163898
rect 126804 128218 126986 128454
rect 127222 128218 127404 128454
rect 126804 128134 127404 128218
rect 126804 127898 126986 128134
rect 127222 127898 127404 128134
rect 126804 92454 127404 127898
rect 126804 92218 126986 92454
rect 127222 92218 127404 92454
rect 126804 92134 127404 92218
rect 126804 91898 126986 92134
rect 127222 91898 127404 92134
rect 126804 56454 127404 91898
rect 126804 56218 126986 56454
rect 127222 56218 127404 56454
rect 126804 56134 127404 56218
rect 126804 55898 126986 56134
rect 127222 55898 127404 56134
rect 126804 20454 127404 55898
rect 126804 20218 126986 20454
rect 127222 20218 127404 20454
rect 126804 20134 127404 20218
rect 126804 19898 126986 20134
rect 127222 19898 127404 20134
rect 126804 -1266 127404 19898
rect 126804 -1502 126986 -1266
rect 127222 -1502 127404 -1266
rect 126804 -1586 127404 -1502
rect 126804 -1822 126986 -1586
rect 127222 -1822 127404 -1586
rect 126804 -1844 127404 -1822
rect 130404 672054 131004 707042
rect 130404 671818 130586 672054
rect 130822 671818 131004 672054
rect 130404 671734 131004 671818
rect 130404 671498 130586 671734
rect 130822 671498 131004 671734
rect 130404 636054 131004 671498
rect 130404 635818 130586 636054
rect 130822 635818 131004 636054
rect 130404 635734 131004 635818
rect 130404 635498 130586 635734
rect 130822 635498 131004 635734
rect 130404 600054 131004 635498
rect 130404 599818 130586 600054
rect 130822 599818 131004 600054
rect 130404 599734 131004 599818
rect 130404 599498 130586 599734
rect 130822 599498 131004 599734
rect 130404 564054 131004 599498
rect 130404 563818 130586 564054
rect 130822 563818 131004 564054
rect 130404 563734 131004 563818
rect 130404 563498 130586 563734
rect 130822 563498 131004 563734
rect 130404 528054 131004 563498
rect 130404 527818 130586 528054
rect 130822 527818 131004 528054
rect 130404 527734 131004 527818
rect 130404 527498 130586 527734
rect 130822 527498 131004 527734
rect 130404 492054 131004 527498
rect 130404 491818 130586 492054
rect 130822 491818 131004 492054
rect 130404 491734 131004 491818
rect 130404 491498 130586 491734
rect 130822 491498 131004 491734
rect 130404 456054 131004 491498
rect 130404 455818 130586 456054
rect 130822 455818 131004 456054
rect 130404 455734 131004 455818
rect 130404 455498 130586 455734
rect 130822 455498 131004 455734
rect 130404 420054 131004 455498
rect 130404 419818 130586 420054
rect 130822 419818 131004 420054
rect 130404 419734 131004 419818
rect 130404 419498 130586 419734
rect 130822 419498 131004 419734
rect 130404 384054 131004 419498
rect 130404 383818 130586 384054
rect 130822 383818 131004 384054
rect 130404 383734 131004 383818
rect 130404 383498 130586 383734
rect 130822 383498 131004 383734
rect 130404 348054 131004 383498
rect 130404 347818 130586 348054
rect 130822 347818 131004 348054
rect 130404 347734 131004 347818
rect 130404 347498 130586 347734
rect 130822 347498 131004 347734
rect 130404 312054 131004 347498
rect 130404 311818 130586 312054
rect 130822 311818 131004 312054
rect 130404 311734 131004 311818
rect 130404 311498 130586 311734
rect 130822 311498 131004 311734
rect 130404 276054 131004 311498
rect 130404 275818 130586 276054
rect 130822 275818 131004 276054
rect 130404 275734 131004 275818
rect 130404 275498 130586 275734
rect 130822 275498 131004 275734
rect 130404 240054 131004 275498
rect 130404 239818 130586 240054
rect 130822 239818 131004 240054
rect 130404 239734 131004 239818
rect 130404 239498 130586 239734
rect 130822 239498 131004 239734
rect 130404 204054 131004 239498
rect 130404 203818 130586 204054
rect 130822 203818 131004 204054
rect 130404 203734 131004 203818
rect 130404 203498 130586 203734
rect 130822 203498 131004 203734
rect 130404 168054 131004 203498
rect 130404 167818 130586 168054
rect 130822 167818 131004 168054
rect 130404 167734 131004 167818
rect 130404 167498 130586 167734
rect 130822 167498 131004 167734
rect 130404 132054 131004 167498
rect 130404 131818 130586 132054
rect 130822 131818 131004 132054
rect 130404 131734 131004 131818
rect 130404 131498 130586 131734
rect 130822 131498 131004 131734
rect 130404 96054 131004 131498
rect 130404 95818 130586 96054
rect 130822 95818 131004 96054
rect 130404 95734 131004 95818
rect 130404 95498 130586 95734
rect 130822 95498 131004 95734
rect 130404 60054 131004 95498
rect 130404 59818 130586 60054
rect 130822 59818 131004 60054
rect 130404 59734 131004 59818
rect 130404 59498 130586 59734
rect 130822 59498 131004 59734
rect 130404 24054 131004 59498
rect 130404 23818 130586 24054
rect 130822 23818 131004 24054
rect 130404 23734 131004 23818
rect 130404 23498 130586 23734
rect 130822 23498 131004 23734
rect 130404 -3106 131004 23498
rect 130404 -3342 130586 -3106
rect 130822 -3342 131004 -3106
rect 130404 -3426 131004 -3342
rect 130404 -3662 130586 -3426
rect 130822 -3662 131004 -3426
rect 130404 -3684 131004 -3662
rect 134004 675654 134604 708882
rect 134004 675418 134186 675654
rect 134422 675418 134604 675654
rect 134004 675334 134604 675418
rect 134004 675098 134186 675334
rect 134422 675098 134604 675334
rect 134004 639654 134604 675098
rect 134004 639418 134186 639654
rect 134422 639418 134604 639654
rect 134004 639334 134604 639418
rect 134004 639098 134186 639334
rect 134422 639098 134604 639334
rect 134004 603654 134604 639098
rect 134004 603418 134186 603654
rect 134422 603418 134604 603654
rect 134004 603334 134604 603418
rect 134004 603098 134186 603334
rect 134422 603098 134604 603334
rect 134004 567654 134604 603098
rect 134004 567418 134186 567654
rect 134422 567418 134604 567654
rect 134004 567334 134604 567418
rect 134004 567098 134186 567334
rect 134422 567098 134604 567334
rect 134004 531654 134604 567098
rect 134004 531418 134186 531654
rect 134422 531418 134604 531654
rect 134004 531334 134604 531418
rect 134004 531098 134186 531334
rect 134422 531098 134604 531334
rect 134004 495654 134604 531098
rect 134004 495418 134186 495654
rect 134422 495418 134604 495654
rect 134004 495334 134604 495418
rect 134004 495098 134186 495334
rect 134422 495098 134604 495334
rect 134004 459654 134604 495098
rect 134004 459418 134186 459654
rect 134422 459418 134604 459654
rect 134004 459334 134604 459418
rect 134004 459098 134186 459334
rect 134422 459098 134604 459334
rect 134004 423654 134604 459098
rect 134004 423418 134186 423654
rect 134422 423418 134604 423654
rect 134004 423334 134604 423418
rect 134004 423098 134186 423334
rect 134422 423098 134604 423334
rect 134004 387654 134604 423098
rect 134004 387418 134186 387654
rect 134422 387418 134604 387654
rect 134004 387334 134604 387418
rect 134004 387098 134186 387334
rect 134422 387098 134604 387334
rect 134004 351654 134604 387098
rect 134004 351418 134186 351654
rect 134422 351418 134604 351654
rect 134004 351334 134604 351418
rect 134004 351098 134186 351334
rect 134422 351098 134604 351334
rect 134004 315654 134604 351098
rect 134004 315418 134186 315654
rect 134422 315418 134604 315654
rect 134004 315334 134604 315418
rect 134004 315098 134186 315334
rect 134422 315098 134604 315334
rect 134004 279654 134604 315098
rect 134004 279418 134186 279654
rect 134422 279418 134604 279654
rect 134004 279334 134604 279418
rect 134004 279098 134186 279334
rect 134422 279098 134604 279334
rect 134004 243654 134604 279098
rect 134004 243418 134186 243654
rect 134422 243418 134604 243654
rect 134004 243334 134604 243418
rect 134004 243098 134186 243334
rect 134422 243098 134604 243334
rect 134004 207654 134604 243098
rect 134004 207418 134186 207654
rect 134422 207418 134604 207654
rect 134004 207334 134604 207418
rect 134004 207098 134186 207334
rect 134422 207098 134604 207334
rect 134004 171654 134604 207098
rect 134004 171418 134186 171654
rect 134422 171418 134604 171654
rect 134004 171334 134604 171418
rect 134004 171098 134186 171334
rect 134422 171098 134604 171334
rect 134004 135654 134604 171098
rect 134004 135418 134186 135654
rect 134422 135418 134604 135654
rect 134004 135334 134604 135418
rect 134004 135098 134186 135334
rect 134422 135098 134604 135334
rect 134004 99654 134604 135098
rect 134004 99418 134186 99654
rect 134422 99418 134604 99654
rect 134004 99334 134604 99418
rect 134004 99098 134186 99334
rect 134422 99098 134604 99334
rect 134004 63654 134604 99098
rect 134004 63418 134186 63654
rect 134422 63418 134604 63654
rect 134004 63334 134604 63418
rect 134004 63098 134186 63334
rect 134422 63098 134604 63334
rect 134004 27654 134604 63098
rect 134004 27418 134186 27654
rect 134422 27418 134604 27654
rect 134004 27334 134604 27418
rect 134004 27098 134186 27334
rect 134422 27098 134604 27334
rect 134004 -4946 134604 27098
rect 134004 -5182 134186 -4946
rect 134422 -5182 134604 -4946
rect 134004 -5266 134604 -5182
rect 134004 -5502 134186 -5266
rect 134422 -5502 134604 -5266
rect 134004 -5524 134604 -5502
rect 137604 679254 138204 710722
rect 155604 710358 156204 711300
rect 155604 710122 155786 710358
rect 156022 710122 156204 710358
rect 155604 710038 156204 710122
rect 155604 709802 155786 710038
rect 156022 709802 156204 710038
rect 152004 708518 152604 709460
rect 152004 708282 152186 708518
rect 152422 708282 152604 708518
rect 152004 708198 152604 708282
rect 152004 707962 152186 708198
rect 152422 707962 152604 708198
rect 148404 706678 149004 707620
rect 148404 706442 148586 706678
rect 148822 706442 149004 706678
rect 148404 706358 149004 706442
rect 148404 706122 148586 706358
rect 148822 706122 149004 706358
rect 137604 679018 137786 679254
rect 138022 679018 138204 679254
rect 137604 678934 138204 679018
rect 137604 678698 137786 678934
rect 138022 678698 138204 678934
rect 137604 643254 138204 678698
rect 137604 643018 137786 643254
rect 138022 643018 138204 643254
rect 137604 642934 138204 643018
rect 137604 642698 137786 642934
rect 138022 642698 138204 642934
rect 137604 607254 138204 642698
rect 137604 607018 137786 607254
rect 138022 607018 138204 607254
rect 137604 606934 138204 607018
rect 137604 606698 137786 606934
rect 138022 606698 138204 606934
rect 137604 571254 138204 606698
rect 137604 571018 137786 571254
rect 138022 571018 138204 571254
rect 137604 570934 138204 571018
rect 137604 570698 137786 570934
rect 138022 570698 138204 570934
rect 137604 535254 138204 570698
rect 137604 535018 137786 535254
rect 138022 535018 138204 535254
rect 137604 534934 138204 535018
rect 137604 534698 137786 534934
rect 138022 534698 138204 534934
rect 137604 499254 138204 534698
rect 137604 499018 137786 499254
rect 138022 499018 138204 499254
rect 137604 498934 138204 499018
rect 137604 498698 137786 498934
rect 138022 498698 138204 498934
rect 137604 463254 138204 498698
rect 137604 463018 137786 463254
rect 138022 463018 138204 463254
rect 137604 462934 138204 463018
rect 137604 462698 137786 462934
rect 138022 462698 138204 462934
rect 137604 427254 138204 462698
rect 137604 427018 137786 427254
rect 138022 427018 138204 427254
rect 137604 426934 138204 427018
rect 137604 426698 137786 426934
rect 138022 426698 138204 426934
rect 137604 391254 138204 426698
rect 137604 391018 137786 391254
rect 138022 391018 138204 391254
rect 137604 390934 138204 391018
rect 137604 390698 137786 390934
rect 138022 390698 138204 390934
rect 137604 355254 138204 390698
rect 137604 355018 137786 355254
rect 138022 355018 138204 355254
rect 137604 354934 138204 355018
rect 137604 354698 137786 354934
rect 138022 354698 138204 354934
rect 137604 319254 138204 354698
rect 137604 319018 137786 319254
rect 138022 319018 138204 319254
rect 137604 318934 138204 319018
rect 137604 318698 137786 318934
rect 138022 318698 138204 318934
rect 137604 283254 138204 318698
rect 137604 283018 137786 283254
rect 138022 283018 138204 283254
rect 137604 282934 138204 283018
rect 137604 282698 137786 282934
rect 138022 282698 138204 282934
rect 137604 247254 138204 282698
rect 137604 247018 137786 247254
rect 138022 247018 138204 247254
rect 137604 246934 138204 247018
rect 137604 246698 137786 246934
rect 138022 246698 138204 246934
rect 137604 211254 138204 246698
rect 137604 211018 137786 211254
rect 138022 211018 138204 211254
rect 137604 210934 138204 211018
rect 137604 210698 137786 210934
rect 138022 210698 138204 210934
rect 137604 175254 138204 210698
rect 137604 175018 137786 175254
rect 138022 175018 138204 175254
rect 137604 174934 138204 175018
rect 137604 174698 137786 174934
rect 138022 174698 138204 174934
rect 137604 139254 138204 174698
rect 137604 139018 137786 139254
rect 138022 139018 138204 139254
rect 137604 138934 138204 139018
rect 137604 138698 137786 138934
rect 138022 138698 138204 138934
rect 137604 103254 138204 138698
rect 137604 103018 137786 103254
rect 138022 103018 138204 103254
rect 137604 102934 138204 103018
rect 137604 102698 137786 102934
rect 138022 102698 138204 102934
rect 137604 67254 138204 102698
rect 137604 67018 137786 67254
rect 138022 67018 138204 67254
rect 137604 66934 138204 67018
rect 137604 66698 137786 66934
rect 138022 66698 138204 66934
rect 137604 31254 138204 66698
rect 137604 31018 137786 31254
rect 138022 31018 138204 31254
rect 137604 30934 138204 31018
rect 137604 30698 137786 30934
rect 138022 30698 138204 30934
rect 119604 -6102 119786 -5866
rect 120022 -6102 120204 -5866
rect 119604 -6186 120204 -6102
rect 119604 -6422 119786 -6186
rect 120022 -6422 120204 -6186
rect 119604 -7364 120204 -6422
rect 137604 -6786 138204 30698
rect 144804 704838 145404 705780
rect 144804 704602 144986 704838
rect 145222 704602 145404 704838
rect 144804 704518 145404 704602
rect 144804 704282 144986 704518
rect 145222 704282 145404 704518
rect 144804 686454 145404 704282
rect 144804 686218 144986 686454
rect 145222 686218 145404 686454
rect 144804 686134 145404 686218
rect 144804 685898 144986 686134
rect 145222 685898 145404 686134
rect 144804 650454 145404 685898
rect 144804 650218 144986 650454
rect 145222 650218 145404 650454
rect 144804 650134 145404 650218
rect 144804 649898 144986 650134
rect 145222 649898 145404 650134
rect 144804 614454 145404 649898
rect 144804 614218 144986 614454
rect 145222 614218 145404 614454
rect 144804 614134 145404 614218
rect 144804 613898 144986 614134
rect 145222 613898 145404 614134
rect 144804 578454 145404 613898
rect 144804 578218 144986 578454
rect 145222 578218 145404 578454
rect 144804 578134 145404 578218
rect 144804 577898 144986 578134
rect 145222 577898 145404 578134
rect 144804 542454 145404 577898
rect 144804 542218 144986 542454
rect 145222 542218 145404 542454
rect 144804 542134 145404 542218
rect 144804 541898 144986 542134
rect 145222 541898 145404 542134
rect 144804 506454 145404 541898
rect 144804 506218 144986 506454
rect 145222 506218 145404 506454
rect 144804 506134 145404 506218
rect 144804 505898 144986 506134
rect 145222 505898 145404 506134
rect 144804 470454 145404 505898
rect 144804 470218 144986 470454
rect 145222 470218 145404 470454
rect 144804 470134 145404 470218
rect 144804 469898 144986 470134
rect 145222 469898 145404 470134
rect 144804 434454 145404 469898
rect 144804 434218 144986 434454
rect 145222 434218 145404 434454
rect 144804 434134 145404 434218
rect 144804 433898 144986 434134
rect 145222 433898 145404 434134
rect 144804 398454 145404 433898
rect 144804 398218 144986 398454
rect 145222 398218 145404 398454
rect 144804 398134 145404 398218
rect 144804 397898 144986 398134
rect 145222 397898 145404 398134
rect 144804 362454 145404 397898
rect 144804 362218 144986 362454
rect 145222 362218 145404 362454
rect 144804 362134 145404 362218
rect 144804 361898 144986 362134
rect 145222 361898 145404 362134
rect 144804 326454 145404 361898
rect 144804 326218 144986 326454
rect 145222 326218 145404 326454
rect 144804 326134 145404 326218
rect 144804 325898 144986 326134
rect 145222 325898 145404 326134
rect 144804 290454 145404 325898
rect 144804 290218 144986 290454
rect 145222 290218 145404 290454
rect 144804 290134 145404 290218
rect 144804 289898 144986 290134
rect 145222 289898 145404 290134
rect 144804 254454 145404 289898
rect 144804 254218 144986 254454
rect 145222 254218 145404 254454
rect 144804 254134 145404 254218
rect 144804 253898 144986 254134
rect 145222 253898 145404 254134
rect 144804 218454 145404 253898
rect 144804 218218 144986 218454
rect 145222 218218 145404 218454
rect 144804 218134 145404 218218
rect 144804 217898 144986 218134
rect 145222 217898 145404 218134
rect 144804 182454 145404 217898
rect 144804 182218 144986 182454
rect 145222 182218 145404 182454
rect 144804 182134 145404 182218
rect 144804 181898 144986 182134
rect 145222 181898 145404 182134
rect 144804 146454 145404 181898
rect 144804 146218 144986 146454
rect 145222 146218 145404 146454
rect 144804 146134 145404 146218
rect 144804 145898 144986 146134
rect 145222 145898 145404 146134
rect 144804 110454 145404 145898
rect 144804 110218 144986 110454
rect 145222 110218 145404 110454
rect 144804 110134 145404 110218
rect 144804 109898 144986 110134
rect 145222 109898 145404 110134
rect 144804 74454 145404 109898
rect 144804 74218 144986 74454
rect 145222 74218 145404 74454
rect 144804 74134 145404 74218
rect 144804 73898 144986 74134
rect 145222 73898 145404 74134
rect 144804 38454 145404 73898
rect 144804 38218 144986 38454
rect 145222 38218 145404 38454
rect 144804 38134 145404 38218
rect 144804 37898 144986 38134
rect 145222 37898 145404 38134
rect 144804 2454 145404 37898
rect 144804 2218 144986 2454
rect 145222 2218 145404 2454
rect 144804 2134 145404 2218
rect 144804 1898 144986 2134
rect 145222 1898 145404 2134
rect 144804 -346 145404 1898
rect 144804 -582 144986 -346
rect 145222 -582 145404 -346
rect 144804 -666 145404 -582
rect 144804 -902 144986 -666
rect 145222 -902 145404 -666
rect 144804 -1844 145404 -902
rect 148404 690054 149004 706122
rect 148404 689818 148586 690054
rect 148822 689818 149004 690054
rect 148404 689734 149004 689818
rect 148404 689498 148586 689734
rect 148822 689498 149004 689734
rect 148404 654054 149004 689498
rect 148404 653818 148586 654054
rect 148822 653818 149004 654054
rect 148404 653734 149004 653818
rect 148404 653498 148586 653734
rect 148822 653498 149004 653734
rect 148404 618054 149004 653498
rect 148404 617818 148586 618054
rect 148822 617818 149004 618054
rect 148404 617734 149004 617818
rect 148404 617498 148586 617734
rect 148822 617498 149004 617734
rect 148404 582054 149004 617498
rect 148404 581818 148586 582054
rect 148822 581818 149004 582054
rect 148404 581734 149004 581818
rect 148404 581498 148586 581734
rect 148822 581498 149004 581734
rect 148404 546054 149004 581498
rect 148404 545818 148586 546054
rect 148822 545818 149004 546054
rect 148404 545734 149004 545818
rect 148404 545498 148586 545734
rect 148822 545498 149004 545734
rect 148404 510054 149004 545498
rect 148404 509818 148586 510054
rect 148822 509818 149004 510054
rect 148404 509734 149004 509818
rect 148404 509498 148586 509734
rect 148822 509498 149004 509734
rect 148404 474054 149004 509498
rect 148404 473818 148586 474054
rect 148822 473818 149004 474054
rect 148404 473734 149004 473818
rect 148404 473498 148586 473734
rect 148822 473498 149004 473734
rect 148404 438054 149004 473498
rect 148404 437818 148586 438054
rect 148822 437818 149004 438054
rect 148404 437734 149004 437818
rect 148404 437498 148586 437734
rect 148822 437498 149004 437734
rect 148404 402054 149004 437498
rect 148404 401818 148586 402054
rect 148822 401818 149004 402054
rect 148404 401734 149004 401818
rect 148404 401498 148586 401734
rect 148822 401498 149004 401734
rect 148404 366054 149004 401498
rect 148404 365818 148586 366054
rect 148822 365818 149004 366054
rect 148404 365734 149004 365818
rect 148404 365498 148586 365734
rect 148822 365498 149004 365734
rect 148404 330054 149004 365498
rect 148404 329818 148586 330054
rect 148822 329818 149004 330054
rect 148404 329734 149004 329818
rect 148404 329498 148586 329734
rect 148822 329498 149004 329734
rect 148404 294054 149004 329498
rect 148404 293818 148586 294054
rect 148822 293818 149004 294054
rect 148404 293734 149004 293818
rect 148404 293498 148586 293734
rect 148822 293498 149004 293734
rect 148404 258054 149004 293498
rect 148404 257818 148586 258054
rect 148822 257818 149004 258054
rect 148404 257734 149004 257818
rect 148404 257498 148586 257734
rect 148822 257498 149004 257734
rect 148404 222054 149004 257498
rect 148404 221818 148586 222054
rect 148822 221818 149004 222054
rect 148404 221734 149004 221818
rect 148404 221498 148586 221734
rect 148822 221498 149004 221734
rect 148404 186054 149004 221498
rect 148404 185818 148586 186054
rect 148822 185818 149004 186054
rect 148404 185734 149004 185818
rect 148404 185498 148586 185734
rect 148822 185498 149004 185734
rect 148404 150054 149004 185498
rect 148404 149818 148586 150054
rect 148822 149818 149004 150054
rect 148404 149734 149004 149818
rect 148404 149498 148586 149734
rect 148822 149498 149004 149734
rect 148404 114054 149004 149498
rect 148404 113818 148586 114054
rect 148822 113818 149004 114054
rect 148404 113734 149004 113818
rect 148404 113498 148586 113734
rect 148822 113498 149004 113734
rect 148404 78054 149004 113498
rect 148404 77818 148586 78054
rect 148822 77818 149004 78054
rect 148404 77734 149004 77818
rect 148404 77498 148586 77734
rect 148822 77498 149004 77734
rect 148404 42054 149004 77498
rect 148404 41818 148586 42054
rect 148822 41818 149004 42054
rect 148404 41734 149004 41818
rect 148404 41498 148586 41734
rect 148822 41498 149004 41734
rect 148404 6054 149004 41498
rect 148404 5818 148586 6054
rect 148822 5818 149004 6054
rect 148404 5734 149004 5818
rect 148404 5498 148586 5734
rect 148822 5498 149004 5734
rect 148404 -2186 149004 5498
rect 148404 -2422 148586 -2186
rect 148822 -2422 149004 -2186
rect 148404 -2506 149004 -2422
rect 148404 -2742 148586 -2506
rect 148822 -2742 149004 -2506
rect 148404 -3684 149004 -2742
rect 152004 693654 152604 707962
rect 152004 693418 152186 693654
rect 152422 693418 152604 693654
rect 152004 693334 152604 693418
rect 152004 693098 152186 693334
rect 152422 693098 152604 693334
rect 152004 657654 152604 693098
rect 152004 657418 152186 657654
rect 152422 657418 152604 657654
rect 152004 657334 152604 657418
rect 152004 657098 152186 657334
rect 152422 657098 152604 657334
rect 152004 621654 152604 657098
rect 152004 621418 152186 621654
rect 152422 621418 152604 621654
rect 152004 621334 152604 621418
rect 152004 621098 152186 621334
rect 152422 621098 152604 621334
rect 152004 585654 152604 621098
rect 152004 585418 152186 585654
rect 152422 585418 152604 585654
rect 152004 585334 152604 585418
rect 152004 585098 152186 585334
rect 152422 585098 152604 585334
rect 152004 549654 152604 585098
rect 152004 549418 152186 549654
rect 152422 549418 152604 549654
rect 152004 549334 152604 549418
rect 152004 549098 152186 549334
rect 152422 549098 152604 549334
rect 152004 513654 152604 549098
rect 152004 513418 152186 513654
rect 152422 513418 152604 513654
rect 152004 513334 152604 513418
rect 152004 513098 152186 513334
rect 152422 513098 152604 513334
rect 152004 477654 152604 513098
rect 152004 477418 152186 477654
rect 152422 477418 152604 477654
rect 152004 477334 152604 477418
rect 152004 477098 152186 477334
rect 152422 477098 152604 477334
rect 152004 441654 152604 477098
rect 152004 441418 152186 441654
rect 152422 441418 152604 441654
rect 152004 441334 152604 441418
rect 152004 441098 152186 441334
rect 152422 441098 152604 441334
rect 152004 405654 152604 441098
rect 152004 405418 152186 405654
rect 152422 405418 152604 405654
rect 152004 405334 152604 405418
rect 152004 405098 152186 405334
rect 152422 405098 152604 405334
rect 152004 369654 152604 405098
rect 152004 369418 152186 369654
rect 152422 369418 152604 369654
rect 152004 369334 152604 369418
rect 152004 369098 152186 369334
rect 152422 369098 152604 369334
rect 152004 333654 152604 369098
rect 152004 333418 152186 333654
rect 152422 333418 152604 333654
rect 152004 333334 152604 333418
rect 152004 333098 152186 333334
rect 152422 333098 152604 333334
rect 152004 297654 152604 333098
rect 152004 297418 152186 297654
rect 152422 297418 152604 297654
rect 152004 297334 152604 297418
rect 152004 297098 152186 297334
rect 152422 297098 152604 297334
rect 152004 261654 152604 297098
rect 152004 261418 152186 261654
rect 152422 261418 152604 261654
rect 152004 261334 152604 261418
rect 152004 261098 152186 261334
rect 152422 261098 152604 261334
rect 152004 225654 152604 261098
rect 152004 225418 152186 225654
rect 152422 225418 152604 225654
rect 152004 225334 152604 225418
rect 152004 225098 152186 225334
rect 152422 225098 152604 225334
rect 152004 189654 152604 225098
rect 152004 189418 152186 189654
rect 152422 189418 152604 189654
rect 152004 189334 152604 189418
rect 152004 189098 152186 189334
rect 152422 189098 152604 189334
rect 152004 153654 152604 189098
rect 152004 153418 152186 153654
rect 152422 153418 152604 153654
rect 152004 153334 152604 153418
rect 152004 153098 152186 153334
rect 152422 153098 152604 153334
rect 152004 117654 152604 153098
rect 152004 117418 152186 117654
rect 152422 117418 152604 117654
rect 152004 117334 152604 117418
rect 152004 117098 152186 117334
rect 152422 117098 152604 117334
rect 152004 81654 152604 117098
rect 152004 81418 152186 81654
rect 152422 81418 152604 81654
rect 152004 81334 152604 81418
rect 152004 81098 152186 81334
rect 152422 81098 152604 81334
rect 152004 45654 152604 81098
rect 152004 45418 152186 45654
rect 152422 45418 152604 45654
rect 152004 45334 152604 45418
rect 152004 45098 152186 45334
rect 152422 45098 152604 45334
rect 152004 9654 152604 45098
rect 152004 9418 152186 9654
rect 152422 9418 152604 9654
rect 152004 9334 152604 9418
rect 152004 9098 152186 9334
rect 152422 9098 152604 9334
rect 152004 -4026 152604 9098
rect 152004 -4262 152186 -4026
rect 152422 -4262 152604 -4026
rect 152004 -4346 152604 -4262
rect 152004 -4582 152186 -4346
rect 152422 -4582 152604 -4346
rect 152004 -5524 152604 -4582
rect 155604 697254 156204 709802
rect 173604 711278 174204 711300
rect 173604 711042 173786 711278
rect 174022 711042 174204 711278
rect 173604 710958 174204 711042
rect 173604 710722 173786 710958
rect 174022 710722 174204 710958
rect 170004 709438 170604 709460
rect 170004 709202 170186 709438
rect 170422 709202 170604 709438
rect 170004 709118 170604 709202
rect 170004 708882 170186 709118
rect 170422 708882 170604 709118
rect 166404 707598 167004 707620
rect 166404 707362 166586 707598
rect 166822 707362 167004 707598
rect 166404 707278 167004 707362
rect 166404 707042 166586 707278
rect 166822 707042 167004 707278
rect 155604 697018 155786 697254
rect 156022 697018 156204 697254
rect 155604 696934 156204 697018
rect 155604 696698 155786 696934
rect 156022 696698 156204 696934
rect 155604 661254 156204 696698
rect 155604 661018 155786 661254
rect 156022 661018 156204 661254
rect 155604 660934 156204 661018
rect 155604 660698 155786 660934
rect 156022 660698 156204 660934
rect 155604 625254 156204 660698
rect 155604 625018 155786 625254
rect 156022 625018 156204 625254
rect 155604 624934 156204 625018
rect 155604 624698 155786 624934
rect 156022 624698 156204 624934
rect 155604 589254 156204 624698
rect 155604 589018 155786 589254
rect 156022 589018 156204 589254
rect 155604 588934 156204 589018
rect 155604 588698 155786 588934
rect 156022 588698 156204 588934
rect 155604 553254 156204 588698
rect 155604 553018 155786 553254
rect 156022 553018 156204 553254
rect 155604 552934 156204 553018
rect 155604 552698 155786 552934
rect 156022 552698 156204 552934
rect 155604 517254 156204 552698
rect 155604 517018 155786 517254
rect 156022 517018 156204 517254
rect 155604 516934 156204 517018
rect 155604 516698 155786 516934
rect 156022 516698 156204 516934
rect 155604 481254 156204 516698
rect 155604 481018 155786 481254
rect 156022 481018 156204 481254
rect 155604 480934 156204 481018
rect 155604 480698 155786 480934
rect 156022 480698 156204 480934
rect 155604 445254 156204 480698
rect 155604 445018 155786 445254
rect 156022 445018 156204 445254
rect 155604 444934 156204 445018
rect 155604 444698 155786 444934
rect 156022 444698 156204 444934
rect 155604 409254 156204 444698
rect 155604 409018 155786 409254
rect 156022 409018 156204 409254
rect 155604 408934 156204 409018
rect 155604 408698 155786 408934
rect 156022 408698 156204 408934
rect 155604 373254 156204 408698
rect 155604 373018 155786 373254
rect 156022 373018 156204 373254
rect 155604 372934 156204 373018
rect 155604 372698 155786 372934
rect 156022 372698 156204 372934
rect 155604 337254 156204 372698
rect 155604 337018 155786 337254
rect 156022 337018 156204 337254
rect 155604 336934 156204 337018
rect 155604 336698 155786 336934
rect 156022 336698 156204 336934
rect 155604 301254 156204 336698
rect 155604 301018 155786 301254
rect 156022 301018 156204 301254
rect 155604 300934 156204 301018
rect 155604 300698 155786 300934
rect 156022 300698 156204 300934
rect 155604 265254 156204 300698
rect 155604 265018 155786 265254
rect 156022 265018 156204 265254
rect 155604 264934 156204 265018
rect 155604 264698 155786 264934
rect 156022 264698 156204 264934
rect 155604 229254 156204 264698
rect 155604 229018 155786 229254
rect 156022 229018 156204 229254
rect 155604 228934 156204 229018
rect 155604 228698 155786 228934
rect 156022 228698 156204 228934
rect 155604 193254 156204 228698
rect 155604 193018 155786 193254
rect 156022 193018 156204 193254
rect 155604 192934 156204 193018
rect 155604 192698 155786 192934
rect 156022 192698 156204 192934
rect 155604 157254 156204 192698
rect 155604 157018 155786 157254
rect 156022 157018 156204 157254
rect 155604 156934 156204 157018
rect 155604 156698 155786 156934
rect 156022 156698 156204 156934
rect 155604 121254 156204 156698
rect 155604 121018 155786 121254
rect 156022 121018 156204 121254
rect 155604 120934 156204 121018
rect 155604 120698 155786 120934
rect 156022 120698 156204 120934
rect 155604 85254 156204 120698
rect 155604 85018 155786 85254
rect 156022 85018 156204 85254
rect 155604 84934 156204 85018
rect 155604 84698 155786 84934
rect 156022 84698 156204 84934
rect 155604 49254 156204 84698
rect 155604 49018 155786 49254
rect 156022 49018 156204 49254
rect 155604 48934 156204 49018
rect 155604 48698 155786 48934
rect 156022 48698 156204 48934
rect 155604 13254 156204 48698
rect 155604 13018 155786 13254
rect 156022 13018 156204 13254
rect 155604 12934 156204 13018
rect 155604 12698 155786 12934
rect 156022 12698 156204 12934
rect 137604 -7022 137786 -6786
rect 138022 -7022 138204 -6786
rect 137604 -7106 138204 -7022
rect 137604 -7342 137786 -7106
rect 138022 -7342 138204 -7106
rect 137604 -7364 138204 -7342
rect 155604 -5866 156204 12698
rect 162804 705758 163404 705780
rect 162804 705522 162986 705758
rect 163222 705522 163404 705758
rect 162804 705438 163404 705522
rect 162804 705202 162986 705438
rect 163222 705202 163404 705438
rect 162804 668454 163404 705202
rect 162804 668218 162986 668454
rect 163222 668218 163404 668454
rect 162804 668134 163404 668218
rect 162804 667898 162986 668134
rect 163222 667898 163404 668134
rect 162804 632454 163404 667898
rect 162804 632218 162986 632454
rect 163222 632218 163404 632454
rect 162804 632134 163404 632218
rect 162804 631898 162986 632134
rect 163222 631898 163404 632134
rect 162804 596454 163404 631898
rect 162804 596218 162986 596454
rect 163222 596218 163404 596454
rect 162804 596134 163404 596218
rect 162804 595898 162986 596134
rect 163222 595898 163404 596134
rect 162804 560454 163404 595898
rect 162804 560218 162986 560454
rect 163222 560218 163404 560454
rect 162804 560134 163404 560218
rect 162804 559898 162986 560134
rect 163222 559898 163404 560134
rect 162804 524454 163404 559898
rect 162804 524218 162986 524454
rect 163222 524218 163404 524454
rect 162804 524134 163404 524218
rect 162804 523898 162986 524134
rect 163222 523898 163404 524134
rect 162804 488454 163404 523898
rect 162804 488218 162986 488454
rect 163222 488218 163404 488454
rect 162804 488134 163404 488218
rect 162804 487898 162986 488134
rect 163222 487898 163404 488134
rect 162804 452454 163404 487898
rect 162804 452218 162986 452454
rect 163222 452218 163404 452454
rect 162804 452134 163404 452218
rect 162804 451898 162986 452134
rect 163222 451898 163404 452134
rect 162804 416454 163404 451898
rect 162804 416218 162986 416454
rect 163222 416218 163404 416454
rect 162804 416134 163404 416218
rect 162804 415898 162986 416134
rect 163222 415898 163404 416134
rect 162804 380454 163404 415898
rect 162804 380218 162986 380454
rect 163222 380218 163404 380454
rect 162804 380134 163404 380218
rect 162804 379898 162986 380134
rect 163222 379898 163404 380134
rect 162804 344454 163404 379898
rect 162804 344218 162986 344454
rect 163222 344218 163404 344454
rect 162804 344134 163404 344218
rect 162804 343898 162986 344134
rect 163222 343898 163404 344134
rect 162804 308454 163404 343898
rect 162804 308218 162986 308454
rect 163222 308218 163404 308454
rect 162804 308134 163404 308218
rect 162804 307898 162986 308134
rect 163222 307898 163404 308134
rect 162804 272454 163404 307898
rect 162804 272218 162986 272454
rect 163222 272218 163404 272454
rect 162804 272134 163404 272218
rect 162804 271898 162986 272134
rect 163222 271898 163404 272134
rect 162804 236454 163404 271898
rect 162804 236218 162986 236454
rect 163222 236218 163404 236454
rect 162804 236134 163404 236218
rect 162804 235898 162986 236134
rect 163222 235898 163404 236134
rect 162804 200454 163404 235898
rect 162804 200218 162986 200454
rect 163222 200218 163404 200454
rect 162804 200134 163404 200218
rect 162804 199898 162986 200134
rect 163222 199898 163404 200134
rect 162804 164454 163404 199898
rect 162804 164218 162986 164454
rect 163222 164218 163404 164454
rect 162804 164134 163404 164218
rect 162804 163898 162986 164134
rect 163222 163898 163404 164134
rect 162804 128454 163404 163898
rect 162804 128218 162986 128454
rect 163222 128218 163404 128454
rect 162804 128134 163404 128218
rect 162804 127898 162986 128134
rect 163222 127898 163404 128134
rect 162804 92454 163404 127898
rect 162804 92218 162986 92454
rect 163222 92218 163404 92454
rect 162804 92134 163404 92218
rect 162804 91898 162986 92134
rect 163222 91898 163404 92134
rect 162804 56454 163404 91898
rect 162804 56218 162986 56454
rect 163222 56218 163404 56454
rect 162804 56134 163404 56218
rect 162804 55898 162986 56134
rect 163222 55898 163404 56134
rect 162804 20454 163404 55898
rect 162804 20218 162986 20454
rect 163222 20218 163404 20454
rect 162804 20134 163404 20218
rect 162804 19898 162986 20134
rect 163222 19898 163404 20134
rect 162804 -1266 163404 19898
rect 162804 -1502 162986 -1266
rect 163222 -1502 163404 -1266
rect 162804 -1586 163404 -1502
rect 162804 -1822 162986 -1586
rect 163222 -1822 163404 -1586
rect 162804 -1844 163404 -1822
rect 166404 672054 167004 707042
rect 166404 671818 166586 672054
rect 166822 671818 167004 672054
rect 166404 671734 167004 671818
rect 166404 671498 166586 671734
rect 166822 671498 167004 671734
rect 166404 636054 167004 671498
rect 166404 635818 166586 636054
rect 166822 635818 167004 636054
rect 166404 635734 167004 635818
rect 166404 635498 166586 635734
rect 166822 635498 167004 635734
rect 166404 600054 167004 635498
rect 166404 599818 166586 600054
rect 166822 599818 167004 600054
rect 166404 599734 167004 599818
rect 166404 599498 166586 599734
rect 166822 599498 167004 599734
rect 166404 564054 167004 599498
rect 166404 563818 166586 564054
rect 166822 563818 167004 564054
rect 166404 563734 167004 563818
rect 166404 563498 166586 563734
rect 166822 563498 167004 563734
rect 166404 528054 167004 563498
rect 166404 527818 166586 528054
rect 166822 527818 167004 528054
rect 166404 527734 167004 527818
rect 166404 527498 166586 527734
rect 166822 527498 167004 527734
rect 166404 492054 167004 527498
rect 166404 491818 166586 492054
rect 166822 491818 167004 492054
rect 166404 491734 167004 491818
rect 166404 491498 166586 491734
rect 166822 491498 167004 491734
rect 166404 456054 167004 491498
rect 166404 455818 166586 456054
rect 166822 455818 167004 456054
rect 166404 455734 167004 455818
rect 166404 455498 166586 455734
rect 166822 455498 167004 455734
rect 166404 420054 167004 455498
rect 166404 419818 166586 420054
rect 166822 419818 167004 420054
rect 166404 419734 167004 419818
rect 166404 419498 166586 419734
rect 166822 419498 167004 419734
rect 166404 384054 167004 419498
rect 166404 383818 166586 384054
rect 166822 383818 167004 384054
rect 166404 383734 167004 383818
rect 166404 383498 166586 383734
rect 166822 383498 167004 383734
rect 166404 348054 167004 383498
rect 166404 347818 166586 348054
rect 166822 347818 167004 348054
rect 166404 347734 167004 347818
rect 166404 347498 166586 347734
rect 166822 347498 167004 347734
rect 166404 312054 167004 347498
rect 166404 311818 166586 312054
rect 166822 311818 167004 312054
rect 166404 311734 167004 311818
rect 166404 311498 166586 311734
rect 166822 311498 167004 311734
rect 166404 276054 167004 311498
rect 166404 275818 166586 276054
rect 166822 275818 167004 276054
rect 166404 275734 167004 275818
rect 166404 275498 166586 275734
rect 166822 275498 167004 275734
rect 166404 240054 167004 275498
rect 166404 239818 166586 240054
rect 166822 239818 167004 240054
rect 166404 239734 167004 239818
rect 166404 239498 166586 239734
rect 166822 239498 167004 239734
rect 166404 204054 167004 239498
rect 166404 203818 166586 204054
rect 166822 203818 167004 204054
rect 166404 203734 167004 203818
rect 166404 203498 166586 203734
rect 166822 203498 167004 203734
rect 166404 168054 167004 203498
rect 166404 167818 166586 168054
rect 166822 167818 167004 168054
rect 166404 167734 167004 167818
rect 166404 167498 166586 167734
rect 166822 167498 167004 167734
rect 166404 132054 167004 167498
rect 166404 131818 166586 132054
rect 166822 131818 167004 132054
rect 166404 131734 167004 131818
rect 166404 131498 166586 131734
rect 166822 131498 167004 131734
rect 166404 96054 167004 131498
rect 166404 95818 166586 96054
rect 166822 95818 167004 96054
rect 166404 95734 167004 95818
rect 166404 95498 166586 95734
rect 166822 95498 167004 95734
rect 166404 60054 167004 95498
rect 166404 59818 166586 60054
rect 166822 59818 167004 60054
rect 166404 59734 167004 59818
rect 166404 59498 166586 59734
rect 166822 59498 167004 59734
rect 166404 24054 167004 59498
rect 166404 23818 166586 24054
rect 166822 23818 167004 24054
rect 166404 23734 167004 23818
rect 166404 23498 166586 23734
rect 166822 23498 167004 23734
rect 166404 -3106 167004 23498
rect 166404 -3342 166586 -3106
rect 166822 -3342 167004 -3106
rect 166404 -3426 167004 -3342
rect 166404 -3662 166586 -3426
rect 166822 -3662 167004 -3426
rect 166404 -3684 167004 -3662
rect 170004 675654 170604 708882
rect 170004 675418 170186 675654
rect 170422 675418 170604 675654
rect 170004 675334 170604 675418
rect 170004 675098 170186 675334
rect 170422 675098 170604 675334
rect 170004 639654 170604 675098
rect 170004 639418 170186 639654
rect 170422 639418 170604 639654
rect 170004 639334 170604 639418
rect 170004 639098 170186 639334
rect 170422 639098 170604 639334
rect 170004 603654 170604 639098
rect 170004 603418 170186 603654
rect 170422 603418 170604 603654
rect 170004 603334 170604 603418
rect 170004 603098 170186 603334
rect 170422 603098 170604 603334
rect 170004 567654 170604 603098
rect 170004 567418 170186 567654
rect 170422 567418 170604 567654
rect 170004 567334 170604 567418
rect 170004 567098 170186 567334
rect 170422 567098 170604 567334
rect 170004 531654 170604 567098
rect 170004 531418 170186 531654
rect 170422 531418 170604 531654
rect 170004 531334 170604 531418
rect 170004 531098 170186 531334
rect 170422 531098 170604 531334
rect 170004 495654 170604 531098
rect 170004 495418 170186 495654
rect 170422 495418 170604 495654
rect 170004 495334 170604 495418
rect 170004 495098 170186 495334
rect 170422 495098 170604 495334
rect 170004 459654 170604 495098
rect 170004 459418 170186 459654
rect 170422 459418 170604 459654
rect 170004 459334 170604 459418
rect 170004 459098 170186 459334
rect 170422 459098 170604 459334
rect 170004 423654 170604 459098
rect 170004 423418 170186 423654
rect 170422 423418 170604 423654
rect 170004 423334 170604 423418
rect 170004 423098 170186 423334
rect 170422 423098 170604 423334
rect 170004 387654 170604 423098
rect 170004 387418 170186 387654
rect 170422 387418 170604 387654
rect 170004 387334 170604 387418
rect 170004 387098 170186 387334
rect 170422 387098 170604 387334
rect 170004 351654 170604 387098
rect 170004 351418 170186 351654
rect 170422 351418 170604 351654
rect 170004 351334 170604 351418
rect 170004 351098 170186 351334
rect 170422 351098 170604 351334
rect 170004 315654 170604 351098
rect 170004 315418 170186 315654
rect 170422 315418 170604 315654
rect 170004 315334 170604 315418
rect 170004 315098 170186 315334
rect 170422 315098 170604 315334
rect 170004 279654 170604 315098
rect 170004 279418 170186 279654
rect 170422 279418 170604 279654
rect 170004 279334 170604 279418
rect 170004 279098 170186 279334
rect 170422 279098 170604 279334
rect 170004 243654 170604 279098
rect 170004 243418 170186 243654
rect 170422 243418 170604 243654
rect 170004 243334 170604 243418
rect 170004 243098 170186 243334
rect 170422 243098 170604 243334
rect 170004 207654 170604 243098
rect 170004 207418 170186 207654
rect 170422 207418 170604 207654
rect 170004 207334 170604 207418
rect 170004 207098 170186 207334
rect 170422 207098 170604 207334
rect 170004 171654 170604 207098
rect 170004 171418 170186 171654
rect 170422 171418 170604 171654
rect 170004 171334 170604 171418
rect 170004 171098 170186 171334
rect 170422 171098 170604 171334
rect 170004 135654 170604 171098
rect 170004 135418 170186 135654
rect 170422 135418 170604 135654
rect 170004 135334 170604 135418
rect 170004 135098 170186 135334
rect 170422 135098 170604 135334
rect 170004 99654 170604 135098
rect 170004 99418 170186 99654
rect 170422 99418 170604 99654
rect 170004 99334 170604 99418
rect 170004 99098 170186 99334
rect 170422 99098 170604 99334
rect 170004 63654 170604 99098
rect 170004 63418 170186 63654
rect 170422 63418 170604 63654
rect 170004 63334 170604 63418
rect 170004 63098 170186 63334
rect 170422 63098 170604 63334
rect 170004 27654 170604 63098
rect 170004 27418 170186 27654
rect 170422 27418 170604 27654
rect 170004 27334 170604 27418
rect 170004 27098 170186 27334
rect 170422 27098 170604 27334
rect 170004 -4946 170604 27098
rect 170004 -5182 170186 -4946
rect 170422 -5182 170604 -4946
rect 170004 -5266 170604 -5182
rect 170004 -5502 170186 -5266
rect 170422 -5502 170604 -5266
rect 170004 -5524 170604 -5502
rect 173604 679254 174204 710722
rect 191604 710358 192204 711300
rect 191604 710122 191786 710358
rect 192022 710122 192204 710358
rect 191604 710038 192204 710122
rect 191604 709802 191786 710038
rect 192022 709802 192204 710038
rect 188004 708518 188604 709460
rect 188004 708282 188186 708518
rect 188422 708282 188604 708518
rect 188004 708198 188604 708282
rect 188004 707962 188186 708198
rect 188422 707962 188604 708198
rect 184404 706678 185004 707620
rect 184404 706442 184586 706678
rect 184822 706442 185004 706678
rect 184404 706358 185004 706442
rect 184404 706122 184586 706358
rect 184822 706122 185004 706358
rect 173604 679018 173786 679254
rect 174022 679018 174204 679254
rect 173604 678934 174204 679018
rect 173604 678698 173786 678934
rect 174022 678698 174204 678934
rect 173604 643254 174204 678698
rect 173604 643018 173786 643254
rect 174022 643018 174204 643254
rect 173604 642934 174204 643018
rect 173604 642698 173786 642934
rect 174022 642698 174204 642934
rect 173604 607254 174204 642698
rect 173604 607018 173786 607254
rect 174022 607018 174204 607254
rect 173604 606934 174204 607018
rect 173604 606698 173786 606934
rect 174022 606698 174204 606934
rect 173604 571254 174204 606698
rect 173604 571018 173786 571254
rect 174022 571018 174204 571254
rect 173604 570934 174204 571018
rect 173604 570698 173786 570934
rect 174022 570698 174204 570934
rect 173604 535254 174204 570698
rect 173604 535018 173786 535254
rect 174022 535018 174204 535254
rect 173604 534934 174204 535018
rect 173604 534698 173786 534934
rect 174022 534698 174204 534934
rect 173604 499254 174204 534698
rect 173604 499018 173786 499254
rect 174022 499018 174204 499254
rect 173604 498934 174204 499018
rect 173604 498698 173786 498934
rect 174022 498698 174204 498934
rect 173604 463254 174204 498698
rect 173604 463018 173786 463254
rect 174022 463018 174204 463254
rect 173604 462934 174204 463018
rect 173604 462698 173786 462934
rect 174022 462698 174204 462934
rect 173604 427254 174204 462698
rect 173604 427018 173786 427254
rect 174022 427018 174204 427254
rect 173604 426934 174204 427018
rect 173604 426698 173786 426934
rect 174022 426698 174204 426934
rect 173604 391254 174204 426698
rect 173604 391018 173786 391254
rect 174022 391018 174204 391254
rect 173604 390934 174204 391018
rect 173604 390698 173786 390934
rect 174022 390698 174204 390934
rect 173604 355254 174204 390698
rect 173604 355018 173786 355254
rect 174022 355018 174204 355254
rect 173604 354934 174204 355018
rect 173604 354698 173786 354934
rect 174022 354698 174204 354934
rect 173604 319254 174204 354698
rect 173604 319018 173786 319254
rect 174022 319018 174204 319254
rect 173604 318934 174204 319018
rect 173604 318698 173786 318934
rect 174022 318698 174204 318934
rect 173604 283254 174204 318698
rect 173604 283018 173786 283254
rect 174022 283018 174204 283254
rect 173604 282934 174204 283018
rect 173604 282698 173786 282934
rect 174022 282698 174204 282934
rect 173604 247254 174204 282698
rect 173604 247018 173786 247254
rect 174022 247018 174204 247254
rect 173604 246934 174204 247018
rect 173604 246698 173786 246934
rect 174022 246698 174204 246934
rect 173604 211254 174204 246698
rect 173604 211018 173786 211254
rect 174022 211018 174204 211254
rect 173604 210934 174204 211018
rect 173604 210698 173786 210934
rect 174022 210698 174204 210934
rect 173604 175254 174204 210698
rect 173604 175018 173786 175254
rect 174022 175018 174204 175254
rect 173604 174934 174204 175018
rect 173604 174698 173786 174934
rect 174022 174698 174204 174934
rect 173604 139254 174204 174698
rect 173604 139018 173786 139254
rect 174022 139018 174204 139254
rect 173604 138934 174204 139018
rect 173604 138698 173786 138934
rect 174022 138698 174204 138934
rect 173604 103254 174204 138698
rect 173604 103018 173786 103254
rect 174022 103018 174204 103254
rect 173604 102934 174204 103018
rect 173604 102698 173786 102934
rect 174022 102698 174204 102934
rect 173604 67254 174204 102698
rect 173604 67018 173786 67254
rect 174022 67018 174204 67254
rect 173604 66934 174204 67018
rect 173604 66698 173786 66934
rect 174022 66698 174204 66934
rect 173604 31254 174204 66698
rect 173604 31018 173786 31254
rect 174022 31018 174204 31254
rect 173604 30934 174204 31018
rect 173604 30698 173786 30934
rect 174022 30698 174204 30934
rect 155604 -6102 155786 -5866
rect 156022 -6102 156204 -5866
rect 155604 -6186 156204 -6102
rect 155604 -6422 155786 -6186
rect 156022 -6422 156204 -6186
rect 155604 -7364 156204 -6422
rect 173604 -6786 174204 30698
rect 180804 704838 181404 705780
rect 180804 704602 180986 704838
rect 181222 704602 181404 704838
rect 180804 704518 181404 704602
rect 180804 704282 180986 704518
rect 181222 704282 181404 704518
rect 180804 686454 181404 704282
rect 180804 686218 180986 686454
rect 181222 686218 181404 686454
rect 180804 686134 181404 686218
rect 180804 685898 180986 686134
rect 181222 685898 181404 686134
rect 180804 650454 181404 685898
rect 180804 650218 180986 650454
rect 181222 650218 181404 650454
rect 180804 650134 181404 650218
rect 180804 649898 180986 650134
rect 181222 649898 181404 650134
rect 180804 614454 181404 649898
rect 180804 614218 180986 614454
rect 181222 614218 181404 614454
rect 180804 614134 181404 614218
rect 180804 613898 180986 614134
rect 181222 613898 181404 614134
rect 180804 578454 181404 613898
rect 180804 578218 180986 578454
rect 181222 578218 181404 578454
rect 180804 578134 181404 578218
rect 180804 577898 180986 578134
rect 181222 577898 181404 578134
rect 180804 542454 181404 577898
rect 180804 542218 180986 542454
rect 181222 542218 181404 542454
rect 180804 542134 181404 542218
rect 180804 541898 180986 542134
rect 181222 541898 181404 542134
rect 180804 506454 181404 541898
rect 180804 506218 180986 506454
rect 181222 506218 181404 506454
rect 180804 506134 181404 506218
rect 180804 505898 180986 506134
rect 181222 505898 181404 506134
rect 180804 470454 181404 505898
rect 180804 470218 180986 470454
rect 181222 470218 181404 470454
rect 180804 470134 181404 470218
rect 180804 469898 180986 470134
rect 181222 469898 181404 470134
rect 180804 434454 181404 469898
rect 180804 434218 180986 434454
rect 181222 434218 181404 434454
rect 180804 434134 181404 434218
rect 180804 433898 180986 434134
rect 181222 433898 181404 434134
rect 180804 398454 181404 433898
rect 180804 398218 180986 398454
rect 181222 398218 181404 398454
rect 180804 398134 181404 398218
rect 180804 397898 180986 398134
rect 181222 397898 181404 398134
rect 180804 362454 181404 397898
rect 180804 362218 180986 362454
rect 181222 362218 181404 362454
rect 180804 362134 181404 362218
rect 180804 361898 180986 362134
rect 181222 361898 181404 362134
rect 180804 326454 181404 361898
rect 180804 326218 180986 326454
rect 181222 326218 181404 326454
rect 180804 326134 181404 326218
rect 180804 325898 180986 326134
rect 181222 325898 181404 326134
rect 180804 290454 181404 325898
rect 180804 290218 180986 290454
rect 181222 290218 181404 290454
rect 180804 290134 181404 290218
rect 180804 289898 180986 290134
rect 181222 289898 181404 290134
rect 180804 254454 181404 289898
rect 180804 254218 180986 254454
rect 181222 254218 181404 254454
rect 180804 254134 181404 254218
rect 180804 253898 180986 254134
rect 181222 253898 181404 254134
rect 180804 218454 181404 253898
rect 180804 218218 180986 218454
rect 181222 218218 181404 218454
rect 180804 218134 181404 218218
rect 180804 217898 180986 218134
rect 181222 217898 181404 218134
rect 180804 182454 181404 217898
rect 180804 182218 180986 182454
rect 181222 182218 181404 182454
rect 180804 182134 181404 182218
rect 180804 181898 180986 182134
rect 181222 181898 181404 182134
rect 180804 146454 181404 181898
rect 180804 146218 180986 146454
rect 181222 146218 181404 146454
rect 180804 146134 181404 146218
rect 180804 145898 180986 146134
rect 181222 145898 181404 146134
rect 180804 110454 181404 145898
rect 180804 110218 180986 110454
rect 181222 110218 181404 110454
rect 180804 110134 181404 110218
rect 180804 109898 180986 110134
rect 181222 109898 181404 110134
rect 180804 74454 181404 109898
rect 180804 74218 180986 74454
rect 181222 74218 181404 74454
rect 180804 74134 181404 74218
rect 180804 73898 180986 74134
rect 181222 73898 181404 74134
rect 180804 38454 181404 73898
rect 180804 38218 180986 38454
rect 181222 38218 181404 38454
rect 180804 38134 181404 38218
rect 180804 37898 180986 38134
rect 181222 37898 181404 38134
rect 180804 2454 181404 37898
rect 180804 2218 180986 2454
rect 181222 2218 181404 2454
rect 180804 2134 181404 2218
rect 180804 1898 180986 2134
rect 181222 1898 181404 2134
rect 180804 -346 181404 1898
rect 180804 -582 180986 -346
rect 181222 -582 181404 -346
rect 180804 -666 181404 -582
rect 180804 -902 180986 -666
rect 181222 -902 181404 -666
rect 180804 -1844 181404 -902
rect 184404 690054 185004 706122
rect 184404 689818 184586 690054
rect 184822 689818 185004 690054
rect 184404 689734 185004 689818
rect 184404 689498 184586 689734
rect 184822 689498 185004 689734
rect 184404 654054 185004 689498
rect 184404 653818 184586 654054
rect 184822 653818 185004 654054
rect 184404 653734 185004 653818
rect 184404 653498 184586 653734
rect 184822 653498 185004 653734
rect 184404 618054 185004 653498
rect 184404 617818 184586 618054
rect 184822 617818 185004 618054
rect 184404 617734 185004 617818
rect 184404 617498 184586 617734
rect 184822 617498 185004 617734
rect 184404 582054 185004 617498
rect 184404 581818 184586 582054
rect 184822 581818 185004 582054
rect 184404 581734 185004 581818
rect 184404 581498 184586 581734
rect 184822 581498 185004 581734
rect 184404 546054 185004 581498
rect 184404 545818 184586 546054
rect 184822 545818 185004 546054
rect 184404 545734 185004 545818
rect 184404 545498 184586 545734
rect 184822 545498 185004 545734
rect 184404 510054 185004 545498
rect 184404 509818 184586 510054
rect 184822 509818 185004 510054
rect 184404 509734 185004 509818
rect 184404 509498 184586 509734
rect 184822 509498 185004 509734
rect 184404 474054 185004 509498
rect 184404 473818 184586 474054
rect 184822 473818 185004 474054
rect 184404 473734 185004 473818
rect 184404 473498 184586 473734
rect 184822 473498 185004 473734
rect 184404 438054 185004 473498
rect 184404 437818 184586 438054
rect 184822 437818 185004 438054
rect 184404 437734 185004 437818
rect 184404 437498 184586 437734
rect 184822 437498 185004 437734
rect 184404 402054 185004 437498
rect 184404 401818 184586 402054
rect 184822 401818 185004 402054
rect 184404 401734 185004 401818
rect 184404 401498 184586 401734
rect 184822 401498 185004 401734
rect 184404 366054 185004 401498
rect 184404 365818 184586 366054
rect 184822 365818 185004 366054
rect 184404 365734 185004 365818
rect 184404 365498 184586 365734
rect 184822 365498 185004 365734
rect 184404 330054 185004 365498
rect 184404 329818 184586 330054
rect 184822 329818 185004 330054
rect 184404 329734 185004 329818
rect 184404 329498 184586 329734
rect 184822 329498 185004 329734
rect 184404 294054 185004 329498
rect 184404 293818 184586 294054
rect 184822 293818 185004 294054
rect 184404 293734 185004 293818
rect 184404 293498 184586 293734
rect 184822 293498 185004 293734
rect 184404 258054 185004 293498
rect 184404 257818 184586 258054
rect 184822 257818 185004 258054
rect 184404 257734 185004 257818
rect 184404 257498 184586 257734
rect 184822 257498 185004 257734
rect 184404 222054 185004 257498
rect 184404 221818 184586 222054
rect 184822 221818 185004 222054
rect 184404 221734 185004 221818
rect 184404 221498 184586 221734
rect 184822 221498 185004 221734
rect 184404 186054 185004 221498
rect 184404 185818 184586 186054
rect 184822 185818 185004 186054
rect 184404 185734 185004 185818
rect 184404 185498 184586 185734
rect 184822 185498 185004 185734
rect 184404 150054 185004 185498
rect 184404 149818 184586 150054
rect 184822 149818 185004 150054
rect 184404 149734 185004 149818
rect 184404 149498 184586 149734
rect 184822 149498 185004 149734
rect 184404 114054 185004 149498
rect 184404 113818 184586 114054
rect 184822 113818 185004 114054
rect 184404 113734 185004 113818
rect 184404 113498 184586 113734
rect 184822 113498 185004 113734
rect 184404 78054 185004 113498
rect 184404 77818 184586 78054
rect 184822 77818 185004 78054
rect 184404 77734 185004 77818
rect 184404 77498 184586 77734
rect 184822 77498 185004 77734
rect 184404 42054 185004 77498
rect 184404 41818 184586 42054
rect 184822 41818 185004 42054
rect 184404 41734 185004 41818
rect 184404 41498 184586 41734
rect 184822 41498 185004 41734
rect 184404 6054 185004 41498
rect 184404 5818 184586 6054
rect 184822 5818 185004 6054
rect 184404 5734 185004 5818
rect 184404 5498 184586 5734
rect 184822 5498 185004 5734
rect 184404 -2186 185004 5498
rect 184404 -2422 184586 -2186
rect 184822 -2422 185004 -2186
rect 184404 -2506 185004 -2422
rect 184404 -2742 184586 -2506
rect 184822 -2742 185004 -2506
rect 184404 -3684 185004 -2742
rect 188004 693654 188604 707962
rect 188004 693418 188186 693654
rect 188422 693418 188604 693654
rect 188004 693334 188604 693418
rect 188004 693098 188186 693334
rect 188422 693098 188604 693334
rect 188004 657654 188604 693098
rect 188004 657418 188186 657654
rect 188422 657418 188604 657654
rect 188004 657334 188604 657418
rect 188004 657098 188186 657334
rect 188422 657098 188604 657334
rect 188004 621654 188604 657098
rect 188004 621418 188186 621654
rect 188422 621418 188604 621654
rect 188004 621334 188604 621418
rect 188004 621098 188186 621334
rect 188422 621098 188604 621334
rect 188004 585654 188604 621098
rect 188004 585418 188186 585654
rect 188422 585418 188604 585654
rect 188004 585334 188604 585418
rect 188004 585098 188186 585334
rect 188422 585098 188604 585334
rect 188004 549654 188604 585098
rect 188004 549418 188186 549654
rect 188422 549418 188604 549654
rect 188004 549334 188604 549418
rect 188004 549098 188186 549334
rect 188422 549098 188604 549334
rect 188004 513654 188604 549098
rect 188004 513418 188186 513654
rect 188422 513418 188604 513654
rect 188004 513334 188604 513418
rect 188004 513098 188186 513334
rect 188422 513098 188604 513334
rect 188004 477654 188604 513098
rect 188004 477418 188186 477654
rect 188422 477418 188604 477654
rect 188004 477334 188604 477418
rect 188004 477098 188186 477334
rect 188422 477098 188604 477334
rect 188004 441654 188604 477098
rect 188004 441418 188186 441654
rect 188422 441418 188604 441654
rect 188004 441334 188604 441418
rect 188004 441098 188186 441334
rect 188422 441098 188604 441334
rect 188004 405654 188604 441098
rect 188004 405418 188186 405654
rect 188422 405418 188604 405654
rect 188004 405334 188604 405418
rect 188004 405098 188186 405334
rect 188422 405098 188604 405334
rect 188004 369654 188604 405098
rect 188004 369418 188186 369654
rect 188422 369418 188604 369654
rect 188004 369334 188604 369418
rect 188004 369098 188186 369334
rect 188422 369098 188604 369334
rect 188004 333654 188604 369098
rect 188004 333418 188186 333654
rect 188422 333418 188604 333654
rect 188004 333334 188604 333418
rect 188004 333098 188186 333334
rect 188422 333098 188604 333334
rect 188004 297654 188604 333098
rect 188004 297418 188186 297654
rect 188422 297418 188604 297654
rect 188004 297334 188604 297418
rect 188004 297098 188186 297334
rect 188422 297098 188604 297334
rect 188004 261654 188604 297098
rect 188004 261418 188186 261654
rect 188422 261418 188604 261654
rect 188004 261334 188604 261418
rect 188004 261098 188186 261334
rect 188422 261098 188604 261334
rect 188004 225654 188604 261098
rect 188004 225418 188186 225654
rect 188422 225418 188604 225654
rect 188004 225334 188604 225418
rect 188004 225098 188186 225334
rect 188422 225098 188604 225334
rect 188004 189654 188604 225098
rect 188004 189418 188186 189654
rect 188422 189418 188604 189654
rect 188004 189334 188604 189418
rect 188004 189098 188186 189334
rect 188422 189098 188604 189334
rect 188004 153654 188604 189098
rect 188004 153418 188186 153654
rect 188422 153418 188604 153654
rect 188004 153334 188604 153418
rect 188004 153098 188186 153334
rect 188422 153098 188604 153334
rect 188004 117654 188604 153098
rect 188004 117418 188186 117654
rect 188422 117418 188604 117654
rect 188004 117334 188604 117418
rect 188004 117098 188186 117334
rect 188422 117098 188604 117334
rect 188004 81654 188604 117098
rect 188004 81418 188186 81654
rect 188422 81418 188604 81654
rect 188004 81334 188604 81418
rect 188004 81098 188186 81334
rect 188422 81098 188604 81334
rect 188004 45654 188604 81098
rect 188004 45418 188186 45654
rect 188422 45418 188604 45654
rect 188004 45334 188604 45418
rect 188004 45098 188186 45334
rect 188422 45098 188604 45334
rect 188004 9654 188604 45098
rect 188004 9418 188186 9654
rect 188422 9418 188604 9654
rect 188004 9334 188604 9418
rect 188004 9098 188186 9334
rect 188422 9098 188604 9334
rect 188004 -4026 188604 9098
rect 188004 -4262 188186 -4026
rect 188422 -4262 188604 -4026
rect 188004 -4346 188604 -4262
rect 188004 -4582 188186 -4346
rect 188422 -4582 188604 -4346
rect 188004 -5524 188604 -4582
rect 191604 697254 192204 709802
rect 209604 711278 210204 711300
rect 209604 711042 209786 711278
rect 210022 711042 210204 711278
rect 209604 710958 210204 711042
rect 209604 710722 209786 710958
rect 210022 710722 210204 710958
rect 206004 709438 206604 709460
rect 206004 709202 206186 709438
rect 206422 709202 206604 709438
rect 206004 709118 206604 709202
rect 206004 708882 206186 709118
rect 206422 708882 206604 709118
rect 202404 707598 203004 707620
rect 202404 707362 202586 707598
rect 202822 707362 203004 707598
rect 202404 707278 203004 707362
rect 202404 707042 202586 707278
rect 202822 707042 203004 707278
rect 191604 697018 191786 697254
rect 192022 697018 192204 697254
rect 191604 696934 192204 697018
rect 191604 696698 191786 696934
rect 192022 696698 192204 696934
rect 191604 661254 192204 696698
rect 191604 661018 191786 661254
rect 192022 661018 192204 661254
rect 191604 660934 192204 661018
rect 191604 660698 191786 660934
rect 192022 660698 192204 660934
rect 191604 625254 192204 660698
rect 191604 625018 191786 625254
rect 192022 625018 192204 625254
rect 191604 624934 192204 625018
rect 191604 624698 191786 624934
rect 192022 624698 192204 624934
rect 191604 589254 192204 624698
rect 191604 589018 191786 589254
rect 192022 589018 192204 589254
rect 191604 588934 192204 589018
rect 191604 588698 191786 588934
rect 192022 588698 192204 588934
rect 191604 553254 192204 588698
rect 191604 553018 191786 553254
rect 192022 553018 192204 553254
rect 191604 552934 192204 553018
rect 191604 552698 191786 552934
rect 192022 552698 192204 552934
rect 191604 517254 192204 552698
rect 191604 517018 191786 517254
rect 192022 517018 192204 517254
rect 191604 516934 192204 517018
rect 191604 516698 191786 516934
rect 192022 516698 192204 516934
rect 191604 481254 192204 516698
rect 191604 481018 191786 481254
rect 192022 481018 192204 481254
rect 191604 480934 192204 481018
rect 191604 480698 191786 480934
rect 192022 480698 192204 480934
rect 191604 445254 192204 480698
rect 191604 445018 191786 445254
rect 192022 445018 192204 445254
rect 191604 444934 192204 445018
rect 191604 444698 191786 444934
rect 192022 444698 192204 444934
rect 191604 409254 192204 444698
rect 191604 409018 191786 409254
rect 192022 409018 192204 409254
rect 191604 408934 192204 409018
rect 191604 408698 191786 408934
rect 192022 408698 192204 408934
rect 191604 373254 192204 408698
rect 191604 373018 191786 373254
rect 192022 373018 192204 373254
rect 191604 372934 192204 373018
rect 191604 372698 191786 372934
rect 192022 372698 192204 372934
rect 191604 337254 192204 372698
rect 191604 337018 191786 337254
rect 192022 337018 192204 337254
rect 191604 336934 192204 337018
rect 191604 336698 191786 336934
rect 192022 336698 192204 336934
rect 191604 301254 192204 336698
rect 191604 301018 191786 301254
rect 192022 301018 192204 301254
rect 191604 300934 192204 301018
rect 191604 300698 191786 300934
rect 192022 300698 192204 300934
rect 191604 265254 192204 300698
rect 191604 265018 191786 265254
rect 192022 265018 192204 265254
rect 191604 264934 192204 265018
rect 191604 264698 191786 264934
rect 192022 264698 192204 264934
rect 191604 229254 192204 264698
rect 191604 229018 191786 229254
rect 192022 229018 192204 229254
rect 191604 228934 192204 229018
rect 191604 228698 191786 228934
rect 192022 228698 192204 228934
rect 191604 193254 192204 228698
rect 191604 193018 191786 193254
rect 192022 193018 192204 193254
rect 191604 192934 192204 193018
rect 191604 192698 191786 192934
rect 192022 192698 192204 192934
rect 191604 157254 192204 192698
rect 191604 157018 191786 157254
rect 192022 157018 192204 157254
rect 191604 156934 192204 157018
rect 191604 156698 191786 156934
rect 192022 156698 192204 156934
rect 191604 121254 192204 156698
rect 191604 121018 191786 121254
rect 192022 121018 192204 121254
rect 191604 120934 192204 121018
rect 191604 120698 191786 120934
rect 192022 120698 192204 120934
rect 191604 85254 192204 120698
rect 191604 85018 191786 85254
rect 192022 85018 192204 85254
rect 191604 84934 192204 85018
rect 191604 84698 191786 84934
rect 192022 84698 192204 84934
rect 191604 49254 192204 84698
rect 191604 49018 191786 49254
rect 192022 49018 192204 49254
rect 191604 48934 192204 49018
rect 191604 48698 191786 48934
rect 192022 48698 192204 48934
rect 191604 13254 192204 48698
rect 191604 13018 191786 13254
rect 192022 13018 192204 13254
rect 191604 12934 192204 13018
rect 191604 12698 191786 12934
rect 192022 12698 192204 12934
rect 173604 -7022 173786 -6786
rect 174022 -7022 174204 -6786
rect 173604 -7106 174204 -7022
rect 173604 -7342 173786 -7106
rect 174022 -7342 174204 -7106
rect 173604 -7364 174204 -7342
rect 191604 -5866 192204 12698
rect 198804 705758 199404 705780
rect 198804 705522 198986 705758
rect 199222 705522 199404 705758
rect 198804 705438 199404 705522
rect 198804 705202 198986 705438
rect 199222 705202 199404 705438
rect 198804 668454 199404 705202
rect 198804 668218 198986 668454
rect 199222 668218 199404 668454
rect 198804 668134 199404 668218
rect 198804 667898 198986 668134
rect 199222 667898 199404 668134
rect 198804 632454 199404 667898
rect 198804 632218 198986 632454
rect 199222 632218 199404 632454
rect 198804 632134 199404 632218
rect 198804 631898 198986 632134
rect 199222 631898 199404 632134
rect 198804 596454 199404 631898
rect 198804 596218 198986 596454
rect 199222 596218 199404 596454
rect 198804 596134 199404 596218
rect 198804 595898 198986 596134
rect 199222 595898 199404 596134
rect 198804 560454 199404 595898
rect 198804 560218 198986 560454
rect 199222 560218 199404 560454
rect 198804 560134 199404 560218
rect 198804 559898 198986 560134
rect 199222 559898 199404 560134
rect 198804 524454 199404 559898
rect 198804 524218 198986 524454
rect 199222 524218 199404 524454
rect 198804 524134 199404 524218
rect 198804 523898 198986 524134
rect 199222 523898 199404 524134
rect 198804 488454 199404 523898
rect 198804 488218 198986 488454
rect 199222 488218 199404 488454
rect 198804 488134 199404 488218
rect 198804 487898 198986 488134
rect 199222 487898 199404 488134
rect 198804 452454 199404 487898
rect 198804 452218 198986 452454
rect 199222 452218 199404 452454
rect 198804 452134 199404 452218
rect 198804 451898 198986 452134
rect 199222 451898 199404 452134
rect 198804 416454 199404 451898
rect 198804 416218 198986 416454
rect 199222 416218 199404 416454
rect 198804 416134 199404 416218
rect 198804 415898 198986 416134
rect 199222 415898 199404 416134
rect 198804 380454 199404 415898
rect 198804 380218 198986 380454
rect 199222 380218 199404 380454
rect 198804 380134 199404 380218
rect 198804 379898 198986 380134
rect 199222 379898 199404 380134
rect 198804 344454 199404 379898
rect 198804 344218 198986 344454
rect 199222 344218 199404 344454
rect 198804 344134 199404 344218
rect 198804 343898 198986 344134
rect 199222 343898 199404 344134
rect 198804 308454 199404 343898
rect 198804 308218 198986 308454
rect 199222 308218 199404 308454
rect 198804 308134 199404 308218
rect 198804 307898 198986 308134
rect 199222 307898 199404 308134
rect 198804 272454 199404 307898
rect 198804 272218 198986 272454
rect 199222 272218 199404 272454
rect 198804 272134 199404 272218
rect 198804 271898 198986 272134
rect 199222 271898 199404 272134
rect 198804 236454 199404 271898
rect 198804 236218 198986 236454
rect 199222 236218 199404 236454
rect 198804 236134 199404 236218
rect 198804 235898 198986 236134
rect 199222 235898 199404 236134
rect 198804 200454 199404 235898
rect 198804 200218 198986 200454
rect 199222 200218 199404 200454
rect 198804 200134 199404 200218
rect 198804 199898 198986 200134
rect 199222 199898 199404 200134
rect 198804 164454 199404 199898
rect 198804 164218 198986 164454
rect 199222 164218 199404 164454
rect 198804 164134 199404 164218
rect 198804 163898 198986 164134
rect 199222 163898 199404 164134
rect 198804 128454 199404 163898
rect 198804 128218 198986 128454
rect 199222 128218 199404 128454
rect 198804 128134 199404 128218
rect 198804 127898 198986 128134
rect 199222 127898 199404 128134
rect 198804 92454 199404 127898
rect 198804 92218 198986 92454
rect 199222 92218 199404 92454
rect 198804 92134 199404 92218
rect 198804 91898 198986 92134
rect 199222 91898 199404 92134
rect 198804 56454 199404 91898
rect 198804 56218 198986 56454
rect 199222 56218 199404 56454
rect 198804 56134 199404 56218
rect 198804 55898 198986 56134
rect 199222 55898 199404 56134
rect 198804 20454 199404 55898
rect 198804 20218 198986 20454
rect 199222 20218 199404 20454
rect 198804 20134 199404 20218
rect 198804 19898 198986 20134
rect 199222 19898 199404 20134
rect 198804 -1266 199404 19898
rect 198804 -1502 198986 -1266
rect 199222 -1502 199404 -1266
rect 198804 -1586 199404 -1502
rect 198804 -1822 198986 -1586
rect 199222 -1822 199404 -1586
rect 198804 -1844 199404 -1822
rect 202404 672054 203004 707042
rect 202404 671818 202586 672054
rect 202822 671818 203004 672054
rect 202404 671734 203004 671818
rect 202404 671498 202586 671734
rect 202822 671498 203004 671734
rect 202404 636054 203004 671498
rect 202404 635818 202586 636054
rect 202822 635818 203004 636054
rect 202404 635734 203004 635818
rect 202404 635498 202586 635734
rect 202822 635498 203004 635734
rect 202404 600054 203004 635498
rect 202404 599818 202586 600054
rect 202822 599818 203004 600054
rect 202404 599734 203004 599818
rect 202404 599498 202586 599734
rect 202822 599498 203004 599734
rect 202404 564054 203004 599498
rect 202404 563818 202586 564054
rect 202822 563818 203004 564054
rect 202404 563734 203004 563818
rect 202404 563498 202586 563734
rect 202822 563498 203004 563734
rect 202404 528054 203004 563498
rect 202404 527818 202586 528054
rect 202822 527818 203004 528054
rect 202404 527734 203004 527818
rect 202404 527498 202586 527734
rect 202822 527498 203004 527734
rect 202404 492054 203004 527498
rect 202404 491818 202586 492054
rect 202822 491818 203004 492054
rect 202404 491734 203004 491818
rect 202404 491498 202586 491734
rect 202822 491498 203004 491734
rect 202404 456054 203004 491498
rect 202404 455818 202586 456054
rect 202822 455818 203004 456054
rect 202404 455734 203004 455818
rect 202404 455498 202586 455734
rect 202822 455498 203004 455734
rect 202404 420054 203004 455498
rect 202404 419818 202586 420054
rect 202822 419818 203004 420054
rect 202404 419734 203004 419818
rect 202404 419498 202586 419734
rect 202822 419498 203004 419734
rect 202404 384054 203004 419498
rect 202404 383818 202586 384054
rect 202822 383818 203004 384054
rect 202404 383734 203004 383818
rect 202404 383498 202586 383734
rect 202822 383498 203004 383734
rect 202404 348054 203004 383498
rect 202404 347818 202586 348054
rect 202822 347818 203004 348054
rect 202404 347734 203004 347818
rect 202404 347498 202586 347734
rect 202822 347498 203004 347734
rect 202404 312054 203004 347498
rect 202404 311818 202586 312054
rect 202822 311818 203004 312054
rect 202404 311734 203004 311818
rect 202404 311498 202586 311734
rect 202822 311498 203004 311734
rect 202404 276054 203004 311498
rect 202404 275818 202586 276054
rect 202822 275818 203004 276054
rect 202404 275734 203004 275818
rect 202404 275498 202586 275734
rect 202822 275498 203004 275734
rect 202404 240054 203004 275498
rect 202404 239818 202586 240054
rect 202822 239818 203004 240054
rect 202404 239734 203004 239818
rect 202404 239498 202586 239734
rect 202822 239498 203004 239734
rect 202404 204054 203004 239498
rect 202404 203818 202586 204054
rect 202822 203818 203004 204054
rect 202404 203734 203004 203818
rect 202404 203498 202586 203734
rect 202822 203498 203004 203734
rect 202404 168054 203004 203498
rect 202404 167818 202586 168054
rect 202822 167818 203004 168054
rect 202404 167734 203004 167818
rect 202404 167498 202586 167734
rect 202822 167498 203004 167734
rect 202404 132054 203004 167498
rect 202404 131818 202586 132054
rect 202822 131818 203004 132054
rect 202404 131734 203004 131818
rect 202404 131498 202586 131734
rect 202822 131498 203004 131734
rect 202404 96054 203004 131498
rect 202404 95818 202586 96054
rect 202822 95818 203004 96054
rect 202404 95734 203004 95818
rect 202404 95498 202586 95734
rect 202822 95498 203004 95734
rect 202404 60054 203004 95498
rect 202404 59818 202586 60054
rect 202822 59818 203004 60054
rect 202404 59734 203004 59818
rect 202404 59498 202586 59734
rect 202822 59498 203004 59734
rect 202404 24054 203004 59498
rect 202404 23818 202586 24054
rect 202822 23818 203004 24054
rect 202404 23734 203004 23818
rect 202404 23498 202586 23734
rect 202822 23498 203004 23734
rect 202404 -3106 203004 23498
rect 202404 -3342 202586 -3106
rect 202822 -3342 203004 -3106
rect 202404 -3426 203004 -3342
rect 202404 -3662 202586 -3426
rect 202822 -3662 203004 -3426
rect 202404 -3684 203004 -3662
rect 206004 675654 206604 708882
rect 206004 675418 206186 675654
rect 206422 675418 206604 675654
rect 206004 675334 206604 675418
rect 206004 675098 206186 675334
rect 206422 675098 206604 675334
rect 206004 639654 206604 675098
rect 206004 639418 206186 639654
rect 206422 639418 206604 639654
rect 206004 639334 206604 639418
rect 206004 639098 206186 639334
rect 206422 639098 206604 639334
rect 206004 603654 206604 639098
rect 206004 603418 206186 603654
rect 206422 603418 206604 603654
rect 206004 603334 206604 603418
rect 206004 603098 206186 603334
rect 206422 603098 206604 603334
rect 206004 567654 206604 603098
rect 206004 567418 206186 567654
rect 206422 567418 206604 567654
rect 206004 567334 206604 567418
rect 206004 567098 206186 567334
rect 206422 567098 206604 567334
rect 206004 531654 206604 567098
rect 206004 531418 206186 531654
rect 206422 531418 206604 531654
rect 206004 531334 206604 531418
rect 206004 531098 206186 531334
rect 206422 531098 206604 531334
rect 206004 495654 206604 531098
rect 206004 495418 206186 495654
rect 206422 495418 206604 495654
rect 206004 495334 206604 495418
rect 206004 495098 206186 495334
rect 206422 495098 206604 495334
rect 206004 459654 206604 495098
rect 206004 459418 206186 459654
rect 206422 459418 206604 459654
rect 206004 459334 206604 459418
rect 206004 459098 206186 459334
rect 206422 459098 206604 459334
rect 206004 423654 206604 459098
rect 206004 423418 206186 423654
rect 206422 423418 206604 423654
rect 206004 423334 206604 423418
rect 206004 423098 206186 423334
rect 206422 423098 206604 423334
rect 206004 387654 206604 423098
rect 206004 387418 206186 387654
rect 206422 387418 206604 387654
rect 206004 387334 206604 387418
rect 206004 387098 206186 387334
rect 206422 387098 206604 387334
rect 206004 351654 206604 387098
rect 206004 351418 206186 351654
rect 206422 351418 206604 351654
rect 206004 351334 206604 351418
rect 206004 351098 206186 351334
rect 206422 351098 206604 351334
rect 206004 315654 206604 351098
rect 206004 315418 206186 315654
rect 206422 315418 206604 315654
rect 206004 315334 206604 315418
rect 206004 315098 206186 315334
rect 206422 315098 206604 315334
rect 206004 279654 206604 315098
rect 206004 279418 206186 279654
rect 206422 279418 206604 279654
rect 206004 279334 206604 279418
rect 206004 279098 206186 279334
rect 206422 279098 206604 279334
rect 206004 243654 206604 279098
rect 206004 243418 206186 243654
rect 206422 243418 206604 243654
rect 206004 243334 206604 243418
rect 206004 243098 206186 243334
rect 206422 243098 206604 243334
rect 206004 207654 206604 243098
rect 206004 207418 206186 207654
rect 206422 207418 206604 207654
rect 206004 207334 206604 207418
rect 206004 207098 206186 207334
rect 206422 207098 206604 207334
rect 206004 171654 206604 207098
rect 206004 171418 206186 171654
rect 206422 171418 206604 171654
rect 206004 171334 206604 171418
rect 206004 171098 206186 171334
rect 206422 171098 206604 171334
rect 206004 135654 206604 171098
rect 206004 135418 206186 135654
rect 206422 135418 206604 135654
rect 206004 135334 206604 135418
rect 206004 135098 206186 135334
rect 206422 135098 206604 135334
rect 206004 99654 206604 135098
rect 206004 99418 206186 99654
rect 206422 99418 206604 99654
rect 206004 99334 206604 99418
rect 206004 99098 206186 99334
rect 206422 99098 206604 99334
rect 206004 63654 206604 99098
rect 206004 63418 206186 63654
rect 206422 63418 206604 63654
rect 206004 63334 206604 63418
rect 206004 63098 206186 63334
rect 206422 63098 206604 63334
rect 206004 27654 206604 63098
rect 206004 27418 206186 27654
rect 206422 27418 206604 27654
rect 206004 27334 206604 27418
rect 206004 27098 206186 27334
rect 206422 27098 206604 27334
rect 206004 -4946 206604 27098
rect 206004 -5182 206186 -4946
rect 206422 -5182 206604 -4946
rect 206004 -5266 206604 -5182
rect 206004 -5502 206186 -5266
rect 206422 -5502 206604 -5266
rect 206004 -5524 206604 -5502
rect 209604 679254 210204 710722
rect 227604 710358 228204 711300
rect 227604 710122 227786 710358
rect 228022 710122 228204 710358
rect 227604 710038 228204 710122
rect 227604 709802 227786 710038
rect 228022 709802 228204 710038
rect 224004 708518 224604 709460
rect 224004 708282 224186 708518
rect 224422 708282 224604 708518
rect 224004 708198 224604 708282
rect 224004 707962 224186 708198
rect 224422 707962 224604 708198
rect 220404 706678 221004 707620
rect 220404 706442 220586 706678
rect 220822 706442 221004 706678
rect 220404 706358 221004 706442
rect 220404 706122 220586 706358
rect 220822 706122 221004 706358
rect 209604 679018 209786 679254
rect 210022 679018 210204 679254
rect 209604 678934 210204 679018
rect 209604 678698 209786 678934
rect 210022 678698 210204 678934
rect 209604 643254 210204 678698
rect 209604 643018 209786 643254
rect 210022 643018 210204 643254
rect 209604 642934 210204 643018
rect 209604 642698 209786 642934
rect 210022 642698 210204 642934
rect 209604 607254 210204 642698
rect 209604 607018 209786 607254
rect 210022 607018 210204 607254
rect 209604 606934 210204 607018
rect 209604 606698 209786 606934
rect 210022 606698 210204 606934
rect 209604 571254 210204 606698
rect 209604 571018 209786 571254
rect 210022 571018 210204 571254
rect 209604 570934 210204 571018
rect 209604 570698 209786 570934
rect 210022 570698 210204 570934
rect 209604 535254 210204 570698
rect 209604 535018 209786 535254
rect 210022 535018 210204 535254
rect 209604 534934 210204 535018
rect 209604 534698 209786 534934
rect 210022 534698 210204 534934
rect 209604 499254 210204 534698
rect 209604 499018 209786 499254
rect 210022 499018 210204 499254
rect 209604 498934 210204 499018
rect 209604 498698 209786 498934
rect 210022 498698 210204 498934
rect 209604 463254 210204 498698
rect 209604 463018 209786 463254
rect 210022 463018 210204 463254
rect 209604 462934 210204 463018
rect 209604 462698 209786 462934
rect 210022 462698 210204 462934
rect 209604 427254 210204 462698
rect 209604 427018 209786 427254
rect 210022 427018 210204 427254
rect 209604 426934 210204 427018
rect 209604 426698 209786 426934
rect 210022 426698 210204 426934
rect 209604 391254 210204 426698
rect 209604 391018 209786 391254
rect 210022 391018 210204 391254
rect 209604 390934 210204 391018
rect 209604 390698 209786 390934
rect 210022 390698 210204 390934
rect 209604 355254 210204 390698
rect 209604 355018 209786 355254
rect 210022 355018 210204 355254
rect 209604 354934 210204 355018
rect 209604 354698 209786 354934
rect 210022 354698 210204 354934
rect 209604 319254 210204 354698
rect 209604 319018 209786 319254
rect 210022 319018 210204 319254
rect 209604 318934 210204 319018
rect 209604 318698 209786 318934
rect 210022 318698 210204 318934
rect 209604 283254 210204 318698
rect 209604 283018 209786 283254
rect 210022 283018 210204 283254
rect 209604 282934 210204 283018
rect 209604 282698 209786 282934
rect 210022 282698 210204 282934
rect 209604 247254 210204 282698
rect 209604 247018 209786 247254
rect 210022 247018 210204 247254
rect 209604 246934 210204 247018
rect 209604 246698 209786 246934
rect 210022 246698 210204 246934
rect 209604 211254 210204 246698
rect 209604 211018 209786 211254
rect 210022 211018 210204 211254
rect 209604 210934 210204 211018
rect 209604 210698 209786 210934
rect 210022 210698 210204 210934
rect 209604 175254 210204 210698
rect 209604 175018 209786 175254
rect 210022 175018 210204 175254
rect 209604 174934 210204 175018
rect 209604 174698 209786 174934
rect 210022 174698 210204 174934
rect 209604 139254 210204 174698
rect 209604 139018 209786 139254
rect 210022 139018 210204 139254
rect 209604 138934 210204 139018
rect 209604 138698 209786 138934
rect 210022 138698 210204 138934
rect 209604 103254 210204 138698
rect 209604 103018 209786 103254
rect 210022 103018 210204 103254
rect 209604 102934 210204 103018
rect 209604 102698 209786 102934
rect 210022 102698 210204 102934
rect 209604 67254 210204 102698
rect 209604 67018 209786 67254
rect 210022 67018 210204 67254
rect 209604 66934 210204 67018
rect 209604 66698 209786 66934
rect 210022 66698 210204 66934
rect 209604 31254 210204 66698
rect 209604 31018 209786 31254
rect 210022 31018 210204 31254
rect 209604 30934 210204 31018
rect 209604 30698 209786 30934
rect 210022 30698 210204 30934
rect 191604 -6102 191786 -5866
rect 192022 -6102 192204 -5866
rect 191604 -6186 192204 -6102
rect 191604 -6422 191786 -6186
rect 192022 -6422 192204 -6186
rect 191604 -7364 192204 -6422
rect 209604 -6786 210204 30698
rect 216804 704838 217404 705780
rect 216804 704602 216986 704838
rect 217222 704602 217404 704838
rect 216804 704518 217404 704602
rect 216804 704282 216986 704518
rect 217222 704282 217404 704518
rect 216804 686454 217404 704282
rect 216804 686218 216986 686454
rect 217222 686218 217404 686454
rect 216804 686134 217404 686218
rect 216804 685898 216986 686134
rect 217222 685898 217404 686134
rect 216804 650454 217404 685898
rect 216804 650218 216986 650454
rect 217222 650218 217404 650454
rect 216804 650134 217404 650218
rect 216804 649898 216986 650134
rect 217222 649898 217404 650134
rect 216804 614454 217404 649898
rect 216804 614218 216986 614454
rect 217222 614218 217404 614454
rect 216804 614134 217404 614218
rect 216804 613898 216986 614134
rect 217222 613898 217404 614134
rect 216804 578454 217404 613898
rect 216804 578218 216986 578454
rect 217222 578218 217404 578454
rect 216804 578134 217404 578218
rect 216804 577898 216986 578134
rect 217222 577898 217404 578134
rect 216804 542454 217404 577898
rect 216804 542218 216986 542454
rect 217222 542218 217404 542454
rect 216804 542134 217404 542218
rect 216804 541898 216986 542134
rect 217222 541898 217404 542134
rect 216804 506454 217404 541898
rect 216804 506218 216986 506454
rect 217222 506218 217404 506454
rect 216804 506134 217404 506218
rect 216804 505898 216986 506134
rect 217222 505898 217404 506134
rect 216804 470454 217404 505898
rect 216804 470218 216986 470454
rect 217222 470218 217404 470454
rect 216804 470134 217404 470218
rect 216804 469898 216986 470134
rect 217222 469898 217404 470134
rect 216804 434454 217404 469898
rect 216804 434218 216986 434454
rect 217222 434218 217404 434454
rect 216804 434134 217404 434218
rect 216804 433898 216986 434134
rect 217222 433898 217404 434134
rect 216804 398454 217404 433898
rect 216804 398218 216986 398454
rect 217222 398218 217404 398454
rect 216804 398134 217404 398218
rect 216804 397898 216986 398134
rect 217222 397898 217404 398134
rect 216804 362454 217404 397898
rect 216804 362218 216986 362454
rect 217222 362218 217404 362454
rect 216804 362134 217404 362218
rect 216804 361898 216986 362134
rect 217222 361898 217404 362134
rect 216804 326454 217404 361898
rect 216804 326218 216986 326454
rect 217222 326218 217404 326454
rect 216804 326134 217404 326218
rect 216804 325898 216986 326134
rect 217222 325898 217404 326134
rect 216804 290454 217404 325898
rect 216804 290218 216986 290454
rect 217222 290218 217404 290454
rect 216804 290134 217404 290218
rect 216804 289898 216986 290134
rect 217222 289898 217404 290134
rect 216804 254454 217404 289898
rect 216804 254218 216986 254454
rect 217222 254218 217404 254454
rect 216804 254134 217404 254218
rect 216804 253898 216986 254134
rect 217222 253898 217404 254134
rect 216804 218454 217404 253898
rect 216804 218218 216986 218454
rect 217222 218218 217404 218454
rect 216804 218134 217404 218218
rect 216804 217898 216986 218134
rect 217222 217898 217404 218134
rect 216804 182454 217404 217898
rect 216804 182218 216986 182454
rect 217222 182218 217404 182454
rect 216804 182134 217404 182218
rect 216804 181898 216986 182134
rect 217222 181898 217404 182134
rect 216804 146454 217404 181898
rect 216804 146218 216986 146454
rect 217222 146218 217404 146454
rect 216804 146134 217404 146218
rect 216804 145898 216986 146134
rect 217222 145898 217404 146134
rect 216804 110454 217404 145898
rect 216804 110218 216986 110454
rect 217222 110218 217404 110454
rect 216804 110134 217404 110218
rect 216804 109898 216986 110134
rect 217222 109898 217404 110134
rect 216804 74454 217404 109898
rect 216804 74218 216986 74454
rect 217222 74218 217404 74454
rect 216804 74134 217404 74218
rect 216804 73898 216986 74134
rect 217222 73898 217404 74134
rect 216804 38454 217404 73898
rect 216804 38218 216986 38454
rect 217222 38218 217404 38454
rect 216804 38134 217404 38218
rect 216804 37898 216986 38134
rect 217222 37898 217404 38134
rect 216804 2454 217404 37898
rect 216804 2218 216986 2454
rect 217222 2218 217404 2454
rect 216804 2134 217404 2218
rect 216804 1898 216986 2134
rect 217222 1898 217404 2134
rect 216804 -346 217404 1898
rect 216804 -582 216986 -346
rect 217222 -582 217404 -346
rect 216804 -666 217404 -582
rect 216804 -902 216986 -666
rect 217222 -902 217404 -666
rect 216804 -1844 217404 -902
rect 220404 690054 221004 706122
rect 220404 689818 220586 690054
rect 220822 689818 221004 690054
rect 220404 689734 221004 689818
rect 220404 689498 220586 689734
rect 220822 689498 221004 689734
rect 220404 654054 221004 689498
rect 220404 653818 220586 654054
rect 220822 653818 221004 654054
rect 220404 653734 221004 653818
rect 220404 653498 220586 653734
rect 220822 653498 221004 653734
rect 220404 618054 221004 653498
rect 220404 617818 220586 618054
rect 220822 617818 221004 618054
rect 220404 617734 221004 617818
rect 220404 617498 220586 617734
rect 220822 617498 221004 617734
rect 220404 582054 221004 617498
rect 220404 581818 220586 582054
rect 220822 581818 221004 582054
rect 220404 581734 221004 581818
rect 220404 581498 220586 581734
rect 220822 581498 221004 581734
rect 220404 546054 221004 581498
rect 220404 545818 220586 546054
rect 220822 545818 221004 546054
rect 220404 545734 221004 545818
rect 220404 545498 220586 545734
rect 220822 545498 221004 545734
rect 220404 510054 221004 545498
rect 220404 509818 220586 510054
rect 220822 509818 221004 510054
rect 220404 509734 221004 509818
rect 220404 509498 220586 509734
rect 220822 509498 221004 509734
rect 220404 474054 221004 509498
rect 220404 473818 220586 474054
rect 220822 473818 221004 474054
rect 220404 473734 221004 473818
rect 220404 473498 220586 473734
rect 220822 473498 221004 473734
rect 220404 438054 221004 473498
rect 220404 437818 220586 438054
rect 220822 437818 221004 438054
rect 220404 437734 221004 437818
rect 220404 437498 220586 437734
rect 220822 437498 221004 437734
rect 220404 402054 221004 437498
rect 220404 401818 220586 402054
rect 220822 401818 221004 402054
rect 220404 401734 221004 401818
rect 220404 401498 220586 401734
rect 220822 401498 221004 401734
rect 220404 366054 221004 401498
rect 220404 365818 220586 366054
rect 220822 365818 221004 366054
rect 220404 365734 221004 365818
rect 220404 365498 220586 365734
rect 220822 365498 221004 365734
rect 220404 330054 221004 365498
rect 220404 329818 220586 330054
rect 220822 329818 221004 330054
rect 220404 329734 221004 329818
rect 220404 329498 220586 329734
rect 220822 329498 221004 329734
rect 220404 294054 221004 329498
rect 220404 293818 220586 294054
rect 220822 293818 221004 294054
rect 220404 293734 221004 293818
rect 220404 293498 220586 293734
rect 220822 293498 221004 293734
rect 220404 258054 221004 293498
rect 220404 257818 220586 258054
rect 220822 257818 221004 258054
rect 220404 257734 221004 257818
rect 220404 257498 220586 257734
rect 220822 257498 221004 257734
rect 220404 222054 221004 257498
rect 220404 221818 220586 222054
rect 220822 221818 221004 222054
rect 220404 221734 221004 221818
rect 220404 221498 220586 221734
rect 220822 221498 221004 221734
rect 220404 186054 221004 221498
rect 220404 185818 220586 186054
rect 220822 185818 221004 186054
rect 220404 185734 221004 185818
rect 220404 185498 220586 185734
rect 220822 185498 221004 185734
rect 220404 150054 221004 185498
rect 220404 149818 220586 150054
rect 220822 149818 221004 150054
rect 220404 149734 221004 149818
rect 220404 149498 220586 149734
rect 220822 149498 221004 149734
rect 220404 114054 221004 149498
rect 220404 113818 220586 114054
rect 220822 113818 221004 114054
rect 220404 113734 221004 113818
rect 220404 113498 220586 113734
rect 220822 113498 221004 113734
rect 220404 78054 221004 113498
rect 220404 77818 220586 78054
rect 220822 77818 221004 78054
rect 220404 77734 221004 77818
rect 220404 77498 220586 77734
rect 220822 77498 221004 77734
rect 220404 42054 221004 77498
rect 220404 41818 220586 42054
rect 220822 41818 221004 42054
rect 220404 41734 221004 41818
rect 220404 41498 220586 41734
rect 220822 41498 221004 41734
rect 220404 6054 221004 41498
rect 220404 5818 220586 6054
rect 220822 5818 221004 6054
rect 220404 5734 221004 5818
rect 220404 5498 220586 5734
rect 220822 5498 221004 5734
rect 220404 -2186 221004 5498
rect 220404 -2422 220586 -2186
rect 220822 -2422 221004 -2186
rect 220404 -2506 221004 -2422
rect 220404 -2742 220586 -2506
rect 220822 -2742 221004 -2506
rect 220404 -3684 221004 -2742
rect 224004 693654 224604 707962
rect 224004 693418 224186 693654
rect 224422 693418 224604 693654
rect 224004 693334 224604 693418
rect 224004 693098 224186 693334
rect 224422 693098 224604 693334
rect 224004 657654 224604 693098
rect 224004 657418 224186 657654
rect 224422 657418 224604 657654
rect 224004 657334 224604 657418
rect 224004 657098 224186 657334
rect 224422 657098 224604 657334
rect 224004 621654 224604 657098
rect 224004 621418 224186 621654
rect 224422 621418 224604 621654
rect 224004 621334 224604 621418
rect 224004 621098 224186 621334
rect 224422 621098 224604 621334
rect 224004 585654 224604 621098
rect 224004 585418 224186 585654
rect 224422 585418 224604 585654
rect 224004 585334 224604 585418
rect 224004 585098 224186 585334
rect 224422 585098 224604 585334
rect 224004 549654 224604 585098
rect 224004 549418 224186 549654
rect 224422 549418 224604 549654
rect 224004 549334 224604 549418
rect 224004 549098 224186 549334
rect 224422 549098 224604 549334
rect 224004 513654 224604 549098
rect 224004 513418 224186 513654
rect 224422 513418 224604 513654
rect 224004 513334 224604 513418
rect 224004 513098 224186 513334
rect 224422 513098 224604 513334
rect 224004 477654 224604 513098
rect 224004 477418 224186 477654
rect 224422 477418 224604 477654
rect 224004 477334 224604 477418
rect 224004 477098 224186 477334
rect 224422 477098 224604 477334
rect 224004 441654 224604 477098
rect 224004 441418 224186 441654
rect 224422 441418 224604 441654
rect 224004 441334 224604 441418
rect 224004 441098 224186 441334
rect 224422 441098 224604 441334
rect 224004 405654 224604 441098
rect 224004 405418 224186 405654
rect 224422 405418 224604 405654
rect 224004 405334 224604 405418
rect 224004 405098 224186 405334
rect 224422 405098 224604 405334
rect 224004 369654 224604 405098
rect 224004 369418 224186 369654
rect 224422 369418 224604 369654
rect 224004 369334 224604 369418
rect 224004 369098 224186 369334
rect 224422 369098 224604 369334
rect 224004 333654 224604 369098
rect 224004 333418 224186 333654
rect 224422 333418 224604 333654
rect 224004 333334 224604 333418
rect 224004 333098 224186 333334
rect 224422 333098 224604 333334
rect 224004 297654 224604 333098
rect 224004 297418 224186 297654
rect 224422 297418 224604 297654
rect 224004 297334 224604 297418
rect 224004 297098 224186 297334
rect 224422 297098 224604 297334
rect 224004 261654 224604 297098
rect 224004 261418 224186 261654
rect 224422 261418 224604 261654
rect 224004 261334 224604 261418
rect 224004 261098 224186 261334
rect 224422 261098 224604 261334
rect 224004 225654 224604 261098
rect 224004 225418 224186 225654
rect 224422 225418 224604 225654
rect 224004 225334 224604 225418
rect 224004 225098 224186 225334
rect 224422 225098 224604 225334
rect 224004 189654 224604 225098
rect 224004 189418 224186 189654
rect 224422 189418 224604 189654
rect 224004 189334 224604 189418
rect 224004 189098 224186 189334
rect 224422 189098 224604 189334
rect 224004 153654 224604 189098
rect 224004 153418 224186 153654
rect 224422 153418 224604 153654
rect 224004 153334 224604 153418
rect 224004 153098 224186 153334
rect 224422 153098 224604 153334
rect 224004 117654 224604 153098
rect 224004 117418 224186 117654
rect 224422 117418 224604 117654
rect 224004 117334 224604 117418
rect 224004 117098 224186 117334
rect 224422 117098 224604 117334
rect 224004 81654 224604 117098
rect 224004 81418 224186 81654
rect 224422 81418 224604 81654
rect 224004 81334 224604 81418
rect 224004 81098 224186 81334
rect 224422 81098 224604 81334
rect 224004 45654 224604 81098
rect 224004 45418 224186 45654
rect 224422 45418 224604 45654
rect 224004 45334 224604 45418
rect 224004 45098 224186 45334
rect 224422 45098 224604 45334
rect 224004 9654 224604 45098
rect 224004 9418 224186 9654
rect 224422 9418 224604 9654
rect 224004 9334 224604 9418
rect 224004 9098 224186 9334
rect 224422 9098 224604 9334
rect 224004 -4026 224604 9098
rect 224004 -4262 224186 -4026
rect 224422 -4262 224604 -4026
rect 224004 -4346 224604 -4262
rect 224004 -4582 224186 -4346
rect 224422 -4582 224604 -4346
rect 224004 -5524 224604 -4582
rect 227604 697254 228204 709802
rect 245604 711278 246204 711300
rect 245604 711042 245786 711278
rect 246022 711042 246204 711278
rect 245604 710958 246204 711042
rect 245604 710722 245786 710958
rect 246022 710722 246204 710958
rect 242004 709438 242604 709460
rect 242004 709202 242186 709438
rect 242422 709202 242604 709438
rect 242004 709118 242604 709202
rect 242004 708882 242186 709118
rect 242422 708882 242604 709118
rect 238404 707598 239004 707620
rect 238404 707362 238586 707598
rect 238822 707362 239004 707598
rect 238404 707278 239004 707362
rect 238404 707042 238586 707278
rect 238822 707042 239004 707278
rect 227604 697018 227786 697254
rect 228022 697018 228204 697254
rect 227604 696934 228204 697018
rect 227604 696698 227786 696934
rect 228022 696698 228204 696934
rect 227604 661254 228204 696698
rect 227604 661018 227786 661254
rect 228022 661018 228204 661254
rect 227604 660934 228204 661018
rect 227604 660698 227786 660934
rect 228022 660698 228204 660934
rect 227604 625254 228204 660698
rect 227604 625018 227786 625254
rect 228022 625018 228204 625254
rect 227604 624934 228204 625018
rect 227604 624698 227786 624934
rect 228022 624698 228204 624934
rect 227604 589254 228204 624698
rect 227604 589018 227786 589254
rect 228022 589018 228204 589254
rect 227604 588934 228204 589018
rect 227604 588698 227786 588934
rect 228022 588698 228204 588934
rect 227604 553254 228204 588698
rect 227604 553018 227786 553254
rect 228022 553018 228204 553254
rect 227604 552934 228204 553018
rect 227604 552698 227786 552934
rect 228022 552698 228204 552934
rect 227604 517254 228204 552698
rect 227604 517018 227786 517254
rect 228022 517018 228204 517254
rect 227604 516934 228204 517018
rect 227604 516698 227786 516934
rect 228022 516698 228204 516934
rect 227604 481254 228204 516698
rect 227604 481018 227786 481254
rect 228022 481018 228204 481254
rect 227604 480934 228204 481018
rect 227604 480698 227786 480934
rect 228022 480698 228204 480934
rect 227604 445254 228204 480698
rect 227604 445018 227786 445254
rect 228022 445018 228204 445254
rect 227604 444934 228204 445018
rect 227604 444698 227786 444934
rect 228022 444698 228204 444934
rect 227604 409254 228204 444698
rect 227604 409018 227786 409254
rect 228022 409018 228204 409254
rect 227604 408934 228204 409018
rect 227604 408698 227786 408934
rect 228022 408698 228204 408934
rect 227604 373254 228204 408698
rect 234804 705758 235404 705780
rect 234804 705522 234986 705758
rect 235222 705522 235404 705758
rect 234804 705438 235404 705522
rect 234804 705202 234986 705438
rect 235222 705202 235404 705438
rect 234804 668454 235404 705202
rect 234804 668218 234986 668454
rect 235222 668218 235404 668454
rect 234804 668134 235404 668218
rect 234804 667898 234986 668134
rect 235222 667898 235404 668134
rect 234804 632454 235404 667898
rect 234804 632218 234986 632454
rect 235222 632218 235404 632454
rect 234804 632134 235404 632218
rect 234804 631898 234986 632134
rect 235222 631898 235404 632134
rect 234804 596454 235404 631898
rect 234804 596218 234986 596454
rect 235222 596218 235404 596454
rect 234804 596134 235404 596218
rect 234804 595898 234986 596134
rect 235222 595898 235404 596134
rect 234804 560454 235404 595898
rect 234804 560218 234986 560454
rect 235222 560218 235404 560454
rect 234804 560134 235404 560218
rect 234804 559898 234986 560134
rect 235222 559898 235404 560134
rect 234804 524454 235404 559898
rect 234804 524218 234986 524454
rect 235222 524218 235404 524454
rect 234804 524134 235404 524218
rect 234804 523898 234986 524134
rect 235222 523898 235404 524134
rect 234804 488454 235404 523898
rect 234804 488218 234986 488454
rect 235222 488218 235404 488454
rect 234804 488134 235404 488218
rect 234804 487898 234986 488134
rect 235222 487898 235404 488134
rect 234804 452454 235404 487898
rect 234804 452218 234986 452454
rect 235222 452218 235404 452454
rect 234804 452134 235404 452218
rect 234804 451898 234986 452134
rect 235222 451898 235404 452134
rect 234804 416454 235404 451898
rect 234804 416218 234986 416454
rect 235222 416218 235404 416454
rect 234804 416134 235404 416218
rect 234804 415898 234986 416134
rect 235222 415898 235404 416134
rect 231715 399396 231781 399397
rect 231715 399332 231716 399396
rect 231780 399332 231781 399396
rect 231715 399331 231781 399332
rect 233003 399396 233069 399397
rect 233003 399332 233004 399396
rect 233068 399332 233069 399396
rect 233003 399331 233069 399332
rect 233923 399396 233989 399397
rect 233923 399332 233924 399396
rect 233988 399332 233989 399396
rect 233923 399331 233989 399332
rect 227604 373018 227786 373254
rect 228022 373018 228204 373254
rect 227604 372934 228204 373018
rect 227604 372698 227786 372934
rect 228022 372698 228204 372934
rect 227604 337254 228204 372698
rect 227604 337018 227786 337254
rect 228022 337018 228204 337254
rect 227604 336934 228204 337018
rect 227604 336698 227786 336934
rect 228022 336698 228204 336934
rect 227604 301254 228204 336698
rect 227604 301018 227786 301254
rect 228022 301018 228204 301254
rect 227604 300934 228204 301018
rect 227604 300698 227786 300934
rect 228022 300698 228204 300934
rect 227604 265254 228204 300698
rect 227604 265018 227786 265254
rect 228022 265018 228204 265254
rect 227604 264934 228204 265018
rect 227604 264698 227786 264934
rect 228022 264698 228204 264934
rect 227604 229254 228204 264698
rect 227604 229018 227786 229254
rect 228022 229018 228204 229254
rect 227604 228934 228204 229018
rect 227604 228698 227786 228934
rect 228022 228698 228204 228934
rect 227604 193254 228204 228698
rect 227604 193018 227786 193254
rect 228022 193018 228204 193254
rect 227604 192934 228204 193018
rect 227604 192698 227786 192934
rect 228022 192698 228204 192934
rect 227604 157254 228204 192698
rect 227604 157018 227786 157254
rect 228022 157018 228204 157254
rect 227604 156934 228204 157018
rect 227604 156698 227786 156934
rect 228022 156698 228204 156934
rect 227604 121254 228204 156698
rect 227604 121018 227786 121254
rect 228022 121018 228204 121254
rect 227604 120934 228204 121018
rect 227604 120698 227786 120934
rect 228022 120698 228204 120934
rect 227604 85254 228204 120698
rect 227604 85018 227786 85254
rect 228022 85018 228204 85254
rect 227604 84934 228204 85018
rect 227604 84698 227786 84934
rect 228022 84698 228204 84934
rect 227604 49254 228204 84698
rect 229507 67556 229573 67557
rect 229507 67492 229508 67556
rect 229572 67492 229573 67556
rect 229507 67491 229573 67492
rect 229510 58170 229570 67491
rect 229510 58110 229754 58170
rect 229694 58037 229754 58110
rect 229691 58036 229757 58037
rect 229691 57972 229692 58036
rect 229756 57972 229757 58036
rect 229691 57971 229757 57972
rect 227604 49018 227786 49254
rect 228022 49018 228204 49254
rect 227604 48934 228204 49018
rect 227604 48698 227786 48934
rect 228022 48698 228204 48934
rect 227604 13254 228204 48698
rect 231718 29205 231778 399331
rect 233006 76261 233066 399331
rect 233926 338741 233986 399331
rect 234804 380454 235404 415898
rect 238404 672054 239004 707042
rect 238404 671818 238586 672054
rect 238822 671818 239004 672054
rect 238404 671734 239004 671818
rect 238404 671498 238586 671734
rect 238822 671498 239004 671734
rect 238404 636054 239004 671498
rect 238404 635818 238586 636054
rect 238822 635818 239004 636054
rect 238404 635734 239004 635818
rect 238404 635498 238586 635734
rect 238822 635498 239004 635734
rect 238404 600054 239004 635498
rect 238404 599818 238586 600054
rect 238822 599818 239004 600054
rect 238404 599734 239004 599818
rect 238404 599498 238586 599734
rect 238822 599498 239004 599734
rect 238404 564054 239004 599498
rect 238404 563818 238586 564054
rect 238822 563818 239004 564054
rect 238404 563734 239004 563818
rect 238404 563498 238586 563734
rect 238822 563498 239004 563734
rect 238404 528054 239004 563498
rect 238404 527818 238586 528054
rect 238822 527818 239004 528054
rect 238404 527734 239004 527818
rect 238404 527498 238586 527734
rect 238822 527498 239004 527734
rect 238404 492054 239004 527498
rect 238404 491818 238586 492054
rect 238822 491818 239004 492054
rect 238404 491734 239004 491818
rect 238404 491498 238586 491734
rect 238822 491498 239004 491734
rect 238404 456054 239004 491498
rect 238404 455818 238586 456054
rect 238822 455818 239004 456054
rect 238404 455734 239004 455818
rect 238404 455498 238586 455734
rect 238822 455498 239004 455734
rect 238404 420054 239004 455498
rect 238404 419818 238586 420054
rect 238822 419818 239004 420054
rect 238404 419734 239004 419818
rect 238404 419498 238586 419734
rect 238822 419498 239004 419734
rect 237235 399396 237301 399397
rect 237235 399332 237236 399396
rect 237300 399332 237301 399396
rect 237235 399331 237301 399332
rect 238155 399396 238221 399397
rect 238155 399332 238156 399396
rect 238220 399332 238221 399396
rect 238155 399331 238221 399332
rect 234804 380218 234986 380454
rect 235222 380218 235404 380454
rect 234804 380134 235404 380218
rect 234804 379898 234986 380134
rect 235222 379898 235404 380134
rect 234804 344454 235404 379898
rect 234804 344218 234986 344454
rect 235222 344218 235404 344454
rect 234804 344134 235404 344218
rect 234804 343898 234986 344134
rect 235222 343898 235404 344134
rect 233923 338740 233989 338741
rect 233923 338676 233924 338740
rect 233988 338676 233989 338740
rect 233923 338675 233989 338676
rect 234804 308454 235404 343898
rect 234804 308218 234986 308454
rect 235222 308218 235404 308454
rect 234804 308134 235404 308218
rect 234804 307898 234986 308134
rect 235222 307898 235404 308134
rect 234804 272454 235404 307898
rect 234804 272218 234986 272454
rect 235222 272218 235404 272454
rect 234804 272134 235404 272218
rect 234804 271898 234986 272134
rect 235222 271898 235404 272134
rect 234804 236454 235404 271898
rect 234804 236218 234986 236454
rect 235222 236218 235404 236454
rect 234804 236134 235404 236218
rect 234804 235898 234986 236134
rect 235222 235898 235404 236134
rect 234804 200454 235404 235898
rect 237238 228173 237298 399331
rect 238158 340101 238218 399331
rect 238404 384054 239004 419498
rect 242004 675654 242604 708882
rect 242004 675418 242186 675654
rect 242422 675418 242604 675654
rect 242004 675334 242604 675418
rect 242004 675098 242186 675334
rect 242422 675098 242604 675334
rect 242004 639654 242604 675098
rect 242004 639418 242186 639654
rect 242422 639418 242604 639654
rect 242004 639334 242604 639418
rect 242004 639098 242186 639334
rect 242422 639098 242604 639334
rect 242004 603654 242604 639098
rect 242004 603418 242186 603654
rect 242422 603418 242604 603654
rect 242004 603334 242604 603418
rect 242004 603098 242186 603334
rect 242422 603098 242604 603334
rect 242004 567654 242604 603098
rect 242004 567418 242186 567654
rect 242422 567418 242604 567654
rect 242004 567334 242604 567418
rect 242004 567098 242186 567334
rect 242422 567098 242604 567334
rect 242004 531654 242604 567098
rect 242004 531418 242186 531654
rect 242422 531418 242604 531654
rect 242004 531334 242604 531418
rect 242004 531098 242186 531334
rect 242422 531098 242604 531334
rect 242004 495654 242604 531098
rect 242004 495418 242186 495654
rect 242422 495418 242604 495654
rect 242004 495334 242604 495418
rect 242004 495098 242186 495334
rect 242422 495098 242604 495334
rect 242004 459654 242604 495098
rect 242004 459418 242186 459654
rect 242422 459418 242604 459654
rect 242004 459334 242604 459418
rect 242004 459098 242186 459334
rect 242422 459098 242604 459334
rect 242004 423654 242604 459098
rect 242004 423418 242186 423654
rect 242422 423418 242604 423654
rect 242004 423334 242604 423418
rect 242004 423098 242186 423334
rect 242422 423098 242604 423334
rect 239995 399396 240061 399397
rect 239995 399332 239996 399396
rect 240060 399332 240061 399396
rect 239995 399331 240061 399332
rect 241283 399396 241349 399397
rect 241283 399332 241284 399396
rect 241348 399332 241349 399396
rect 241283 399331 241349 399332
rect 238404 383818 238586 384054
rect 238822 383818 239004 384054
rect 238404 383734 239004 383818
rect 238404 383498 238586 383734
rect 238822 383498 239004 383734
rect 238404 348054 239004 383498
rect 238404 347818 238586 348054
rect 238822 347818 239004 348054
rect 238404 347734 239004 347818
rect 238404 347498 238586 347734
rect 238822 347498 239004 347734
rect 238155 340100 238221 340101
rect 238155 340036 238156 340100
rect 238220 340036 238221 340100
rect 238155 340035 238221 340036
rect 238404 312054 239004 347498
rect 239998 338877 240058 399331
rect 239995 338876 240061 338877
rect 239995 338812 239996 338876
rect 240060 338812 240061 338876
rect 239995 338811 240061 338812
rect 238404 311818 238586 312054
rect 238822 311818 239004 312054
rect 238404 311734 239004 311818
rect 238404 311498 238586 311734
rect 238822 311498 239004 311734
rect 237787 278764 237853 278765
rect 237787 278700 237788 278764
rect 237852 278700 237853 278764
rect 237787 278699 237853 278700
rect 237790 264349 237850 278699
rect 238404 276054 239004 311498
rect 241286 310997 241346 399331
rect 242004 387654 242604 423098
rect 245604 679254 246204 710722
rect 263604 710358 264204 711300
rect 263604 710122 263786 710358
rect 264022 710122 264204 710358
rect 263604 710038 264204 710122
rect 263604 709802 263786 710038
rect 264022 709802 264204 710038
rect 260004 708518 260604 709460
rect 260004 708282 260186 708518
rect 260422 708282 260604 708518
rect 260004 708198 260604 708282
rect 260004 707962 260186 708198
rect 260422 707962 260604 708198
rect 256404 706678 257004 707620
rect 256404 706442 256586 706678
rect 256822 706442 257004 706678
rect 256404 706358 257004 706442
rect 256404 706122 256586 706358
rect 256822 706122 257004 706358
rect 245604 679018 245786 679254
rect 246022 679018 246204 679254
rect 245604 678934 246204 679018
rect 245604 678698 245786 678934
rect 246022 678698 246204 678934
rect 245604 643254 246204 678698
rect 245604 643018 245786 643254
rect 246022 643018 246204 643254
rect 245604 642934 246204 643018
rect 245604 642698 245786 642934
rect 246022 642698 246204 642934
rect 245604 607254 246204 642698
rect 245604 607018 245786 607254
rect 246022 607018 246204 607254
rect 245604 606934 246204 607018
rect 245604 606698 245786 606934
rect 246022 606698 246204 606934
rect 245604 571254 246204 606698
rect 245604 571018 245786 571254
rect 246022 571018 246204 571254
rect 245604 570934 246204 571018
rect 245604 570698 245786 570934
rect 246022 570698 246204 570934
rect 245604 535254 246204 570698
rect 245604 535018 245786 535254
rect 246022 535018 246204 535254
rect 245604 534934 246204 535018
rect 245604 534698 245786 534934
rect 246022 534698 246204 534934
rect 245604 499254 246204 534698
rect 245604 499018 245786 499254
rect 246022 499018 246204 499254
rect 245604 498934 246204 499018
rect 245604 498698 245786 498934
rect 246022 498698 246204 498934
rect 245604 463254 246204 498698
rect 245604 463018 245786 463254
rect 246022 463018 246204 463254
rect 245604 462934 246204 463018
rect 245604 462698 245786 462934
rect 246022 462698 246204 462934
rect 245604 427254 246204 462698
rect 245604 427018 245786 427254
rect 246022 427018 246204 427254
rect 245604 426934 246204 427018
rect 245604 426698 245786 426934
rect 246022 426698 246204 426934
rect 243491 399532 243557 399533
rect 243491 399468 243492 399532
rect 243556 399468 243557 399532
rect 243491 399467 243557 399468
rect 242004 387418 242186 387654
rect 242422 387418 242604 387654
rect 242004 387334 242604 387418
rect 242004 387098 242186 387334
rect 242422 387098 242604 387334
rect 242004 351654 242604 387098
rect 242004 351418 242186 351654
rect 242422 351418 242604 351654
rect 242004 351334 242604 351418
rect 242004 351098 242186 351334
rect 242422 351098 242604 351334
rect 242004 315654 242604 351098
rect 243494 321605 243554 399467
rect 245604 391254 246204 426698
rect 245604 391018 245786 391254
rect 246022 391018 246204 391254
rect 245604 390934 246204 391018
rect 245604 390698 245786 390934
rect 246022 390698 246204 390934
rect 245604 355254 246204 390698
rect 245604 355018 245786 355254
rect 246022 355018 246204 355254
rect 245604 354934 246204 355018
rect 245604 354698 245786 354934
rect 246022 354698 246204 354934
rect 243491 321604 243557 321605
rect 243491 321540 243492 321604
rect 243556 321540 243557 321604
rect 243491 321539 243557 321540
rect 242004 315418 242186 315654
rect 242422 315418 242604 315654
rect 242004 315334 242604 315418
rect 242004 315098 242186 315334
rect 242422 315098 242604 315334
rect 241283 310996 241349 310997
rect 241283 310932 241284 310996
rect 241348 310932 241349 310996
rect 241283 310931 241349 310932
rect 238404 275818 238586 276054
rect 238822 275818 239004 276054
rect 238404 275734 239004 275818
rect 238404 275498 238586 275734
rect 238822 275498 239004 275734
rect 237787 264348 237853 264349
rect 237787 264284 237788 264348
rect 237852 264284 237853 264348
rect 237787 264283 237853 264284
rect 238404 240054 239004 275498
rect 238404 239818 238586 240054
rect 238822 239818 239004 240054
rect 238404 239734 239004 239818
rect 238404 239498 238586 239734
rect 238822 239498 239004 239734
rect 237235 228172 237301 228173
rect 237235 228108 237236 228172
rect 237300 228108 237301 228172
rect 237235 228107 237301 228108
rect 234804 200218 234986 200454
rect 235222 200218 235404 200454
rect 234804 200134 235404 200218
rect 234804 199898 234986 200134
rect 235222 199898 235404 200134
rect 234804 164454 235404 199898
rect 234804 164218 234986 164454
rect 235222 164218 235404 164454
rect 234804 164134 235404 164218
rect 234804 163898 234986 164134
rect 235222 163898 235404 164134
rect 234804 128454 235404 163898
rect 234804 128218 234986 128454
rect 235222 128218 235404 128454
rect 234804 128134 235404 128218
rect 234804 127898 234986 128134
rect 235222 127898 235404 128134
rect 234804 92454 235404 127898
rect 234804 92218 234986 92454
rect 235222 92218 235404 92454
rect 234804 92134 235404 92218
rect 234804 91898 234986 92134
rect 235222 91898 235404 92134
rect 233003 76260 233069 76261
rect 233003 76196 233004 76260
rect 233068 76196 233069 76260
rect 233003 76195 233069 76196
rect 234804 56454 235404 91898
rect 234804 56218 234986 56454
rect 235222 56218 235404 56454
rect 234804 56134 235404 56218
rect 234804 55898 234986 56134
rect 235222 55898 235404 56134
rect 231715 29204 231781 29205
rect 231715 29140 231716 29204
rect 231780 29140 231781 29204
rect 231715 29139 231781 29140
rect 227604 13018 227786 13254
rect 228022 13018 228204 13254
rect 227604 12934 228204 13018
rect 227604 12698 227786 12934
rect 228022 12698 228204 12934
rect 209604 -7022 209786 -6786
rect 210022 -7022 210204 -6786
rect 209604 -7106 210204 -7022
rect 209604 -7342 209786 -7106
rect 210022 -7342 210204 -7106
rect 209604 -7364 210204 -7342
rect 227604 -5866 228204 12698
rect 234804 20454 235404 55898
rect 234804 20218 234986 20454
rect 235222 20218 235404 20454
rect 234804 20134 235404 20218
rect 234804 19898 234986 20134
rect 235222 19898 235404 20134
rect 234804 -1266 235404 19898
rect 234804 -1502 234986 -1266
rect 235222 -1502 235404 -1266
rect 234804 -1586 235404 -1502
rect 234804 -1822 234986 -1586
rect 235222 -1822 235404 -1586
rect 234804 -1844 235404 -1822
rect 238404 204054 239004 239498
rect 238404 203818 238586 204054
rect 238822 203818 239004 204054
rect 238404 203734 239004 203818
rect 238404 203498 238586 203734
rect 238822 203498 239004 203734
rect 238404 168054 239004 203498
rect 238404 167818 238586 168054
rect 238822 167818 239004 168054
rect 238404 167734 239004 167818
rect 238404 167498 238586 167734
rect 238822 167498 239004 167734
rect 238404 132054 239004 167498
rect 238404 131818 238586 132054
rect 238822 131818 239004 132054
rect 238404 131734 239004 131818
rect 238404 131498 238586 131734
rect 238822 131498 239004 131734
rect 238404 96054 239004 131498
rect 238404 95818 238586 96054
rect 238822 95818 239004 96054
rect 238404 95734 239004 95818
rect 238404 95498 238586 95734
rect 238822 95498 239004 95734
rect 238404 60054 239004 95498
rect 242004 279654 242604 315098
rect 242004 279418 242186 279654
rect 242422 279418 242604 279654
rect 242004 279334 242604 279418
rect 242004 279098 242186 279334
rect 242422 279098 242604 279334
rect 242004 243654 242604 279098
rect 242004 243418 242186 243654
rect 242422 243418 242604 243654
rect 242004 243334 242604 243418
rect 242004 243098 242186 243334
rect 242422 243098 242604 243334
rect 242004 207654 242604 243098
rect 242004 207418 242186 207654
rect 242422 207418 242604 207654
rect 242004 207334 242604 207418
rect 242004 207098 242186 207334
rect 242422 207098 242604 207334
rect 242004 171654 242604 207098
rect 242004 171418 242186 171654
rect 242422 171418 242604 171654
rect 242004 171334 242604 171418
rect 242004 171098 242186 171334
rect 242422 171098 242604 171334
rect 242004 135654 242604 171098
rect 242004 135418 242186 135654
rect 242422 135418 242604 135654
rect 242004 135334 242604 135418
rect 242004 135098 242186 135334
rect 242422 135098 242604 135334
rect 242004 99654 242604 135098
rect 242004 99418 242186 99654
rect 242422 99418 242604 99654
rect 242004 99334 242604 99418
rect 242004 99098 242186 99334
rect 242422 99098 242604 99334
rect 241467 76260 241533 76261
rect 241467 76196 241468 76260
rect 241532 76196 241533 76260
rect 241467 76195 241533 76196
rect 241470 75989 241530 76195
rect 241467 75988 241533 75989
rect 241467 75924 241468 75988
rect 241532 75924 241533 75988
rect 241467 75923 241533 75924
rect 238404 59818 238586 60054
rect 238822 59818 239004 60054
rect 238404 59734 239004 59818
rect 238404 59498 238586 59734
rect 238822 59498 239004 59734
rect 238404 24054 239004 59498
rect 238404 23818 238586 24054
rect 238822 23818 239004 24054
rect 238404 23734 239004 23818
rect 238404 23498 238586 23734
rect 238822 23498 239004 23734
rect 238404 -3106 239004 23498
rect 238404 -3342 238586 -3106
rect 238822 -3342 239004 -3106
rect 238404 -3426 239004 -3342
rect 238404 -3662 238586 -3426
rect 238822 -3662 239004 -3426
rect 238404 -3684 239004 -3662
rect 242004 63654 242604 99098
rect 242004 63418 242186 63654
rect 242422 63418 242604 63654
rect 242004 63334 242604 63418
rect 242004 63098 242186 63334
rect 242422 63098 242604 63334
rect 242004 27654 242604 63098
rect 242004 27418 242186 27654
rect 242422 27418 242604 27654
rect 242004 27334 242604 27418
rect 242004 27098 242186 27334
rect 242422 27098 242604 27334
rect 242004 -4946 242604 27098
rect 242004 -5182 242186 -4946
rect 242422 -5182 242604 -4946
rect 242004 -5266 242604 -5182
rect 242004 -5502 242186 -5266
rect 242422 -5502 242604 -5266
rect 242004 -5524 242604 -5502
rect 245604 319254 246204 354698
rect 245604 319018 245786 319254
rect 246022 319018 246204 319254
rect 245604 318934 246204 319018
rect 245604 318698 245786 318934
rect 246022 318698 246204 318934
rect 245604 283254 246204 318698
rect 245604 283018 245786 283254
rect 246022 283018 246204 283254
rect 245604 282934 246204 283018
rect 245604 282698 245786 282934
rect 246022 282698 246204 282934
rect 245604 247254 246204 282698
rect 245604 247018 245786 247254
rect 246022 247018 246204 247254
rect 245604 246934 246204 247018
rect 245604 246698 245786 246934
rect 246022 246698 246204 246934
rect 245604 211254 246204 246698
rect 245604 211018 245786 211254
rect 246022 211018 246204 211254
rect 245604 210934 246204 211018
rect 245604 210698 245786 210934
rect 246022 210698 246204 210934
rect 245604 175254 246204 210698
rect 245604 175018 245786 175254
rect 246022 175018 246204 175254
rect 245604 174934 246204 175018
rect 245604 174698 245786 174934
rect 246022 174698 246204 174934
rect 245604 139254 246204 174698
rect 245604 139018 245786 139254
rect 246022 139018 246204 139254
rect 245604 138934 246204 139018
rect 245604 138698 245786 138934
rect 246022 138698 246204 138934
rect 245604 103254 246204 138698
rect 245604 103018 245786 103254
rect 246022 103018 246204 103254
rect 245604 102934 246204 103018
rect 245604 102698 245786 102934
rect 246022 102698 246204 102934
rect 245604 67254 246204 102698
rect 245604 67018 245786 67254
rect 246022 67018 246204 67254
rect 245604 66934 246204 67018
rect 245604 66698 245786 66934
rect 246022 66698 246204 66934
rect 245604 31254 246204 66698
rect 245604 31018 245786 31254
rect 246022 31018 246204 31254
rect 245604 30934 246204 31018
rect 245604 30698 245786 30934
rect 246022 30698 246204 30934
rect 227604 -6102 227786 -5866
rect 228022 -6102 228204 -5866
rect 227604 -6186 228204 -6102
rect 227604 -6422 227786 -6186
rect 228022 -6422 228204 -6186
rect 227604 -7364 228204 -6422
rect 245604 -6786 246204 30698
rect 252804 704838 253404 705780
rect 252804 704602 252986 704838
rect 253222 704602 253404 704838
rect 252804 704518 253404 704602
rect 252804 704282 252986 704518
rect 253222 704282 253404 704518
rect 252804 686454 253404 704282
rect 252804 686218 252986 686454
rect 253222 686218 253404 686454
rect 252804 686134 253404 686218
rect 252804 685898 252986 686134
rect 253222 685898 253404 686134
rect 252804 650454 253404 685898
rect 252804 650218 252986 650454
rect 253222 650218 253404 650454
rect 252804 650134 253404 650218
rect 252804 649898 252986 650134
rect 253222 649898 253404 650134
rect 252804 614454 253404 649898
rect 252804 614218 252986 614454
rect 253222 614218 253404 614454
rect 252804 614134 253404 614218
rect 252804 613898 252986 614134
rect 253222 613898 253404 614134
rect 252804 578454 253404 613898
rect 252804 578218 252986 578454
rect 253222 578218 253404 578454
rect 252804 578134 253404 578218
rect 252804 577898 252986 578134
rect 253222 577898 253404 578134
rect 252804 542454 253404 577898
rect 252804 542218 252986 542454
rect 253222 542218 253404 542454
rect 252804 542134 253404 542218
rect 252804 541898 252986 542134
rect 253222 541898 253404 542134
rect 252804 506454 253404 541898
rect 252804 506218 252986 506454
rect 253222 506218 253404 506454
rect 252804 506134 253404 506218
rect 252804 505898 252986 506134
rect 253222 505898 253404 506134
rect 252804 470454 253404 505898
rect 252804 470218 252986 470454
rect 253222 470218 253404 470454
rect 252804 470134 253404 470218
rect 252804 469898 252986 470134
rect 253222 469898 253404 470134
rect 252804 434454 253404 469898
rect 252804 434218 252986 434454
rect 253222 434218 253404 434454
rect 252804 434134 253404 434218
rect 252804 433898 252986 434134
rect 253222 433898 253404 434134
rect 252804 398454 253404 433898
rect 252804 398218 252986 398454
rect 253222 398218 253404 398454
rect 252804 398134 253404 398218
rect 252804 397898 252986 398134
rect 253222 397898 253404 398134
rect 252804 362454 253404 397898
rect 252804 362218 252986 362454
rect 253222 362218 253404 362454
rect 252804 362134 253404 362218
rect 252804 361898 252986 362134
rect 253222 361898 253404 362134
rect 252804 326454 253404 361898
rect 252804 326218 252986 326454
rect 253222 326218 253404 326454
rect 252804 326134 253404 326218
rect 252804 325898 252986 326134
rect 253222 325898 253404 326134
rect 252804 290454 253404 325898
rect 252804 290218 252986 290454
rect 253222 290218 253404 290454
rect 252804 290134 253404 290218
rect 252804 289898 252986 290134
rect 253222 289898 253404 290134
rect 252804 254454 253404 289898
rect 252804 254218 252986 254454
rect 253222 254218 253404 254454
rect 252804 254134 253404 254218
rect 252804 253898 252986 254134
rect 253222 253898 253404 254134
rect 252804 218454 253404 253898
rect 252804 218218 252986 218454
rect 253222 218218 253404 218454
rect 252804 218134 253404 218218
rect 252804 217898 252986 218134
rect 253222 217898 253404 218134
rect 252804 182454 253404 217898
rect 252804 182218 252986 182454
rect 253222 182218 253404 182454
rect 252804 182134 253404 182218
rect 252804 181898 252986 182134
rect 253222 181898 253404 182134
rect 252804 146454 253404 181898
rect 252804 146218 252986 146454
rect 253222 146218 253404 146454
rect 252804 146134 253404 146218
rect 252804 145898 252986 146134
rect 253222 145898 253404 146134
rect 252804 110454 253404 145898
rect 252804 110218 252986 110454
rect 253222 110218 253404 110454
rect 252804 110134 253404 110218
rect 252804 109898 252986 110134
rect 253222 109898 253404 110134
rect 252804 74454 253404 109898
rect 252804 74218 252986 74454
rect 253222 74218 253404 74454
rect 252804 74134 253404 74218
rect 252804 73898 252986 74134
rect 253222 73898 253404 74134
rect 252804 38454 253404 73898
rect 252804 38218 252986 38454
rect 253222 38218 253404 38454
rect 252804 38134 253404 38218
rect 252804 37898 252986 38134
rect 253222 37898 253404 38134
rect 249747 29204 249813 29205
rect 249747 29140 249748 29204
rect 249812 29202 249813 29204
rect 249812 29142 249994 29202
rect 249812 29140 249813 29142
rect 249747 29139 249813 29140
rect 249934 29069 249994 29142
rect 249931 29068 249997 29069
rect 249931 29004 249932 29068
rect 249996 29004 249997 29068
rect 249931 29003 249997 29004
rect 252804 2454 253404 37898
rect 252804 2218 252986 2454
rect 253222 2218 253404 2454
rect 252804 2134 253404 2218
rect 252804 1898 252986 2134
rect 253222 1898 253404 2134
rect 252804 -346 253404 1898
rect 252804 -582 252986 -346
rect 253222 -582 253404 -346
rect 252804 -666 253404 -582
rect 252804 -902 252986 -666
rect 253222 -902 253404 -666
rect 252804 -1844 253404 -902
rect 256404 690054 257004 706122
rect 256404 689818 256586 690054
rect 256822 689818 257004 690054
rect 256404 689734 257004 689818
rect 256404 689498 256586 689734
rect 256822 689498 257004 689734
rect 256404 654054 257004 689498
rect 256404 653818 256586 654054
rect 256822 653818 257004 654054
rect 256404 653734 257004 653818
rect 256404 653498 256586 653734
rect 256822 653498 257004 653734
rect 256404 618054 257004 653498
rect 256404 617818 256586 618054
rect 256822 617818 257004 618054
rect 256404 617734 257004 617818
rect 256404 617498 256586 617734
rect 256822 617498 257004 617734
rect 256404 582054 257004 617498
rect 256404 581818 256586 582054
rect 256822 581818 257004 582054
rect 256404 581734 257004 581818
rect 256404 581498 256586 581734
rect 256822 581498 257004 581734
rect 256404 546054 257004 581498
rect 256404 545818 256586 546054
rect 256822 545818 257004 546054
rect 256404 545734 257004 545818
rect 256404 545498 256586 545734
rect 256822 545498 257004 545734
rect 256404 510054 257004 545498
rect 256404 509818 256586 510054
rect 256822 509818 257004 510054
rect 256404 509734 257004 509818
rect 256404 509498 256586 509734
rect 256822 509498 257004 509734
rect 256404 474054 257004 509498
rect 256404 473818 256586 474054
rect 256822 473818 257004 474054
rect 256404 473734 257004 473818
rect 256404 473498 256586 473734
rect 256822 473498 257004 473734
rect 256404 438054 257004 473498
rect 256404 437818 256586 438054
rect 256822 437818 257004 438054
rect 256404 437734 257004 437818
rect 256404 437498 256586 437734
rect 256822 437498 257004 437734
rect 256404 402054 257004 437498
rect 256404 401818 256586 402054
rect 256822 401818 257004 402054
rect 256404 401734 257004 401818
rect 256404 401498 256586 401734
rect 256822 401498 257004 401734
rect 256404 366054 257004 401498
rect 256404 365818 256586 366054
rect 256822 365818 257004 366054
rect 256404 365734 257004 365818
rect 256404 365498 256586 365734
rect 256822 365498 257004 365734
rect 256404 330054 257004 365498
rect 256404 329818 256586 330054
rect 256822 329818 257004 330054
rect 256404 329734 257004 329818
rect 256404 329498 256586 329734
rect 256822 329498 257004 329734
rect 256404 294054 257004 329498
rect 260004 693654 260604 707962
rect 260004 693418 260186 693654
rect 260422 693418 260604 693654
rect 260004 693334 260604 693418
rect 260004 693098 260186 693334
rect 260422 693098 260604 693334
rect 260004 657654 260604 693098
rect 260004 657418 260186 657654
rect 260422 657418 260604 657654
rect 260004 657334 260604 657418
rect 260004 657098 260186 657334
rect 260422 657098 260604 657334
rect 260004 621654 260604 657098
rect 260004 621418 260186 621654
rect 260422 621418 260604 621654
rect 260004 621334 260604 621418
rect 260004 621098 260186 621334
rect 260422 621098 260604 621334
rect 260004 585654 260604 621098
rect 260004 585418 260186 585654
rect 260422 585418 260604 585654
rect 260004 585334 260604 585418
rect 260004 585098 260186 585334
rect 260422 585098 260604 585334
rect 260004 549654 260604 585098
rect 260004 549418 260186 549654
rect 260422 549418 260604 549654
rect 260004 549334 260604 549418
rect 260004 549098 260186 549334
rect 260422 549098 260604 549334
rect 260004 513654 260604 549098
rect 260004 513418 260186 513654
rect 260422 513418 260604 513654
rect 260004 513334 260604 513418
rect 260004 513098 260186 513334
rect 260422 513098 260604 513334
rect 260004 477654 260604 513098
rect 260004 477418 260186 477654
rect 260422 477418 260604 477654
rect 260004 477334 260604 477418
rect 260004 477098 260186 477334
rect 260422 477098 260604 477334
rect 260004 441654 260604 477098
rect 260004 441418 260186 441654
rect 260422 441418 260604 441654
rect 260004 441334 260604 441418
rect 260004 441098 260186 441334
rect 260422 441098 260604 441334
rect 260004 405654 260604 441098
rect 260004 405418 260186 405654
rect 260422 405418 260604 405654
rect 260004 405334 260604 405418
rect 260004 405098 260186 405334
rect 260422 405098 260604 405334
rect 260004 369654 260604 405098
rect 263604 697254 264204 709802
rect 281604 711278 282204 711300
rect 281604 711042 281786 711278
rect 282022 711042 282204 711278
rect 281604 710958 282204 711042
rect 281604 710722 281786 710958
rect 282022 710722 282204 710958
rect 278004 709438 278604 709460
rect 278004 709202 278186 709438
rect 278422 709202 278604 709438
rect 278004 709118 278604 709202
rect 278004 708882 278186 709118
rect 278422 708882 278604 709118
rect 274404 707598 275004 707620
rect 274404 707362 274586 707598
rect 274822 707362 275004 707598
rect 274404 707278 275004 707362
rect 274404 707042 274586 707278
rect 274822 707042 275004 707278
rect 263604 697018 263786 697254
rect 264022 697018 264204 697254
rect 263604 696934 264204 697018
rect 263604 696698 263786 696934
rect 264022 696698 264204 696934
rect 263604 661254 264204 696698
rect 263604 661018 263786 661254
rect 264022 661018 264204 661254
rect 263604 660934 264204 661018
rect 263604 660698 263786 660934
rect 264022 660698 264204 660934
rect 263604 625254 264204 660698
rect 263604 625018 263786 625254
rect 264022 625018 264204 625254
rect 263604 624934 264204 625018
rect 263604 624698 263786 624934
rect 264022 624698 264204 624934
rect 263604 589254 264204 624698
rect 263604 589018 263786 589254
rect 264022 589018 264204 589254
rect 263604 588934 264204 589018
rect 263604 588698 263786 588934
rect 264022 588698 264204 588934
rect 263604 553254 264204 588698
rect 263604 553018 263786 553254
rect 264022 553018 264204 553254
rect 263604 552934 264204 553018
rect 263604 552698 263786 552934
rect 264022 552698 264204 552934
rect 263604 517254 264204 552698
rect 263604 517018 263786 517254
rect 264022 517018 264204 517254
rect 263604 516934 264204 517018
rect 263604 516698 263786 516934
rect 264022 516698 264204 516934
rect 263604 481254 264204 516698
rect 263604 481018 263786 481254
rect 264022 481018 264204 481254
rect 263604 480934 264204 481018
rect 263604 480698 263786 480934
rect 264022 480698 264204 480934
rect 263604 445254 264204 480698
rect 263604 445018 263786 445254
rect 264022 445018 264204 445254
rect 263604 444934 264204 445018
rect 263604 444698 263786 444934
rect 264022 444698 264204 444934
rect 263604 409254 264204 444698
rect 263604 409018 263786 409254
rect 264022 409018 264204 409254
rect 263604 408934 264204 409018
rect 263604 408698 263786 408934
rect 264022 408698 264204 408934
rect 262811 401844 262877 401845
rect 262811 401780 262812 401844
rect 262876 401780 262877 401844
rect 262811 401779 262877 401780
rect 260004 369418 260186 369654
rect 260422 369418 260604 369654
rect 260004 369334 260604 369418
rect 260004 369098 260186 369334
rect 260422 369098 260604 369334
rect 260004 333654 260604 369098
rect 262814 336021 262874 401779
rect 263604 373254 264204 408698
rect 263604 373018 263786 373254
rect 264022 373018 264204 373254
rect 263604 372934 264204 373018
rect 263604 372698 263786 372934
rect 264022 372698 264204 372934
rect 263604 337254 264204 372698
rect 263604 337018 263786 337254
rect 264022 337018 264204 337254
rect 263604 336934 264204 337018
rect 263604 336698 263786 336934
rect 264022 336698 264204 336934
rect 262811 336020 262877 336021
rect 262811 335956 262812 336020
rect 262876 335956 262877 336020
rect 262811 335955 262877 335956
rect 260004 333418 260186 333654
rect 260422 333418 260604 333654
rect 260004 333334 260604 333418
rect 260004 333098 260186 333334
rect 260422 333098 260604 333334
rect 257843 310996 257909 310997
rect 257843 310932 257844 310996
rect 257908 310932 257909 310996
rect 257843 310931 257909 310932
rect 258027 310996 258093 310997
rect 258027 310932 258028 310996
rect 258092 310932 258093 310996
rect 258027 310931 258093 310932
rect 257846 310725 257906 310931
rect 258030 310725 258090 310931
rect 257843 310724 257909 310725
rect 257843 310660 257844 310724
rect 257908 310660 257909 310724
rect 257843 310659 257909 310660
rect 258027 310724 258093 310725
rect 258027 310660 258028 310724
rect 258092 310660 258093 310724
rect 258027 310659 258093 310660
rect 256404 293818 256586 294054
rect 256822 293818 257004 294054
rect 256404 293734 257004 293818
rect 256404 293498 256586 293734
rect 256822 293498 257004 293734
rect 256404 258054 257004 293498
rect 256404 257818 256586 258054
rect 256822 257818 257004 258054
rect 256404 257734 257004 257818
rect 256404 257498 256586 257734
rect 256822 257498 257004 257734
rect 256404 222054 257004 257498
rect 260004 297654 260604 333098
rect 260004 297418 260186 297654
rect 260422 297418 260604 297654
rect 260004 297334 260604 297418
rect 260004 297098 260186 297334
rect 260422 297098 260604 297334
rect 260004 261654 260604 297098
rect 260004 261418 260186 261654
rect 260422 261418 260604 261654
rect 260004 261334 260604 261418
rect 260004 261098 260186 261334
rect 260422 261098 260604 261334
rect 257843 228036 257909 228037
rect 257843 227972 257844 228036
rect 257908 227972 257909 228036
rect 257843 227971 257909 227972
rect 257846 227629 257906 227971
rect 257843 227628 257909 227629
rect 257843 227564 257844 227628
rect 257908 227564 257909 227628
rect 257843 227563 257909 227564
rect 256404 221818 256586 222054
rect 256822 221818 257004 222054
rect 256404 221734 257004 221818
rect 256404 221498 256586 221734
rect 256822 221498 257004 221734
rect 256404 186054 257004 221498
rect 256404 185818 256586 186054
rect 256822 185818 257004 186054
rect 256404 185734 257004 185818
rect 256404 185498 256586 185734
rect 256822 185498 257004 185734
rect 256404 150054 257004 185498
rect 256404 149818 256586 150054
rect 256822 149818 257004 150054
rect 256404 149734 257004 149818
rect 256404 149498 256586 149734
rect 256822 149498 257004 149734
rect 256404 114054 257004 149498
rect 256404 113818 256586 114054
rect 256822 113818 257004 114054
rect 256404 113734 257004 113818
rect 256404 113498 256586 113734
rect 256822 113498 257004 113734
rect 256404 78054 257004 113498
rect 256404 77818 256586 78054
rect 256822 77818 257004 78054
rect 256404 77734 257004 77818
rect 256404 77498 256586 77734
rect 256822 77498 257004 77734
rect 256404 42054 257004 77498
rect 256404 41818 256586 42054
rect 256822 41818 257004 42054
rect 256404 41734 257004 41818
rect 256404 41498 256586 41734
rect 256822 41498 257004 41734
rect 256404 6054 257004 41498
rect 256404 5818 256586 6054
rect 256822 5818 257004 6054
rect 256404 5734 257004 5818
rect 256404 5498 256586 5734
rect 256822 5498 257004 5734
rect 256404 -2186 257004 5498
rect 256404 -2422 256586 -2186
rect 256822 -2422 257004 -2186
rect 256404 -2506 257004 -2422
rect 256404 -2742 256586 -2506
rect 256822 -2742 257004 -2506
rect 256404 -3684 257004 -2742
rect 260004 225654 260604 261098
rect 260004 225418 260186 225654
rect 260422 225418 260604 225654
rect 260004 225334 260604 225418
rect 260004 225098 260186 225334
rect 260422 225098 260604 225334
rect 260004 189654 260604 225098
rect 260004 189418 260186 189654
rect 260422 189418 260604 189654
rect 260004 189334 260604 189418
rect 260004 189098 260186 189334
rect 260422 189098 260604 189334
rect 260004 153654 260604 189098
rect 260004 153418 260186 153654
rect 260422 153418 260604 153654
rect 260004 153334 260604 153418
rect 260004 153098 260186 153334
rect 260422 153098 260604 153334
rect 260004 117654 260604 153098
rect 260004 117418 260186 117654
rect 260422 117418 260604 117654
rect 260004 117334 260604 117418
rect 260004 117098 260186 117334
rect 260422 117098 260604 117334
rect 260004 81654 260604 117098
rect 260004 81418 260186 81654
rect 260422 81418 260604 81654
rect 260004 81334 260604 81418
rect 260004 81098 260186 81334
rect 260422 81098 260604 81334
rect 260004 45654 260604 81098
rect 263604 301254 264204 336698
rect 263604 301018 263786 301254
rect 264022 301018 264204 301254
rect 263604 300934 264204 301018
rect 263604 300698 263786 300934
rect 264022 300698 264204 300934
rect 263604 265254 264204 300698
rect 263604 265018 263786 265254
rect 264022 265018 264204 265254
rect 263604 264934 264204 265018
rect 263604 264698 263786 264934
rect 264022 264698 264204 264934
rect 263604 229254 264204 264698
rect 263604 229018 263786 229254
rect 264022 229018 264204 229254
rect 263604 228934 264204 229018
rect 263604 228698 263786 228934
rect 264022 228698 264204 228934
rect 263604 193254 264204 228698
rect 263604 193018 263786 193254
rect 264022 193018 264204 193254
rect 263604 192934 264204 193018
rect 263604 192698 263786 192934
rect 264022 192698 264204 192934
rect 263604 157254 264204 192698
rect 263604 157018 263786 157254
rect 264022 157018 264204 157254
rect 263604 156934 264204 157018
rect 263604 156698 263786 156934
rect 264022 156698 264204 156934
rect 263604 121254 264204 156698
rect 263604 121018 263786 121254
rect 264022 121018 264204 121254
rect 263604 120934 264204 121018
rect 263604 120698 263786 120934
rect 264022 120698 264204 120934
rect 263604 85254 264204 120698
rect 263604 85018 263786 85254
rect 264022 85018 264204 85254
rect 263604 84934 264204 85018
rect 263604 84698 263786 84934
rect 264022 84698 264204 84934
rect 260971 76124 261037 76125
rect 260971 76060 260972 76124
rect 261036 76060 261037 76124
rect 260971 76059 261037 76060
rect 260787 75988 260853 75989
rect 260787 75924 260788 75988
rect 260852 75924 260853 75988
rect 260787 75923 260853 75924
rect 260790 75850 260850 75923
rect 260974 75850 261034 76059
rect 260790 75790 261034 75850
rect 260004 45418 260186 45654
rect 260422 45418 260604 45654
rect 260004 45334 260604 45418
rect 260004 45098 260186 45334
rect 260422 45098 260604 45334
rect 260004 9654 260604 45098
rect 260004 9418 260186 9654
rect 260422 9418 260604 9654
rect 260004 9334 260604 9418
rect 260004 9098 260186 9334
rect 260422 9098 260604 9334
rect 260004 -4026 260604 9098
rect 260004 -4262 260186 -4026
rect 260422 -4262 260604 -4026
rect 260004 -4346 260604 -4262
rect 260004 -4582 260186 -4346
rect 260422 -4582 260604 -4346
rect 260004 -5524 260604 -4582
rect 263604 49254 264204 84698
rect 263604 49018 263786 49254
rect 264022 49018 264204 49254
rect 263604 48934 264204 49018
rect 263604 48698 263786 48934
rect 264022 48698 264204 48934
rect 263604 13254 264204 48698
rect 270804 705758 271404 705780
rect 270804 705522 270986 705758
rect 271222 705522 271404 705758
rect 270804 705438 271404 705522
rect 270804 705202 270986 705438
rect 271222 705202 271404 705438
rect 270804 668454 271404 705202
rect 270804 668218 270986 668454
rect 271222 668218 271404 668454
rect 270804 668134 271404 668218
rect 270804 667898 270986 668134
rect 271222 667898 271404 668134
rect 270804 632454 271404 667898
rect 270804 632218 270986 632454
rect 271222 632218 271404 632454
rect 270804 632134 271404 632218
rect 270804 631898 270986 632134
rect 271222 631898 271404 632134
rect 270804 596454 271404 631898
rect 270804 596218 270986 596454
rect 271222 596218 271404 596454
rect 270804 596134 271404 596218
rect 270804 595898 270986 596134
rect 271222 595898 271404 596134
rect 270804 560454 271404 595898
rect 270804 560218 270986 560454
rect 271222 560218 271404 560454
rect 270804 560134 271404 560218
rect 270804 559898 270986 560134
rect 271222 559898 271404 560134
rect 270804 524454 271404 559898
rect 270804 524218 270986 524454
rect 271222 524218 271404 524454
rect 270804 524134 271404 524218
rect 270804 523898 270986 524134
rect 271222 523898 271404 524134
rect 270804 488454 271404 523898
rect 270804 488218 270986 488454
rect 271222 488218 271404 488454
rect 270804 488134 271404 488218
rect 270804 487898 270986 488134
rect 271222 487898 271404 488134
rect 270804 452454 271404 487898
rect 270804 452218 270986 452454
rect 271222 452218 271404 452454
rect 270804 452134 271404 452218
rect 270804 451898 270986 452134
rect 271222 451898 271404 452134
rect 270804 416454 271404 451898
rect 270804 416218 270986 416454
rect 271222 416218 271404 416454
rect 270804 416134 271404 416218
rect 270804 415898 270986 416134
rect 271222 415898 271404 416134
rect 270804 380454 271404 415898
rect 270804 380218 270986 380454
rect 271222 380218 271404 380454
rect 270804 380134 271404 380218
rect 270804 379898 270986 380134
rect 271222 379898 271404 380134
rect 270804 344454 271404 379898
rect 270804 344218 270986 344454
rect 271222 344218 271404 344454
rect 270804 344134 271404 344218
rect 270804 343898 270986 344134
rect 271222 343898 271404 344134
rect 270804 308454 271404 343898
rect 270804 308218 270986 308454
rect 271222 308218 271404 308454
rect 270804 308134 271404 308218
rect 270804 307898 270986 308134
rect 271222 307898 271404 308134
rect 270804 272454 271404 307898
rect 270804 272218 270986 272454
rect 271222 272218 271404 272454
rect 270804 272134 271404 272218
rect 270804 271898 270986 272134
rect 271222 271898 271404 272134
rect 270804 236454 271404 271898
rect 270804 236218 270986 236454
rect 271222 236218 271404 236454
rect 270804 236134 271404 236218
rect 270804 235898 270986 236134
rect 271222 235898 271404 236134
rect 270804 200454 271404 235898
rect 270804 200218 270986 200454
rect 271222 200218 271404 200454
rect 270804 200134 271404 200218
rect 270804 199898 270986 200134
rect 271222 199898 271404 200134
rect 270804 164454 271404 199898
rect 270804 164218 270986 164454
rect 271222 164218 271404 164454
rect 270804 164134 271404 164218
rect 270804 163898 270986 164134
rect 271222 163898 271404 164134
rect 270804 128454 271404 163898
rect 270804 128218 270986 128454
rect 271222 128218 271404 128454
rect 270804 128134 271404 128218
rect 270804 127898 270986 128134
rect 271222 127898 271404 128134
rect 270804 92454 271404 127898
rect 270804 92218 270986 92454
rect 271222 92218 271404 92454
rect 270804 92134 271404 92218
rect 270804 91898 270986 92134
rect 271222 91898 271404 92134
rect 270804 56454 271404 91898
rect 270804 56218 270986 56454
rect 271222 56218 271404 56454
rect 270804 56134 271404 56218
rect 270804 55898 270986 56134
rect 271222 55898 271404 56134
rect 269067 29340 269133 29341
rect 269067 29276 269068 29340
rect 269132 29276 269133 29340
rect 269067 29275 269133 29276
rect 269070 29069 269130 29275
rect 269067 29068 269133 29069
rect 269067 29004 269068 29068
rect 269132 29004 269133 29068
rect 269067 29003 269133 29004
rect 263604 13018 263786 13254
rect 264022 13018 264204 13254
rect 263604 12934 264204 13018
rect 263604 12698 263786 12934
rect 264022 12698 264204 12934
rect 245604 -7022 245786 -6786
rect 246022 -7022 246204 -6786
rect 245604 -7106 246204 -7022
rect 245604 -7342 245786 -7106
rect 246022 -7342 246204 -7106
rect 245604 -7364 246204 -7342
rect 263604 -5866 264204 12698
rect 270804 20454 271404 55898
rect 270804 20218 270986 20454
rect 271222 20218 271404 20454
rect 270804 20134 271404 20218
rect 270804 19898 270986 20134
rect 271222 19898 271404 20134
rect 270804 -1266 271404 19898
rect 270804 -1502 270986 -1266
rect 271222 -1502 271404 -1266
rect 270804 -1586 271404 -1502
rect 270804 -1822 270986 -1586
rect 271222 -1822 271404 -1586
rect 270804 -1844 271404 -1822
rect 274404 672054 275004 707042
rect 274404 671818 274586 672054
rect 274822 671818 275004 672054
rect 274404 671734 275004 671818
rect 274404 671498 274586 671734
rect 274822 671498 275004 671734
rect 274404 636054 275004 671498
rect 274404 635818 274586 636054
rect 274822 635818 275004 636054
rect 274404 635734 275004 635818
rect 274404 635498 274586 635734
rect 274822 635498 275004 635734
rect 274404 600054 275004 635498
rect 274404 599818 274586 600054
rect 274822 599818 275004 600054
rect 274404 599734 275004 599818
rect 274404 599498 274586 599734
rect 274822 599498 275004 599734
rect 274404 564054 275004 599498
rect 274404 563818 274586 564054
rect 274822 563818 275004 564054
rect 274404 563734 275004 563818
rect 274404 563498 274586 563734
rect 274822 563498 275004 563734
rect 274404 528054 275004 563498
rect 274404 527818 274586 528054
rect 274822 527818 275004 528054
rect 274404 527734 275004 527818
rect 274404 527498 274586 527734
rect 274822 527498 275004 527734
rect 274404 492054 275004 527498
rect 274404 491818 274586 492054
rect 274822 491818 275004 492054
rect 274404 491734 275004 491818
rect 274404 491498 274586 491734
rect 274822 491498 275004 491734
rect 274404 456054 275004 491498
rect 274404 455818 274586 456054
rect 274822 455818 275004 456054
rect 274404 455734 275004 455818
rect 274404 455498 274586 455734
rect 274822 455498 275004 455734
rect 274404 420054 275004 455498
rect 274404 419818 274586 420054
rect 274822 419818 275004 420054
rect 274404 419734 275004 419818
rect 274404 419498 274586 419734
rect 274822 419498 275004 419734
rect 274404 384054 275004 419498
rect 274404 383818 274586 384054
rect 274822 383818 275004 384054
rect 274404 383734 275004 383818
rect 274404 383498 274586 383734
rect 274822 383498 275004 383734
rect 274404 348054 275004 383498
rect 274404 347818 274586 348054
rect 274822 347818 275004 348054
rect 274404 347734 275004 347818
rect 274404 347498 274586 347734
rect 274822 347498 275004 347734
rect 274404 312054 275004 347498
rect 278004 675654 278604 708882
rect 278004 675418 278186 675654
rect 278422 675418 278604 675654
rect 278004 675334 278604 675418
rect 278004 675098 278186 675334
rect 278422 675098 278604 675334
rect 278004 639654 278604 675098
rect 278004 639418 278186 639654
rect 278422 639418 278604 639654
rect 278004 639334 278604 639418
rect 278004 639098 278186 639334
rect 278422 639098 278604 639334
rect 278004 603654 278604 639098
rect 278004 603418 278186 603654
rect 278422 603418 278604 603654
rect 278004 603334 278604 603418
rect 278004 603098 278186 603334
rect 278422 603098 278604 603334
rect 278004 567654 278604 603098
rect 278004 567418 278186 567654
rect 278422 567418 278604 567654
rect 278004 567334 278604 567418
rect 278004 567098 278186 567334
rect 278422 567098 278604 567334
rect 278004 531654 278604 567098
rect 278004 531418 278186 531654
rect 278422 531418 278604 531654
rect 278004 531334 278604 531418
rect 278004 531098 278186 531334
rect 278422 531098 278604 531334
rect 278004 495654 278604 531098
rect 278004 495418 278186 495654
rect 278422 495418 278604 495654
rect 278004 495334 278604 495418
rect 278004 495098 278186 495334
rect 278422 495098 278604 495334
rect 278004 459654 278604 495098
rect 278004 459418 278186 459654
rect 278422 459418 278604 459654
rect 278004 459334 278604 459418
rect 278004 459098 278186 459334
rect 278422 459098 278604 459334
rect 278004 423654 278604 459098
rect 278004 423418 278186 423654
rect 278422 423418 278604 423654
rect 278004 423334 278604 423418
rect 278004 423098 278186 423334
rect 278422 423098 278604 423334
rect 278004 387654 278604 423098
rect 278004 387418 278186 387654
rect 278422 387418 278604 387654
rect 278004 387334 278604 387418
rect 278004 387098 278186 387334
rect 278422 387098 278604 387334
rect 278004 351654 278604 387098
rect 278004 351418 278186 351654
rect 278422 351418 278604 351654
rect 278004 351334 278604 351418
rect 278004 351098 278186 351334
rect 278422 351098 278604 351334
rect 275323 325684 275389 325685
rect 275323 325620 275324 325684
rect 275388 325620 275389 325684
rect 275323 325619 275389 325620
rect 275326 314941 275386 325619
rect 278004 315654 278604 351098
rect 278004 315418 278186 315654
rect 278422 315418 278604 315654
rect 278004 315334 278604 315418
rect 278004 315098 278186 315334
rect 278422 315098 278604 315334
rect 275323 314940 275389 314941
rect 275323 314876 275324 314940
rect 275388 314876 275389 314940
rect 275323 314875 275389 314876
rect 274404 311818 274586 312054
rect 274822 311818 275004 312054
rect 274404 311734 275004 311818
rect 274404 311498 274586 311734
rect 274822 311498 275004 311734
rect 274404 276054 275004 311498
rect 274404 275818 274586 276054
rect 274822 275818 275004 276054
rect 274404 275734 275004 275818
rect 274404 275498 274586 275734
rect 274822 275498 275004 275734
rect 274404 240054 275004 275498
rect 274404 239818 274586 240054
rect 274822 239818 275004 240054
rect 274404 239734 275004 239818
rect 274404 239498 274586 239734
rect 274822 239498 275004 239734
rect 274404 204054 275004 239498
rect 274404 203818 274586 204054
rect 274822 203818 275004 204054
rect 274404 203734 275004 203818
rect 274404 203498 274586 203734
rect 274822 203498 275004 203734
rect 274404 168054 275004 203498
rect 274404 167818 274586 168054
rect 274822 167818 275004 168054
rect 274404 167734 275004 167818
rect 274404 167498 274586 167734
rect 274822 167498 275004 167734
rect 274404 132054 275004 167498
rect 274404 131818 274586 132054
rect 274822 131818 275004 132054
rect 274404 131734 275004 131818
rect 274404 131498 274586 131734
rect 274822 131498 275004 131734
rect 274404 96054 275004 131498
rect 274404 95818 274586 96054
rect 274822 95818 275004 96054
rect 274404 95734 275004 95818
rect 274404 95498 274586 95734
rect 274822 95498 275004 95734
rect 274404 60054 275004 95498
rect 274404 59818 274586 60054
rect 274822 59818 275004 60054
rect 274404 59734 275004 59818
rect 274404 59498 274586 59734
rect 274822 59498 275004 59734
rect 274404 24054 275004 59498
rect 274404 23818 274586 24054
rect 274822 23818 275004 24054
rect 274404 23734 275004 23818
rect 274404 23498 274586 23734
rect 274822 23498 275004 23734
rect 274404 -3106 275004 23498
rect 274404 -3342 274586 -3106
rect 274822 -3342 275004 -3106
rect 274404 -3426 275004 -3342
rect 274404 -3662 274586 -3426
rect 274822 -3662 275004 -3426
rect 274404 -3684 275004 -3662
rect 278004 279654 278604 315098
rect 278004 279418 278186 279654
rect 278422 279418 278604 279654
rect 278004 279334 278604 279418
rect 278004 279098 278186 279334
rect 278422 279098 278604 279334
rect 278004 243654 278604 279098
rect 278004 243418 278186 243654
rect 278422 243418 278604 243654
rect 278004 243334 278604 243418
rect 278004 243098 278186 243334
rect 278422 243098 278604 243334
rect 278004 207654 278604 243098
rect 278004 207418 278186 207654
rect 278422 207418 278604 207654
rect 278004 207334 278604 207418
rect 278004 207098 278186 207334
rect 278422 207098 278604 207334
rect 278004 171654 278604 207098
rect 278004 171418 278186 171654
rect 278422 171418 278604 171654
rect 278004 171334 278604 171418
rect 278004 171098 278186 171334
rect 278422 171098 278604 171334
rect 278004 135654 278604 171098
rect 278004 135418 278186 135654
rect 278422 135418 278604 135654
rect 278004 135334 278604 135418
rect 278004 135098 278186 135334
rect 278422 135098 278604 135334
rect 278004 99654 278604 135098
rect 278004 99418 278186 99654
rect 278422 99418 278604 99654
rect 278004 99334 278604 99418
rect 278004 99098 278186 99334
rect 278422 99098 278604 99334
rect 278004 63654 278604 99098
rect 278004 63418 278186 63654
rect 278422 63418 278604 63654
rect 278004 63334 278604 63418
rect 278004 63098 278186 63334
rect 278422 63098 278604 63334
rect 278004 27654 278604 63098
rect 278004 27418 278186 27654
rect 278422 27418 278604 27654
rect 278004 27334 278604 27418
rect 278004 27098 278186 27334
rect 278422 27098 278604 27334
rect 278004 -4946 278604 27098
rect 278004 -5182 278186 -4946
rect 278422 -5182 278604 -4946
rect 278004 -5266 278604 -5182
rect 278004 -5502 278186 -5266
rect 278422 -5502 278604 -5266
rect 278004 -5524 278604 -5502
rect 281604 679254 282204 710722
rect 299604 710358 300204 711300
rect 299604 710122 299786 710358
rect 300022 710122 300204 710358
rect 299604 710038 300204 710122
rect 299604 709802 299786 710038
rect 300022 709802 300204 710038
rect 296004 708518 296604 709460
rect 296004 708282 296186 708518
rect 296422 708282 296604 708518
rect 296004 708198 296604 708282
rect 296004 707962 296186 708198
rect 296422 707962 296604 708198
rect 292404 706678 293004 707620
rect 292404 706442 292586 706678
rect 292822 706442 293004 706678
rect 292404 706358 293004 706442
rect 292404 706122 292586 706358
rect 292822 706122 293004 706358
rect 281604 679018 281786 679254
rect 282022 679018 282204 679254
rect 281604 678934 282204 679018
rect 281604 678698 281786 678934
rect 282022 678698 282204 678934
rect 281604 643254 282204 678698
rect 281604 643018 281786 643254
rect 282022 643018 282204 643254
rect 281604 642934 282204 643018
rect 281604 642698 281786 642934
rect 282022 642698 282204 642934
rect 281604 607254 282204 642698
rect 281604 607018 281786 607254
rect 282022 607018 282204 607254
rect 281604 606934 282204 607018
rect 281604 606698 281786 606934
rect 282022 606698 282204 606934
rect 281604 571254 282204 606698
rect 281604 571018 281786 571254
rect 282022 571018 282204 571254
rect 281604 570934 282204 571018
rect 281604 570698 281786 570934
rect 282022 570698 282204 570934
rect 281604 535254 282204 570698
rect 281604 535018 281786 535254
rect 282022 535018 282204 535254
rect 281604 534934 282204 535018
rect 281604 534698 281786 534934
rect 282022 534698 282204 534934
rect 281604 499254 282204 534698
rect 281604 499018 281786 499254
rect 282022 499018 282204 499254
rect 281604 498934 282204 499018
rect 281604 498698 281786 498934
rect 282022 498698 282204 498934
rect 281604 463254 282204 498698
rect 281604 463018 281786 463254
rect 282022 463018 282204 463254
rect 281604 462934 282204 463018
rect 281604 462698 281786 462934
rect 282022 462698 282204 462934
rect 281604 427254 282204 462698
rect 281604 427018 281786 427254
rect 282022 427018 282204 427254
rect 281604 426934 282204 427018
rect 281604 426698 281786 426934
rect 282022 426698 282204 426934
rect 281604 391254 282204 426698
rect 288804 704838 289404 705780
rect 288804 704602 288986 704838
rect 289222 704602 289404 704838
rect 288804 704518 289404 704602
rect 288804 704282 288986 704518
rect 289222 704282 289404 704518
rect 288804 686454 289404 704282
rect 288804 686218 288986 686454
rect 289222 686218 289404 686454
rect 288804 686134 289404 686218
rect 288804 685898 288986 686134
rect 289222 685898 289404 686134
rect 288804 650454 289404 685898
rect 288804 650218 288986 650454
rect 289222 650218 289404 650454
rect 288804 650134 289404 650218
rect 288804 649898 288986 650134
rect 289222 649898 289404 650134
rect 288804 614454 289404 649898
rect 288804 614218 288986 614454
rect 289222 614218 289404 614454
rect 288804 614134 289404 614218
rect 288804 613898 288986 614134
rect 289222 613898 289404 614134
rect 288804 578454 289404 613898
rect 288804 578218 288986 578454
rect 289222 578218 289404 578454
rect 288804 578134 289404 578218
rect 288804 577898 288986 578134
rect 289222 577898 289404 578134
rect 288804 542454 289404 577898
rect 288804 542218 288986 542454
rect 289222 542218 289404 542454
rect 288804 542134 289404 542218
rect 288804 541898 288986 542134
rect 289222 541898 289404 542134
rect 288804 506454 289404 541898
rect 288804 506218 288986 506454
rect 289222 506218 289404 506454
rect 288804 506134 289404 506218
rect 288804 505898 288986 506134
rect 289222 505898 289404 506134
rect 288804 470454 289404 505898
rect 288804 470218 288986 470454
rect 289222 470218 289404 470454
rect 288804 470134 289404 470218
rect 288804 469898 288986 470134
rect 289222 469898 289404 470134
rect 288804 434454 289404 469898
rect 288804 434218 288986 434454
rect 289222 434218 289404 434454
rect 288804 434134 289404 434218
rect 288804 433898 288986 434134
rect 289222 433898 289404 434134
rect 282867 399396 282933 399397
rect 282867 399332 282868 399396
rect 282932 399332 282933 399396
rect 282867 399331 282933 399332
rect 284339 399396 284405 399397
rect 284339 399332 284340 399396
rect 284404 399332 284405 399396
rect 284339 399331 284405 399332
rect 285627 399396 285693 399397
rect 285627 399332 285628 399396
rect 285692 399332 285693 399396
rect 285627 399331 285693 399332
rect 287099 399396 287165 399397
rect 287099 399332 287100 399396
rect 287164 399332 287165 399396
rect 287099 399331 287165 399332
rect 281604 391018 281786 391254
rect 282022 391018 282204 391254
rect 281604 390934 282204 391018
rect 281604 390698 281786 390934
rect 282022 390698 282204 390934
rect 281604 355254 282204 390698
rect 281604 355018 281786 355254
rect 282022 355018 282204 355254
rect 281604 354934 282204 355018
rect 281604 354698 281786 354934
rect 282022 354698 282204 354934
rect 281604 319254 282204 354698
rect 281604 319018 281786 319254
rect 282022 319018 282204 319254
rect 281604 318934 282204 319018
rect 281604 318698 281786 318934
rect 282022 318698 282204 318934
rect 281604 283254 282204 318698
rect 281604 283018 281786 283254
rect 282022 283018 282204 283254
rect 281604 282934 282204 283018
rect 281604 282698 281786 282934
rect 282022 282698 282204 282934
rect 281604 247254 282204 282698
rect 281604 247018 281786 247254
rect 282022 247018 282204 247254
rect 281604 246934 282204 247018
rect 281604 246698 281786 246934
rect 282022 246698 282204 246934
rect 281604 211254 282204 246698
rect 281604 211018 281786 211254
rect 282022 211018 282204 211254
rect 281604 210934 282204 211018
rect 281604 210698 281786 210934
rect 282022 210698 282204 210934
rect 281604 175254 282204 210698
rect 282870 194581 282930 399331
rect 282867 194580 282933 194581
rect 282867 194516 282868 194580
rect 282932 194516 282933 194580
rect 282867 194515 282933 194516
rect 281604 175018 281786 175254
rect 282022 175018 282204 175254
rect 281604 174934 282204 175018
rect 281604 174698 281786 174934
rect 282022 174698 282204 174934
rect 281604 139254 282204 174698
rect 284342 151741 284402 399331
rect 284339 151740 284405 151741
rect 284339 151676 284340 151740
rect 284404 151676 284405 151740
rect 284339 151675 284405 151676
rect 281604 139018 281786 139254
rect 282022 139018 282204 139254
rect 281604 138934 282204 139018
rect 281604 138698 281786 138934
rect 282022 138698 282204 138934
rect 281604 103254 282204 138698
rect 285630 109037 285690 399331
rect 285627 109036 285693 109037
rect 285627 108972 285628 109036
rect 285692 108972 285693 109036
rect 285627 108971 285693 108972
rect 281604 103018 281786 103254
rect 282022 103018 282204 103254
rect 281604 102934 282204 103018
rect 281604 102698 281786 102934
rect 282022 102698 282204 102934
rect 281604 67254 282204 102698
rect 281604 67018 281786 67254
rect 282022 67018 282204 67254
rect 281604 66934 282204 67018
rect 281604 66698 281786 66934
rect 282022 66698 282204 66934
rect 281604 31254 282204 66698
rect 287102 64837 287162 399331
rect 288804 398454 289404 433898
rect 288804 398218 288986 398454
rect 289222 398218 289404 398454
rect 288804 398134 289404 398218
rect 288804 397898 288986 398134
rect 289222 397898 289404 398134
rect 288804 362454 289404 397898
rect 288804 362218 288986 362454
rect 289222 362218 289404 362454
rect 288804 362134 289404 362218
rect 288804 361898 288986 362134
rect 289222 361898 289404 362134
rect 288804 326454 289404 361898
rect 288804 326218 288986 326454
rect 289222 326218 289404 326454
rect 288804 326134 289404 326218
rect 288804 325898 288986 326134
rect 289222 325898 289404 326134
rect 288804 290454 289404 325898
rect 288804 290218 288986 290454
rect 289222 290218 289404 290454
rect 288804 290134 289404 290218
rect 288804 289898 288986 290134
rect 289222 289898 289404 290134
rect 288804 254454 289404 289898
rect 288804 254218 288986 254454
rect 289222 254218 289404 254454
rect 288804 254134 289404 254218
rect 288804 253898 288986 254134
rect 289222 253898 289404 254134
rect 288804 218454 289404 253898
rect 288804 218218 288986 218454
rect 289222 218218 289404 218454
rect 288804 218134 289404 218218
rect 288804 217898 288986 218134
rect 289222 217898 289404 218134
rect 288804 182454 289404 217898
rect 288804 182218 288986 182454
rect 289222 182218 289404 182454
rect 288804 182134 289404 182218
rect 288804 181898 288986 182134
rect 289222 181898 289404 182134
rect 288804 146454 289404 181898
rect 288804 146218 288986 146454
rect 289222 146218 289404 146454
rect 288804 146134 289404 146218
rect 288804 145898 288986 146134
rect 289222 145898 289404 146134
rect 288804 110454 289404 145898
rect 288804 110218 288986 110454
rect 289222 110218 289404 110454
rect 288804 110134 289404 110218
rect 288804 109898 288986 110134
rect 289222 109898 289404 110134
rect 288804 74454 289404 109898
rect 288804 74218 288986 74454
rect 289222 74218 289404 74454
rect 288804 74134 289404 74218
rect 288804 73898 288986 74134
rect 289222 73898 289404 74134
rect 287099 64836 287165 64837
rect 287099 64772 287100 64836
rect 287164 64772 287165 64836
rect 287099 64771 287165 64772
rect 281604 31018 281786 31254
rect 282022 31018 282204 31254
rect 281604 30934 282204 31018
rect 281604 30698 281786 30934
rect 282022 30698 282204 30934
rect 263604 -6102 263786 -5866
rect 264022 -6102 264204 -5866
rect 263604 -6186 264204 -6102
rect 263604 -6422 263786 -6186
rect 264022 -6422 264204 -6186
rect 263604 -7364 264204 -6422
rect 281604 -6786 282204 30698
rect 288804 38454 289404 73898
rect 288804 38218 288986 38454
rect 289222 38218 289404 38454
rect 288804 38134 289404 38218
rect 288804 37898 288986 38134
rect 289222 37898 289404 38134
rect 288804 2454 289404 37898
rect 288804 2218 288986 2454
rect 289222 2218 289404 2454
rect 288804 2134 289404 2218
rect 288804 1898 288986 2134
rect 289222 1898 289404 2134
rect 288804 -346 289404 1898
rect 288804 -582 288986 -346
rect 289222 -582 289404 -346
rect 288804 -666 289404 -582
rect 288804 -902 288986 -666
rect 289222 -902 289404 -666
rect 288804 -1844 289404 -902
rect 292404 690054 293004 706122
rect 292404 689818 292586 690054
rect 292822 689818 293004 690054
rect 292404 689734 293004 689818
rect 292404 689498 292586 689734
rect 292822 689498 293004 689734
rect 292404 654054 293004 689498
rect 292404 653818 292586 654054
rect 292822 653818 293004 654054
rect 292404 653734 293004 653818
rect 292404 653498 292586 653734
rect 292822 653498 293004 653734
rect 292404 618054 293004 653498
rect 292404 617818 292586 618054
rect 292822 617818 293004 618054
rect 292404 617734 293004 617818
rect 292404 617498 292586 617734
rect 292822 617498 293004 617734
rect 292404 582054 293004 617498
rect 292404 581818 292586 582054
rect 292822 581818 293004 582054
rect 292404 581734 293004 581818
rect 292404 581498 292586 581734
rect 292822 581498 293004 581734
rect 292404 546054 293004 581498
rect 292404 545818 292586 546054
rect 292822 545818 293004 546054
rect 292404 545734 293004 545818
rect 292404 545498 292586 545734
rect 292822 545498 293004 545734
rect 292404 510054 293004 545498
rect 292404 509818 292586 510054
rect 292822 509818 293004 510054
rect 292404 509734 293004 509818
rect 292404 509498 292586 509734
rect 292822 509498 293004 509734
rect 292404 474054 293004 509498
rect 292404 473818 292586 474054
rect 292822 473818 293004 474054
rect 292404 473734 293004 473818
rect 292404 473498 292586 473734
rect 292822 473498 293004 473734
rect 292404 438054 293004 473498
rect 292404 437818 292586 438054
rect 292822 437818 293004 438054
rect 292404 437734 293004 437818
rect 292404 437498 292586 437734
rect 292822 437498 293004 437734
rect 292404 402054 293004 437498
rect 292404 401818 292586 402054
rect 292822 401818 293004 402054
rect 292404 401734 293004 401818
rect 292404 401498 292586 401734
rect 292822 401498 293004 401734
rect 292404 366054 293004 401498
rect 292404 365818 292586 366054
rect 292822 365818 293004 366054
rect 292404 365734 293004 365818
rect 292404 365498 292586 365734
rect 292822 365498 293004 365734
rect 292404 330054 293004 365498
rect 292404 329818 292586 330054
rect 292822 329818 293004 330054
rect 292404 329734 293004 329818
rect 292404 329498 292586 329734
rect 292822 329498 293004 329734
rect 292404 294054 293004 329498
rect 292404 293818 292586 294054
rect 292822 293818 293004 294054
rect 292404 293734 293004 293818
rect 292404 293498 292586 293734
rect 292822 293498 293004 293734
rect 292404 258054 293004 293498
rect 292404 257818 292586 258054
rect 292822 257818 293004 258054
rect 292404 257734 293004 257818
rect 292404 257498 292586 257734
rect 292822 257498 293004 257734
rect 292404 222054 293004 257498
rect 292404 221818 292586 222054
rect 292822 221818 293004 222054
rect 292404 221734 293004 221818
rect 292404 221498 292586 221734
rect 292822 221498 293004 221734
rect 292404 186054 293004 221498
rect 292404 185818 292586 186054
rect 292822 185818 293004 186054
rect 292404 185734 293004 185818
rect 292404 185498 292586 185734
rect 292822 185498 293004 185734
rect 292404 150054 293004 185498
rect 292404 149818 292586 150054
rect 292822 149818 293004 150054
rect 292404 149734 293004 149818
rect 292404 149498 292586 149734
rect 292822 149498 293004 149734
rect 292404 114054 293004 149498
rect 292404 113818 292586 114054
rect 292822 113818 293004 114054
rect 292404 113734 293004 113818
rect 292404 113498 292586 113734
rect 292822 113498 293004 113734
rect 292404 78054 293004 113498
rect 292404 77818 292586 78054
rect 292822 77818 293004 78054
rect 292404 77734 293004 77818
rect 292404 77498 292586 77734
rect 292822 77498 293004 77734
rect 292404 42054 293004 77498
rect 292404 41818 292586 42054
rect 292822 41818 293004 42054
rect 292404 41734 293004 41818
rect 292404 41498 292586 41734
rect 292822 41498 293004 41734
rect 292404 6054 293004 41498
rect 292404 5818 292586 6054
rect 292822 5818 293004 6054
rect 292404 5734 293004 5818
rect 292404 5498 292586 5734
rect 292822 5498 293004 5734
rect 292404 -2186 293004 5498
rect 292404 -2422 292586 -2186
rect 292822 -2422 293004 -2186
rect 292404 -2506 293004 -2422
rect 292404 -2742 292586 -2506
rect 292822 -2742 293004 -2506
rect 292404 -3684 293004 -2742
rect 296004 693654 296604 707962
rect 296004 693418 296186 693654
rect 296422 693418 296604 693654
rect 296004 693334 296604 693418
rect 296004 693098 296186 693334
rect 296422 693098 296604 693334
rect 296004 657654 296604 693098
rect 296004 657418 296186 657654
rect 296422 657418 296604 657654
rect 296004 657334 296604 657418
rect 296004 657098 296186 657334
rect 296422 657098 296604 657334
rect 296004 621654 296604 657098
rect 296004 621418 296186 621654
rect 296422 621418 296604 621654
rect 296004 621334 296604 621418
rect 296004 621098 296186 621334
rect 296422 621098 296604 621334
rect 296004 585654 296604 621098
rect 296004 585418 296186 585654
rect 296422 585418 296604 585654
rect 296004 585334 296604 585418
rect 296004 585098 296186 585334
rect 296422 585098 296604 585334
rect 296004 549654 296604 585098
rect 296004 549418 296186 549654
rect 296422 549418 296604 549654
rect 296004 549334 296604 549418
rect 296004 549098 296186 549334
rect 296422 549098 296604 549334
rect 296004 513654 296604 549098
rect 296004 513418 296186 513654
rect 296422 513418 296604 513654
rect 296004 513334 296604 513418
rect 296004 513098 296186 513334
rect 296422 513098 296604 513334
rect 296004 477654 296604 513098
rect 296004 477418 296186 477654
rect 296422 477418 296604 477654
rect 296004 477334 296604 477418
rect 296004 477098 296186 477334
rect 296422 477098 296604 477334
rect 296004 441654 296604 477098
rect 296004 441418 296186 441654
rect 296422 441418 296604 441654
rect 296004 441334 296604 441418
rect 296004 441098 296186 441334
rect 296422 441098 296604 441334
rect 296004 405654 296604 441098
rect 296004 405418 296186 405654
rect 296422 405418 296604 405654
rect 296004 405334 296604 405418
rect 296004 405098 296186 405334
rect 296422 405098 296604 405334
rect 296004 369654 296604 405098
rect 296004 369418 296186 369654
rect 296422 369418 296604 369654
rect 296004 369334 296604 369418
rect 296004 369098 296186 369334
rect 296422 369098 296604 369334
rect 296004 333654 296604 369098
rect 296004 333418 296186 333654
rect 296422 333418 296604 333654
rect 296004 333334 296604 333418
rect 296004 333098 296186 333334
rect 296422 333098 296604 333334
rect 296004 297654 296604 333098
rect 299604 697254 300204 709802
rect 317604 711278 318204 711300
rect 317604 711042 317786 711278
rect 318022 711042 318204 711278
rect 317604 710958 318204 711042
rect 317604 710722 317786 710958
rect 318022 710722 318204 710958
rect 314004 709438 314604 709460
rect 314004 709202 314186 709438
rect 314422 709202 314604 709438
rect 314004 709118 314604 709202
rect 314004 708882 314186 709118
rect 314422 708882 314604 709118
rect 310404 707598 311004 707620
rect 310404 707362 310586 707598
rect 310822 707362 311004 707598
rect 310404 707278 311004 707362
rect 310404 707042 310586 707278
rect 310822 707042 311004 707278
rect 299604 697018 299786 697254
rect 300022 697018 300204 697254
rect 299604 696934 300204 697018
rect 299604 696698 299786 696934
rect 300022 696698 300204 696934
rect 299604 661254 300204 696698
rect 299604 661018 299786 661254
rect 300022 661018 300204 661254
rect 299604 660934 300204 661018
rect 299604 660698 299786 660934
rect 300022 660698 300204 660934
rect 299604 625254 300204 660698
rect 299604 625018 299786 625254
rect 300022 625018 300204 625254
rect 299604 624934 300204 625018
rect 299604 624698 299786 624934
rect 300022 624698 300204 624934
rect 299604 589254 300204 624698
rect 299604 589018 299786 589254
rect 300022 589018 300204 589254
rect 299604 588934 300204 589018
rect 299604 588698 299786 588934
rect 300022 588698 300204 588934
rect 299604 553254 300204 588698
rect 299604 553018 299786 553254
rect 300022 553018 300204 553254
rect 299604 552934 300204 553018
rect 299604 552698 299786 552934
rect 300022 552698 300204 552934
rect 299604 517254 300204 552698
rect 299604 517018 299786 517254
rect 300022 517018 300204 517254
rect 299604 516934 300204 517018
rect 299604 516698 299786 516934
rect 300022 516698 300204 516934
rect 299604 481254 300204 516698
rect 299604 481018 299786 481254
rect 300022 481018 300204 481254
rect 299604 480934 300204 481018
rect 299604 480698 299786 480934
rect 300022 480698 300204 480934
rect 299604 445254 300204 480698
rect 299604 445018 299786 445254
rect 300022 445018 300204 445254
rect 299604 444934 300204 445018
rect 299604 444698 299786 444934
rect 300022 444698 300204 444934
rect 299604 409254 300204 444698
rect 299604 409018 299786 409254
rect 300022 409018 300204 409254
rect 299604 408934 300204 409018
rect 299604 408698 299786 408934
rect 300022 408698 300204 408934
rect 299604 373254 300204 408698
rect 299604 373018 299786 373254
rect 300022 373018 300204 373254
rect 299604 372934 300204 373018
rect 299604 372698 299786 372934
rect 300022 372698 300204 372934
rect 299604 337254 300204 372698
rect 299604 337018 299786 337254
rect 300022 337018 300204 337254
rect 299604 336934 300204 337018
rect 299604 336698 299786 336934
rect 300022 336698 300204 336934
rect 299427 322148 299493 322149
rect 299427 322084 299428 322148
rect 299492 322084 299493 322148
rect 299427 322083 299493 322084
rect 299430 321741 299490 322083
rect 299427 321740 299493 321741
rect 299427 321676 299428 321740
rect 299492 321676 299493 321740
rect 299427 321675 299493 321676
rect 296004 297418 296186 297654
rect 296422 297418 296604 297654
rect 296004 297334 296604 297418
rect 296004 297098 296186 297334
rect 296422 297098 296604 297334
rect 296004 261654 296604 297098
rect 296004 261418 296186 261654
rect 296422 261418 296604 261654
rect 296004 261334 296604 261418
rect 296004 261098 296186 261334
rect 296422 261098 296604 261334
rect 296004 225654 296604 261098
rect 296004 225418 296186 225654
rect 296422 225418 296604 225654
rect 296004 225334 296604 225418
rect 296004 225098 296186 225334
rect 296422 225098 296604 225334
rect 296004 189654 296604 225098
rect 296004 189418 296186 189654
rect 296422 189418 296604 189654
rect 296004 189334 296604 189418
rect 296004 189098 296186 189334
rect 296422 189098 296604 189334
rect 296004 153654 296604 189098
rect 296004 153418 296186 153654
rect 296422 153418 296604 153654
rect 296004 153334 296604 153418
rect 296004 153098 296186 153334
rect 296422 153098 296604 153334
rect 296004 117654 296604 153098
rect 296004 117418 296186 117654
rect 296422 117418 296604 117654
rect 296004 117334 296604 117418
rect 296004 117098 296186 117334
rect 296422 117098 296604 117334
rect 296004 81654 296604 117098
rect 296004 81418 296186 81654
rect 296422 81418 296604 81654
rect 296004 81334 296604 81418
rect 296004 81098 296186 81334
rect 296422 81098 296604 81334
rect 296004 45654 296604 81098
rect 296004 45418 296186 45654
rect 296422 45418 296604 45654
rect 296004 45334 296604 45418
rect 296004 45098 296186 45334
rect 296422 45098 296604 45334
rect 296004 9654 296604 45098
rect 296004 9418 296186 9654
rect 296422 9418 296604 9654
rect 296004 9334 296604 9418
rect 296004 9098 296186 9334
rect 296422 9098 296604 9334
rect 296004 -4026 296604 9098
rect 296004 -4262 296186 -4026
rect 296422 -4262 296604 -4026
rect 296004 -4346 296604 -4262
rect 296004 -4582 296186 -4346
rect 296422 -4582 296604 -4346
rect 296004 -5524 296604 -4582
rect 299604 301254 300204 336698
rect 299604 301018 299786 301254
rect 300022 301018 300204 301254
rect 299604 300934 300204 301018
rect 299604 300698 299786 300934
rect 300022 300698 300204 300934
rect 299604 265254 300204 300698
rect 299604 265018 299786 265254
rect 300022 265018 300204 265254
rect 299604 264934 300204 265018
rect 299604 264698 299786 264934
rect 300022 264698 300204 264934
rect 299604 229254 300204 264698
rect 299604 229018 299786 229254
rect 300022 229018 300204 229254
rect 299604 228934 300204 229018
rect 299604 228698 299786 228934
rect 300022 228698 300204 228934
rect 299604 193254 300204 228698
rect 299604 193018 299786 193254
rect 300022 193018 300204 193254
rect 299604 192934 300204 193018
rect 299604 192698 299786 192934
rect 300022 192698 300204 192934
rect 299604 157254 300204 192698
rect 299604 157018 299786 157254
rect 300022 157018 300204 157254
rect 299604 156934 300204 157018
rect 299604 156698 299786 156934
rect 300022 156698 300204 156934
rect 299604 121254 300204 156698
rect 299604 121018 299786 121254
rect 300022 121018 300204 121254
rect 299604 120934 300204 121018
rect 299604 120698 299786 120934
rect 300022 120698 300204 120934
rect 299604 85254 300204 120698
rect 299604 85018 299786 85254
rect 300022 85018 300204 85254
rect 299604 84934 300204 85018
rect 299604 84698 299786 84934
rect 300022 84698 300204 84934
rect 299604 49254 300204 84698
rect 299604 49018 299786 49254
rect 300022 49018 300204 49254
rect 299604 48934 300204 49018
rect 299604 48698 299786 48934
rect 300022 48698 300204 48934
rect 299604 13254 300204 48698
rect 299604 13018 299786 13254
rect 300022 13018 300204 13254
rect 299604 12934 300204 13018
rect 299604 12698 299786 12934
rect 300022 12698 300204 12934
rect 281604 -7022 281786 -6786
rect 282022 -7022 282204 -6786
rect 281604 -7106 282204 -7022
rect 281604 -7342 281786 -7106
rect 282022 -7342 282204 -7106
rect 281604 -7364 282204 -7342
rect 299604 -5866 300204 12698
rect 306804 705758 307404 705780
rect 306804 705522 306986 705758
rect 307222 705522 307404 705758
rect 306804 705438 307404 705522
rect 306804 705202 306986 705438
rect 307222 705202 307404 705438
rect 306804 668454 307404 705202
rect 306804 668218 306986 668454
rect 307222 668218 307404 668454
rect 306804 668134 307404 668218
rect 306804 667898 306986 668134
rect 307222 667898 307404 668134
rect 306804 632454 307404 667898
rect 306804 632218 306986 632454
rect 307222 632218 307404 632454
rect 306804 632134 307404 632218
rect 306804 631898 306986 632134
rect 307222 631898 307404 632134
rect 306804 596454 307404 631898
rect 306804 596218 306986 596454
rect 307222 596218 307404 596454
rect 306804 596134 307404 596218
rect 306804 595898 306986 596134
rect 307222 595898 307404 596134
rect 306804 560454 307404 595898
rect 306804 560218 306986 560454
rect 307222 560218 307404 560454
rect 306804 560134 307404 560218
rect 306804 559898 306986 560134
rect 307222 559898 307404 560134
rect 306804 524454 307404 559898
rect 306804 524218 306986 524454
rect 307222 524218 307404 524454
rect 306804 524134 307404 524218
rect 306804 523898 306986 524134
rect 307222 523898 307404 524134
rect 306804 488454 307404 523898
rect 306804 488218 306986 488454
rect 307222 488218 307404 488454
rect 306804 488134 307404 488218
rect 306804 487898 306986 488134
rect 307222 487898 307404 488134
rect 306804 452454 307404 487898
rect 306804 452218 306986 452454
rect 307222 452218 307404 452454
rect 306804 452134 307404 452218
rect 306804 451898 306986 452134
rect 307222 451898 307404 452134
rect 306804 416454 307404 451898
rect 306804 416218 306986 416454
rect 307222 416218 307404 416454
rect 306804 416134 307404 416218
rect 306804 415898 306986 416134
rect 307222 415898 307404 416134
rect 306804 380454 307404 415898
rect 306804 380218 306986 380454
rect 307222 380218 307404 380454
rect 306804 380134 307404 380218
rect 306804 379898 306986 380134
rect 307222 379898 307404 380134
rect 306804 344454 307404 379898
rect 306804 344218 306986 344454
rect 307222 344218 307404 344454
rect 306804 344134 307404 344218
rect 306804 343898 306986 344134
rect 307222 343898 307404 344134
rect 306804 308454 307404 343898
rect 306804 308218 306986 308454
rect 307222 308218 307404 308454
rect 306804 308134 307404 308218
rect 306804 307898 306986 308134
rect 307222 307898 307404 308134
rect 306804 272454 307404 307898
rect 306804 272218 306986 272454
rect 307222 272218 307404 272454
rect 306804 272134 307404 272218
rect 306804 271898 306986 272134
rect 307222 271898 307404 272134
rect 306804 236454 307404 271898
rect 306804 236218 306986 236454
rect 307222 236218 307404 236454
rect 306804 236134 307404 236218
rect 306804 235898 306986 236134
rect 307222 235898 307404 236134
rect 306804 200454 307404 235898
rect 306804 200218 306986 200454
rect 307222 200218 307404 200454
rect 306804 200134 307404 200218
rect 306804 199898 306986 200134
rect 307222 199898 307404 200134
rect 306804 164454 307404 199898
rect 306804 164218 306986 164454
rect 307222 164218 307404 164454
rect 306804 164134 307404 164218
rect 306804 163898 306986 164134
rect 307222 163898 307404 164134
rect 306804 128454 307404 163898
rect 306804 128218 306986 128454
rect 307222 128218 307404 128454
rect 306804 128134 307404 128218
rect 306804 127898 306986 128134
rect 307222 127898 307404 128134
rect 306804 92454 307404 127898
rect 306804 92218 306986 92454
rect 307222 92218 307404 92454
rect 306804 92134 307404 92218
rect 306804 91898 306986 92134
rect 307222 91898 307404 92134
rect 306804 56454 307404 91898
rect 306804 56218 306986 56454
rect 307222 56218 307404 56454
rect 306804 56134 307404 56218
rect 306804 55898 306986 56134
rect 307222 55898 307404 56134
rect 306804 20454 307404 55898
rect 306804 20218 306986 20454
rect 307222 20218 307404 20454
rect 306804 20134 307404 20218
rect 306804 19898 306986 20134
rect 307222 19898 307404 20134
rect 306804 -1266 307404 19898
rect 306804 -1502 306986 -1266
rect 307222 -1502 307404 -1266
rect 306804 -1586 307404 -1502
rect 306804 -1822 306986 -1586
rect 307222 -1822 307404 -1586
rect 306804 -1844 307404 -1822
rect 310404 672054 311004 707042
rect 310404 671818 310586 672054
rect 310822 671818 311004 672054
rect 310404 671734 311004 671818
rect 310404 671498 310586 671734
rect 310822 671498 311004 671734
rect 310404 636054 311004 671498
rect 310404 635818 310586 636054
rect 310822 635818 311004 636054
rect 310404 635734 311004 635818
rect 310404 635498 310586 635734
rect 310822 635498 311004 635734
rect 310404 600054 311004 635498
rect 310404 599818 310586 600054
rect 310822 599818 311004 600054
rect 310404 599734 311004 599818
rect 310404 599498 310586 599734
rect 310822 599498 311004 599734
rect 310404 564054 311004 599498
rect 310404 563818 310586 564054
rect 310822 563818 311004 564054
rect 310404 563734 311004 563818
rect 310404 563498 310586 563734
rect 310822 563498 311004 563734
rect 310404 528054 311004 563498
rect 310404 527818 310586 528054
rect 310822 527818 311004 528054
rect 310404 527734 311004 527818
rect 310404 527498 310586 527734
rect 310822 527498 311004 527734
rect 310404 492054 311004 527498
rect 310404 491818 310586 492054
rect 310822 491818 311004 492054
rect 310404 491734 311004 491818
rect 310404 491498 310586 491734
rect 310822 491498 311004 491734
rect 310404 456054 311004 491498
rect 310404 455818 310586 456054
rect 310822 455818 311004 456054
rect 310404 455734 311004 455818
rect 310404 455498 310586 455734
rect 310822 455498 311004 455734
rect 310404 420054 311004 455498
rect 310404 419818 310586 420054
rect 310822 419818 311004 420054
rect 310404 419734 311004 419818
rect 310404 419498 310586 419734
rect 310822 419498 311004 419734
rect 310404 384054 311004 419498
rect 310404 383818 310586 384054
rect 310822 383818 311004 384054
rect 310404 383734 311004 383818
rect 310404 383498 310586 383734
rect 310822 383498 311004 383734
rect 310404 348054 311004 383498
rect 310404 347818 310586 348054
rect 310822 347818 311004 348054
rect 310404 347734 311004 347818
rect 310404 347498 310586 347734
rect 310822 347498 311004 347734
rect 310404 312054 311004 347498
rect 310404 311818 310586 312054
rect 310822 311818 311004 312054
rect 310404 311734 311004 311818
rect 310404 311498 310586 311734
rect 310822 311498 311004 311734
rect 310404 276054 311004 311498
rect 310404 275818 310586 276054
rect 310822 275818 311004 276054
rect 310404 275734 311004 275818
rect 310404 275498 310586 275734
rect 310822 275498 311004 275734
rect 310404 240054 311004 275498
rect 310404 239818 310586 240054
rect 310822 239818 311004 240054
rect 310404 239734 311004 239818
rect 310404 239498 310586 239734
rect 310822 239498 311004 239734
rect 310404 204054 311004 239498
rect 310404 203818 310586 204054
rect 310822 203818 311004 204054
rect 310404 203734 311004 203818
rect 310404 203498 310586 203734
rect 310822 203498 311004 203734
rect 310404 168054 311004 203498
rect 310404 167818 310586 168054
rect 310822 167818 311004 168054
rect 310404 167734 311004 167818
rect 310404 167498 310586 167734
rect 310822 167498 311004 167734
rect 310404 132054 311004 167498
rect 310404 131818 310586 132054
rect 310822 131818 311004 132054
rect 310404 131734 311004 131818
rect 310404 131498 310586 131734
rect 310822 131498 311004 131734
rect 310404 96054 311004 131498
rect 310404 95818 310586 96054
rect 310822 95818 311004 96054
rect 310404 95734 311004 95818
rect 310404 95498 310586 95734
rect 310822 95498 311004 95734
rect 310404 60054 311004 95498
rect 310404 59818 310586 60054
rect 310822 59818 311004 60054
rect 310404 59734 311004 59818
rect 310404 59498 310586 59734
rect 310822 59498 311004 59734
rect 310404 24054 311004 59498
rect 310404 23818 310586 24054
rect 310822 23818 311004 24054
rect 310404 23734 311004 23818
rect 310404 23498 310586 23734
rect 310822 23498 311004 23734
rect 310404 -3106 311004 23498
rect 310404 -3342 310586 -3106
rect 310822 -3342 311004 -3106
rect 310404 -3426 311004 -3342
rect 310404 -3662 310586 -3426
rect 310822 -3662 311004 -3426
rect 310404 -3684 311004 -3662
rect 314004 675654 314604 708882
rect 314004 675418 314186 675654
rect 314422 675418 314604 675654
rect 314004 675334 314604 675418
rect 314004 675098 314186 675334
rect 314422 675098 314604 675334
rect 314004 639654 314604 675098
rect 314004 639418 314186 639654
rect 314422 639418 314604 639654
rect 314004 639334 314604 639418
rect 314004 639098 314186 639334
rect 314422 639098 314604 639334
rect 314004 603654 314604 639098
rect 314004 603418 314186 603654
rect 314422 603418 314604 603654
rect 314004 603334 314604 603418
rect 314004 603098 314186 603334
rect 314422 603098 314604 603334
rect 314004 567654 314604 603098
rect 314004 567418 314186 567654
rect 314422 567418 314604 567654
rect 314004 567334 314604 567418
rect 314004 567098 314186 567334
rect 314422 567098 314604 567334
rect 314004 531654 314604 567098
rect 314004 531418 314186 531654
rect 314422 531418 314604 531654
rect 314004 531334 314604 531418
rect 314004 531098 314186 531334
rect 314422 531098 314604 531334
rect 314004 495654 314604 531098
rect 314004 495418 314186 495654
rect 314422 495418 314604 495654
rect 314004 495334 314604 495418
rect 314004 495098 314186 495334
rect 314422 495098 314604 495334
rect 314004 459654 314604 495098
rect 314004 459418 314186 459654
rect 314422 459418 314604 459654
rect 314004 459334 314604 459418
rect 314004 459098 314186 459334
rect 314422 459098 314604 459334
rect 314004 423654 314604 459098
rect 314004 423418 314186 423654
rect 314422 423418 314604 423654
rect 314004 423334 314604 423418
rect 314004 423098 314186 423334
rect 314422 423098 314604 423334
rect 314004 387654 314604 423098
rect 314004 387418 314186 387654
rect 314422 387418 314604 387654
rect 314004 387334 314604 387418
rect 314004 387098 314186 387334
rect 314422 387098 314604 387334
rect 314004 351654 314604 387098
rect 314004 351418 314186 351654
rect 314422 351418 314604 351654
rect 314004 351334 314604 351418
rect 314004 351098 314186 351334
rect 314422 351098 314604 351334
rect 314004 315654 314604 351098
rect 314004 315418 314186 315654
rect 314422 315418 314604 315654
rect 314004 315334 314604 315418
rect 314004 315098 314186 315334
rect 314422 315098 314604 315334
rect 314004 279654 314604 315098
rect 314004 279418 314186 279654
rect 314422 279418 314604 279654
rect 314004 279334 314604 279418
rect 314004 279098 314186 279334
rect 314422 279098 314604 279334
rect 314004 243654 314604 279098
rect 314004 243418 314186 243654
rect 314422 243418 314604 243654
rect 314004 243334 314604 243418
rect 314004 243098 314186 243334
rect 314422 243098 314604 243334
rect 314004 207654 314604 243098
rect 314004 207418 314186 207654
rect 314422 207418 314604 207654
rect 314004 207334 314604 207418
rect 314004 207098 314186 207334
rect 314422 207098 314604 207334
rect 314004 171654 314604 207098
rect 314004 171418 314186 171654
rect 314422 171418 314604 171654
rect 314004 171334 314604 171418
rect 314004 171098 314186 171334
rect 314422 171098 314604 171334
rect 314004 135654 314604 171098
rect 314004 135418 314186 135654
rect 314422 135418 314604 135654
rect 314004 135334 314604 135418
rect 314004 135098 314186 135334
rect 314422 135098 314604 135334
rect 314004 99654 314604 135098
rect 314004 99418 314186 99654
rect 314422 99418 314604 99654
rect 314004 99334 314604 99418
rect 314004 99098 314186 99334
rect 314422 99098 314604 99334
rect 314004 63654 314604 99098
rect 314004 63418 314186 63654
rect 314422 63418 314604 63654
rect 314004 63334 314604 63418
rect 314004 63098 314186 63334
rect 314422 63098 314604 63334
rect 314004 27654 314604 63098
rect 314004 27418 314186 27654
rect 314422 27418 314604 27654
rect 314004 27334 314604 27418
rect 314004 27098 314186 27334
rect 314422 27098 314604 27334
rect 314004 -4946 314604 27098
rect 314004 -5182 314186 -4946
rect 314422 -5182 314604 -4946
rect 314004 -5266 314604 -5182
rect 314004 -5502 314186 -5266
rect 314422 -5502 314604 -5266
rect 314004 -5524 314604 -5502
rect 317604 679254 318204 710722
rect 335604 710358 336204 711300
rect 335604 710122 335786 710358
rect 336022 710122 336204 710358
rect 335604 710038 336204 710122
rect 335604 709802 335786 710038
rect 336022 709802 336204 710038
rect 332004 708518 332604 709460
rect 332004 708282 332186 708518
rect 332422 708282 332604 708518
rect 332004 708198 332604 708282
rect 332004 707962 332186 708198
rect 332422 707962 332604 708198
rect 328404 706678 329004 707620
rect 328404 706442 328586 706678
rect 328822 706442 329004 706678
rect 328404 706358 329004 706442
rect 328404 706122 328586 706358
rect 328822 706122 329004 706358
rect 317604 679018 317786 679254
rect 318022 679018 318204 679254
rect 317604 678934 318204 679018
rect 317604 678698 317786 678934
rect 318022 678698 318204 678934
rect 317604 643254 318204 678698
rect 317604 643018 317786 643254
rect 318022 643018 318204 643254
rect 317604 642934 318204 643018
rect 317604 642698 317786 642934
rect 318022 642698 318204 642934
rect 317604 607254 318204 642698
rect 317604 607018 317786 607254
rect 318022 607018 318204 607254
rect 317604 606934 318204 607018
rect 317604 606698 317786 606934
rect 318022 606698 318204 606934
rect 317604 571254 318204 606698
rect 317604 571018 317786 571254
rect 318022 571018 318204 571254
rect 317604 570934 318204 571018
rect 317604 570698 317786 570934
rect 318022 570698 318204 570934
rect 317604 535254 318204 570698
rect 317604 535018 317786 535254
rect 318022 535018 318204 535254
rect 317604 534934 318204 535018
rect 317604 534698 317786 534934
rect 318022 534698 318204 534934
rect 317604 499254 318204 534698
rect 317604 499018 317786 499254
rect 318022 499018 318204 499254
rect 317604 498934 318204 499018
rect 317604 498698 317786 498934
rect 318022 498698 318204 498934
rect 317604 463254 318204 498698
rect 317604 463018 317786 463254
rect 318022 463018 318204 463254
rect 317604 462934 318204 463018
rect 317604 462698 317786 462934
rect 318022 462698 318204 462934
rect 317604 427254 318204 462698
rect 317604 427018 317786 427254
rect 318022 427018 318204 427254
rect 317604 426934 318204 427018
rect 317604 426698 317786 426934
rect 318022 426698 318204 426934
rect 317604 391254 318204 426698
rect 317604 391018 317786 391254
rect 318022 391018 318204 391254
rect 317604 390934 318204 391018
rect 317604 390698 317786 390934
rect 318022 390698 318204 390934
rect 317604 355254 318204 390698
rect 317604 355018 317786 355254
rect 318022 355018 318204 355254
rect 317604 354934 318204 355018
rect 317604 354698 317786 354934
rect 318022 354698 318204 354934
rect 317604 319254 318204 354698
rect 317604 319018 317786 319254
rect 318022 319018 318204 319254
rect 317604 318934 318204 319018
rect 317604 318698 317786 318934
rect 318022 318698 318204 318934
rect 317604 283254 318204 318698
rect 317604 283018 317786 283254
rect 318022 283018 318204 283254
rect 317604 282934 318204 283018
rect 317604 282698 317786 282934
rect 318022 282698 318204 282934
rect 317604 247254 318204 282698
rect 317604 247018 317786 247254
rect 318022 247018 318204 247254
rect 317604 246934 318204 247018
rect 317604 246698 317786 246934
rect 318022 246698 318204 246934
rect 317604 211254 318204 246698
rect 317604 211018 317786 211254
rect 318022 211018 318204 211254
rect 317604 210934 318204 211018
rect 317604 210698 317786 210934
rect 318022 210698 318204 210934
rect 317604 175254 318204 210698
rect 317604 175018 317786 175254
rect 318022 175018 318204 175254
rect 317604 174934 318204 175018
rect 317604 174698 317786 174934
rect 318022 174698 318204 174934
rect 317604 139254 318204 174698
rect 317604 139018 317786 139254
rect 318022 139018 318204 139254
rect 317604 138934 318204 139018
rect 317604 138698 317786 138934
rect 318022 138698 318204 138934
rect 317604 103254 318204 138698
rect 317604 103018 317786 103254
rect 318022 103018 318204 103254
rect 317604 102934 318204 103018
rect 317604 102698 317786 102934
rect 318022 102698 318204 102934
rect 317604 67254 318204 102698
rect 317604 67018 317786 67254
rect 318022 67018 318204 67254
rect 317604 66934 318204 67018
rect 317604 66698 317786 66934
rect 318022 66698 318204 66934
rect 317604 31254 318204 66698
rect 317604 31018 317786 31254
rect 318022 31018 318204 31254
rect 317604 30934 318204 31018
rect 317604 30698 317786 30934
rect 318022 30698 318204 30934
rect 299604 -6102 299786 -5866
rect 300022 -6102 300204 -5866
rect 299604 -6186 300204 -6102
rect 299604 -6422 299786 -6186
rect 300022 -6422 300204 -6186
rect 299604 -7364 300204 -6422
rect 317604 -6786 318204 30698
rect 324804 704838 325404 705780
rect 324804 704602 324986 704838
rect 325222 704602 325404 704838
rect 324804 704518 325404 704602
rect 324804 704282 324986 704518
rect 325222 704282 325404 704518
rect 324804 686454 325404 704282
rect 324804 686218 324986 686454
rect 325222 686218 325404 686454
rect 324804 686134 325404 686218
rect 324804 685898 324986 686134
rect 325222 685898 325404 686134
rect 324804 650454 325404 685898
rect 324804 650218 324986 650454
rect 325222 650218 325404 650454
rect 324804 650134 325404 650218
rect 324804 649898 324986 650134
rect 325222 649898 325404 650134
rect 324804 614454 325404 649898
rect 324804 614218 324986 614454
rect 325222 614218 325404 614454
rect 324804 614134 325404 614218
rect 324804 613898 324986 614134
rect 325222 613898 325404 614134
rect 324804 578454 325404 613898
rect 324804 578218 324986 578454
rect 325222 578218 325404 578454
rect 324804 578134 325404 578218
rect 324804 577898 324986 578134
rect 325222 577898 325404 578134
rect 324804 542454 325404 577898
rect 324804 542218 324986 542454
rect 325222 542218 325404 542454
rect 324804 542134 325404 542218
rect 324804 541898 324986 542134
rect 325222 541898 325404 542134
rect 324804 506454 325404 541898
rect 324804 506218 324986 506454
rect 325222 506218 325404 506454
rect 324804 506134 325404 506218
rect 324804 505898 324986 506134
rect 325222 505898 325404 506134
rect 324804 470454 325404 505898
rect 324804 470218 324986 470454
rect 325222 470218 325404 470454
rect 324804 470134 325404 470218
rect 324804 469898 324986 470134
rect 325222 469898 325404 470134
rect 324804 434454 325404 469898
rect 324804 434218 324986 434454
rect 325222 434218 325404 434454
rect 324804 434134 325404 434218
rect 324804 433898 324986 434134
rect 325222 433898 325404 434134
rect 324804 398454 325404 433898
rect 324804 398218 324986 398454
rect 325222 398218 325404 398454
rect 324804 398134 325404 398218
rect 324804 397898 324986 398134
rect 325222 397898 325404 398134
rect 324804 362454 325404 397898
rect 324804 362218 324986 362454
rect 325222 362218 325404 362454
rect 324804 362134 325404 362218
rect 324804 361898 324986 362134
rect 325222 361898 325404 362134
rect 324804 326454 325404 361898
rect 324804 326218 324986 326454
rect 325222 326218 325404 326454
rect 324804 326134 325404 326218
rect 324804 325898 324986 326134
rect 325222 325898 325404 326134
rect 324804 290454 325404 325898
rect 324804 290218 324986 290454
rect 325222 290218 325404 290454
rect 324804 290134 325404 290218
rect 324804 289898 324986 290134
rect 325222 289898 325404 290134
rect 324804 254454 325404 289898
rect 324804 254218 324986 254454
rect 325222 254218 325404 254454
rect 324804 254134 325404 254218
rect 324804 253898 324986 254134
rect 325222 253898 325404 254134
rect 324804 218454 325404 253898
rect 324804 218218 324986 218454
rect 325222 218218 325404 218454
rect 324804 218134 325404 218218
rect 324804 217898 324986 218134
rect 325222 217898 325404 218134
rect 324804 182454 325404 217898
rect 324804 182218 324986 182454
rect 325222 182218 325404 182454
rect 324804 182134 325404 182218
rect 324804 181898 324986 182134
rect 325222 181898 325404 182134
rect 324804 146454 325404 181898
rect 324804 146218 324986 146454
rect 325222 146218 325404 146454
rect 324804 146134 325404 146218
rect 324804 145898 324986 146134
rect 325222 145898 325404 146134
rect 324804 110454 325404 145898
rect 324804 110218 324986 110454
rect 325222 110218 325404 110454
rect 324804 110134 325404 110218
rect 324804 109898 324986 110134
rect 325222 109898 325404 110134
rect 324804 74454 325404 109898
rect 324804 74218 324986 74454
rect 325222 74218 325404 74454
rect 324804 74134 325404 74218
rect 324804 73898 324986 74134
rect 325222 73898 325404 74134
rect 324804 38454 325404 73898
rect 324804 38218 324986 38454
rect 325222 38218 325404 38454
rect 324804 38134 325404 38218
rect 324804 37898 324986 38134
rect 325222 37898 325404 38134
rect 324804 2454 325404 37898
rect 324804 2218 324986 2454
rect 325222 2218 325404 2454
rect 324804 2134 325404 2218
rect 324804 1898 324986 2134
rect 325222 1898 325404 2134
rect 324804 -346 325404 1898
rect 324804 -582 324986 -346
rect 325222 -582 325404 -346
rect 324804 -666 325404 -582
rect 324804 -902 324986 -666
rect 325222 -902 325404 -666
rect 324804 -1844 325404 -902
rect 328404 690054 329004 706122
rect 328404 689818 328586 690054
rect 328822 689818 329004 690054
rect 328404 689734 329004 689818
rect 328404 689498 328586 689734
rect 328822 689498 329004 689734
rect 328404 654054 329004 689498
rect 328404 653818 328586 654054
rect 328822 653818 329004 654054
rect 328404 653734 329004 653818
rect 328404 653498 328586 653734
rect 328822 653498 329004 653734
rect 328404 618054 329004 653498
rect 328404 617818 328586 618054
rect 328822 617818 329004 618054
rect 328404 617734 329004 617818
rect 328404 617498 328586 617734
rect 328822 617498 329004 617734
rect 328404 582054 329004 617498
rect 328404 581818 328586 582054
rect 328822 581818 329004 582054
rect 328404 581734 329004 581818
rect 328404 581498 328586 581734
rect 328822 581498 329004 581734
rect 328404 546054 329004 581498
rect 328404 545818 328586 546054
rect 328822 545818 329004 546054
rect 328404 545734 329004 545818
rect 328404 545498 328586 545734
rect 328822 545498 329004 545734
rect 328404 510054 329004 545498
rect 328404 509818 328586 510054
rect 328822 509818 329004 510054
rect 328404 509734 329004 509818
rect 328404 509498 328586 509734
rect 328822 509498 329004 509734
rect 328404 474054 329004 509498
rect 328404 473818 328586 474054
rect 328822 473818 329004 474054
rect 328404 473734 329004 473818
rect 328404 473498 328586 473734
rect 328822 473498 329004 473734
rect 328404 438054 329004 473498
rect 328404 437818 328586 438054
rect 328822 437818 329004 438054
rect 328404 437734 329004 437818
rect 328404 437498 328586 437734
rect 328822 437498 329004 437734
rect 328404 402054 329004 437498
rect 328404 401818 328586 402054
rect 328822 401818 329004 402054
rect 328404 401734 329004 401818
rect 328404 401498 328586 401734
rect 328822 401498 329004 401734
rect 328404 366054 329004 401498
rect 328404 365818 328586 366054
rect 328822 365818 329004 366054
rect 328404 365734 329004 365818
rect 328404 365498 328586 365734
rect 328822 365498 329004 365734
rect 328404 330054 329004 365498
rect 328404 329818 328586 330054
rect 328822 329818 329004 330054
rect 328404 329734 329004 329818
rect 328404 329498 328586 329734
rect 328822 329498 329004 329734
rect 328404 294054 329004 329498
rect 328404 293818 328586 294054
rect 328822 293818 329004 294054
rect 328404 293734 329004 293818
rect 328404 293498 328586 293734
rect 328822 293498 329004 293734
rect 328404 258054 329004 293498
rect 328404 257818 328586 258054
rect 328822 257818 329004 258054
rect 328404 257734 329004 257818
rect 328404 257498 328586 257734
rect 328822 257498 329004 257734
rect 328404 222054 329004 257498
rect 328404 221818 328586 222054
rect 328822 221818 329004 222054
rect 328404 221734 329004 221818
rect 328404 221498 328586 221734
rect 328822 221498 329004 221734
rect 328404 186054 329004 221498
rect 328404 185818 328586 186054
rect 328822 185818 329004 186054
rect 328404 185734 329004 185818
rect 328404 185498 328586 185734
rect 328822 185498 329004 185734
rect 328404 150054 329004 185498
rect 328404 149818 328586 150054
rect 328822 149818 329004 150054
rect 328404 149734 329004 149818
rect 328404 149498 328586 149734
rect 328822 149498 329004 149734
rect 328404 114054 329004 149498
rect 328404 113818 328586 114054
rect 328822 113818 329004 114054
rect 328404 113734 329004 113818
rect 328404 113498 328586 113734
rect 328822 113498 329004 113734
rect 328404 78054 329004 113498
rect 328404 77818 328586 78054
rect 328822 77818 329004 78054
rect 328404 77734 329004 77818
rect 328404 77498 328586 77734
rect 328822 77498 329004 77734
rect 328404 42054 329004 77498
rect 328404 41818 328586 42054
rect 328822 41818 329004 42054
rect 328404 41734 329004 41818
rect 328404 41498 328586 41734
rect 328822 41498 329004 41734
rect 328404 6054 329004 41498
rect 328404 5818 328586 6054
rect 328822 5818 329004 6054
rect 328404 5734 329004 5818
rect 328404 5498 328586 5734
rect 328822 5498 329004 5734
rect 328404 -2186 329004 5498
rect 328404 -2422 328586 -2186
rect 328822 -2422 329004 -2186
rect 328404 -2506 329004 -2422
rect 328404 -2742 328586 -2506
rect 328822 -2742 329004 -2506
rect 328404 -3684 329004 -2742
rect 332004 693654 332604 707962
rect 332004 693418 332186 693654
rect 332422 693418 332604 693654
rect 332004 693334 332604 693418
rect 332004 693098 332186 693334
rect 332422 693098 332604 693334
rect 332004 657654 332604 693098
rect 332004 657418 332186 657654
rect 332422 657418 332604 657654
rect 332004 657334 332604 657418
rect 332004 657098 332186 657334
rect 332422 657098 332604 657334
rect 332004 621654 332604 657098
rect 332004 621418 332186 621654
rect 332422 621418 332604 621654
rect 332004 621334 332604 621418
rect 332004 621098 332186 621334
rect 332422 621098 332604 621334
rect 332004 585654 332604 621098
rect 332004 585418 332186 585654
rect 332422 585418 332604 585654
rect 332004 585334 332604 585418
rect 332004 585098 332186 585334
rect 332422 585098 332604 585334
rect 332004 549654 332604 585098
rect 332004 549418 332186 549654
rect 332422 549418 332604 549654
rect 332004 549334 332604 549418
rect 332004 549098 332186 549334
rect 332422 549098 332604 549334
rect 332004 513654 332604 549098
rect 332004 513418 332186 513654
rect 332422 513418 332604 513654
rect 332004 513334 332604 513418
rect 332004 513098 332186 513334
rect 332422 513098 332604 513334
rect 332004 477654 332604 513098
rect 332004 477418 332186 477654
rect 332422 477418 332604 477654
rect 332004 477334 332604 477418
rect 332004 477098 332186 477334
rect 332422 477098 332604 477334
rect 332004 441654 332604 477098
rect 332004 441418 332186 441654
rect 332422 441418 332604 441654
rect 332004 441334 332604 441418
rect 332004 441098 332186 441334
rect 332422 441098 332604 441334
rect 332004 405654 332604 441098
rect 332004 405418 332186 405654
rect 332422 405418 332604 405654
rect 332004 405334 332604 405418
rect 332004 405098 332186 405334
rect 332422 405098 332604 405334
rect 332004 369654 332604 405098
rect 332004 369418 332186 369654
rect 332422 369418 332604 369654
rect 332004 369334 332604 369418
rect 332004 369098 332186 369334
rect 332422 369098 332604 369334
rect 332004 333654 332604 369098
rect 332004 333418 332186 333654
rect 332422 333418 332604 333654
rect 332004 333334 332604 333418
rect 332004 333098 332186 333334
rect 332422 333098 332604 333334
rect 332004 297654 332604 333098
rect 332004 297418 332186 297654
rect 332422 297418 332604 297654
rect 332004 297334 332604 297418
rect 332004 297098 332186 297334
rect 332422 297098 332604 297334
rect 332004 261654 332604 297098
rect 332004 261418 332186 261654
rect 332422 261418 332604 261654
rect 332004 261334 332604 261418
rect 332004 261098 332186 261334
rect 332422 261098 332604 261334
rect 332004 225654 332604 261098
rect 332004 225418 332186 225654
rect 332422 225418 332604 225654
rect 332004 225334 332604 225418
rect 332004 225098 332186 225334
rect 332422 225098 332604 225334
rect 332004 189654 332604 225098
rect 332004 189418 332186 189654
rect 332422 189418 332604 189654
rect 332004 189334 332604 189418
rect 332004 189098 332186 189334
rect 332422 189098 332604 189334
rect 332004 153654 332604 189098
rect 332004 153418 332186 153654
rect 332422 153418 332604 153654
rect 332004 153334 332604 153418
rect 332004 153098 332186 153334
rect 332422 153098 332604 153334
rect 332004 117654 332604 153098
rect 332004 117418 332186 117654
rect 332422 117418 332604 117654
rect 332004 117334 332604 117418
rect 332004 117098 332186 117334
rect 332422 117098 332604 117334
rect 332004 81654 332604 117098
rect 332004 81418 332186 81654
rect 332422 81418 332604 81654
rect 332004 81334 332604 81418
rect 332004 81098 332186 81334
rect 332422 81098 332604 81334
rect 332004 45654 332604 81098
rect 332004 45418 332186 45654
rect 332422 45418 332604 45654
rect 332004 45334 332604 45418
rect 332004 45098 332186 45334
rect 332422 45098 332604 45334
rect 332004 9654 332604 45098
rect 332004 9418 332186 9654
rect 332422 9418 332604 9654
rect 332004 9334 332604 9418
rect 332004 9098 332186 9334
rect 332422 9098 332604 9334
rect 332004 -4026 332604 9098
rect 332004 -4262 332186 -4026
rect 332422 -4262 332604 -4026
rect 332004 -4346 332604 -4262
rect 332004 -4582 332186 -4346
rect 332422 -4582 332604 -4346
rect 332004 -5524 332604 -4582
rect 335604 697254 336204 709802
rect 353604 711278 354204 711300
rect 353604 711042 353786 711278
rect 354022 711042 354204 711278
rect 353604 710958 354204 711042
rect 353604 710722 353786 710958
rect 354022 710722 354204 710958
rect 350004 709438 350604 709460
rect 350004 709202 350186 709438
rect 350422 709202 350604 709438
rect 350004 709118 350604 709202
rect 350004 708882 350186 709118
rect 350422 708882 350604 709118
rect 346404 707598 347004 707620
rect 346404 707362 346586 707598
rect 346822 707362 347004 707598
rect 346404 707278 347004 707362
rect 346404 707042 346586 707278
rect 346822 707042 347004 707278
rect 335604 697018 335786 697254
rect 336022 697018 336204 697254
rect 335604 696934 336204 697018
rect 335604 696698 335786 696934
rect 336022 696698 336204 696934
rect 335604 661254 336204 696698
rect 335604 661018 335786 661254
rect 336022 661018 336204 661254
rect 335604 660934 336204 661018
rect 335604 660698 335786 660934
rect 336022 660698 336204 660934
rect 335604 625254 336204 660698
rect 335604 625018 335786 625254
rect 336022 625018 336204 625254
rect 335604 624934 336204 625018
rect 335604 624698 335786 624934
rect 336022 624698 336204 624934
rect 335604 589254 336204 624698
rect 335604 589018 335786 589254
rect 336022 589018 336204 589254
rect 335604 588934 336204 589018
rect 335604 588698 335786 588934
rect 336022 588698 336204 588934
rect 335604 553254 336204 588698
rect 335604 553018 335786 553254
rect 336022 553018 336204 553254
rect 335604 552934 336204 553018
rect 335604 552698 335786 552934
rect 336022 552698 336204 552934
rect 335604 517254 336204 552698
rect 335604 517018 335786 517254
rect 336022 517018 336204 517254
rect 335604 516934 336204 517018
rect 335604 516698 335786 516934
rect 336022 516698 336204 516934
rect 335604 481254 336204 516698
rect 335604 481018 335786 481254
rect 336022 481018 336204 481254
rect 335604 480934 336204 481018
rect 335604 480698 335786 480934
rect 336022 480698 336204 480934
rect 335604 445254 336204 480698
rect 335604 445018 335786 445254
rect 336022 445018 336204 445254
rect 335604 444934 336204 445018
rect 335604 444698 335786 444934
rect 336022 444698 336204 444934
rect 335604 409254 336204 444698
rect 335604 409018 335786 409254
rect 336022 409018 336204 409254
rect 335604 408934 336204 409018
rect 335604 408698 335786 408934
rect 336022 408698 336204 408934
rect 335604 373254 336204 408698
rect 335604 373018 335786 373254
rect 336022 373018 336204 373254
rect 335604 372934 336204 373018
rect 335604 372698 335786 372934
rect 336022 372698 336204 372934
rect 335604 337254 336204 372698
rect 335604 337018 335786 337254
rect 336022 337018 336204 337254
rect 335604 336934 336204 337018
rect 335604 336698 335786 336934
rect 336022 336698 336204 336934
rect 335604 301254 336204 336698
rect 335604 301018 335786 301254
rect 336022 301018 336204 301254
rect 335604 300934 336204 301018
rect 335604 300698 335786 300934
rect 336022 300698 336204 300934
rect 335604 265254 336204 300698
rect 335604 265018 335786 265254
rect 336022 265018 336204 265254
rect 335604 264934 336204 265018
rect 335604 264698 335786 264934
rect 336022 264698 336204 264934
rect 335604 229254 336204 264698
rect 335604 229018 335786 229254
rect 336022 229018 336204 229254
rect 335604 228934 336204 229018
rect 335604 228698 335786 228934
rect 336022 228698 336204 228934
rect 335604 193254 336204 228698
rect 335604 193018 335786 193254
rect 336022 193018 336204 193254
rect 335604 192934 336204 193018
rect 335604 192698 335786 192934
rect 336022 192698 336204 192934
rect 335604 157254 336204 192698
rect 335604 157018 335786 157254
rect 336022 157018 336204 157254
rect 335604 156934 336204 157018
rect 335604 156698 335786 156934
rect 336022 156698 336204 156934
rect 335604 121254 336204 156698
rect 335604 121018 335786 121254
rect 336022 121018 336204 121254
rect 335604 120934 336204 121018
rect 335604 120698 335786 120934
rect 336022 120698 336204 120934
rect 335604 85254 336204 120698
rect 335604 85018 335786 85254
rect 336022 85018 336204 85254
rect 335604 84934 336204 85018
rect 335604 84698 335786 84934
rect 336022 84698 336204 84934
rect 335604 49254 336204 84698
rect 335604 49018 335786 49254
rect 336022 49018 336204 49254
rect 335604 48934 336204 49018
rect 335604 48698 335786 48934
rect 336022 48698 336204 48934
rect 335604 13254 336204 48698
rect 335604 13018 335786 13254
rect 336022 13018 336204 13254
rect 335604 12934 336204 13018
rect 335604 12698 335786 12934
rect 336022 12698 336204 12934
rect 317604 -7022 317786 -6786
rect 318022 -7022 318204 -6786
rect 317604 -7106 318204 -7022
rect 317604 -7342 317786 -7106
rect 318022 -7342 318204 -7106
rect 317604 -7364 318204 -7342
rect 335604 -5866 336204 12698
rect 342804 705758 343404 705780
rect 342804 705522 342986 705758
rect 343222 705522 343404 705758
rect 342804 705438 343404 705522
rect 342804 705202 342986 705438
rect 343222 705202 343404 705438
rect 342804 668454 343404 705202
rect 342804 668218 342986 668454
rect 343222 668218 343404 668454
rect 342804 668134 343404 668218
rect 342804 667898 342986 668134
rect 343222 667898 343404 668134
rect 342804 632454 343404 667898
rect 342804 632218 342986 632454
rect 343222 632218 343404 632454
rect 342804 632134 343404 632218
rect 342804 631898 342986 632134
rect 343222 631898 343404 632134
rect 342804 596454 343404 631898
rect 342804 596218 342986 596454
rect 343222 596218 343404 596454
rect 342804 596134 343404 596218
rect 342804 595898 342986 596134
rect 343222 595898 343404 596134
rect 342804 560454 343404 595898
rect 342804 560218 342986 560454
rect 343222 560218 343404 560454
rect 342804 560134 343404 560218
rect 342804 559898 342986 560134
rect 343222 559898 343404 560134
rect 342804 524454 343404 559898
rect 342804 524218 342986 524454
rect 343222 524218 343404 524454
rect 342804 524134 343404 524218
rect 342804 523898 342986 524134
rect 343222 523898 343404 524134
rect 342804 488454 343404 523898
rect 342804 488218 342986 488454
rect 343222 488218 343404 488454
rect 342804 488134 343404 488218
rect 342804 487898 342986 488134
rect 343222 487898 343404 488134
rect 342804 452454 343404 487898
rect 342804 452218 342986 452454
rect 343222 452218 343404 452454
rect 342804 452134 343404 452218
rect 342804 451898 342986 452134
rect 343222 451898 343404 452134
rect 342804 416454 343404 451898
rect 342804 416218 342986 416454
rect 343222 416218 343404 416454
rect 342804 416134 343404 416218
rect 342804 415898 342986 416134
rect 343222 415898 343404 416134
rect 342804 380454 343404 415898
rect 342804 380218 342986 380454
rect 343222 380218 343404 380454
rect 342804 380134 343404 380218
rect 342804 379898 342986 380134
rect 343222 379898 343404 380134
rect 342804 344454 343404 379898
rect 342804 344218 342986 344454
rect 343222 344218 343404 344454
rect 342804 344134 343404 344218
rect 342804 343898 342986 344134
rect 343222 343898 343404 344134
rect 342804 308454 343404 343898
rect 342804 308218 342986 308454
rect 343222 308218 343404 308454
rect 342804 308134 343404 308218
rect 342804 307898 342986 308134
rect 343222 307898 343404 308134
rect 342804 272454 343404 307898
rect 342804 272218 342986 272454
rect 343222 272218 343404 272454
rect 342804 272134 343404 272218
rect 342804 271898 342986 272134
rect 343222 271898 343404 272134
rect 342804 236454 343404 271898
rect 342804 236218 342986 236454
rect 343222 236218 343404 236454
rect 342804 236134 343404 236218
rect 342804 235898 342986 236134
rect 343222 235898 343404 236134
rect 342804 200454 343404 235898
rect 342804 200218 342986 200454
rect 343222 200218 343404 200454
rect 342804 200134 343404 200218
rect 342804 199898 342986 200134
rect 343222 199898 343404 200134
rect 342804 164454 343404 199898
rect 342804 164218 342986 164454
rect 343222 164218 343404 164454
rect 342804 164134 343404 164218
rect 342804 163898 342986 164134
rect 343222 163898 343404 164134
rect 342804 128454 343404 163898
rect 342804 128218 342986 128454
rect 343222 128218 343404 128454
rect 342804 128134 343404 128218
rect 342804 127898 342986 128134
rect 343222 127898 343404 128134
rect 342804 92454 343404 127898
rect 342804 92218 342986 92454
rect 343222 92218 343404 92454
rect 342804 92134 343404 92218
rect 342804 91898 342986 92134
rect 343222 91898 343404 92134
rect 342804 56454 343404 91898
rect 342804 56218 342986 56454
rect 343222 56218 343404 56454
rect 342804 56134 343404 56218
rect 342804 55898 342986 56134
rect 343222 55898 343404 56134
rect 342804 20454 343404 55898
rect 342804 20218 342986 20454
rect 343222 20218 343404 20454
rect 342804 20134 343404 20218
rect 342804 19898 342986 20134
rect 343222 19898 343404 20134
rect 342804 -1266 343404 19898
rect 342804 -1502 342986 -1266
rect 343222 -1502 343404 -1266
rect 342804 -1586 343404 -1502
rect 342804 -1822 342986 -1586
rect 343222 -1822 343404 -1586
rect 342804 -1844 343404 -1822
rect 346404 672054 347004 707042
rect 346404 671818 346586 672054
rect 346822 671818 347004 672054
rect 346404 671734 347004 671818
rect 346404 671498 346586 671734
rect 346822 671498 347004 671734
rect 346404 636054 347004 671498
rect 346404 635818 346586 636054
rect 346822 635818 347004 636054
rect 346404 635734 347004 635818
rect 346404 635498 346586 635734
rect 346822 635498 347004 635734
rect 346404 600054 347004 635498
rect 346404 599818 346586 600054
rect 346822 599818 347004 600054
rect 346404 599734 347004 599818
rect 346404 599498 346586 599734
rect 346822 599498 347004 599734
rect 346404 564054 347004 599498
rect 346404 563818 346586 564054
rect 346822 563818 347004 564054
rect 346404 563734 347004 563818
rect 346404 563498 346586 563734
rect 346822 563498 347004 563734
rect 346404 528054 347004 563498
rect 346404 527818 346586 528054
rect 346822 527818 347004 528054
rect 346404 527734 347004 527818
rect 346404 527498 346586 527734
rect 346822 527498 347004 527734
rect 346404 492054 347004 527498
rect 346404 491818 346586 492054
rect 346822 491818 347004 492054
rect 346404 491734 347004 491818
rect 346404 491498 346586 491734
rect 346822 491498 347004 491734
rect 346404 456054 347004 491498
rect 346404 455818 346586 456054
rect 346822 455818 347004 456054
rect 346404 455734 347004 455818
rect 346404 455498 346586 455734
rect 346822 455498 347004 455734
rect 346404 420054 347004 455498
rect 346404 419818 346586 420054
rect 346822 419818 347004 420054
rect 346404 419734 347004 419818
rect 346404 419498 346586 419734
rect 346822 419498 347004 419734
rect 346404 384054 347004 419498
rect 346404 383818 346586 384054
rect 346822 383818 347004 384054
rect 346404 383734 347004 383818
rect 346404 383498 346586 383734
rect 346822 383498 347004 383734
rect 346404 348054 347004 383498
rect 346404 347818 346586 348054
rect 346822 347818 347004 348054
rect 346404 347734 347004 347818
rect 346404 347498 346586 347734
rect 346822 347498 347004 347734
rect 346404 312054 347004 347498
rect 346404 311818 346586 312054
rect 346822 311818 347004 312054
rect 346404 311734 347004 311818
rect 346404 311498 346586 311734
rect 346822 311498 347004 311734
rect 346404 276054 347004 311498
rect 346404 275818 346586 276054
rect 346822 275818 347004 276054
rect 346404 275734 347004 275818
rect 346404 275498 346586 275734
rect 346822 275498 347004 275734
rect 346404 240054 347004 275498
rect 346404 239818 346586 240054
rect 346822 239818 347004 240054
rect 346404 239734 347004 239818
rect 346404 239498 346586 239734
rect 346822 239498 347004 239734
rect 346404 204054 347004 239498
rect 346404 203818 346586 204054
rect 346822 203818 347004 204054
rect 346404 203734 347004 203818
rect 346404 203498 346586 203734
rect 346822 203498 347004 203734
rect 346404 168054 347004 203498
rect 346404 167818 346586 168054
rect 346822 167818 347004 168054
rect 346404 167734 347004 167818
rect 346404 167498 346586 167734
rect 346822 167498 347004 167734
rect 346404 132054 347004 167498
rect 346404 131818 346586 132054
rect 346822 131818 347004 132054
rect 346404 131734 347004 131818
rect 346404 131498 346586 131734
rect 346822 131498 347004 131734
rect 346404 96054 347004 131498
rect 346404 95818 346586 96054
rect 346822 95818 347004 96054
rect 346404 95734 347004 95818
rect 346404 95498 346586 95734
rect 346822 95498 347004 95734
rect 346404 60054 347004 95498
rect 346404 59818 346586 60054
rect 346822 59818 347004 60054
rect 346404 59734 347004 59818
rect 346404 59498 346586 59734
rect 346822 59498 347004 59734
rect 346404 24054 347004 59498
rect 346404 23818 346586 24054
rect 346822 23818 347004 24054
rect 346404 23734 347004 23818
rect 346404 23498 346586 23734
rect 346822 23498 347004 23734
rect 346404 -3106 347004 23498
rect 346404 -3342 346586 -3106
rect 346822 -3342 347004 -3106
rect 346404 -3426 347004 -3342
rect 346404 -3662 346586 -3426
rect 346822 -3662 347004 -3426
rect 346404 -3684 347004 -3662
rect 350004 675654 350604 708882
rect 350004 675418 350186 675654
rect 350422 675418 350604 675654
rect 350004 675334 350604 675418
rect 350004 675098 350186 675334
rect 350422 675098 350604 675334
rect 350004 639654 350604 675098
rect 350004 639418 350186 639654
rect 350422 639418 350604 639654
rect 350004 639334 350604 639418
rect 350004 639098 350186 639334
rect 350422 639098 350604 639334
rect 350004 603654 350604 639098
rect 350004 603418 350186 603654
rect 350422 603418 350604 603654
rect 350004 603334 350604 603418
rect 350004 603098 350186 603334
rect 350422 603098 350604 603334
rect 350004 567654 350604 603098
rect 350004 567418 350186 567654
rect 350422 567418 350604 567654
rect 350004 567334 350604 567418
rect 350004 567098 350186 567334
rect 350422 567098 350604 567334
rect 350004 531654 350604 567098
rect 350004 531418 350186 531654
rect 350422 531418 350604 531654
rect 350004 531334 350604 531418
rect 350004 531098 350186 531334
rect 350422 531098 350604 531334
rect 350004 495654 350604 531098
rect 350004 495418 350186 495654
rect 350422 495418 350604 495654
rect 350004 495334 350604 495418
rect 350004 495098 350186 495334
rect 350422 495098 350604 495334
rect 350004 459654 350604 495098
rect 350004 459418 350186 459654
rect 350422 459418 350604 459654
rect 350004 459334 350604 459418
rect 350004 459098 350186 459334
rect 350422 459098 350604 459334
rect 350004 423654 350604 459098
rect 350004 423418 350186 423654
rect 350422 423418 350604 423654
rect 350004 423334 350604 423418
rect 350004 423098 350186 423334
rect 350422 423098 350604 423334
rect 350004 387654 350604 423098
rect 350004 387418 350186 387654
rect 350422 387418 350604 387654
rect 350004 387334 350604 387418
rect 350004 387098 350186 387334
rect 350422 387098 350604 387334
rect 350004 351654 350604 387098
rect 350004 351418 350186 351654
rect 350422 351418 350604 351654
rect 350004 351334 350604 351418
rect 350004 351098 350186 351334
rect 350422 351098 350604 351334
rect 350004 315654 350604 351098
rect 350004 315418 350186 315654
rect 350422 315418 350604 315654
rect 350004 315334 350604 315418
rect 350004 315098 350186 315334
rect 350422 315098 350604 315334
rect 350004 279654 350604 315098
rect 350004 279418 350186 279654
rect 350422 279418 350604 279654
rect 350004 279334 350604 279418
rect 350004 279098 350186 279334
rect 350422 279098 350604 279334
rect 350004 243654 350604 279098
rect 350004 243418 350186 243654
rect 350422 243418 350604 243654
rect 350004 243334 350604 243418
rect 350004 243098 350186 243334
rect 350422 243098 350604 243334
rect 350004 207654 350604 243098
rect 350004 207418 350186 207654
rect 350422 207418 350604 207654
rect 350004 207334 350604 207418
rect 350004 207098 350186 207334
rect 350422 207098 350604 207334
rect 350004 171654 350604 207098
rect 350004 171418 350186 171654
rect 350422 171418 350604 171654
rect 350004 171334 350604 171418
rect 350004 171098 350186 171334
rect 350422 171098 350604 171334
rect 350004 135654 350604 171098
rect 350004 135418 350186 135654
rect 350422 135418 350604 135654
rect 350004 135334 350604 135418
rect 350004 135098 350186 135334
rect 350422 135098 350604 135334
rect 350004 99654 350604 135098
rect 350004 99418 350186 99654
rect 350422 99418 350604 99654
rect 350004 99334 350604 99418
rect 350004 99098 350186 99334
rect 350422 99098 350604 99334
rect 350004 63654 350604 99098
rect 350004 63418 350186 63654
rect 350422 63418 350604 63654
rect 350004 63334 350604 63418
rect 350004 63098 350186 63334
rect 350422 63098 350604 63334
rect 350004 27654 350604 63098
rect 350004 27418 350186 27654
rect 350422 27418 350604 27654
rect 350004 27334 350604 27418
rect 350004 27098 350186 27334
rect 350422 27098 350604 27334
rect 350004 -4946 350604 27098
rect 350004 -5182 350186 -4946
rect 350422 -5182 350604 -4946
rect 350004 -5266 350604 -5182
rect 350004 -5502 350186 -5266
rect 350422 -5502 350604 -5266
rect 350004 -5524 350604 -5502
rect 353604 679254 354204 710722
rect 371604 710358 372204 711300
rect 371604 710122 371786 710358
rect 372022 710122 372204 710358
rect 371604 710038 372204 710122
rect 371604 709802 371786 710038
rect 372022 709802 372204 710038
rect 368004 708518 368604 709460
rect 368004 708282 368186 708518
rect 368422 708282 368604 708518
rect 368004 708198 368604 708282
rect 368004 707962 368186 708198
rect 368422 707962 368604 708198
rect 364404 706678 365004 707620
rect 364404 706442 364586 706678
rect 364822 706442 365004 706678
rect 364404 706358 365004 706442
rect 364404 706122 364586 706358
rect 364822 706122 365004 706358
rect 353604 679018 353786 679254
rect 354022 679018 354204 679254
rect 353604 678934 354204 679018
rect 353604 678698 353786 678934
rect 354022 678698 354204 678934
rect 353604 643254 354204 678698
rect 353604 643018 353786 643254
rect 354022 643018 354204 643254
rect 353604 642934 354204 643018
rect 353604 642698 353786 642934
rect 354022 642698 354204 642934
rect 353604 607254 354204 642698
rect 353604 607018 353786 607254
rect 354022 607018 354204 607254
rect 353604 606934 354204 607018
rect 353604 606698 353786 606934
rect 354022 606698 354204 606934
rect 353604 571254 354204 606698
rect 353604 571018 353786 571254
rect 354022 571018 354204 571254
rect 353604 570934 354204 571018
rect 353604 570698 353786 570934
rect 354022 570698 354204 570934
rect 353604 535254 354204 570698
rect 353604 535018 353786 535254
rect 354022 535018 354204 535254
rect 353604 534934 354204 535018
rect 353604 534698 353786 534934
rect 354022 534698 354204 534934
rect 353604 499254 354204 534698
rect 353604 499018 353786 499254
rect 354022 499018 354204 499254
rect 353604 498934 354204 499018
rect 353604 498698 353786 498934
rect 354022 498698 354204 498934
rect 353604 463254 354204 498698
rect 353604 463018 353786 463254
rect 354022 463018 354204 463254
rect 353604 462934 354204 463018
rect 353604 462698 353786 462934
rect 354022 462698 354204 462934
rect 353604 427254 354204 462698
rect 353604 427018 353786 427254
rect 354022 427018 354204 427254
rect 353604 426934 354204 427018
rect 353604 426698 353786 426934
rect 354022 426698 354204 426934
rect 353604 391254 354204 426698
rect 353604 391018 353786 391254
rect 354022 391018 354204 391254
rect 353604 390934 354204 391018
rect 353604 390698 353786 390934
rect 354022 390698 354204 390934
rect 353604 355254 354204 390698
rect 353604 355018 353786 355254
rect 354022 355018 354204 355254
rect 353604 354934 354204 355018
rect 353604 354698 353786 354934
rect 354022 354698 354204 354934
rect 353604 319254 354204 354698
rect 360804 704838 361404 705780
rect 360804 704602 360986 704838
rect 361222 704602 361404 704838
rect 360804 704518 361404 704602
rect 360804 704282 360986 704518
rect 361222 704282 361404 704518
rect 360804 686454 361404 704282
rect 360804 686218 360986 686454
rect 361222 686218 361404 686454
rect 360804 686134 361404 686218
rect 360804 685898 360986 686134
rect 361222 685898 361404 686134
rect 360804 650454 361404 685898
rect 360804 650218 360986 650454
rect 361222 650218 361404 650454
rect 360804 650134 361404 650218
rect 360804 649898 360986 650134
rect 361222 649898 361404 650134
rect 360804 614454 361404 649898
rect 360804 614218 360986 614454
rect 361222 614218 361404 614454
rect 360804 614134 361404 614218
rect 360804 613898 360986 614134
rect 361222 613898 361404 614134
rect 360804 578454 361404 613898
rect 360804 578218 360986 578454
rect 361222 578218 361404 578454
rect 360804 578134 361404 578218
rect 360804 577898 360986 578134
rect 361222 577898 361404 578134
rect 360804 542454 361404 577898
rect 360804 542218 360986 542454
rect 361222 542218 361404 542454
rect 360804 542134 361404 542218
rect 360804 541898 360986 542134
rect 361222 541898 361404 542134
rect 360804 506454 361404 541898
rect 360804 506218 360986 506454
rect 361222 506218 361404 506454
rect 360804 506134 361404 506218
rect 360804 505898 360986 506134
rect 361222 505898 361404 506134
rect 360804 470454 361404 505898
rect 360804 470218 360986 470454
rect 361222 470218 361404 470454
rect 360804 470134 361404 470218
rect 360804 469898 360986 470134
rect 361222 469898 361404 470134
rect 360804 434454 361404 469898
rect 360804 434218 360986 434454
rect 361222 434218 361404 434454
rect 360804 434134 361404 434218
rect 360804 433898 360986 434134
rect 361222 433898 361404 434134
rect 360804 398454 361404 433898
rect 360804 398218 360986 398454
rect 361222 398218 361404 398454
rect 360804 398134 361404 398218
rect 360804 397898 360986 398134
rect 361222 397898 361404 398134
rect 360804 362454 361404 397898
rect 360804 362218 360986 362454
rect 361222 362218 361404 362454
rect 360804 362134 361404 362218
rect 360804 361898 360986 362134
rect 361222 361898 361404 362134
rect 360804 326454 361404 361898
rect 360804 326218 360986 326454
rect 361222 326218 361404 326454
rect 360804 326134 361404 326218
rect 360804 325898 360986 326134
rect 361222 325898 361404 326134
rect 357387 322148 357453 322149
rect 357387 322084 357388 322148
rect 357452 322084 357453 322148
rect 357387 322083 357453 322084
rect 357390 321741 357450 322083
rect 357387 321740 357453 321741
rect 357387 321676 357388 321740
rect 357452 321676 357453 321740
rect 357387 321675 357453 321676
rect 353604 319018 353786 319254
rect 354022 319018 354204 319254
rect 353604 318934 354204 319018
rect 353604 318698 353786 318934
rect 354022 318698 354204 318934
rect 353604 283254 354204 318698
rect 353604 283018 353786 283254
rect 354022 283018 354204 283254
rect 353604 282934 354204 283018
rect 353604 282698 353786 282934
rect 354022 282698 354204 282934
rect 353604 247254 354204 282698
rect 353604 247018 353786 247254
rect 354022 247018 354204 247254
rect 353604 246934 354204 247018
rect 353604 246698 353786 246934
rect 354022 246698 354204 246934
rect 353604 211254 354204 246698
rect 353604 211018 353786 211254
rect 354022 211018 354204 211254
rect 353604 210934 354204 211018
rect 353604 210698 353786 210934
rect 354022 210698 354204 210934
rect 353604 175254 354204 210698
rect 353604 175018 353786 175254
rect 354022 175018 354204 175254
rect 353604 174934 354204 175018
rect 353604 174698 353786 174934
rect 354022 174698 354204 174934
rect 353604 139254 354204 174698
rect 353604 139018 353786 139254
rect 354022 139018 354204 139254
rect 353604 138934 354204 139018
rect 353604 138698 353786 138934
rect 354022 138698 354204 138934
rect 353604 103254 354204 138698
rect 353604 103018 353786 103254
rect 354022 103018 354204 103254
rect 353604 102934 354204 103018
rect 353604 102698 353786 102934
rect 354022 102698 354204 102934
rect 353604 67254 354204 102698
rect 353604 67018 353786 67254
rect 354022 67018 354204 67254
rect 353604 66934 354204 67018
rect 353604 66698 353786 66934
rect 354022 66698 354204 66934
rect 353604 31254 354204 66698
rect 353604 31018 353786 31254
rect 354022 31018 354204 31254
rect 353604 30934 354204 31018
rect 353604 30698 353786 30934
rect 354022 30698 354204 30934
rect 335604 -6102 335786 -5866
rect 336022 -6102 336204 -5866
rect 335604 -6186 336204 -6102
rect 335604 -6422 335786 -6186
rect 336022 -6422 336204 -6186
rect 335604 -7364 336204 -6422
rect 353604 -6786 354204 30698
rect 360804 290454 361404 325898
rect 360804 290218 360986 290454
rect 361222 290218 361404 290454
rect 360804 290134 361404 290218
rect 360804 289898 360986 290134
rect 361222 289898 361404 290134
rect 360804 254454 361404 289898
rect 360804 254218 360986 254454
rect 361222 254218 361404 254454
rect 360804 254134 361404 254218
rect 360804 253898 360986 254134
rect 361222 253898 361404 254134
rect 360804 218454 361404 253898
rect 360804 218218 360986 218454
rect 361222 218218 361404 218454
rect 360804 218134 361404 218218
rect 360804 217898 360986 218134
rect 361222 217898 361404 218134
rect 360804 182454 361404 217898
rect 360804 182218 360986 182454
rect 361222 182218 361404 182454
rect 360804 182134 361404 182218
rect 360804 181898 360986 182134
rect 361222 181898 361404 182134
rect 360804 146454 361404 181898
rect 360804 146218 360986 146454
rect 361222 146218 361404 146454
rect 360804 146134 361404 146218
rect 360804 145898 360986 146134
rect 361222 145898 361404 146134
rect 360804 110454 361404 145898
rect 360804 110218 360986 110454
rect 361222 110218 361404 110454
rect 360804 110134 361404 110218
rect 360804 109898 360986 110134
rect 361222 109898 361404 110134
rect 360804 74454 361404 109898
rect 360804 74218 360986 74454
rect 361222 74218 361404 74454
rect 360804 74134 361404 74218
rect 360804 73898 360986 74134
rect 361222 73898 361404 74134
rect 360804 38454 361404 73898
rect 360804 38218 360986 38454
rect 361222 38218 361404 38454
rect 360804 38134 361404 38218
rect 360804 37898 360986 38134
rect 361222 37898 361404 38134
rect 360804 2454 361404 37898
rect 360804 2218 360986 2454
rect 361222 2218 361404 2454
rect 360804 2134 361404 2218
rect 360804 1898 360986 2134
rect 361222 1898 361404 2134
rect 360804 -346 361404 1898
rect 360804 -582 360986 -346
rect 361222 -582 361404 -346
rect 360804 -666 361404 -582
rect 360804 -902 360986 -666
rect 361222 -902 361404 -666
rect 360804 -1844 361404 -902
rect 364404 690054 365004 706122
rect 364404 689818 364586 690054
rect 364822 689818 365004 690054
rect 364404 689734 365004 689818
rect 364404 689498 364586 689734
rect 364822 689498 365004 689734
rect 364404 654054 365004 689498
rect 364404 653818 364586 654054
rect 364822 653818 365004 654054
rect 364404 653734 365004 653818
rect 364404 653498 364586 653734
rect 364822 653498 365004 653734
rect 364404 618054 365004 653498
rect 364404 617818 364586 618054
rect 364822 617818 365004 618054
rect 364404 617734 365004 617818
rect 364404 617498 364586 617734
rect 364822 617498 365004 617734
rect 364404 582054 365004 617498
rect 364404 581818 364586 582054
rect 364822 581818 365004 582054
rect 364404 581734 365004 581818
rect 364404 581498 364586 581734
rect 364822 581498 365004 581734
rect 364404 546054 365004 581498
rect 364404 545818 364586 546054
rect 364822 545818 365004 546054
rect 364404 545734 365004 545818
rect 364404 545498 364586 545734
rect 364822 545498 365004 545734
rect 364404 510054 365004 545498
rect 364404 509818 364586 510054
rect 364822 509818 365004 510054
rect 364404 509734 365004 509818
rect 364404 509498 364586 509734
rect 364822 509498 365004 509734
rect 364404 474054 365004 509498
rect 364404 473818 364586 474054
rect 364822 473818 365004 474054
rect 364404 473734 365004 473818
rect 364404 473498 364586 473734
rect 364822 473498 365004 473734
rect 364404 438054 365004 473498
rect 364404 437818 364586 438054
rect 364822 437818 365004 438054
rect 364404 437734 365004 437818
rect 364404 437498 364586 437734
rect 364822 437498 365004 437734
rect 364404 402054 365004 437498
rect 364404 401818 364586 402054
rect 364822 401818 365004 402054
rect 364404 401734 365004 401818
rect 364404 401498 364586 401734
rect 364822 401498 365004 401734
rect 364404 366054 365004 401498
rect 364404 365818 364586 366054
rect 364822 365818 365004 366054
rect 364404 365734 365004 365818
rect 364404 365498 364586 365734
rect 364822 365498 365004 365734
rect 364404 330054 365004 365498
rect 364404 329818 364586 330054
rect 364822 329818 365004 330054
rect 364404 329734 365004 329818
rect 364404 329498 364586 329734
rect 364822 329498 365004 329734
rect 364404 294054 365004 329498
rect 364404 293818 364586 294054
rect 364822 293818 365004 294054
rect 364404 293734 365004 293818
rect 364404 293498 364586 293734
rect 364822 293498 365004 293734
rect 364404 258054 365004 293498
rect 364404 257818 364586 258054
rect 364822 257818 365004 258054
rect 364404 257734 365004 257818
rect 364404 257498 364586 257734
rect 364822 257498 365004 257734
rect 364404 222054 365004 257498
rect 364404 221818 364586 222054
rect 364822 221818 365004 222054
rect 364404 221734 365004 221818
rect 364404 221498 364586 221734
rect 364822 221498 365004 221734
rect 364404 186054 365004 221498
rect 364404 185818 364586 186054
rect 364822 185818 365004 186054
rect 364404 185734 365004 185818
rect 364404 185498 364586 185734
rect 364822 185498 365004 185734
rect 364404 150054 365004 185498
rect 364404 149818 364586 150054
rect 364822 149818 365004 150054
rect 364404 149734 365004 149818
rect 364404 149498 364586 149734
rect 364822 149498 365004 149734
rect 364404 114054 365004 149498
rect 364404 113818 364586 114054
rect 364822 113818 365004 114054
rect 364404 113734 365004 113818
rect 364404 113498 364586 113734
rect 364822 113498 365004 113734
rect 364404 78054 365004 113498
rect 364404 77818 364586 78054
rect 364822 77818 365004 78054
rect 364404 77734 365004 77818
rect 364404 77498 364586 77734
rect 364822 77498 365004 77734
rect 364404 42054 365004 77498
rect 364404 41818 364586 42054
rect 364822 41818 365004 42054
rect 364404 41734 365004 41818
rect 364404 41498 364586 41734
rect 364822 41498 365004 41734
rect 364404 6054 365004 41498
rect 364404 5818 364586 6054
rect 364822 5818 365004 6054
rect 364404 5734 365004 5818
rect 364404 5498 364586 5734
rect 364822 5498 365004 5734
rect 364404 -2186 365004 5498
rect 364404 -2422 364586 -2186
rect 364822 -2422 365004 -2186
rect 364404 -2506 365004 -2422
rect 364404 -2742 364586 -2506
rect 364822 -2742 365004 -2506
rect 364404 -3684 365004 -2742
rect 368004 693654 368604 707962
rect 368004 693418 368186 693654
rect 368422 693418 368604 693654
rect 368004 693334 368604 693418
rect 368004 693098 368186 693334
rect 368422 693098 368604 693334
rect 368004 657654 368604 693098
rect 368004 657418 368186 657654
rect 368422 657418 368604 657654
rect 368004 657334 368604 657418
rect 368004 657098 368186 657334
rect 368422 657098 368604 657334
rect 368004 621654 368604 657098
rect 368004 621418 368186 621654
rect 368422 621418 368604 621654
rect 368004 621334 368604 621418
rect 368004 621098 368186 621334
rect 368422 621098 368604 621334
rect 368004 585654 368604 621098
rect 368004 585418 368186 585654
rect 368422 585418 368604 585654
rect 368004 585334 368604 585418
rect 368004 585098 368186 585334
rect 368422 585098 368604 585334
rect 368004 549654 368604 585098
rect 368004 549418 368186 549654
rect 368422 549418 368604 549654
rect 368004 549334 368604 549418
rect 368004 549098 368186 549334
rect 368422 549098 368604 549334
rect 368004 513654 368604 549098
rect 368004 513418 368186 513654
rect 368422 513418 368604 513654
rect 368004 513334 368604 513418
rect 368004 513098 368186 513334
rect 368422 513098 368604 513334
rect 368004 477654 368604 513098
rect 368004 477418 368186 477654
rect 368422 477418 368604 477654
rect 368004 477334 368604 477418
rect 368004 477098 368186 477334
rect 368422 477098 368604 477334
rect 368004 441654 368604 477098
rect 368004 441418 368186 441654
rect 368422 441418 368604 441654
rect 368004 441334 368604 441418
rect 368004 441098 368186 441334
rect 368422 441098 368604 441334
rect 368004 405654 368604 441098
rect 368004 405418 368186 405654
rect 368422 405418 368604 405654
rect 368004 405334 368604 405418
rect 368004 405098 368186 405334
rect 368422 405098 368604 405334
rect 368004 369654 368604 405098
rect 368004 369418 368186 369654
rect 368422 369418 368604 369654
rect 368004 369334 368604 369418
rect 368004 369098 368186 369334
rect 368422 369098 368604 369334
rect 368004 333654 368604 369098
rect 368004 333418 368186 333654
rect 368422 333418 368604 333654
rect 368004 333334 368604 333418
rect 368004 333098 368186 333334
rect 368422 333098 368604 333334
rect 368004 297654 368604 333098
rect 368004 297418 368186 297654
rect 368422 297418 368604 297654
rect 368004 297334 368604 297418
rect 368004 297098 368186 297334
rect 368422 297098 368604 297334
rect 368004 261654 368604 297098
rect 368004 261418 368186 261654
rect 368422 261418 368604 261654
rect 368004 261334 368604 261418
rect 368004 261098 368186 261334
rect 368422 261098 368604 261334
rect 368004 225654 368604 261098
rect 368004 225418 368186 225654
rect 368422 225418 368604 225654
rect 368004 225334 368604 225418
rect 368004 225098 368186 225334
rect 368422 225098 368604 225334
rect 368004 189654 368604 225098
rect 368004 189418 368186 189654
rect 368422 189418 368604 189654
rect 368004 189334 368604 189418
rect 368004 189098 368186 189334
rect 368422 189098 368604 189334
rect 368004 153654 368604 189098
rect 368004 153418 368186 153654
rect 368422 153418 368604 153654
rect 368004 153334 368604 153418
rect 368004 153098 368186 153334
rect 368422 153098 368604 153334
rect 368004 117654 368604 153098
rect 368004 117418 368186 117654
rect 368422 117418 368604 117654
rect 368004 117334 368604 117418
rect 368004 117098 368186 117334
rect 368422 117098 368604 117334
rect 368004 81654 368604 117098
rect 368004 81418 368186 81654
rect 368422 81418 368604 81654
rect 368004 81334 368604 81418
rect 368004 81098 368186 81334
rect 368422 81098 368604 81334
rect 368004 45654 368604 81098
rect 368004 45418 368186 45654
rect 368422 45418 368604 45654
rect 368004 45334 368604 45418
rect 368004 45098 368186 45334
rect 368422 45098 368604 45334
rect 368004 9654 368604 45098
rect 368004 9418 368186 9654
rect 368422 9418 368604 9654
rect 368004 9334 368604 9418
rect 368004 9098 368186 9334
rect 368422 9098 368604 9334
rect 368004 -4026 368604 9098
rect 368004 -4262 368186 -4026
rect 368422 -4262 368604 -4026
rect 368004 -4346 368604 -4262
rect 368004 -4582 368186 -4346
rect 368422 -4582 368604 -4346
rect 368004 -5524 368604 -4582
rect 371604 697254 372204 709802
rect 389604 711278 390204 711300
rect 389604 711042 389786 711278
rect 390022 711042 390204 711278
rect 389604 710958 390204 711042
rect 389604 710722 389786 710958
rect 390022 710722 390204 710958
rect 386004 709438 386604 709460
rect 386004 709202 386186 709438
rect 386422 709202 386604 709438
rect 386004 709118 386604 709202
rect 386004 708882 386186 709118
rect 386422 708882 386604 709118
rect 382404 707598 383004 707620
rect 382404 707362 382586 707598
rect 382822 707362 383004 707598
rect 382404 707278 383004 707362
rect 382404 707042 382586 707278
rect 382822 707042 383004 707278
rect 371604 697018 371786 697254
rect 372022 697018 372204 697254
rect 371604 696934 372204 697018
rect 371604 696698 371786 696934
rect 372022 696698 372204 696934
rect 371604 661254 372204 696698
rect 371604 661018 371786 661254
rect 372022 661018 372204 661254
rect 371604 660934 372204 661018
rect 371604 660698 371786 660934
rect 372022 660698 372204 660934
rect 371604 625254 372204 660698
rect 371604 625018 371786 625254
rect 372022 625018 372204 625254
rect 371604 624934 372204 625018
rect 371604 624698 371786 624934
rect 372022 624698 372204 624934
rect 371604 589254 372204 624698
rect 371604 589018 371786 589254
rect 372022 589018 372204 589254
rect 371604 588934 372204 589018
rect 371604 588698 371786 588934
rect 372022 588698 372204 588934
rect 371604 553254 372204 588698
rect 371604 553018 371786 553254
rect 372022 553018 372204 553254
rect 371604 552934 372204 553018
rect 371604 552698 371786 552934
rect 372022 552698 372204 552934
rect 371604 517254 372204 552698
rect 371604 517018 371786 517254
rect 372022 517018 372204 517254
rect 371604 516934 372204 517018
rect 371604 516698 371786 516934
rect 372022 516698 372204 516934
rect 371604 481254 372204 516698
rect 371604 481018 371786 481254
rect 372022 481018 372204 481254
rect 371604 480934 372204 481018
rect 371604 480698 371786 480934
rect 372022 480698 372204 480934
rect 371604 445254 372204 480698
rect 371604 445018 371786 445254
rect 372022 445018 372204 445254
rect 371604 444934 372204 445018
rect 371604 444698 371786 444934
rect 372022 444698 372204 444934
rect 371604 409254 372204 444698
rect 371604 409018 371786 409254
rect 372022 409018 372204 409254
rect 371604 408934 372204 409018
rect 371604 408698 371786 408934
rect 372022 408698 372204 408934
rect 371604 373254 372204 408698
rect 371604 373018 371786 373254
rect 372022 373018 372204 373254
rect 371604 372934 372204 373018
rect 371604 372698 371786 372934
rect 372022 372698 372204 372934
rect 371604 337254 372204 372698
rect 371604 337018 371786 337254
rect 372022 337018 372204 337254
rect 371604 336934 372204 337018
rect 371604 336698 371786 336934
rect 372022 336698 372204 336934
rect 371604 301254 372204 336698
rect 371604 301018 371786 301254
rect 372022 301018 372204 301254
rect 371604 300934 372204 301018
rect 371604 300698 371786 300934
rect 372022 300698 372204 300934
rect 371604 265254 372204 300698
rect 371604 265018 371786 265254
rect 372022 265018 372204 265254
rect 371604 264934 372204 265018
rect 371604 264698 371786 264934
rect 372022 264698 372204 264934
rect 371604 229254 372204 264698
rect 371604 229018 371786 229254
rect 372022 229018 372204 229254
rect 371604 228934 372204 229018
rect 371604 228698 371786 228934
rect 372022 228698 372204 228934
rect 371604 193254 372204 228698
rect 371604 193018 371786 193254
rect 372022 193018 372204 193254
rect 371604 192934 372204 193018
rect 371604 192698 371786 192934
rect 372022 192698 372204 192934
rect 371604 157254 372204 192698
rect 371604 157018 371786 157254
rect 372022 157018 372204 157254
rect 371604 156934 372204 157018
rect 371604 156698 371786 156934
rect 372022 156698 372204 156934
rect 371604 121254 372204 156698
rect 371604 121018 371786 121254
rect 372022 121018 372204 121254
rect 371604 120934 372204 121018
rect 371604 120698 371786 120934
rect 372022 120698 372204 120934
rect 371604 85254 372204 120698
rect 371604 85018 371786 85254
rect 372022 85018 372204 85254
rect 371604 84934 372204 85018
rect 371604 84698 371786 84934
rect 372022 84698 372204 84934
rect 371604 49254 372204 84698
rect 371604 49018 371786 49254
rect 372022 49018 372204 49254
rect 371604 48934 372204 49018
rect 371604 48698 371786 48934
rect 372022 48698 372204 48934
rect 371604 13254 372204 48698
rect 371604 13018 371786 13254
rect 372022 13018 372204 13254
rect 371604 12934 372204 13018
rect 371604 12698 371786 12934
rect 372022 12698 372204 12934
rect 353604 -7022 353786 -6786
rect 354022 -7022 354204 -6786
rect 353604 -7106 354204 -7022
rect 353604 -7342 353786 -7106
rect 354022 -7342 354204 -7106
rect 353604 -7364 354204 -7342
rect 371604 -5866 372204 12698
rect 378804 705758 379404 705780
rect 378804 705522 378986 705758
rect 379222 705522 379404 705758
rect 378804 705438 379404 705522
rect 378804 705202 378986 705438
rect 379222 705202 379404 705438
rect 378804 668454 379404 705202
rect 378804 668218 378986 668454
rect 379222 668218 379404 668454
rect 378804 668134 379404 668218
rect 378804 667898 378986 668134
rect 379222 667898 379404 668134
rect 378804 632454 379404 667898
rect 378804 632218 378986 632454
rect 379222 632218 379404 632454
rect 378804 632134 379404 632218
rect 378804 631898 378986 632134
rect 379222 631898 379404 632134
rect 378804 596454 379404 631898
rect 378804 596218 378986 596454
rect 379222 596218 379404 596454
rect 378804 596134 379404 596218
rect 378804 595898 378986 596134
rect 379222 595898 379404 596134
rect 378804 560454 379404 595898
rect 378804 560218 378986 560454
rect 379222 560218 379404 560454
rect 378804 560134 379404 560218
rect 378804 559898 378986 560134
rect 379222 559898 379404 560134
rect 378804 524454 379404 559898
rect 378804 524218 378986 524454
rect 379222 524218 379404 524454
rect 378804 524134 379404 524218
rect 378804 523898 378986 524134
rect 379222 523898 379404 524134
rect 378804 488454 379404 523898
rect 378804 488218 378986 488454
rect 379222 488218 379404 488454
rect 378804 488134 379404 488218
rect 378804 487898 378986 488134
rect 379222 487898 379404 488134
rect 378804 452454 379404 487898
rect 378804 452218 378986 452454
rect 379222 452218 379404 452454
rect 378804 452134 379404 452218
rect 378804 451898 378986 452134
rect 379222 451898 379404 452134
rect 378804 416454 379404 451898
rect 378804 416218 378986 416454
rect 379222 416218 379404 416454
rect 378804 416134 379404 416218
rect 378804 415898 378986 416134
rect 379222 415898 379404 416134
rect 378804 380454 379404 415898
rect 378804 380218 378986 380454
rect 379222 380218 379404 380454
rect 378804 380134 379404 380218
rect 378804 379898 378986 380134
rect 379222 379898 379404 380134
rect 378804 344454 379404 379898
rect 378804 344218 378986 344454
rect 379222 344218 379404 344454
rect 378804 344134 379404 344218
rect 378804 343898 378986 344134
rect 379222 343898 379404 344134
rect 378804 308454 379404 343898
rect 378804 308218 378986 308454
rect 379222 308218 379404 308454
rect 378804 308134 379404 308218
rect 378804 307898 378986 308134
rect 379222 307898 379404 308134
rect 378804 272454 379404 307898
rect 378804 272218 378986 272454
rect 379222 272218 379404 272454
rect 378804 272134 379404 272218
rect 378804 271898 378986 272134
rect 379222 271898 379404 272134
rect 378804 236454 379404 271898
rect 378804 236218 378986 236454
rect 379222 236218 379404 236454
rect 378804 236134 379404 236218
rect 378804 235898 378986 236134
rect 379222 235898 379404 236134
rect 378804 200454 379404 235898
rect 378804 200218 378986 200454
rect 379222 200218 379404 200454
rect 378804 200134 379404 200218
rect 378804 199898 378986 200134
rect 379222 199898 379404 200134
rect 378804 164454 379404 199898
rect 378804 164218 378986 164454
rect 379222 164218 379404 164454
rect 378804 164134 379404 164218
rect 378804 163898 378986 164134
rect 379222 163898 379404 164134
rect 378804 128454 379404 163898
rect 378804 128218 378986 128454
rect 379222 128218 379404 128454
rect 378804 128134 379404 128218
rect 378804 127898 378986 128134
rect 379222 127898 379404 128134
rect 378804 92454 379404 127898
rect 378804 92218 378986 92454
rect 379222 92218 379404 92454
rect 378804 92134 379404 92218
rect 378804 91898 378986 92134
rect 379222 91898 379404 92134
rect 378804 56454 379404 91898
rect 378804 56218 378986 56454
rect 379222 56218 379404 56454
rect 378804 56134 379404 56218
rect 378804 55898 378986 56134
rect 379222 55898 379404 56134
rect 378804 20454 379404 55898
rect 378804 20218 378986 20454
rect 379222 20218 379404 20454
rect 378804 20134 379404 20218
rect 378804 19898 378986 20134
rect 379222 19898 379404 20134
rect 378804 -1266 379404 19898
rect 378804 -1502 378986 -1266
rect 379222 -1502 379404 -1266
rect 378804 -1586 379404 -1502
rect 378804 -1822 378986 -1586
rect 379222 -1822 379404 -1586
rect 378804 -1844 379404 -1822
rect 382404 672054 383004 707042
rect 382404 671818 382586 672054
rect 382822 671818 383004 672054
rect 382404 671734 383004 671818
rect 382404 671498 382586 671734
rect 382822 671498 383004 671734
rect 382404 636054 383004 671498
rect 382404 635818 382586 636054
rect 382822 635818 383004 636054
rect 382404 635734 383004 635818
rect 382404 635498 382586 635734
rect 382822 635498 383004 635734
rect 382404 600054 383004 635498
rect 382404 599818 382586 600054
rect 382822 599818 383004 600054
rect 382404 599734 383004 599818
rect 382404 599498 382586 599734
rect 382822 599498 383004 599734
rect 382404 564054 383004 599498
rect 382404 563818 382586 564054
rect 382822 563818 383004 564054
rect 382404 563734 383004 563818
rect 382404 563498 382586 563734
rect 382822 563498 383004 563734
rect 382404 528054 383004 563498
rect 382404 527818 382586 528054
rect 382822 527818 383004 528054
rect 382404 527734 383004 527818
rect 382404 527498 382586 527734
rect 382822 527498 383004 527734
rect 382404 492054 383004 527498
rect 382404 491818 382586 492054
rect 382822 491818 383004 492054
rect 382404 491734 383004 491818
rect 382404 491498 382586 491734
rect 382822 491498 383004 491734
rect 382404 456054 383004 491498
rect 382404 455818 382586 456054
rect 382822 455818 383004 456054
rect 382404 455734 383004 455818
rect 382404 455498 382586 455734
rect 382822 455498 383004 455734
rect 382404 420054 383004 455498
rect 382404 419818 382586 420054
rect 382822 419818 383004 420054
rect 382404 419734 383004 419818
rect 382404 419498 382586 419734
rect 382822 419498 383004 419734
rect 382404 384054 383004 419498
rect 382404 383818 382586 384054
rect 382822 383818 383004 384054
rect 382404 383734 383004 383818
rect 382404 383498 382586 383734
rect 382822 383498 383004 383734
rect 382404 348054 383004 383498
rect 382404 347818 382586 348054
rect 382822 347818 383004 348054
rect 382404 347734 383004 347818
rect 382404 347498 382586 347734
rect 382822 347498 383004 347734
rect 382404 312054 383004 347498
rect 382404 311818 382586 312054
rect 382822 311818 383004 312054
rect 382404 311734 383004 311818
rect 382404 311498 382586 311734
rect 382822 311498 383004 311734
rect 382404 276054 383004 311498
rect 382404 275818 382586 276054
rect 382822 275818 383004 276054
rect 382404 275734 383004 275818
rect 382404 275498 382586 275734
rect 382822 275498 383004 275734
rect 382404 240054 383004 275498
rect 382404 239818 382586 240054
rect 382822 239818 383004 240054
rect 382404 239734 383004 239818
rect 382404 239498 382586 239734
rect 382822 239498 383004 239734
rect 382404 204054 383004 239498
rect 382404 203818 382586 204054
rect 382822 203818 383004 204054
rect 382404 203734 383004 203818
rect 382404 203498 382586 203734
rect 382822 203498 383004 203734
rect 382404 168054 383004 203498
rect 382404 167818 382586 168054
rect 382822 167818 383004 168054
rect 382404 167734 383004 167818
rect 382404 167498 382586 167734
rect 382822 167498 383004 167734
rect 382404 132054 383004 167498
rect 382404 131818 382586 132054
rect 382822 131818 383004 132054
rect 382404 131734 383004 131818
rect 382404 131498 382586 131734
rect 382822 131498 383004 131734
rect 382404 96054 383004 131498
rect 382404 95818 382586 96054
rect 382822 95818 383004 96054
rect 382404 95734 383004 95818
rect 382404 95498 382586 95734
rect 382822 95498 383004 95734
rect 382404 60054 383004 95498
rect 382404 59818 382586 60054
rect 382822 59818 383004 60054
rect 382404 59734 383004 59818
rect 382404 59498 382586 59734
rect 382822 59498 383004 59734
rect 382404 24054 383004 59498
rect 382404 23818 382586 24054
rect 382822 23818 383004 24054
rect 382404 23734 383004 23818
rect 382404 23498 382586 23734
rect 382822 23498 383004 23734
rect 382404 -3106 383004 23498
rect 382404 -3342 382586 -3106
rect 382822 -3342 383004 -3106
rect 382404 -3426 383004 -3342
rect 382404 -3662 382586 -3426
rect 382822 -3662 383004 -3426
rect 382404 -3684 383004 -3662
rect 386004 675654 386604 708882
rect 386004 675418 386186 675654
rect 386422 675418 386604 675654
rect 386004 675334 386604 675418
rect 386004 675098 386186 675334
rect 386422 675098 386604 675334
rect 386004 639654 386604 675098
rect 386004 639418 386186 639654
rect 386422 639418 386604 639654
rect 386004 639334 386604 639418
rect 386004 639098 386186 639334
rect 386422 639098 386604 639334
rect 386004 603654 386604 639098
rect 386004 603418 386186 603654
rect 386422 603418 386604 603654
rect 386004 603334 386604 603418
rect 386004 603098 386186 603334
rect 386422 603098 386604 603334
rect 386004 567654 386604 603098
rect 386004 567418 386186 567654
rect 386422 567418 386604 567654
rect 386004 567334 386604 567418
rect 386004 567098 386186 567334
rect 386422 567098 386604 567334
rect 386004 531654 386604 567098
rect 386004 531418 386186 531654
rect 386422 531418 386604 531654
rect 386004 531334 386604 531418
rect 386004 531098 386186 531334
rect 386422 531098 386604 531334
rect 386004 495654 386604 531098
rect 386004 495418 386186 495654
rect 386422 495418 386604 495654
rect 386004 495334 386604 495418
rect 386004 495098 386186 495334
rect 386422 495098 386604 495334
rect 386004 459654 386604 495098
rect 386004 459418 386186 459654
rect 386422 459418 386604 459654
rect 386004 459334 386604 459418
rect 386004 459098 386186 459334
rect 386422 459098 386604 459334
rect 386004 423654 386604 459098
rect 386004 423418 386186 423654
rect 386422 423418 386604 423654
rect 386004 423334 386604 423418
rect 386004 423098 386186 423334
rect 386422 423098 386604 423334
rect 386004 387654 386604 423098
rect 386004 387418 386186 387654
rect 386422 387418 386604 387654
rect 386004 387334 386604 387418
rect 386004 387098 386186 387334
rect 386422 387098 386604 387334
rect 386004 351654 386604 387098
rect 386004 351418 386186 351654
rect 386422 351418 386604 351654
rect 386004 351334 386604 351418
rect 386004 351098 386186 351334
rect 386422 351098 386604 351334
rect 386004 315654 386604 351098
rect 386004 315418 386186 315654
rect 386422 315418 386604 315654
rect 386004 315334 386604 315418
rect 386004 315098 386186 315334
rect 386422 315098 386604 315334
rect 386004 279654 386604 315098
rect 386004 279418 386186 279654
rect 386422 279418 386604 279654
rect 386004 279334 386604 279418
rect 386004 279098 386186 279334
rect 386422 279098 386604 279334
rect 386004 243654 386604 279098
rect 386004 243418 386186 243654
rect 386422 243418 386604 243654
rect 386004 243334 386604 243418
rect 386004 243098 386186 243334
rect 386422 243098 386604 243334
rect 386004 207654 386604 243098
rect 386004 207418 386186 207654
rect 386422 207418 386604 207654
rect 386004 207334 386604 207418
rect 386004 207098 386186 207334
rect 386422 207098 386604 207334
rect 386004 171654 386604 207098
rect 386004 171418 386186 171654
rect 386422 171418 386604 171654
rect 386004 171334 386604 171418
rect 386004 171098 386186 171334
rect 386422 171098 386604 171334
rect 386004 135654 386604 171098
rect 386004 135418 386186 135654
rect 386422 135418 386604 135654
rect 386004 135334 386604 135418
rect 386004 135098 386186 135334
rect 386422 135098 386604 135334
rect 386004 99654 386604 135098
rect 386004 99418 386186 99654
rect 386422 99418 386604 99654
rect 386004 99334 386604 99418
rect 386004 99098 386186 99334
rect 386422 99098 386604 99334
rect 386004 63654 386604 99098
rect 386004 63418 386186 63654
rect 386422 63418 386604 63654
rect 386004 63334 386604 63418
rect 386004 63098 386186 63334
rect 386422 63098 386604 63334
rect 386004 27654 386604 63098
rect 386004 27418 386186 27654
rect 386422 27418 386604 27654
rect 386004 27334 386604 27418
rect 386004 27098 386186 27334
rect 386422 27098 386604 27334
rect 386004 -4946 386604 27098
rect 386004 -5182 386186 -4946
rect 386422 -5182 386604 -4946
rect 386004 -5266 386604 -5182
rect 386004 -5502 386186 -5266
rect 386422 -5502 386604 -5266
rect 386004 -5524 386604 -5502
rect 389604 679254 390204 710722
rect 407604 710358 408204 711300
rect 407604 710122 407786 710358
rect 408022 710122 408204 710358
rect 407604 710038 408204 710122
rect 407604 709802 407786 710038
rect 408022 709802 408204 710038
rect 404004 708518 404604 709460
rect 404004 708282 404186 708518
rect 404422 708282 404604 708518
rect 404004 708198 404604 708282
rect 404004 707962 404186 708198
rect 404422 707962 404604 708198
rect 400404 706678 401004 707620
rect 400404 706442 400586 706678
rect 400822 706442 401004 706678
rect 400404 706358 401004 706442
rect 400404 706122 400586 706358
rect 400822 706122 401004 706358
rect 389604 679018 389786 679254
rect 390022 679018 390204 679254
rect 389604 678934 390204 679018
rect 389604 678698 389786 678934
rect 390022 678698 390204 678934
rect 389604 643254 390204 678698
rect 389604 643018 389786 643254
rect 390022 643018 390204 643254
rect 389604 642934 390204 643018
rect 389604 642698 389786 642934
rect 390022 642698 390204 642934
rect 389604 607254 390204 642698
rect 389604 607018 389786 607254
rect 390022 607018 390204 607254
rect 389604 606934 390204 607018
rect 389604 606698 389786 606934
rect 390022 606698 390204 606934
rect 389604 571254 390204 606698
rect 389604 571018 389786 571254
rect 390022 571018 390204 571254
rect 389604 570934 390204 571018
rect 389604 570698 389786 570934
rect 390022 570698 390204 570934
rect 389604 535254 390204 570698
rect 389604 535018 389786 535254
rect 390022 535018 390204 535254
rect 389604 534934 390204 535018
rect 389604 534698 389786 534934
rect 390022 534698 390204 534934
rect 389604 499254 390204 534698
rect 389604 499018 389786 499254
rect 390022 499018 390204 499254
rect 389604 498934 390204 499018
rect 389604 498698 389786 498934
rect 390022 498698 390204 498934
rect 389604 463254 390204 498698
rect 389604 463018 389786 463254
rect 390022 463018 390204 463254
rect 389604 462934 390204 463018
rect 389604 462698 389786 462934
rect 390022 462698 390204 462934
rect 389604 427254 390204 462698
rect 389604 427018 389786 427254
rect 390022 427018 390204 427254
rect 389604 426934 390204 427018
rect 389604 426698 389786 426934
rect 390022 426698 390204 426934
rect 389604 391254 390204 426698
rect 389604 391018 389786 391254
rect 390022 391018 390204 391254
rect 389604 390934 390204 391018
rect 389604 390698 389786 390934
rect 390022 390698 390204 390934
rect 389604 355254 390204 390698
rect 389604 355018 389786 355254
rect 390022 355018 390204 355254
rect 389604 354934 390204 355018
rect 389604 354698 389786 354934
rect 390022 354698 390204 354934
rect 389604 319254 390204 354698
rect 396804 704838 397404 705780
rect 396804 704602 396986 704838
rect 397222 704602 397404 704838
rect 396804 704518 397404 704602
rect 396804 704282 396986 704518
rect 397222 704282 397404 704518
rect 396804 686454 397404 704282
rect 396804 686218 396986 686454
rect 397222 686218 397404 686454
rect 396804 686134 397404 686218
rect 396804 685898 396986 686134
rect 397222 685898 397404 686134
rect 396804 650454 397404 685898
rect 396804 650218 396986 650454
rect 397222 650218 397404 650454
rect 396804 650134 397404 650218
rect 396804 649898 396986 650134
rect 397222 649898 397404 650134
rect 396804 614454 397404 649898
rect 396804 614218 396986 614454
rect 397222 614218 397404 614454
rect 396804 614134 397404 614218
rect 396804 613898 396986 614134
rect 397222 613898 397404 614134
rect 396804 578454 397404 613898
rect 396804 578218 396986 578454
rect 397222 578218 397404 578454
rect 396804 578134 397404 578218
rect 396804 577898 396986 578134
rect 397222 577898 397404 578134
rect 396804 542454 397404 577898
rect 396804 542218 396986 542454
rect 397222 542218 397404 542454
rect 396804 542134 397404 542218
rect 396804 541898 396986 542134
rect 397222 541898 397404 542134
rect 396804 506454 397404 541898
rect 396804 506218 396986 506454
rect 397222 506218 397404 506454
rect 396804 506134 397404 506218
rect 396804 505898 396986 506134
rect 397222 505898 397404 506134
rect 396804 470454 397404 505898
rect 396804 470218 396986 470454
rect 397222 470218 397404 470454
rect 396804 470134 397404 470218
rect 396804 469898 396986 470134
rect 397222 469898 397404 470134
rect 396804 434454 397404 469898
rect 396804 434218 396986 434454
rect 397222 434218 397404 434454
rect 396804 434134 397404 434218
rect 396804 433898 396986 434134
rect 397222 433898 397404 434134
rect 396804 398454 397404 433898
rect 396804 398218 396986 398454
rect 397222 398218 397404 398454
rect 396804 398134 397404 398218
rect 396804 397898 396986 398134
rect 397222 397898 397404 398134
rect 396804 362454 397404 397898
rect 396804 362218 396986 362454
rect 397222 362218 397404 362454
rect 396804 362134 397404 362218
rect 396804 361898 396986 362134
rect 397222 361898 397404 362134
rect 396804 326454 397404 361898
rect 396804 326218 396986 326454
rect 397222 326218 397404 326454
rect 396804 326134 397404 326218
rect 396804 325898 396986 326134
rect 397222 325898 397404 326134
rect 396027 322148 396093 322149
rect 396027 322084 396028 322148
rect 396092 322084 396093 322148
rect 396027 322083 396093 322084
rect 396030 321741 396090 322083
rect 396027 321740 396093 321741
rect 396027 321676 396028 321740
rect 396092 321676 396093 321740
rect 396027 321675 396093 321676
rect 389604 319018 389786 319254
rect 390022 319018 390204 319254
rect 389604 318934 390204 319018
rect 389604 318698 389786 318934
rect 390022 318698 390204 318934
rect 389604 283254 390204 318698
rect 389604 283018 389786 283254
rect 390022 283018 390204 283254
rect 389604 282934 390204 283018
rect 389604 282698 389786 282934
rect 390022 282698 390204 282934
rect 389604 247254 390204 282698
rect 389604 247018 389786 247254
rect 390022 247018 390204 247254
rect 389604 246934 390204 247018
rect 389604 246698 389786 246934
rect 390022 246698 390204 246934
rect 389604 211254 390204 246698
rect 389604 211018 389786 211254
rect 390022 211018 390204 211254
rect 389604 210934 390204 211018
rect 389604 210698 389786 210934
rect 390022 210698 390204 210934
rect 389604 175254 390204 210698
rect 389604 175018 389786 175254
rect 390022 175018 390204 175254
rect 389604 174934 390204 175018
rect 389604 174698 389786 174934
rect 390022 174698 390204 174934
rect 389604 139254 390204 174698
rect 389604 139018 389786 139254
rect 390022 139018 390204 139254
rect 389604 138934 390204 139018
rect 389604 138698 389786 138934
rect 390022 138698 390204 138934
rect 389604 103254 390204 138698
rect 389604 103018 389786 103254
rect 390022 103018 390204 103254
rect 389604 102934 390204 103018
rect 389604 102698 389786 102934
rect 390022 102698 390204 102934
rect 389604 67254 390204 102698
rect 389604 67018 389786 67254
rect 390022 67018 390204 67254
rect 389604 66934 390204 67018
rect 389604 66698 389786 66934
rect 390022 66698 390204 66934
rect 389604 31254 390204 66698
rect 389604 31018 389786 31254
rect 390022 31018 390204 31254
rect 389604 30934 390204 31018
rect 389604 30698 389786 30934
rect 390022 30698 390204 30934
rect 371604 -6102 371786 -5866
rect 372022 -6102 372204 -5866
rect 371604 -6186 372204 -6102
rect 371604 -6422 371786 -6186
rect 372022 -6422 372204 -6186
rect 371604 -7364 372204 -6422
rect 389604 -6786 390204 30698
rect 396804 290454 397404 325898
rect 396804 290218 396986 290454
rect 397222 290218 397404 290454
rect 396804 290134 397404 290218
rect 396804 289898 396986 290134
rect 397222 289898 397404 290134
rect 396804 254454 397404 289898
rect 396804 254218 396986 254454
rect 397222 254218 397404 254454
rect 396804 254134 397404 254218
rect 396804 253898 396986 254134
rect 397222 253898 397404 254134
rect 396804 218454 397404 253898
rect 396804 218218 396986 218454
rect 397222 218218 397404 218454
rect 396804 218134 397404 218218
rect 396804 217898 396986 218134
rect 397222 217898 397404 218134
rect 396804 182454 397404 217898
rect 396804 182218 396986 182454
rect 397222 182218 397404 182454
rect 396804 182134 397404 182218
rect 396804 181898 396986 182134
rect 397222 181898 397404 182134
rect 396804 146454 397404 181898
rect 396804 146218 396986 146454
rect 397222 146218 397404 146454
rect 396804 146134 397404 146218
rect 396804 145898 396986 146134
rect 397222 145898 397404 146134
rect 396804 110454 397404 145898
rect 396804 110218 396986 110454
rect 397222 110218 397404 110454
rect 396804 110134 397404 110218
rect 396804 109898 396986 110134
rect 397222 109898 397404 110134
rect 396804 74454 397404 109898
rect 396804 74218 396986 74454
rect 397222 74218 397404 74454
rect 396804 74134 397404 74218
rect 396804 73898 396986 74134
rect 397222 73898 397404 74134
rect 396804 38454 397404 73898
rect 396804 38218 396986 38454
rect 397222 38218 397404 38454
rect 396804 38134 397404 38218
rect 396804 37898 396986 38134
rect 397222 37898 397404 38134
rect 396804 2454 397404 37898
rect 396804 2218 396986 2454
rect 397222 2218 397404 2454
rect 396804 2134 397404 2218
rect 396804 1898 396986 2134
rect 397222 1898 397404 2134
rect 396804 -346 397404 1898
rect 396804 -582 396986 -346
rect 397222 -582 397404 -346
rect 396804 -666 397404 -582
rect 396804 -902 396986 -666
rect 397222 -902 397404 -666
rect 396804 -1844 397404 -902
rect 400404 690054 401004 706122
rect 400404 689818 400586 690054
rect 400822 689818 401004 690054
rect 400404 689734 401004 689818
rect 400404 689498 400586 689734
rect 400822 689498 401004 689734
rect 400404 654054 401004 689498
rect 400404 653818 400586 654054
rect 400822 653818 401004 654054
rect 400404 653734 401004 653818
rect 400404 653498 400586 653734
rect 400822 653498 401004 653734
rect 400404 618054 401004 653498
rect 400404 617818 400586 618054
rect 400822 617818 401004 618054
rect 400404 617734 401004 617818
rect 400404 617498 400586 617734
rect 400822 617498 401004 617734
rect 400404 582054 401004 617498
rect 400404 581818 400586 582054
rect 400822 581818 401004 582054
rect 400404 581734 401004 581818
rect 400404 581498 400586 581734
rect 400822 581498 401004 581734
rect 400404 546054 401004 581498
rect 400404 545818 400586 546054
rect 400822 545818 401004 546054
rect 400404 545734 401004 545818
rect 400404 545498 400586 545734
rect 400822 545498 401004 545734
rect 400404 510054 401004 545498
rect 400404 509818 400586 510054
rect 400822 509818 401004 510054
rect 400404 509734 401004 509818
rect 400404 509498 400586 509734
rect 400822 509498 401004 509734
rect 400404 474054 401004 509498
rect 400404 473818 400586 474054
rect 400822 473818 401004 474054
rect 400404 473734 401004 473818
rect 400404 473498 400586 473734
rect 400822 473498 401004 473734
rect 400404 438054 401004 473498
rect 400404 437818 400586 438054
rect 400822 437818 401004 438054
rect 400404 437734 401004 437818
rect 400404 437498 400586 437734
rect 400822 437498 401004 437734
rect 400404 402054 401004 437498
rect 400404 401818 400586 402054
rect 400822 401818 401004 402054
rect 400404 401734 401004 401818
rect 400404 401498 400586 401734
rect 400822 401498 401004 401734
rect 400404 366054 401004 401498
rect 400404 365818 400586 366054
rect 400822 365818 401004 366054
rect 400404 365734 401004 365818
rect 400404 365498 400586 365734
rect 400822 365498 401004 365734
rect 400404 330054 401004 365498
rect 400404 329818 400586 330054
rect 400822 329818 401004 330054
rect 400404 329734 401004 329818
rect 400404 329498 400586 329734
rect 400822 329498 401004 329734
rect 400404 294054 401004 329498
rect 400404 293818 400586 294054
rect 400822 293818 401004 294054
rect 400404 293734 401004 293818
rect 400404 293498 400586 293734
rect 400822 293498 401004 293734
rect 400404 258054 401004 293498
rect 400404 257818 400586 258054
rect 400822 257818 401004 258054
rect 400404 257734 401004 257818
rect 400404 257498 400586 257734
rect 400822 257498 401004 257734
rect 400404 222054 401004 257498
rect 400404 221818 400586 222054
rect 400822 221818 401004 222054
rect 400404 221734 401004 221818
rect 400404 221498 400586 221734
rect 400822 221498 401004 221734
rect 400404 186054 401004 221498
rect 400404 185818 400586 186054
rect 400822 185818 401004 186054
rect 400404 185734 401004 185818
rect 400404 185498 400586 185734
rect 400822 185498 401004 185734
rect 400404 150054 401004 185498
rect 400404 149818 400586 150054
rect 400822 149818 401004 150054
rect 400404 149734 401004 149818
rect 400404 149498 400586 149734
rect 400822 149498 401004 149734
rect 400404 114054 401004 149498
rect 400404 113818 400586 114054
rect 400822 113818 401004 114054
rect 400404 113734 401004 113818
rect 400404 113498 400586 113734
rect 400822 113498 401004 113734
rect 400404 78054 401004 113498
rect 400404 77818 400586 78054
rect 400822 77818 401004 78054
rect 400404 77734 401004 77818
rect 400404 77498 400586 77734
rect 400822 77498 401004 77734
rect 400404 42054 401004 77498
rect 400404 41818 400586 42054
rect 400822 41818 401004 42054
rect 400404 41734 401004 41818
rect 400404 41498 400586 41734
rect 400822 41498 401004 41734
rect 400404 6054 401004 41498
rect 400404 5818 400586 6054
rect 400822 5818 401004 6054
rect 400404 5734 401004 5818
rect 400404 5498 400586 5734
rect 400822 5498 401004 5734
rect 400404 -2186 401004 5498
rect 400404 -2422 400586 -2186
rect 400822 -2422 401004 -2186
rect 400404 -2506 401004 -2422
rect 400404 -2742 400586 -2506
rect 400822 -2742 401004 -2506
rect 400404 -3684 401004 -2742
rect 404004 693654 404604 707962
rect 404004 693418 404186 693654
rect 404422 693418 404604 693654
rect 404004 693334 404604 693418
rect 404004 693098 404186 693334
rect 404422 693098 404604 693334
rect 404004 657654 404604 693098
rect 404004 657418 404186 657654
rect 404422 657418 404604 657654
rect 404004 657334 404604 657418
rect 404004 657098 404186 657334
rect 404422 657098 404604 657334
rect 404004 621654 404604 657098
rect 404004 621418 404186 621654
rect 404422 621418 404604 621654
rect 404004 621334 404604 621418
rect 404004 621098 404186 621334
rect 404422 621098 404604 621334
rect 404004 585654 404604 621098
rect 404004 585418 404186 585654
rect 404422 585418 404604 585654
rect 404004 585334 404604 585418
rect 404004 585098 404186 585334
rect 404422 585098 404604 585334
rect 404004 549654 404604 585098
rect 404004 549418 404186 549654
rect 404422 549418 404604 549654
rect 404004 549334 404604 549418
rect 404004 549098 404186 549334
rect 404422 549098 404604 549334
rect 404004 513654 404604 549098
rect 404004 513418 404186 513654
rect 404422 513418 404604 513654
rect 404004 513334 404604 513418
rect 404004 513098 404186 513334
rect 404422 513098 404604 513334
rect 404004 477654 404604 513098
rect 404004 477418 404186 477654
rect 404422 477418 404604 477654
rect 404004 477334 404604 477418
rect 404004 477098 404186 477334
rect 404422 477098 404604 477334
rect 404004 441654 404604 477098
rect 404004 441418 404186 441654
rect 404422 441418 404604 441654
rect 404004 441334 404604 441418
rect 404004 441098 404186 441334
rect 404422 441098 404604 441334
rect 404004 405654 404604 441098
rect 404004 405418 404186 405654
rect 404422 405418 404604 405654
rect 404004 405334 404604 405418
rect 404004 405098 404186 405334
rect 404422 405098 404604 405334
rect 404004 369654 404604 405098
rect 404004 369418 404186 369654
rect 404422 369418 404604 369654
rect 404004 369334 404604 369418
rect 404004 369098 404186 369334
rect 404422 369098 404604 369334
rect 404004 333654 404604 369098
rect 404004 333418 404186 333654
rect 404422 333418 404604 333654
rect 404004 333334 404604 333418
rect 404004 333098 404186 333334
rect 404422 333098 404604 333334
rect 404004 297654 404604 333098
rect 404004 297418 404186 297654
rect 404422 297418 404604 297654
rect 404004 297334 404604 297418
rect 404004 297098 404186 297334
rect 404422 297098 404604 297334
rect 404004 261654 404604 297098
rect 404004 261418 404186 261654
rect 404422 261418 404604 261654
rect 404004 261334 404604 261418
rect 404004 261098 404186 261334
rect 404422 261098 404604 261334
rect 404004 225654 404604 261098
rect 404004 225418 404186 225654
rect 404422 225418 404604 225654
rect 404004 225334 404604 225418
rect 404004 225098 404186 225334
rect 404422 225098 404604 225334
rect 404004 189654 404604 225098
rect 404004 189418 404186 189654
rect 404422 189418 404604 189654
rect 404004 189334 404604 189418
rect 404004 189098 404186 189334
rect 404422 189098 404604 189334
rect 404004 153654 404604 189098
rect 404004 153418 404186 153654
rect 404422 153418 404604 153654
rect 404004 153334 404604 153418
rect 404004 153098 404186 153334
rect 404422 153098 404604 153334
rect 404004 117654 404604 153098
rect 404004 117418 404186 117654
rect 404422 117418 404604 117654
rect 404004 117334 404604 117418
rect 404004 117098 404186 117334
rect 404422 117098 404604 117334
rect 404004 81654 404604 117098
rect 404004 81418 404186 81654
rect 404422 81418 404604 81654
rect 404004 81334 404604 81418
rect 404004 81098 404186 81334
rect 404422 81098 404604 81334
rect 404004 45654 404604 81098
rect 404004 45418 404186 45654
rect 404422 45418 404604 45654
rect 404004 45334 404604 45418
rect 404004 45098 404186 45334
rect 404422 45098 404604 45334
rect 404004 9654 404604 45098
rect 404004 9418 404186 9654
rect 404422 9418 404604 9654
rect 404004 9334 404604 9418
rect 404004 9098 404186 9334
rect 404422 9098 404604 9334
rect 404004 -4026 404604 9098
rect 404004 -4262 404186 -4026
rect 404422 -4262 404604 -4026
rect 404004 -4346 404604 -4262
rect 404004 -4582 404186 -4346
rect 404422 -4582 404604 -4346
rect 404004 -5524 404604 -4582
rect 407604 697254 408204 709802
rect 425604 711278 426204 711300
rect 425604 711042 425786 711278
rect 426022 711042 426204 711278
rect 425604 710958 426204 711042
rect 425604 710722 425786 710958
rect 426022 710722 426204 710958
rect 422004 709438 422604 709460
rect 422004 709202 422186 709438
rect 422422 709202 422604 709438
rect 422004 709118 422604 709202
rect 422004 708882 422186 709118
rect 422422 708882 422604 709118
rect 418404 707598 419004 707620
rect 418404 707362 418586 707598
rect 418822 707362 419004 707598
rect 418404 707278 419004 707362
rect 418404 707042 418586 707278
rect 418822 707042 419004 707278
rect 407604 697018 407786 697254
rect 408022 697018 408204 697254
rect 407604 696934 408204 697018
rect 407604 696698 407786 696934
rect 408022 696698 408204 696934
rect 407604 661254 408204 696698
rect 407604 661018 407786 661254
rect 408022 661018 408204 661254
rect 407604 660934 408204 661018
rect 407604 660698 407786 660934
rect 408022 660698 408204 660934
rect 407604 625254 408204 660698
rect 407604 625018 407786 625254
rect 408022 625018 408204 625254
rect 407604 624934 408204 625018
rect 407604 624698 407786 624934
rect 408022 624698 408204 624934
rect 407604 589254 408204 624698
rect 407604 589018 407786 589254
rect 408022 589018 408204 589254
rect 407604 588934 408204 589018
rect 407604 588698 407786 588934
rect 408022 588698 408204 588934
rect 407604 553254 408204 588698
rect 407604 553018 407786 553254
rect 408022 553018 408204 553254
rect 407604 552934 408204 553018
rect 407604 552698 407786 552934
rect 408022 552698 408204 552934
rect 407604 517254 408204 552698
rect 407604 517018 407786 517254
rect 408022 517018 408204 517254
rect 407604 516934 408204 517018
rect 407604 516698 407786 516934
rect 408022 516698 408204 516934
rect 407604 481254 408204 516698
rect 407604 481018 407786 481254
rect 408022 481018 408204 481254
rect 407604 480934 408204 481018
rect 407604 480698 407786 480934
rect 408022 480698 408204 480934
rect 407604 445254 408204 480698
rect 407604 445018 407786 445254
rect 408022 445018 408204 445254
rect 407604 444934 408204 445018
rect 407604 444698 407786 444934
rect 408022 444698 408204 444934
rect 407604 409254 408204 444698
rect 407604 409018 407786 409254
rect 408022 409018 408204 409254
rect 407604 408934 408204 409018
rect 407604 408698 407786 408934
rect 408022 408698 408204 408934
rect 407604 373254 408204 408698
rect 407604 373018 407786 373254
rect 408022 373018 408204 373254
rect 407604 372934 408204 373018
rect 407604 372698 407786 372934
rect 408022 372698 408204 372934
rect 407604 337254 408204 372698
rect 407604 337018 407786 337254
rect 408022 337018 408204 337254
rect 407604 336934 408204 337018
rect 407604 336698 407786 336934
rect 408022 336698 408204 336934
rect 407604 301254 408204 336698
rect 407604 301018 407786 301254
rect 408022 301018 408204 301254
rect 407604 300934 408204 301018
rect 407604 300698 407786 300934
rect 408022 300698 408204 300934
rect 407604 265254 408204 300698
rect 407604 265018 407786 265254
rect 408022 265018 408204 265254
rect 407604 264934 408204 265018
rect 407604 264698 407786 264934
rect 408022 264698 408204 264934
rect 407604 229254 408204 264698
rect 407604 229018 407786 229254
rect 408022 229018 408204 229254
rect 407604 228934 408204 229018
rect 407604 228698 407786 228934
rect 408022 228698 408204 228934
rect 407604 193254 408204 228698
rect 407604 193018 407786 193254
rect 408022 193018 408204 193254
rect 407604 192934 408204 193018
rect 407604 192698 407786 192934
rect 408022 192698 408204 192934
rect 407604 157254 408204 192698
rect 407604 157018 407786 157254
rect 408022 157018 408204 157254
rect 407604 156934 408204 157018
rect 407604 156698 407786 156934
rect 408022 156698 408204 156934
rect 407604 121254 408204 156698
rect 407604 121018 407786 121254
rect 408022 121018 408204 121254
rect 407604 120934 408204 121018
rect 407604 120698 407786 120934
rect 408022 120698 408204 120934
rect 407604 85254 408204 120698
rect 407604 85018 407786 85254
rect 408022 85018 408204 85254
rect 407604 84934 408204 85018
rect 407604 84698 407786 84934
rect 408022 84698 408204 84934
rect 407604 49254 408204 84698
rect 407604 49018 407786 49254
rect 408022 49018 408204 49254
rect 407604 48934 408204 49018
rect 407604 48698 407786 48934
rect 408022 48698 408204 48934
rect 407604 13254 408204 48698
rect 407604 13018 407786 13254
rect 408022 13018 408204 13254
rect 407604 12934 408204 13018
rect 407604 12698 407786 12934
rect 408022 12698 408204 12934
rect 389604 -7022 389786 -6786
rect 390022 -7022 390204 -6786
rect 389604 -7106 390204 -7022
rect 389604 -7342 389786 -7106
rect 390022 -7342 390204 -7106
rect 389604 -7364 390204 -7342
rect 407604 -5866 408204 12698
rect 414804 705758 415404 705780
rect 414804 705522 414986 705758
rect 415222 705522 415404 705758
rect 414804 705438 415404 705522
rect 414804 705202 414986 705438
rect 415222 705202 415404 705438
rect 414804 668454 415404 705202
rect 414804 668218 414986 668454
rect 415222 668218 415404 668454
rect 414804 668134 415404 668218
rect 414804 667898 414986 668134
rect 415222 667898 415404 668134
rect 414804 632454 415404 667898
rect 414804 632218 414986 632454
rect 415222 632218 415404 632454
rect 414804 632134 415404 632218
rect 414804 631898 414986 632134
rect 415222 631898 415404 632134
rect 414804 596454 415404 631898
rect 414804 596218 414986 596454
rect 415222 596218 415404 596454
rect 414804 596134 415404 596218
rect 414804 595898 414986 596134
rect 415222 595898 415404 596134
rect 414804 560454 415404 595898
rect 414804 560218 414986 560454
rect 415222 560218 415404 560454
rect 414804 560134 415404 560218
rect 414804 559898 414986 560134
rect 415222 559898 415404 560134
rect 414804 524454 415404 559898
rect 414804 524218 414986 524454
rect 415222 524218 415404 524454
rect 414804 524134 415404 524218
rect 414804 523898 414986 524134
rect 415222 523898 415404 524134
rect 414804 488454 415404 523898
rect 414804 488218 414986 488454
rect 415222 488218 415404 488454
rect 414804 488134 415404 488218
rect 414804 487898 414986 488134
rect 415222 487898 415404 488134
rect 414804 452454 415404 487898
rect 414804 452218 414986 452454
rect 415222 452218 415404 452454
rect 414804 452134 415404 452218
rect 414804 451898 414986 452134
rect 415222 451898 415404 452134
rect 414804 416454 415404 451898
rect 414804 416218 414986 416454
rect 415222 416218 415404 416454
rect 414804 416134 415404 416218
rect 414804 415898 414986 416134
rect 415222 415898 415404 416134
rect 414804 380454 415404 415898
rect 414804 380218 414986 380454
rect 415222 380218 415404 380454
rect 414804 380134 415404 380218
rect 414804 379898 414986 380134
rect 415222 379898 415404 380134
rect 414804 344454 415404 379898
rect 414804 344218 414986 344454
rect 415222 344218 415404 344454
rect 414804 344134 415404 344218
rect 414804 343898 414986 344134
rect 415222 343898 415404 344134
rect 414804 308454 415404 343898
rect 414804 308218 414986 308454
rect 415222 308218 415404 308454
rect 414804 308134 415404 308218
rect 414804 307898 414986 308134
rect 415222 307898 415404 308134
rect 414804 272454 415404 307898
rect 414804 272218 414986 272454
rect 415222 272218 415404 272454
rect 414804 272134 415404 272218
rect 414804 271898 414986 272134
rect 415222 271898 415404 272134
rect 414804 236454 415404 271898
rect 414804 236218 414986 236454
rect 415222 236218 415404 236454
rect 414804 236134 415404 236218
rect 414804 235898 414986 236134
rect 415222 235898 415404 236134
rect 414804 200454 415404 235898
rect 414804 200218 414986 200454
rect 415222 200218 415404 200454
rect 414804 200134 415404 200218
rect 414804 199898 414986 200134
rect 415222 199898 415404 200134
rect 414804 164454 415404 199898
rect 414804 164218 414986 164454
rect 415222 164218 415404 164454
rect 414804 164134 415404 164218
rect 414804 163898 414986 164134
rect 415222 163898 415404 164134
rect 414804 128454 415404 163898
rect 414804 128218 414986 128454
rect 415222 128218 415404 128454
rect 414804 128134 415404 128218
rect 414804 127898 414986 128134
rect 415222 127898 415404 128134
rect 414804 92454 415404 127898
rect 414804 92218 414986 92454
rect 415222 92218 415404 92454
rect 414804 92134 415404 92218
rect 414804 91898 414986 92134
rect 415222 91898 415404 92134
rect 414804 56454 415404 91898
rect 414804 56218 414986 56454
rect 415222 56218 415404 56454
rect 414804 56134 415404 56218
rect 414804 55898 414986 56134
rect 415222 55898 415404 56134
rect 414804 20454 415404 55898
rect 414804 20218 414986 20454
rect 415222 20218 415404 20454
rect 414804 20134 415404 20218
rect 414804 19898 414986 20134
rect 415222 19898 415404 20134
rect 414804 -1266 415404 19898
rect 414804 -1502 414986 -1266
rect 415222 -1502 415404 -1266
rect 414804 -1586 415404 -1502
rect 414804 -1822 414986 -1586
rect 415222 -1822 415404 -1586
rect 414804 -1844 415404 -1822
rect 418404 672054 419004 707042
rect 418404 671818 418586 672054
rect 418822 671818 419004 672054
rect 418404 671734 419004 671818
rect 418404 671498 418586 671734
rect 418822 671498 419004 671734
rect 418404 636054 419004 671498
rect 418404 635818 418586 636054
rect 418822 635818 419004 636054
rect 418404 635734 419004 635818
rect 418404 635498 418586 635734
rect 418822 635498 419004 635734
rect 418404 600054 419004 635498
rect 418404 599818 418586 600054
rect 418822 599818 419004 600054
rect 418404 599734 419004 599818
rect 418404 599498 418586 599734
rect 418822 599498 419004 599734
rect 418404 564054 419004 599498
rect 418404 563818 418586 564054
rect 418822 563818 419004 564054
rect 418404 563734 419004 563818
rect 418404 563498 418586 563734
rect 418822 563498 419004 563734
rect 418404 528054 419004 563498
rect 418404 527818 418586 528054
rect 418822 527818 419004 528054
rect 418404 527734 419004 527818
rect 418404 527498 418586 527734
rect 418822 527498 419004 527734
rect 418404 492054 419004 527498
rect 418404 491818 418586 492054
rect 418822 491818 419004 492054
rect 418404 491734 419004 491818
rect 418404 491498 418586 491734
rect 418822 491498 419004 491734
rect 418404 456054 419004 491498
rect 418404 455818 418586 456054
rect 418822 455818 419004 456054
rect 418404 455734 419004 455818
rect 418404 455498 418586 455734
rect 418822 455498 419004 455734
rect 418404 420054 419004 455498
rect 418404 419818 418586 420054
rect 418822 419818 419004 420054
rect 418404 419734 419004 419818
rect 418404 419498 418586 419734
rect 418822 419498 419004 419734
rect 418404 384054 419004 419498
rect 418404 383818 418586 384054
rect 418822 383818 419004 384054
rect 418404 383734 419004 383818
rect 418404 383498 418586 383734
rect 418822 383498 419004 383734
rect 418404 348054 419004 383498
rect 418404 347818 418586 348054
rect 418822 347818 419004 348054
rect 418404 347734 419004 347818
rect 418404 347498 418586 347734
rect 418822 347498 419004 347734
rect 418404 312054 419004 347498
rect 418404 311818 418586 312054
rect 418822 311818 419004 312054
rect 418404 311734 419004 311818
rect 418404 311498 418586 311734
rect 418822 311498 419004 311734
rect 418404 276054 419004 311498
rect 418404 275818 418586 276054
rect 418822 275818 419004 276054
rect 418404 275734 419004 275818
rect 418404 275498 418586 275734
rect 418822 275498 419004 275734
rect 418404 240054 419004 275498
rect 418404 239818 418586 240054
rect 418822 239818 419004 240054
rect 418404 239734 419004 239818
rect 418404 239498 418586 239734
rect 418822 239498 419004 239734
rect 418404 204054 419004 239498
rect 418404 203818 418586 204054
rect 418822 203818 419004 204054
rect 418404 203734 419004 203818
rect 418404 203498 418586 203734
rect 418822 203498 419004 203734
rect 418404 168054 419004 203498
rect 418404 167818 418586 168054
rect 418822 167818 419004 168054
rect 418404 167734 419004 167818
rect 418404 167498 418586 167734
rect 418822 167498 419004 167734
rect 418404 132054 419004 167498
rect 418404 131818 418586 132054
rect 418822 131818 419004 132054
rect 418404 131734 419004 131818
rect 418404 131498 418586 131734
rect 418822 131498 419004 131734
rect 418404 96054 419004 131498
rect 418404 95818 418586 96054
rect 418822 95818 419004 96054
rect 418404 95734 419004 95818
rect 418404 95498 418586 95734
rect 418822 95498 419004 95734
rect 418404 60054 419004 95498
rect 418404 59818 418586 60054
rect 418822 59818 419004 60054
rect 418404 59734 419004 59818
rect 418404 59498 418586 59734
rect 418822 59498 419004 59734
rect 418404 24054 419004 59498
rect 418404 23818 418586 24054
rect 418822 23818 419004 24054
rect 418404 23734 419004 23818
rect 418404 23498 418586 23734
rect 418822 23498 419004 23734
rect 418404 -3106 419004 23498
rect 418404 -3342 418586 -3106
rect 418822 -3342 419004 -3106
rect 418404 -3426 419004 -3342
rect 418404 -3662 418586 -3426
rect 418822 -3662 419004 -3426
rect 418404 -3684 419004 -3662
rect 422004 675654 422604 708882
rect 422004 675418 422186 675654
rect 422422 675418 422604 675654
rect 422004 675334 422604 675418
rect 422004 675098 422186 675334
rect 422422 675098 422604 675334
rect 422004 639654 422604 675098
rect 422004 639418 422186 639654
rect 422422 639418 422604 639654
rect 422004 639334 422604 639418
rect 422004 639098 422186 639334
rect 422422 639098 422604 639334
rect 422004 603654 422604 639098
rect 422004 603418 422186 603654
rect 422422 603418 422604 603654
rect 422004 603334 422604 603418
rect 422004 603098 422186 603334
rect 422422 603098 422604 603334
rect 422004 567654 422604 603098
rect 422004 567418 422186 567654
rect 422422 567418 422604 567654
rect 422004 567334 422604 567418
rect 422004 567098 422186 567334
rect 422422 567098 422604 567334
rect 422004 531654 422604 567098
rect 422004 531418 422186 531654
rect 422422 531418 422604 531654
rect 422004 531334 422604 531418
rect 422004 531098 422186 531334
rect 422422 531098 422604 531334
rect 422004 495654 422604 531098
rect 422004 495418 422186 495654
rect 422422 495418 422604 495654
rect 422004 495334 422604 495418
rect 422004 495098 422186 495334
rect 422422 495098 422604 495334
rect 422004 459654 422604 495098
rect 422004 459418 422186 459654
rect 422422 459418 422604 459654
rect 422004 459334 422604 459418
rect 422004 459098 422186 459334
rect 422422 459098 422604 459334
rect 422004 423654 422604 459098
rect 422004 423418 422186 423654
rect 422422 423418 422604 423654
rect 422004 423334 422604 423418
rect 422004 423098 422186 423334
rect 422422 423098 422604 423334
rect 422004 387654 422604 423098
rect 422004 387418 422186 387654
rect 422422 387418 422604 387654
rect 422004 387334 422604 387418
rect 422004 387098 422186 387334
rect 422422 387098 422604 387334
rect 422004 351654 422604 387098
rect 422004 351418 422186 351654
rect 422422 351418 422604 351654
rect 422004 351334 422604 351418
rect 422004 351098 422186 351334
rect 422422 351098 422604 351334
rect 422004 315654 422604 351098
rect 422004 315418 422186 315654
rect 422422 315418 422604 315654
rect 422004 315334 422604 315418
rect 422004 315098 422186 315334
rect 422422 315098 422604 315334
rect 422004 279654 422604 315098
rect 422004 279418 422186 279654
rect 422422 279418 422604 279654
rect 422004 279334 422604 279418
rect 422004 279098 422186 279334
rect 422422 279098 422604 279334
rect 422004 243654 422604 279098
rect 422004 243418 422186 243654
rect 422422 243418 422604 243654
rect 422004 243334 422604 243418
rect 422004 243098 422186 243334
rect 422422 243098 422604 243334
rect 422004 207654 422604 243098
rect 422004 207418 422186 207654
rect 422422 207418 422604 207654
rect 422004 207334 422604 207418
rect 422004 207098 422186 207334
rect 422422 207098 422604 207334
rect 422004 171654 422604 207098
rect 422004 171418 422186 171654
rect 422422 171418 422604 171654
rect 422004 171334 422604 171418
rect 422004 171098 422186 171334
rect 422422 171098 422604 171334
rect 422004 135654 422604 171098
rect 422004 135418 422186 135654
rect 422422 135418 422604 135654
rect 422004 135334 422604 135418
rect 422004 135098 422186 135334
rect 422422 135098 422604 135334
rect 422004 99654 422604 135098
rect 422004 99418 422186 99654
rect 422422 99418 422604 99654
rect 422004 99334 422604 99418
rect 422004 99098 422186 99334
rect 422422 99098 422604 99334
rect 422004 63654 422604 99098
rect 422004 63418 422186 63654
rect 422422 63418 422604 63654
rect 422004 63334 422604 63418
rect 422004 63098 422186 63334
rect 422422 63098 422604 63334
rect 422004 27654 422604 63098
rect 422004 27418 422186 27654
rect 422422 27418 422604 27654
rect 422004 27334 422604 27418
rect 422004 27098 422186 27334
rect 422422 27098 422604 27334
rect 422004 -4946 422604 27098
rect 422004 -5182 422186 -4946
rect 422422 -5182 422604 -4946
rect 422004 -5266 422604 -5182
rect 422004 -5502 422186 -5266
rect 422422 -5502 422604 -5266
rect 422004 -5524 422604 -5502
rect 425604 679254 426204 710722
rect 443604 710358 444204 711300
rect 443604 710122 443786 710358
rect 444022 710122 444204 710358
rect 443604 710038 444204 710122
rect 443604 709802 443786 710038
rect 444022 709802 444204 710038
rect 440004 708518 440604 709460
rect 440004 708282 440186 708518
rect 440422 708282 440604 708518
rect 440004 708198 440604 708282
rect 440004 707962 440186 708198
rect 440422 707962 440604 708198
rect 436404 706678 437004 707620
rect 436404 706442 436586 706678
rect 436822 706442 437004 706678
rect 436404 706358 437004 706442
rect 436404 706122 436586 706358
rect 436822 706122 437004 706358
rect 425604 679018 425786 679254
rect 426022 679018 426204 679254
rect 425604 678934 426204 679018
rect 425604 678698 425786 678934
rect 426022 678698 426204 678934
rect 425604 643254 426204 678698
rect 425604 643018 425786 643254
rect 426022 643018 426204 643254
rect 425604 642934 426204 643018
rect 425604 642698 425786 642934
rect 426022 642698 426204 642934
rect 425604 607254 426204 642698
rect 425604 607018 425786 607254
rect 426022 607018 426204 607254
rect 425604 606934 426204 607018
rect 425604 606698 425786 606934
rect 426022 606698 426204 606934
rect 425604 571254 426204 606698
rect 425604 571018 425786 571254
rect 426022 571018 426204 571254
rect 425604 570934 426204 571018
rect 425604 570698 425786 570934
rect 426022 570698 426204 570934
rect 425604 535254 426204 570698
rect 425604 535018 425786 535254
rect 426022 535018 426204 535254
rect 425604 534934 426204 535018
rect 425604 534698 425786 534934
rect 426022 534698 426204 534934
rect 425604 499254 426204 534698
rect 425604 499018 425786 499254
rect 426022 499018 426204 499254
rect 425604 498934 426204 499018
rect 425604 498698 425786 498934
rect 426022 498698 426204 498934
rect 425604 463254 426204 498698
rect 425604 463018 425786 463254
rect 426022 463018 426204 463254
rect 425604 462934 426204 463018
rect 425604 462698 425786 462934
rect 426022 462698 426204 462934
rect 425604 427254 426204 462698
rect 425604 427018 425786 427254
rect 426022 427018 426204 427254
rect 425604 426934 426204 427018
rect 425604 426698 425786 426934
rect 426022 426698 426204 426934
rect 425604 391254 426204 426698
rect 425604 391018 425786 391254
rect 426022 391018 426204 391254
rect 425604 390934 426204 391018
rect 425604 390698 425786 390934
rect 426022 390698 426204 390934
rect 425604 355254 426204 390698
rect 425604 355018 425786 355254
rect 426022 355018 426204 355254
rect 425604 354934 426204 355018
rect 425604 354698 425786 354934
rect 426022 354698 426204 354934
rect 425604 319254 426204 354698
rect 425604 319018 425786 319254
rect 426022 319018 426204 319254
rect 425604 318934 426204 319018
rect 425604 318698 425786 318934
rect 426022 318698 426204 318934
rect 425604 283254 426204 318698
rect 425604 283018 425786 283254
rect 426022 283018 426204 283254
rect 425604 282934 426204 283018
rect 425604 282698 425786 282934
rect 426022 282698 426204 282934
rect 425604 247254 426204 282698
rect 425604 247018 425786 247254
rect 426022 247018 426204 247254
rect 425604 246934 426204 247018
rect 425604 246698 425786 246934
rect 426022 246698 426204 246934
rect 425604 211254 426204 246698
rect 425604 211018 425786 211254
rect 426022 211018 426204 211254
rect 425604 210934 426204 211018
rect 425604 210698 425786 210934
rect 426022 210698 426204 210934
rect 425604 175254 426204 210698
rect 425604 175018 425786 175254
rect 426022 175018 426204 175254
rect 425604 174934 426204 175018
rect 425604 174698 425786 174934
rect 426022 174698 426204 174934
rect 425604 139254 426204 174698
rect 425604 139018 425786 139254
rect 426022 139018 426204 139254
rect 425604 138934 426204 139018
rect 425604 138698 425786 138934
rect 426022 138698 426204 138934
rect 425604 103254 426204 138698
rect 425604 103018 425786 103254
rect 426022 103018 426204 103254
rect 425604 102934 426204 103018
rect 425604 102698 425786 102934
rect 426022 102698 426204 102934
rect 425604 67254 426204 102698
rect 425604 67018 425786 67254
rect 426022 67018 426204 67254
rect 425604 66934 426204 67018
rect 425604 66698 425786 66934
rect 426022 66698 426204 66934
rect 425604 31254 426204 66698
rect 425604 31018 425786 31254
rect 426022 31018 426204 31254
rect 425604 30934 426204 31018
rect 425604 30698 425786 30934
rect 426022 30698 426204 30934
rect 407604 -6102 407786 -5866
rect 408022 -6102 408204 -5866
rect 407604 -6186 408204 -6102
rect 407604 -6422 407786 -6186
rect 408022 -6422 408204 -6186
rect 407604 -7364 408204 -6422
rect 425604 -6786 426204 30698
rect 432804 704838 433404 705780
rect 432804 704602 432986 704838
rect 433222 704602 433404 704838
rect 432804 704518 433404 704602
rect 432804 704282 432986 704518
rect 433222 704282 433404 704518
rect 432804 686454 433404 704282
rect 432804 686218 432986 686454
rect 433222 686218 433404 686454
rect 432804 686134 433404 686218
rect 432804 685898 432986 686134
rect 433222 685898 433404 686134
rect 432804 650454 433404 685898
rect 432804 650218 432986 650454
rect 433222 650218 433404 650454
rect 432804 650134 433404 650218
rect 432804 649898 432986 650134
rect 433222 649898 433404 650134
rect 432804 614454 433404 649898
rect 432804 614218 432986 614454
rect 433222 614218 433404 614454
rect 432804 614134 433404 614218
rect 432804 613898 432986 614134
rect 433222 613898 433404 614134
rect 432804 578454 433404 613898
rect 432804 578218 432986 578454
rect 433222 578218 433404 578454
rect 432804 578134 433404 578218
rect 432804 577898 432986 578134
rect 433222 577898 433404 578134
rect 432804 542454 433404 577898
rect 432804 542218 432986 542454
rect 433222 542218 433404 542454
rect 432804 542134 433404 542218
rect 432804 541898 432986 542134
rect 433222 541898 433404 542134
rect 432804 506454 433404 541898
rect 432804 506218 432986 506454
rect 433222 506218 433404 506454
rect 432804 506134 433404 506218
rect 432804 505898 432986 506134
rect 433222 505898 433404 506134
rect 432804 470454 433404 505898
rect 432804 470218 432986 470454
rect 433222 470218 433404 470454
rect 432804 470134 433404 470218
rect 432804 469898 432986 470134
rect 433222 469898 433404 470134
rect 432804 434454 433404 469898
rect 432804 434218 432986 434454
rect 433222 434218 433404 434454
rect 432804 434134 433404 434218
rect 432804 433898 432986 434134
rect 433222 433898 433404 434134
rect 432804 398454 433404 433898
rect 432804 398218 432986 398454
rect 433222 398218 433404 398454
rect 432804 398134 433404 398218
rect 432804 397898 432986 398134
rect 433222 397898 433404 398134
rect 432804 362454 433404 397898
rect 432804 362218 432986 362454
rect 433222 362218 433404 362454
rect 432804 362134 433404 362218
rect 432804 361898 432986 362134
rect 433222 361898 433404 362134
rect 432804 326454 433404 361898
rect 432804 326218 432986 326454
rect 433222 326218 433404 326454
rect 432804 326134 433404 326218
rect 432804 325898 432986 326134
rect 433222 325898 433404 326134
rect 432804 290454 433404 325898
rect 432804 290218 432986 290454
rect 433222 290218 433404 290454
rect 432804 290134 433404 290218
rect 432804 289898 432986 290134
rect 433222 289898 433404 290134
rect 432804 254454 433404 289898
rect 432804 254218 432986 254454
rect 433222 254218 433404 254454
rect 432804 254134 433404 254218
rect 432804 253898 432986 254134
rect 433222 253898 433404 254134
rect 432804 218454 433404 253898
rect 432804 218218 432986 218454
rect 433222 218218 433404 218454
rect 432804 218134 433404 218218
rect 432804 217898 432986 218134
rect 433222 217898 433404 218134
rect 432804 182454 433404 217898
rect 432804 182218 432986 182454
rect 433222 182218 433404 182454
rect 432804 182134 433404 182218
rect 432804 181898 432986 182134
rect 433222 181898 433404 182134
rect 432804 146454 433404 181898
rect 432804 146218 432986 146454
rect 433222 146218 433404 146454
rect 432804 146134 433404 146218
rect 432804 145898 432986 146134
rect 433222 145898 433404 146134
rect 432804 110454 433404 145898
rect 432804 110218 432986 110454
rect 433222 110218 433404 110454
rect 432804 110134 433404 110218
rect 432804 109898 432986 110134
rect 433222 109898 433404 110134
rect 432804 74454 433404 109898
rect 432804 74218 432986 74454
rect 433222 74218 433404 74454
rect 432804 74134 433404 74218
rect 432804 73898 432986 74134
rect 433222 73898 433404 74134
rect 432804 38454 433404 73898
rect 432804 38218 432986 38454
rect 433222 38218 433404 38454
rect 432804 38134 433404 38218
rect 432804 37898 432986 38134
rect 433222 37898 433404 38134
rect 432804 2454 433404 37898
rect 432804 2218 432986 2454
rect 433222 2218 433404 2454
rect 432804 2134 433404 2218
rect 432804 1898 432986 2134
rect 433222 1898 433404 2134
rect 432804 -346 433404 1898
rect 432804 -582 432986 -346
rect 433222 -582 433404 -346
rect 432804 -666 433404 -582
rect 432804 -902 432986 -666
rect 433222 -902 433404 -666
rect 432804 -1844 433404 -902
rect 436404 690054 437004 706122
rect 436404 689818 436586 690054
rect 436822 689818 437004 690054
rect 436404 689734 437004 689818
rect 436404 689498 436586 689734
rect 436822 689498 437004 689734
rect 436404 654054 437004 689498
rect 436404 653818 436586 654054
rect 436822 653818 437004 654054
rect 436404 653734 437004 653818
rect 436404 653498 436586 653734
rect 436822 653498 437004 653734
rect 436404 618054 437004 653498
rect 436404 617818 436586 618054
rect 436822 617818 437004 618054
rect 436404 617734 437004 617818
rect 436404 617498 436586 617734
rect 436822 617498 437004 617734
rect 436404 582054 437004 617498
rect 436404 581818 436586 582054
rect 436822 581818 437004 582054
rect 436404 581734 437004 581818
rect 436404 581498 436586 581734
rect 436822 581498 437004 581734
rect 436404 546054 437004 581498
rect 436404 545818 436586 546054
rect 436822 545818 437004 546054
rect 436404 545734 437004 545818
rect 436404 545498 436586 545734
rect 436822 545498 437004 545734
rect 436404 510054 437004 545498
rect 436404 509818 436586 510054
rect 436822 509818 437004 510054
rect 436404 509734 437004 509818
rect 436404 509498 436586 509734
rect 436822 509498 437004 509734
rect 436404 474054 437004 509498
rect 436404 473818 436586 474054
rect 436822 473818 437004 474054
rect 436404 473734 437004 473818
rect 436404 473498 436586 473734
rect 436822 473498 437004 473734
rect 436404 438054 437004 473498
rect 436404 437818 436586 438054
rect 436822 437818 437004 438054
rect 436404 437734 437004 437818
rect 436404 437498 436586 437734
rect 436822 437498 437004 437734
rect 436404 402054 437004 437498
rect 436404 401818 436586 402054
rect 436822 401818 437004 402054
rect 436404 401734 437004 401818
rect 436404 401498 436586 401734
rect 436822 401498 437004 401734
rect 436404 366054 437004 401498
rect 436404 365818 436586 366054
rect 436822 365818 437004 366054
rect 436404 365734 437004 365818
rect 436404 365498 436586 365734
rect 436822 365498 437004 365734
rect 436404 330054 437004 365498
rect 436404 329818 436586 330054
rect 436822 329818 437004 330054
rect 436404 329734 437004 329818
rect 436404 329498 436586 329734
rect 436822 329498 437004 329734
rect 436404 294054 437004 329498
rect 436404 293818 436586 294054
rect 436822 293818 437004 294054
rect 436404 293734 437004 293818
rect 436404 293498 436586 293734
rect 436822 293498 437004 293734
rect 436404 258054 437004 293498
rect 436404 257818 436586 258054
rect 436822 257818 437004 258054
rect 436404 257734 437004 257818
rect 436404 257498 436586 257734
rect 436822 257498 437004 257734
rect 436404 222054 437004 257498
rect 436404 221818 436586 222054
rect 436822 221818 437004 222054
rect 436404 221734 437004 221818
rect 436404 221498 436586 221734
rect 436822 221498 437004 221734
rect 436404 186054 437004 221498
rect 436404 185818 436586 186054
rect 436822 185818 437004 186054
rect 436404 185734 437004 185818
rect 436404 185498 436586 185734
rect 436822 185498 437004 185734
rect 436404 150054 437004 185498
rect 436404 149818 436586 150054
rect 436822 149818 437004 150054
rect 436404 149734 437004 149818
rect 436404 149498 436586 149734
rect 436822 149498 437004 149734
rect 436404 114054 437004 149498
rect 436404 113818 436586 114054
rect 436822 113818 437004 114054
rect 436404 113734 437004 113818
rect 436404 113498 436586 113734
rect 436822 113498 437004 113734
rect 436404 78054 437004 113498
rect 436404 77818 436586 78054
rect 436822 77818 437004 78054
rect 436404 77734 437004 77818
rect 436404 77498 436586 77734
rect 436822 77498 437004 77734
rect 436404 42054 437004 77498
rect 436404 41818 436586 42054
rect 436822 41818 437004 42054
rect 436404 41734 437004 41818
rect 436404 41498 436586 41734
rect 436822 41498 437004 41734
rect 436404 6054 437004 41498
rect 436404 5818 436586 6054
rect 436822 5818 437004 6054
rect 436404 5734 437004 5818
rect 436404 5498 436586 5734
rect 436822 5498 437004 5734
rect 436404 -2186 437004 5498
rect 436404 -2422 436586 -2186
rect 436822 -2422 437004 -2186
rect 436404 -2506 437004 -2422
rect 436404 -2742 436586 -2506
rect 436822 -2742 437004 -2506
rect 436404 -3684 437004 -2742
rect 440004 693654 440604 707962
rect 440004 693418 440186 693654
rect 440422 693418 440604 693654
rect 440004 693334 440604 693418
rect 440004 693098 440186 693334
rect 440422 693098 440604 693334
rect 440004 657654 440604 693098
rect 440004 657418 440186 657654
rect 440422 657418 440604 657654
rect 440004 657334 440604 657418
rect 440004 657098 440186 657334
rect 440422 657098 440604 657334
rect 440004 621654 440604 657098
rect 440004 621418 440186 621654
rect 440422 621418 440604 621654
rect 440004 621334 440604 621418
rect 440004 621098 440186 621334
rect 440422 621098 440604 621334
rect 440004 585654 440604 621098
rect 440004 585418 440186 585654
rect 440422 585418 440604 585654
rect 440004 585334 440604 585418
rect 440004 585098 440186 585334
rect 440422 585098 440604 585334
rect 440004 549654 440604 585098
rect 440004 549418 440186 549654
rect 440422 549418 440604 549654
rect 440004 549334 440604 549418
rect 440004 549098 440186 549334
rect 440422 549098 440604 549334
rect 440004 513654 440604 549098
rect 440004 513418 440186 513654
rect 440422 513418 440604 513654
rect 440004 513334 440604 513418
rect 440004 513098 440186 513334
rect 440422 513098 440604 513334
rect 440004 477654 440604 513098
rect 440004 477418 440186 477654
rect 440422 477418 440604 477654
rect 440004 477334 440604 477418
rect 440004 477098 440186 477334
rect 440422 477098 440604 477334
rect 440004 441654 440604 477098
rect 440004 441418 440186 441654
rect 440422 441418 440604 441654
rect 440004 441334 440604 441418
rect 440004 441098 440186 441334
rect 440422 441098 440604 441334
rect 440004 405654 440604 441098
rect 440004 405418 440186 405654
rect 440422 405418 440604 405654
rect 440004 405334 440604 405418
rect 440004 405098 440186 405334
rect 440422 405098 440604 405334
rect 440004 369654 440604 405098
rect 440004 369418 440186 369654
rect 440422 369418 440604 369654
rect 440004 369334 440604 369418
rect 440004 369098 440186 369334
rect 440422 369098 440604 369334
rect 440004 333654 440604 369098
rect 440004 333418 440186 333654
rect 440422 333418 440604 333654
rect 440004 333334 440604 333418
rect 440004 333098 440186 333334
rect 440422 333098 440604 333334
rect 440004 297654 440604 333098
rect 440004 297418 440186 297654
rect 440422 297418 440604 297654
rect 440004 297334 440604 297418
rect 440004 297098 440186 297334
rect 440422 297098 440604 297334
rect 440004 261654 440604 297098
rect 440004 261418 440186 261654
rect 440422 261418 440604 261654
rect 440004 261334 440604 261418
rect 440004 261098 440186 261334
rect 440422 261098 440604 261334
rect 440004 225654 440604 261098
rect 440004 225418 440186 225654
rect 440422 225418 440604 225654
rect 440004 225334 440604 225418
rect 440004 225098 440186 225334
rect 440422 225098 440604 225334
rect 440004 189654 440604 225098
rect 440004 189418 440186 189654
rect 440422 189418 440604 189654
rect 440004 189334 440604 189418
rect 440004 189098 440186 189334
rect 440422 189098 440604 189334
rect 440004 153654 440604 189098
rect 440004 153418 440186 153654
rect 440422 153418 440604 153654
rect 440004 153334 440604 153418
rect 440004 153098 440186 153334
rect 440422 153098 440604 153334
rect 440004 117654 440604 153098
rect 440004 117418 440186 117654
rect 440422 117418 440604 117654
rect 440004 117334 440604 117418
rect 440004 117098 440186 117334
rect 440422 117098 440604 117334
rect 440004 81654 440604 117098
rect 440004 81418 440186 81654
rect 440422 81418 440604 81654
rect 440004 81334 440604 81418
rect 440004 81098 440186 81334
rect 440422 81098 440604 81334
rect 440004 45654 440604 81098
rect 440004 45418 440186 45654
rect 440422 45418 440604 45654
rect 440004 45334 440604 45418
rect 440004 45098 440186 45334
rect 440422 45098 440604 45334
rect 440004 9654 440604 45098
rect 440004 9418 440186 9654
rect 440422 9418 440604 9654
rect 440004 9334 440604 9418
rect 440004 9098 440186 9334
rect 440422 9098 440604 9334
rect 440004 -4026 440604 9098
rect 440004 -4262 440186 -4026
rect 440422 -4262 440604 -4026
rect 440004 -4346 440604 -4262
rect 440004 -4582 440186 -4346
rect 440422 -4582 440604 -4346
rect 440004 -5524 440604 -4582
rect 443604 697254 444204 709802
rect 461604 711278 462204 711300
rect 461604 711042 461786 711278
rect 462022 711042 462204 711278
rect 461604 710958 462204 711042
rect 461604 710722 461786 710958
rect 462022 710722 462204 710958
rect 458004 709438 458604 709460
rect 458004 709202 458186 709438
rect 458422 709202 458604 709438
rect 458004 709118 458604 709202
rect 458004 708882 458186 709118
rect 458422 708882 458604 709118
rect 454404 707598 455004 707620
rect 454404 707362 454586 707598
rect 454822 707362 455004 707598
rect 454404 707278 455004 707362
rect 454404 707042 454586 707278
rect 454822 707042 455004 707278
rect 443604 697018 443786 697254
rect 444022 697018 444204 697254
rect 443604 696934 444204 697018
rect 443604 696698 443786 696934
rect 444022 696698 444204 696934
rect 443604 661254 444204 696698
rect 443604 661018 443786 661254
rect 444022 661018 444204 661254
rect 443604 660934 444204 661018
rect 443604 660698 443786 660934
rect 444022 660698 444204 660934
rect 443604 625254 444204 660698
rect 443604 625018 443786 625254
rect 444022 625018 444204 625254
rect 443604 624934 444204 625018
rect 443604 624698 443786 624934
rect 444022 624698 444204 624934
rect 443604 589254 444204 624698
rect 443604 589018 443786 589254
rect 444022 589018 444204 589254
rect 443604 588934 444204 589018
rect 443604 588698 443786 588934
rect 444022 588698 444204 588934
rect 443604 553254 444204 588698
rect 443604 553018 443786 553254
rect 444022 553018 444204 553254
rect 443604 552934 444204 553018
rect 443604 552698 443786 552934
rect 444022 552698 444204 552934
rect 443604 517254 444204 552698
rect 443604 517018 443786 517254
rect 444022 517018 444204 517254
rect 443604 516934 444204 517018
rect 443604 516698 443786 516934
rect 444022 516698 444204 516934
rect 443604 481254 444204 516698
rect 443604 481018 443786 481254
rect 444022 481018 444204 481254
rect 443604 480934 444204 481018
rect 443604 480698 443786 480934
rect 444022 480698 444204 480934
rect 443604 445254 444204 480698
rect 443604 445018 443786 445254
rect 444022 445018 444204 445254
rect 443604 444934 444204 445018
rect 443604 444698 443786 444934
rect 444022 444698 444204 444934
rect 443604 409254 444204 444698
rect 443604 409018 443786 409254
rect 444022 409018 444204 409254
rect 443604 408934 444204 409018
rect 443604 408698 443786 408934
rect 444022 408698 444204 408934
rect 443604 373254 444204 408698
rect 443604 373018 443786 373254
rect 444022 373018 444204 373254
rect 443604 372934 444204 373018
rect 443604 372698 443786 372934
rect 444022 372698 444204 372934
rect 443604 337254 444204 372698
rect 443604 337018 443786 337254
rect 444022 337018 444204 337254
rect 443604 336934 444204 337018
rect 443604 336698 443786 336934
rect 444022 336698 444204 336934
rect 443604 301254 444204 336698
rect 443604 301018 443786 301254
rect 444022 301018 444204 301254
rect 443604 300934 444204 301018
rect 443604 300698 443786 300934
rect 444022 300698 444204 300934
rect 443604 265254 444204 300698
rect 443604 265018 443786 265254
rect 444022 265018 444204 265254
rect 443604 264934 444204 265018
rect 443604 264698 443786 264934
rect 444022 264698 444204 264934
rect 443604 229254 444204 264698
rect 443604 229018 443786 229254
rect 444022 229018 444204 229254
rect 443604 228934 444204 229018
rect 443604 228698 443786 228934
rect 444022 228698 444204 228934
rect 443604 193254 444204 228698
rect 443604 193018 443786 193254
rect 444022 193018 444204 193254
rect 443604 192934 444204 193018
rect 443604 192698 443786 192934
rect 444022 192698 444204 192934
rect 443604 157254 444204 192698
rect 443604 157018 443786 157254
rect 444022 157018 444204 157254
rect 443604 156934 444204 157018
rect 443604 156698 443786 156934
rect 444022 156698 444204 156934
rect 443604 121254 444204 156698
rect 443604 121018 443786 121254
rect 444022 121018 444204 121254
rect 443604 120934 444204 121018
rect 443604 120698 443786 120934
rect 444022 120698 444204 120934
rect 443604 85254 444204 120698
rect 443604 85018 443786 85254
rect 444022 85018 444204 85254
rect 443604 84934 444204 85018
rect 443604 84698 443786 84934
rect 444022 84698 444204 84934
rect 443604 49254 444204 84698
rect 443604 49018 443786 49254
rect 444022 49018 444204 49254
rect 443604 48934 444204 49018
rect 443604 48698 443786 48934
rect 444022 48698 444204 48934
rect 443604 13254 444204 48698
rect 443604 13018 443786 13254
rect 444022 13018 444204 13254
rect 443604 12934 444204 13018
rect 443604 12698 443786 12934
rect 444022 12698 444204 12934
rect 425604 -7022 425786 -6786
rect 426022 -7022 426204 -6786
rect 425604 -7106 426204 -7022
rect 425604 -7342 425786 -7106
rect 426022 -7342 426204 -7106
rect 425604 -7364 426204 -7342
rect 443604 -5866 444204 12698
rect 450804 705758 451404 705780
rect 450804 705522 450986 705758
rect 451222 705522 451404 705758
rect 450804 705438 451404 705522
rect 450804 705202 450986 705438
rect 451222 705202 451404 705438
rect 450804 668454 451404 705202
rect 450804 668218 450986 668454
rect 451222 668218 451404 668454
rect 450804 668134 451404 668218
rect 450804 667898 450986 668134
rect 451222 667898 451404 668134
rect 450804 632454 451404 667898
rect 450804 632218 450986 632454
rect 451222 632218 451404 632454
rect 450804 632134 451404 632218
rect 450804 631898 450986 632134
rect 451222 631898 451404 632134
rect 450804 596454 451404 631898
rect 450804 596218 450986 596454
rect 451222 596218 451404 596454
rect 450804 596134 451404 596218
rect 450804 595898 450986 596134
rect 451222 595898 451404 596134
rect 450804 560454 451404 595898
rect 450804 560218 450986 560454
rect 451222 560218 451404 560454
rect 450804 560134 451404 560218
rect 450804 559898 450986 560134
rect 451222 559898 451404 560134
rect 450804 524454 451404 559898
rect 450804 524218 450986 524454
rect 451222 524218 451404 524454
rect 450804 524134 451404 524218
rect 450804 523898 450986 524134
rect 451222 523898 451404 524134
rect 450804 488454 451404 523898
rect 450804 488218 450986 488454
rect 451222 488218 451404 488454
rect 450804 488134 451404 488218
rect 450804 487898 450986 488134
rect 451222 487898 451404 488134
rect 450804 452454 451404 487898
rect 450804 452218 450986 452454
rect 451222 452218 451404 452454
rect 450804 452134 451404 452218
rect 450804 451898 450986 452134
rect 451222 451898 451404 452134
rect 450804 416454 451404 451898
rect 450804 416218 450986 416454
rect 451222 416218 451404 416454
rect 450804 416134 451404 416218
rect 450804 415898 450986 416134
rect 451222 415898 451404 416134
rect 450804 380454 451404 415898
rect 450804 380218 450986 380454
rect 451222 380218 451404 380454
rect 450804 380134 451404 380218
rect 450804 379898 450986 380134
rect 451222 379898 451404 380134
rect 450804 344454 451404 379898
rect 450804 344218 450986 344454
rect 451222 344218 451404 344454
rect 450804 344134 451404 344218
rect 450804 343898 450986 344134
rect 451222 343898 451404 344134
rect 450804 308454 451404 343898
rect 450804 308218 450986 308454
rect 451222 308218 451404 308454
rect 450804 308134 451404 308218
rect 450804 307898 450986 308134
rect 451222 307898 451404 308134
rect 450804 272454 451404 307898
rect 450804 272218 450986 272454
rect 451222 272218 451404 272454
rect 450804 272134 451404 272218
rect 450804 271898 450986 272134
rect 451222 271898 451404 272134
rect 450804 236454 451404 271898
rect 450804 236218 450986 236454
rect 451222 236218 451404 236454
rect 450804 236134 451404 236218
rect 450804 235898 450986 236134
rect 451222 235898 451404 236134
rect 450804 200454 451404 235898
rect 450804 200218 450986 200454
rect 451222 200218 451404 200454
rect 450804 200134 451404 200218
rect 450804 199898 450986 200134
rect 451222 199898 451404 200134
rect 450804 164454 451404 199898
rect 450804 164218 450986 164454
rect 451222 164218 451404 164454
rect 450804 164134 451404 164218
rect 450804 163898 450986 164134
rect 451222 163898 451404 164134
rect 450804 128454 451404 163898
rect 450804 128218 450986 128454
rect 451222 128218 451404 128454
rect 450804 128134 451404 128218
rect 450804 127898 450986 128134
rect 451222 127898 451404 128134
rect 450804 92454 451404 127898
rect 450804 92218 450986 92454
rect 451222 92218 451404 92454
rect 450804 92134 451404 92218
rect 450804 91898 450986 92134
rect 451222 91898 451404 92134
rect 450804 56454 451404 91898
rect 450804 56218 450986 56454
rect 451222 56218 451404 56454
rect 450804 56134 451404 56218
rect 450804 55898 450986 56134
rect 451222 55898 451404 56134
rect 450804 20454 451404 55898
rect 450804 20218 450986 20454
rect 451222 20218 451404 20454
rect 450804 20134 451404 20218
rect 450804 19898 450986 20134
rect 451222 19898 451404 20134
rect 450804 -1266 451404 19898
rect 450804 -1502 450986 -1266
rect 451222 -1502 451404 -1266
rect 450804 -1586 451404 -1502
rect 450804 -1822 450986 -1586
rect 451222 -1822 451404 -1586
rect 450804 -1844 451404 -1822
rect 454404 672054 455004 707042
rect 454404 671818 454586 672054
rect 454822 671818 455004 672054
rect 454404 671734 455004 671818
rect 454404 671498 454586 671734
rect 454822 671498 455004 671734
rect 454404 636054 455004 671498
rect 454404 635818 454586 636054
rect 454822 635818 455004 636054
rect 454404 635734 455004 635818
rect 454404 635498 454586 635734
rect 454822 635498 455004 635734
rect 454404 600054 455004 635498
rect 454404 599818 454586 600054
rect 454822 599818 455004 600054
rect 454404 599734 455004 599818
rect 454404 599498 454586 599734
rect 454822 599498 455004 599734
rect 454404 564054 455004 599498
rect 454404 563818 454586 564054
rect 454822 563818 455004 564054
rect 454404 563734 455004 563818
rect 454404 563498 454586 563734
rect 454822 563498 455004 563734
rect 454404 528054 455004 563498
rect 454404 527818 454586 528054
rect 454822 527818 455004 528054
rect 454404 527734 455004 527818
rect 454404 527498 454586 527734
rect 454822 527498 455004 527734
rect 454404 492054 455004 527498
rect 454404 491818 454586 492054
rect 454822 491818 455004 492054
rect 454404 491734 455004 491818
rect 454404 491498 454586 491734
rect 454822 491498 455004 491734
rect 454404 456054 455004 491498
rect 454404 455818 454586 456054
rect 454822 455818 455004 456054
rect 454404 455734 455004 455818
rect 454404 455498 454586 455734
rect 454822 455498 455004 455734
rect 454404 420054 455004 455498
rect 454404 419818 454586 420054
rect 454822 419818 455004 420054
rect 454404 419734 455004 419818
rect 454404 419498 454586 419734
rect 454822 419498 455004 419734
rect 454404 384054 455004 419498
rect 454404 383818 454586 384054
rect 454822 383818 455004 384054
rect 454404 383734 455004 383818
rect 454404 383498 454586 383734
rect 454822 383498 455004 383734
rect 454404 348054 455004 383498
rect 454404 347818 454586 348054
rect 454822 347818 455004 348054
rect 454404 347734 455004 347818
rect 454404 347498 454586 347734
rect 454822 347498 455004 347734
rect 454404 312054 455004 347498
rect 454404 311818 454586 312054
rect 454822 311818 455004 312054
rect 454404 311734 455004 311818
rect 454404 311498 454586 311734
rect 454822 311498 455004 311734
rect 454404 276054 455004 311498
rect 454404 275818 454586 276054
rect 454822 275818 455004 276054
rect 454404 275734 455004 275818
rect 454404 275498 454586 275734
rect 454822 275498 455004 275734
rect 454404 240054 455004 275498
rect 454404 239818 454586 240054
rect 454822 239818 455004 240054
rect 454404 239734 455004 239818
rect 454404 239498 454586 239734
rect 454822 239498 455004 239734
rect 454404 204054 455004 239498
rect 454404 203818 454586 204054
rect 454822 203818 455004 204054
rect 454404 203734 455004 203818
rect 454404 203498 454586 203734
rect 454822 203498 455004 203734
rect 454404 168054 455004 203498
rect 454404 167818 454586 168054
rect 454822 167818 455004 168054
rect 454404 167734 455004 167818
rect 454404 167498 454586 167734
rect 454822 167498 455004 167734
rect 454404 132054 455004 167498
rect 454404 131818 454586 132054
rect 454822 131818 455004 132054
rect 454404 131734 455004 131818
rect 454404 131498 454586 131734
rect 454822 131498 455004 131734
rect 454404 96054 455004 131498
rect 454404 95818 454586 96054
rect 454822 95818 455004 96054
rect 454404 95734 455004 95818
rect 454404 95498 454586 95734
rect 454822 95498 455004 95734
rect 454404 60054 455004 95498
rect 454404 59818 454586 60054
rect 454822 59818 455004 60054
rect 454404 59734 455004 59818
rect 454404 59498 454586 59734
rect 454822 59498 455004 59734
rect 454404 24054 455004 59498
rect 454404 23818 454586 24054
rect 454822 23818 455004 24054
rect 454404 23734 455004 23818
rect 454404 23498 454586 23734
rect 454822 23498 455004 23734
rect 454404 -3106 455004 23498
rect 454404 -3342 454586 -3106
rect 454822 -3342 455004 -3106
rect 454404 -3426 455004 -3342
rect 454404 -3662 454586 -3426
rect 454822 -3662 455004 -3426
rect 454404 -3684 455004 -3662
rect 458004 675654 458604 708882
rect 458004 675418 458186 675654
rect 458422 675418 458604 675654
rect 458004 675334 458604 675418
rect 458004 675098 458186 675334
rect 458422 675098 458604 675334
rect 458004 639654 458604 675098
rect 458004 639418 458186 639654
rect 458422 639418 458604 639654
rect 458004 639334 458604 639418
rect 458004 639098 458186 639334
rect 458422 639098 458604 639334
rect 458004 603654 458604 639098
rect 458004 603418 458186 603654
rect 458422 603418 458604 603654
rect 458004 603334 458604 603418
rect 458004 603098 458186 603334
rect 458422 603098 458604 603334
rect 458004 567654 458604 603098
rect 458004 567418 458186 567654
rect 458422 567418 458604 567654
rect 458004 567334 458604 567418
rect 458004 567098 458186 567334
rect 458422 567098 458604 567334
rect 458004 531654 458604 567098
rect 458004 531418 458186 531654
rect 458422 531418 458604 531654
rect 458004 531334 458604 531418
rect 458004 531098 458186 531334
rect 458422 531098 458604 531334
rect 458004 495654 458604 531098
rect 458004 495418 458186 495654
rect 458422 495418 458604 495654
rect 458004 495334 458604 495418
rect 458004 495098 458186 495334
rect 458422 495098 458604 495334
rect 458004 459654 458604 495098
rect 458004 459418 458186 459654
rect 458422 459418 458604 459654
rect 458004 459334 458604 459418
rect 458004 459098 458186 459334
rect 458422 459098 458604 459334
rect 458004 423654 458604 459098
rect 458004 423418 458186 423654
rect 458422 423418 458604 423654
rect 458004 423334 458604 423418
rect 458004 423098 458186 423334
rect 458422 423098 458604 423334
rect 458004 387654 458604 423098
rect 458004 387418 458186 387654
rect 458422 387418 458604 387654
rect 458004 387334 458604 387418
rect 458004 387098 458186 387334
rect 458422 387098 458604 387334
rect 458004 351654 458604 387098
rect 458004 351418 458186 351654
rect 458422 351418 458604 351654
rect 458004 351334 458604 351418
rect 458004 351098 458186 351334
rect 458422 351098 458604 351334
rect 458004 315654 458604 351098
rect 458004 315418 458186 315654
rect 458422 315418 458604 315654
rect 458004 315334 458604 315418
rect 458004 315098 458186 315334
rect 458422 315098 458604 315334
rect 458004 279654 458604 315098
rect 458004 279418 458186 279654
rect 458422 279418 458604 279654
rect 458004 279334 458604 279418
rect 458004 279098 458186 279334
rect 458422 279098 458604 279334
rect 458004 243654 458604 279098
rect 458004 243418 458186 243654
rect 458422 243418 458604 243654
rect 458004 243334 458604 243418
rect 458004 243098 458186 243334
rect 458422 243098 458604 243334
rect 458004 207654 458604 243098
rect 458004 207418 458186 207654
rect 458422 207418 458604 207654
rect 458004 207334 458604 207418
rect 458004 207098 458186 207334
rect 458422 207098 458604 207334
rect 458004 171654 458604 207098
rect 458004 171418 458186 171654
rect 458422 171418 458604 171654
rect 458004 171334 458604 171418
rect 458004 171098 458186 171334
rect 458422 171098 458604 171334
rect 458004 135654 458604 171098
rect 458004 135418 458186 135654
rect 458422 135418 458604 135654
rect 458004 135334 458604 135418
rect 458004 135098 458186 135334
rect 458422 135098 458604 135334
rect 458004 99654 458604 135098
rect 458004 99418 458186 99654
rect 458422 99418 458604 99654
rect 458004 99334 458604 99418
rect 458004 99098 458186 99334
rect 458422 99098 458604 99334
rect 458004 63654 458604 99098
rect 458004 63418 458186 63654
rect 458422 63418 458604 63654
rect 458004 63334 458604 63418
rect 458004 63098 458186 63334
rect 458422 63098 458604 63334
rect 458004 27654 458604 63098
rect 458004 27418 458186 27654
rect 458422 27418 458604 27654
rect 458004 27334 458604 27418
rect 458004 27098 458186 27334
rect 458422 27098 458604 27334
rect 458004 -4946 458604 27098
rect 458004 -5182 458186 -4946
rect 458422 -5182 458604 -4946
rect 458004 -5266 458604 -5182
rect 458004 -5502 458186 -5266
rect 458422 -5502 458604 -5266
rect 458004 -5524 458604 -5502
rect 461604 679254 462204 710722
rect 479604 710358 480204 711300
rect 479604 710122 479786 710358
rect 480022 710122 480204 710358
rect 479604 710038 480204 710122
rect 479604 709802 479786 710038
rect 480022 709802 480204 710038
rect 476004 708518 476604 709460
rect 476004 708282 476186 708518
rect 476422 708282 476604 708518
rect 476004 708198 476604 708282
rect 476004 707962 476186 708198
rect 476422 707962 476604 708198
rect 472404 706678 473004 707620
rect 472404 706442 472586 706678
rect 472822 706442 473004 706678
rect 472404 706358 473004 706442
rect 472404 706122 472586 706358
rect 472822 706122 473004 706358
rect 461604 679018 461786 679254
rect 462022 679018 462204 679254
rect 461604 678934 462204 679018
rect 461604 678698 461786 678934
rect 462022 678698 462204 678934
rect 461604 643254 462204 678698
rect 461604 643018 461786 643254
rect 462022 643018 462204 643254
rect 461604 642934 462204 643018
rect 461604 642698 461786 642934
rect 462022 642698 462204 642934
rect 461604 607254 462204 642698
rect 461604 607018 461786 607254
rect 462022 607018 462204 607254
rect 461604 606934 462204 607018
rect 461604 606698 461786 606934
rect 462022 606698 462204 606934
rect 461604 571254 462204 606698
rect 461604 571018 461786 571254
rect 462022 571018 462204 571254
rect 461604 570934 462204 571018
rect 461604 570698 461786 570934
rect 462022 570698 462204 570934
rect 461604 535254 462204 570698
rect 461604 535018 461786 535254
rect 462022 535018 462204 535254
rect 461604 534934 462204 535018
rect 461604 534698 461786 534934
rect 462022 534698 462204 534934
rect 461604 499254 462204 534698
rect 461604 499018 461786 499254
rect 462022 499018 462204 499254
rect 461604 498934 462204 499018
rect 461604 498698 461786 498934
rect 462022 498698 462204 498934
rect 461604 463254 462204 498698
rect 461604 463018 461786 463254
rect 462022 463018 462204 463254
rect 461604 462934 462204 463018
rect 461604 462698 461786 462934
rect 462022 462698 462204 462934
rect 461604 427254 462204 462698
rect 461604 427018 461786 427254
rect 462022 427018 462204 427254
rect 461604 426934 462204 427018
rect 461604 426698 461786 426934
rect 462022 426698 462204 426934
rect 461604 391254 462204 426698
rect 461604 391018 461786 391254
rect 462022 391018 462204 391254
rect 461604 390934 462204 391018
rect 461604 390698 461786 390934
rect 462022 390698 462204 390934
rect 461604 355254 462204 390698
rect 461604 355018 461786 355254
rect 462022 355018 462204 355254
rect 461604 354934 462204 355018
rect 461604 354698 461786 354934
rect 462022 354698 462204 354934
rect 461604 319254 462204 354698
rect 461604 319018 461786 319254
rect 462022 319018 462204 319254
rect 461604 318934 462204 319018
rect 461604 318698 461786 318934
rect 462022 318698 462204 318934
rect 461604 283254 462204 318698
rect 461604 283018 461786 283254
rect 462022 283018 462204 283254
rect 461604 282934 462204 283018
rect 461604 282698 461786 282934
rect 462022 282698 462204 282934
rect 461604 247254 462204 282698
rect 461604 247018 461786 247254
rect 462022 247018 462204 247254
rect 461604 246934 462204 247018
rect 461604 246698 461786 246934
rect 462022 246698 462204 246934
rect 461604 211254 462204 246698
rect 461604 211018 461786 211254
rect 462022 211018 462204 211254
rect 461604 210934 462204 211018
rect 461604 210698 461786 210934
rect 462022 210698 462204 210934
rect 461604 175254 462204 210698
rect 461604 175018 461786 175254
rect 462022 175018 462204 175254
rect 461604 174934 462204 175018
rect 461604 174698 461786 174934
rect 462022 174698 462204 174934
rect 461604 139254 462204 174698
rect 461604 139018 461786 139254
rect 462022 139018 462204 139254
rect 461604 138934 462204 139018
rect 461604 138698 461786 138934
rect 462022 138698 462204 138934
rect 461604 103254 462204 138698
rect 461604 103018 461786 103254
rect 462022 103018 462204 103254
rect 461604 102934 462204 103018
rect 461604 102698 461786 102934
rect 462022 102698 462204 102934
rect 461604 67254 462204 102698
rect 461604 67018 461786 67254
rect 462022 67018 462204 67254
rect 461604 66934 462204 67018
rect 461604 66698 461786 66934
rect 462022 66698 462204 66934
rect 461604 31254 462204 66698
rect 461604 31018 461786 31254
rect 462022 31018 462204 31254
rect 461604 30934 462204 31018
rect 461604 30698 461786 30934
rect 462022 30698 462204 30934
rect 443604 -6102 443786 -5866
rect 444022 -6102 444204 -5866
rect 443604 -6186 444204 -6102
rect 443604 -6422 443786 -6186
rect 444022 -6422 444204 -6186
rect 443604 -7364 444204 -6422
rect 461604 -6786 462204 30698
rect 468804 704838 469404 705780
rect 468804 704602 468986 704838
rect 469222 704602 469404 704838
rect 468804 704518 469404 704602
rect 468804 704282 468986 704518
rect 469222 704282 469404 704518
rect 468804 686454 469404 704282
rect 468804 686218 468986 686454
rect 469222 686218 469404 686454
rect 468804 686134 469404 686218
rect 468804 685898 468986 686134
rect 469222 685898 469404 686134
rect 468804 650454 469404 685898
rect 468804 650218 468986 650454
rect 469222 650218 469404 650454
rect 468804 650134 469404 650218
rect 468804 649898 468986 650134
rect 469222 649898 469404 650134
rect 468804 614454 469404 649898
rect 468804 614218 468986 614454
rect 469222 614218 469404 614454
rect 468804 614134 469404 614218
rect 468804 613898 468986 614134
rect 469222 613898 469404 614134
rect 468804 578454 469404 613898
rect 468804 578218 468986 578454
rect 469222 578218 469404 578454
rect 468804 578134 469404 578218
rect 468804 577898 468986 578134
rect 469222 577898 469404 578134
rect 468804 542454 469404 577898
rect 468804 542218 468986 542454
rect 469222 542218 469404 542454
rect 468804 542134 469404 542218
rect 468804 541898 468986 542134
rect 469222 541898 469404 542134
rect 468804 506454 469404 541898
rect 468804 506218 468986 506454
rect 469222 506218 469404 506454
rect 468804 506134 469404 506218
rect 468804 505898 468986 506134
rect 469222 505898 469404 506134
rect 468804 470454 469404 505898
rect 468804 470218 468986 470454
rect 469222 470218 469404 470454
rect 468804 470134 469404 470218
rect 468804 469898 468986 470134
rect 469222 469898 469404 470134
rect 468804 434454 469404 469898
rect 468804 434218 468986 434454
rect 469222 434218 469404 434454
rect 468804 434134 469404 434218
rect 468804 433898 468986 434134
rect 469222 433898 469404 434134
rect 468804 398454 469404 433898
rect 468804 398218 468986 398454
rect 469222 398218 469404 398454
rect 468804 398134 469404 398218
rect 468804 397898 468986 398134
rect 469222 397898 469404 398134
rect 468804 362454 469404 397898
rect 468804 362218 468986 362454
rect 469222 362218 469404 362454
rect 468804 362134 469404 362218
rect 468804 361898 468986 362134
rect 469222 361898 469404 362134
rect 468804 326454 469404 361898
rect 468804 326218 468986 326454
rect 469222 326218 469404 326454
rect 468804 326134 469404 326218
rect 468804 325898 468986 326134
rect 469222 325898 469404 326134
rect 468804 290454 469404 325898
rect 468804 290218 468986 290454
rect 469222 290218 469404 290454
rect 468804 290134 469404 290218
rect 468804 289898 468986 290134
rect 469222 289898 469404 290134
rect 468804 254454 469404 289898
rect 468804 254218 468986 254454
rect 469222 254218 469404 254454
rect 468804 254134 469404 254218
rect 468804 253898 468986 254134
rect 469222 253898 469404 254134
rect 468804 218454 469404 253898
rect 468804 218218 468986 218454
rect 469222 218218 469404 218454
rect 468804 218134 469404 218218
rect 468804 217898 468986 218134
rect 469222 217898 469404 218134
rect 468804 182454 469404 217898
rect 468804 182218 468986 182454
rect 469222 182218 469404 182454
rect 468804 182134 469404 182218
rect 468804 181898 468986 182134
rect 469222 181898 469404 182134
rect 468804 146454 469404 181898
rect 468804 146218 468986 146454
rect 469222 146218 469404 146454
rect 468804 146134 469404 146218
rect 468804 145898 468986 146134
rect 469222 145898 469404 146134
rect 468804 110454 469404 145898
rect 468804 110218 468986 110454
rect 469222 110218 469404 110454
rect 468804 110134 469404 110218
rect 468804 109898 468986 110134
rect 469222 109898 469404 110134
rect 468804 74454 469404 109898
rect 468804 74218 468986 74454
rect 469222 74218 469404 74454
rect 468804 74134 469404 74218
rect 468804 73898 468986 74134
rect 469222 73898 469404 74134
rect 468804 38454 469404 73898
rect 468804 38218 468986 38454
rect 469222 38218 469404 38454
rect 468804 38134 469404 38218
rect 468804 37898 468986 38134
rect 469222 37898 469404 38134
rect 468804 2454 469404 37898
rect 468804 2218 468986 2454
rect 469222 2218 469404 2454
rect 468804 2134 469404 2218
rect 468804 1898 468986 2134
rect 469222 1898 469404 2134
rect 468804 -346 469404 1898
rect 468804 -582 468986 -346
rect 469222 -582 469404 -346
rect 468804 -666 469404 -582
rect 468804 -902 468986 -666
rect 469222 -902 469404 -666
rect 468804 -1844 469404 -902
rect 472404 690054 473004 706122
rect 472404 689818 472586 690054
rect 472822 689818 473004 690054
rect 472404 689734 473004 689818
rect 472404 689498 472586 689734
rect 472822 689498 473004 689734
rect 472404 654054 473004 689498
rect 472404 653818 472586 654054
rect 472822 653818 473004 654054
rect 472404 653734 473004 653818
rect 472404 653498 472586 653734
rect 472822 653498 473004 653734
rect 472404 618054 473004 653498
rect 472404 617818 472586 618054
rect 472822 617818 473004 618054
rect 472404 617734 473004 617818
rect 472404 617498 472586 617734
rect 472822 617498 473004 617734
rect 472404 582054 473004 617498
rect 472404 581818 472586 582054
rect 472822 581818 473004 582054
rect 472404 581734 473004 581818
rect 472404 581498 472586 581734
rect 472822 581498 473004 581734
rect 472404 546054 473004 581498
rect 472404 545818 472586 546054
rect 472822 545818 473004 546054
rect 472404 545734 473004 545818
rect 472404 545498 472586 545734
rect 472822 545498 473004 545734
rect 472404 510054 473004 545498
rect 472404 509818 472586 510054
rect 472822 509818 473004 510054
rect 472404 509734 473004 509818
rect 472404 509498 472586 509734
rect 472822 509498 473004 509734
rect 472404 474054 473004 509498
rect 472404 473818 472586 474054
rect 472822 473818 473004 474054
rect 472404 473734 473004 473818
rect 472404 473498 472586 473734
rect 472822 473498 473004 473734
rect 472404 438054 473004 473498
rect 472404 437818 472586 438054
rect 472822 437818 473004 438054
rect 472404 437734 473004 437818
rect 472404 437498 472586 437734
rect 472822 437498 473004 437734
rect 472404 402054 473004 437498
rect 472404 401818 472586 402054
rect 472822 401818 473004 402054
rect 472404 401734 473004 401818
rect 472404 401498 472586 401734
rect 472822 401498 473004 401734
rect 472404 366054 473004 401498
rect 472404 365818 472586 366054
rect 472822 365818 473004 366054
rect 472404 365734 473004 365818
rect 472404 365498 472586 365734
rect 472822 365498 473004 365734
rect 472404 330054 473004 365498
rect 472404 329818 472586 330054
rect 472822 329818 473004 330054
rect 472404 329734 473004 329818
rect 472404 329498 472586 329734
rect 472822 329498 473004 329734
rect 472404 294054 473004 329498
rect 472404 293818 472586 294054
rect 472822 293818 473004 294054
rect 472404 293734 473004 293818
rect 472404 293498 472586 293734
rect 472822 293498 473004 293734
rect 472404 258054 473004 293498
rect 472404 257818 472586 258054
rect 472822 257818 473004 258054
rect 472404 257734 473004 257818
rect 472404 257498 472586 257734
rect 472822 257498 473004 257734
rect 472404 222054 473004 257498
rect 472404 221818 472586 222054
rect 472822 221818 473004 222054
rect 472404 221734 473004 221818
rect 472404 221498 472586 221734
rect 472822 221498 473004 221734
rect 472404 186054 473004 221498
rect 472404 185818 472586 186054
rect 472822 185818 473004 186054
rect 472404 185734 473004 185818
rect 472404 185498 472586 185734
rect 472822 185498 473004 185734
rect 472404 150054 473004 185498
rect 472404 149818 472586 150054
rect 472822 149818 473004 150054
rect 472404 149734 473004 149818
rect 472404 149498 472586 149734
rect 472822 149498 473004 149734
rect 472404 114054 473004 149498
rect 472404 113818 472586 114054
rect 472822 113818 473004 114054
rect 472404 113734 473004 113818
rect 472404 113498 472586 113734
rect 472822 113498 473004 113734
rect 472404 78054 473004 113498
rect 472404 77818 472586 78054
rect 472822 77818 473004 78054
rect 472404 77734 473004 77818
rect 472404 77498 472586 77734
rect 472822 77498 473004 77734
rect 472404 42054 473004 77498
rect 472404 41818 472586 42054
rect 472822 41818 473004 42054
rect 472404 41734 473004 41818
rect 472404 41498 472586 41734
rect 472822 41498 473004 41734
rect 472404 6054 473004 41498
rect 472404 5818 472586 6054
rect 472822 5818 473004 6054
rect 472404 5734 473004 5818
rect 472404 5498 472586 5734
rect 472822 5498 473004 5734
rect 472404 -2186 473004 5498
rect 472404 -2422 472586 -2186
rect 472822 -2422 473004 -2186
rect 472404 -2506 473004 -2422
rect 472404 -2742 472586 -2506
rect 472822 -2742 473004 -2506
rect 472404 -3684 473004 -2742
rect 476004 693654 476604 707962
rect 476004 693418 476186 693654
rect 476422 693418 476604 693654
rect 476004 693334 476604 693418
rect 476004 693098 476186 693334
rect 476422 693098 476604 693334
rect 476004 657654 476604 693098
rect 476004 657418 476186 657654
rect 476422 657418 476604 657654
rect 476004 657334 476604 657418
rect 476004 657098 476186 657334
rect 476422 657098 476604 657334
rect 476004 621654 476604 657098
rect 476004 621418 476186 621654
rect 476422 621418 476604 621654
rect 476004 621334 476604 621418
rect 476004 621098 476186 621334
rect 476422 621098 476604 621334
rect 476004 585654 476604 621098
rect 476004 585418 476186 585654
rect 476422 585418 476604 585654
rect 476004 585334 476604 585418
rect 476004 585098 476186 585334
rect 476422 585098 476604 585334
rect 476004 549654 476604 585098
rect 476004 549418 476186 549654
rect 476422 549418 476604 549654
rect 476004 549334 476604 549418
rect 476004 549098 476186 549334
rect 476422 549098 476604 549334
rect 476004 513654 476604 549098
rect 476004 513418 476186 513654
rect 476422 513418 476604 513654
rect 476004 513334 476604 513418
rect 476004 513098 476186 513334
rect 476422 513098 476604 513334
rect 476004 477654 476604 513098
rect 476004 477418 476186 477654
rect 476422 477418 476604 477654
rect 476004 477334 476604 477418
rect 476004 477098 476186 477334
rect 476422 477098 476604 477334
rect 476004 441654 476604 477098
rect 476004 441418 476186 441654
rect 476422 441418 476604 441654
rect 476004 441334 476604 441418
rect 476004 441098 476186 441334
rect 476422 441098 476604 441334
rect 476004 405654 476604 441098
rect 476004 405418 476186 405654
rect 476422 405418 476604 405654
rect 476004 405334 476604 405418
rect 476004 405098 476186 405334
rect 476422 405098 476604 405334
rect 476004 369654 476604 405098
rect 476004 369418 476186 369654
rect 476422 369418 476604 369654
rect 476004 369334 476604 369418
rect 476004 369098 476186 369334
rect 476422 369098 476604 369334
rect 476004 333654 476604 369098
rect 476004 333418 476186 333654
rect 476422 333418 476604 333654
rect 476004 333334 476604 333418
rect 476004 333098 476186 333334
rect 476422 333098 476604 333334
rect 476004 297654 476604 333098
rect 476004 297418 476186 297654
rect 476422 297418 476604 297654
rect 476004 297334 476604 297418
rect 476004 297098 476186 297334
rect 476422 297098 476604 297334
rect 476004 261654 476604 297098
rect 476004 261418 476186 261654
rect 476422 261418 476604 261654
rect 476004 261334 476604 261418
rect 476004 261098 476186 261334
rect 476422 261098 476604 261334
rect 476004 225654 476604 261098
rect 476004 225418 476186 225654
rect 476422 225418 476604 225654
rect 476004 225334 476604 225418
rect 476004 225098 476186 225334
rect 476422 225098 476604 225334
rect 476004 189654 476604 225098
rect 476004 189418 476186 189654
rect 476422 189418 476604 189654
rect 476004 189334 476604 189418
rect 476004 189098 476186 189334
rect 476422 189098 476604 189334
rect 476004 153654 476604 189098
rect 476004 153418 476186 153654
rect 476422 153418 476604 153654
rect 476004 153334 476604 153418
rect 476004 153098 476186 153334
rect 476422 153098 476604 153334
rect 476004 117654 476604 153098
rect 476004 117418 476186 117654
rect 476422 117418 476604 117654
rect 476004 117334 476604 117418
rect 476004 117098 476186 117334
rect 476422 117098 476604 117334
rect 476004 81654 476604 117098
rect 476004 81418 476186 81654
rect 476422 81418 476604 81654
rect 476004 81334 476604 81418
rect 476004 81098 476186 81334
rect 476422 81098 476604 81334
rect 476004 45654 476604 81098
rect 476004 45418 476186 45654
rect 476422 45418 476604 45654
rect 476004 45334 476604 45418
rect 476004 45098 476186 45334
rect 476422 45098 476604 45334
rect 476004 9654 476604 45098
rect 476004 9418 476186 9654
rect 476422 9418 476604 9654
rect 476004 9334 476604 9418
rect 476004 9098 476186 9334
rect 476422 9098 476604 9334
rect 476004 -4026 476604 9098
rect 476004 -4262 476186 -4026
rect 476422 -4262 476604 -4026
rect 476004 -4346 476604 -4262
rect 476004 -4582 476186 -4346
rect 476422 -4582 476604 -4346
rect 476004 -5524 476604 -4582
rect 479604 697254 480204 709802
rect 497604 711278 498204 711300
rect 497604 711042 497786 711278
rect 498022 711042 498204 711278
rect 497604 710958 498204 711042
rect 497604 710722 497786 710958
rect 498022 710722 498204 710958
rect 494004 709438 494604 709460
rect 494004 709202 494186 709438
rect 494422 709202 494604 709438
rect 494004 709118 494604 709202
rect 494004 708882 494186 709118
rect 494422 708882 494604 709118
rect 490404 707598 491004 707620
rect 490404 707362 490586 707598
rect 490822 707362 491004 707598
rect 490404 707278 491004 707362
rect 490404 707042 490586 707278
rect 490822 707042 491004 707278
rect 479604 697018 479786 697254
rect 480022 697018 480204 697254
rect 479604 696934 480204 697018
rect 479604 696698 479786 696934
rect 480022 696698 480204 696934
rect 479604 661254 480204 696698
rect 479604 661018 479786 661254
rect 480022 661018 480204 661254
rect 479604 660934 480204 661018
rect 479604 660698 479786 660934
rect 480022 660698 480204 660934
rect 479604 625254 480204 660698
rect 479604 625018 479786 625254
rect 480022 625018 480204 625254
rect 479604 624934 480204 625018
rect 479604 624698 479786 624934
rect 480022 624698 480204 624934
rect 479604 589254 480204 624698
rect 479604 589018 479786 589254
rect 480022 589018 480204 589254
rect 479604 588934 480204 589018
rect 479604 588698 479786 588934
rect 480022 588698 480204 588934
rect 479604 553254 480204 588698
rect 479604 553018 479786 553254
rect 480022 553018 480204 553254
rect 479604 552934 480204 553018
rect 479604 552698 479786 552934
rect 480022 552698 480204 552934
rect 479604 517254 480204 552698
rect 479604 517018 479786 517254
rect 480022 517018 480204 517254
rect 479604 516934 480204 517018
rect 479604 516698 479786 516934
rect 480022 516698 480204 516934
rect 479604 481254 480204 516698
rect 479604 481018 479786 481254
rect 480022 481018 480204 481254
rect 479604 480934 480204 481018
rect 479604 480698 479786 480934
rect 480022 480698 480204 480934
rect 479604 445254 480204 480698
rect 479604 445018 479786 445254
rect 480022 445018 480204 445254
rect 479604 444934 480204 445018
rect 479604 444698 479786 444934
rect 480022 444698 480204 444934
rect 479604 409254 480204 444698
rect 479604 409018 479786 409254
rect 480022 409018 480204 409254
rect 479604 408934 480204 409018
rect 479604 408698 479786 408934
rect 480022 408698 480204 408934
rect 479604 373254 480204 408698
rect 479604 373018 479786 373254
rect 480022 373018 480204 373254
rect 479604 372934 480204 373018
rect 479604 372698 479786 372934
rect 480022 372698 480204 372934
rect 479604 337254 480204 372698
rect 479604 337018 479786 337254
rect 480022 337018 480204 337254
rect 479604 336934 480204 337018
rect 479604 336698 479786 336934
rect 480022 336698 480204 336934
rect 479604 301254 480204 336698
rect 479604 301018 479786 301254
rect 480022 301018 480204 301254
rect 479604 300934 480204 301018
rect 479604 300698 479786 300934
rect 480022 300698 480204 300934
rect 479604 265254 480204 300698
rect 479604 265018 479786 265254
rect 480022 265018 480204 265254
rect 479604 264934 480204 265018
rect 479604 264698 479786 264934
rect 480022 264698 480204 264934
rect 479604 229254 480204 264698
rect 479604 229018 479786 229254
rect 480022 229018 480204 229254
rect 479604 228934 480204 229018
rect 479604 228698 479786 228934
rect 480022 228698 480204 228934
rect 479604 193254 480204 228698
rect 479604 193018 479786 193254
rect 480022 193018 480204 193254
rect 479604 192934 480204 193018
rect 479604 192698 479786 192934
rect 480022 192698 480204 192934
rect 479604 157254 480204 192698
rect 479604 157018 479786 157254
rect 480022 157018 480204 157254
rect 479604 156934 480204 157018
rect 479604 156698 479786 156934
rect 480022 156698 480204 156934
rect 479604 121254 480204 156698
rect 479604 121018 479786 121254
rect 480022 121018 480204 121254
rect 479604 120934 480204 121018
rect 479604 120698 479786 120934
rect 480022 120698 480204 120934
rect 479604 85254 480204 120698
rect 479604 85018 479786 85254
rect 480022 85018 480204 85254
rect 479604 84934 480204 85018
rect 479604 84698 479786 84934
rect 480022 84698 480204 84934
rect 479604 49254 480204 84698
rect 479604 49018 479786 49254
rect 480022 49018 480204 49254
rect 479604 48934 480204 49018
rect 479604 48698 479786 48934
rect 480022 48698 480204 48934
rect 479604 13254 480204 48698
rect 486804 705758 487404 705780
rect 486804 705522 486986 705758
rect 487222 705522 487404 705758
rect 486804 705438 487404 705522
rect 486804 705202 486986 705438
rect 487222 705202 487404 705438
rect 486804 668454 487404 705202
rect 486804 668218 486986 668454
rect 487222 668218 487404 668454
rect 486804 668134 487404 668218
rect 486804 667898 486986 668134
rect 487222 667898 487404 668134
rect 486804 632454 487404 667898
rect 486804 632218 486986 632454
rect 487222 632218 487404 632454
rect 486804 632134 487404 632218
rect 486804 631898 486986 632134
rect 487222 631898 487404 632134
rect 486804 596454 487404 631898
rect 486804 596218 486986 596454
rect 487222 596218 487404 596454
rect 486804 596134 487404 596218
rect 486804 595898 486986 596134
rect 487222 595898 487404 596134
rect 486804 560454 487404 595898
rect 486804 560218 486986 560454
rect 487222 560218 487404 560454
rect 486804 560134 487404 560218
rect 486804 559898 486986 560134
rect 487222 559898 487404 560134
rect 486804 524454 487404 559898
rect 486804 524218 486986 524454
rect 487222 524218 487404 524454
rect 486804 524134 487404 524218
rect 486804 523898 486986 524134
rect 487222 523898 487404 524134
rect 486804 488454 487404 523898
rect 486804 488218 486986 488454
rect 487222 488218 487404 488454
rect 486804 488134 487404 488218
rect 486804 487898 486986 488134
rect 487222 487898 487404 488134
rect 486804 452454 487404 487898
rect 486804 452218 486986 452454
rect 487222 452218 487404 452454
rect 486804 452134 487404 452218
rect 486804 451898 486986 452134
rect 487222 451898 487404 452134
rect 486804 416454 487404 451898
rect 486804 416218 486986 416454
rect 487222 416218 487404 416454
rect 486804 416134 487404 416218
rect 486804 415898 486986 416134
rect 487222 415898 487404 416134
rect 486804 380454 487404 415898
rect 486804 380218 486986 380454
rect 487222 380218 487404 380454
rect 486804 380134 487404 380218
rect 486804 379898 486986 380134
rect 487222 379898 487404 380134
rect 486804 344454 487404 379898
rect 486804 344218 486986 344454
rect 487222 344218 487404 344454
rect 486804 344134 487404 344218
rect 486804 343898 486986 344134
rect 487222 343898 487404 344134
rect 486804 308454 487404 343898
rect 486804 308218 486986 308454
rect 487222 308218 487404 308454
rect 486804 308134 487404 308218
rect 486804 307898 486986 308134
rect 487222 307898 487404 308134
rect 486804 272454 487404 307898
rect 486804 272218 486986 272454
rect 487222 272218 487404 272454
rect 486804 272134 487404 272218
rect 486804 271898 486986 272134
rect 487222 271898 487404 272134
rect 486804 236454 487404 271898
rect 486804 236218 486986 236454
rect 487222 236218 487404 236454
rect 486804 236134 487404 236218
rect 486804 235898 486986 236134
rect 487222 235898 487404 236134
rect 486804 200454 487404 235898
rect 486804 200218 486986 200454
rect 487222 200218 487404 200454
rect 486804 200134 487404 200218
rect 486804 199898 486986 200134
rect 487222 199898 487404 200134
rect 486804 164454 487404 199898
rect 486804 164218 486986 164454
rect 487222 164218 487404 164454
rect 486804 164134 487404 164218
rect 486804 163898 486986 164134
rect 487222 163898 487404 164134
rect 486804 128454 487404 163898
rect 486804 128218 486986 128454
rect 487222 128218 487404 128454
rect 486804 128134 487404 128218
rect 486804 127898 486986 128134
rect 487222 127898 487404 128134
rect 486804 92454 487404 127898
rect 486804 92218 486986 92454
rect 487222 92218 487404 92454
rect 486804 92134 487404 92218
rect 486804 91898 486986 92134
rect 487222 91898 487404 92134
rect 486804 56454 487404 91898
rect 486804 56218 486986 56454
rect 487222 56218 487404 56454
rect 486804 56134 487404 56218
rect 486804 55898 486986 56134
rect 487222 55898 487404 56134
rect 481587 29068 481653 29069
rect 481587 29004 481588 29068
rect 481652 29004 481653 29068
rect 481587 29003 481653 29004
rect 481590 28797 481650 29003
rect 481587 28796 481653 28797
rect 481587 28732 481588 28796
rect 481652 28732 481653 28796
rect 481587 28731 481653 28732
rect 479604 13018 479786 13254
rect 480022 13018 480204 13254
rect 479604 12934 480204 13018
rect 479604 12698 479786 12934
rect 480022 12698 480204 12934
rect 461604 -7022 461786 -6786
rect 462022 -7022 462204 -6786
rect 461604 -7106 462204 -7022
rect 461604 -7342 461786 -7106
rect 462022 -7342 462204 -7106
rect 461604 -7364 462204 -7342
rect 479604 -5866 480204 12698
rect 486804 20454 487404 55898
rect 486804 20218 486986 20454
rect 487222 20218 487404 20454
rect 486804 20134 487404 20218
rect 486804 19898 486986 20134
rect 487222 19898 487404 20134
rect 486804 -1266 487404 19898
rect 486804 -1502 486986 -1266
rect 487222 -1502 487404 -1266
rect 486804 -1586 487404 -1502
rect 486804 -1822 486986 -1586
rect 487222 -1822 487404 -1586
rect 486804 -1844 487404 -1822
rect 490404 672054 491004 707042
rect 490404 671818 490586 672054
rect 490822 671818 491004 672054
rect 490404 671734 491004 671818
rect 490404 671498 490586 671734
rect 490822 671498 491004 671734
rect 490404 636054 491004 671498
rect 490404 635818 490586 636054
rect 490822 635818 491004 636054
rect 490404 635734 491004 635818
rect 490404 635498 490586 635734
rect 490822 635498 491004 635734
rect 490404 600054 491004 635498
rect 490404 599818 490586 600054
rect 490822 599818 491004 600054
rect 490404 599734 491004 599818
rect 490404 599498 490586 599734
rect 490822 599498 491004 599734
rect 490404 564054 491004 599498
rect 490404 563818 490586 564054
rect 490822 563818 491004 564054
rect 490404 563734 491004 563818
rect 490404 563498 490586 563734
rect 490822 563498 491004 563734
rect 490404 528054 491004 563498
rect 490404 527818 490586 528054
rect 490822 527818 491004 528054
rect 490404 527734 491004 527818
rect 490404 527498 490586 527734
rect 490822 527498 491004 527734
rect 490404 492054 491004 527498
rect 490404 491818 490586 492054
rect 490822 491818 491004 492054
rect 490404 491734 491004 491818
rect 490404 491498 490586 491734
rect 490822 491498 491004 491734
rect 490404 456054 491004 491498
rect 490404 455818 490586 456054
rect 490822 455818 491004 456054
rect 490404 455734 491004 455818
rect 490404 455498 490586 455734
rect 490822 455498 491004 455734
rect 490404 420054 491004 455498
rect 490404 419818 490586 420054
rect 490822 419818 491004 420054
rect 490404 419734 491004 419818
rect 490404 419498 490586 419734
rect 490822 419498 491004 419734
rect 490404 384054 491004 419498
rect 490404 383818 490586 384054
rect 490822 383818 491004 384054
rect 490404 383734 491004 383818
rect 490404 383498 490586 383734
rect 490822 383498 491004 383734
rect 490404 348054 491004 383498
rect 490404 347818 490586 348054
rect 490822 347818 491004 348054
rect 490404 347734 491004 347818
rect 490404 347498 490586 347734
rect 490822 347498 491004 347734
rect 490404 312054 491004 347498
rect 490404 311818 490586 312054
rect 490822 311818 491004 312054
rect 490404 311734 491004 311818
rect 490404 311498 490586 311734
rect 490822 311498 491004 311734
rect 490404 276054 491004 311498
rect 490404 275818 490586 276054
rect 490822 275818 491004 276054
rect 490404 275734 491004 275818
rect 490404 275498 490586 275734
rect 490822 275498 491004 275734
rect 490404 240054 491004 275498
rect 490404 239818 490586 240054
rect 490822 239818 491004 240054
rect 490404 239734 491004 239818
rect 490404 239498 490586 239734
rect 490822 239498 491004 239734
rect 490404 204054 491004 239498
rect 490404 203818 490586 204054
rect 490822 203818 491004 204054
rect 490404 203734 491004 203818
rect 490404 203498 490586 203734
rect 490822 203498 491004 203734
rect 490404 168054 491004 203498
rect 490404 167818 490586 168054
rect 490822 167818 491004 168054
rect 490404 167734 491004 167818
rect 490404 167498 490586 167734
rect 490822 167498 491004 167734
rect 490404 132054 491004 167498
rect 490404 131818 490586 132054
rect 490822 131818 491004 132054
rect 490404 131734 491004 131818
rect 490404 131498 490586 131734
rect 490822 131498 491004 131734
rect 490404 96054 491004 131498
rect 490404 95818 490586 96054
rect 490822 95818 491004 96054
rect 490404 95734 491004 95818
rect 490404 95498 490586 95734
rect 490822 95498 491004 95734
rect 490404 60054 491004 95498
rect 494004 675654 494604 708882
rect 494004 675418 494186 675654
rect 494422 675418 494604 675654
rect 494004 675334 494604 675418
rect 494004 675098 494186 675334
rect 494422 675098 494604 675334
rect 494004 639654 494604 675098
rect 494004 639418 494186 639654
rect 494422 639418 494604 639654
rect 494004 639334 494604 639418
rect 494004 639098 494186 639334
rect 494422 639098 494604 639334
rect 494004 603654 494604 639098
rect 494004 603418 494186 603654
rect 494422 603418 494604 603654
rect 494004 603334 494604 603418
rect 494004 603098 494186 603334
rect 494422 603098 494604 603334
rect 494004 567654 494604 603098
rect 494004 567418 494186 567654
rect 494422 567418 494604 567654
rect 494004 567334 494604 567418
rect 494004 567098 494186 567334
rect 494422 567098 494604 567334
rect 494004 531654 494604 567098
rect 494004 531418 494186 531654
rect 494422 531418 494604 531654
rect 494004 531334 494604 531418
rect 494004 531098 494186 531334
rect 494422 531098 494604 531334
rect 494004 495654 494604 531098
rect 494004 495418 494186 495654
rect 494422 495418 494604 495654
rect 494004 495334 494604 495418
rect 494004 495098 494186 495334
rect 494422 495098 494604 495334
rect 494004 459654 494604 495098
rect 494004 459418 494186 459654
rect 494422 459418 494604 459654
rect 494004 459334 494604 459418
rect 494004 459098 494186 459334
rect 494422 459098 494604 459334
rect 494004 423654 494604 459098
rect 494004 423418 494186 423654
rect 494422 423418 494604 423654
rect 494004 423334 494604 423418
rect 494004 423098 494186 423334
rect 494422 423098 494604 423334
rect 494004 387654 494604 423098
rect 494004 387418 494186 387654
rect 494422 387418 494604 387654
rect 494004 387334 494604 387418
rect 494004 387098 494186 387334
rect 494422 387098 494604 387334
rect 494004 351654 494604 387098
rect 494004 351418 494186 351654
rect 494422 351418 494604 351654
rect 494004 351334 494604 351418
rect 494004 351098 494186 351334
rect 494422 351098 494604 351334
rect 494004 315654 494604 351098
rect 494004 315418 494186 315654
rect 494422 315418 494604 315654
rect 494004 315334 494604 315418
rect 494004 315098 494186 315334
rect 494422 315098 494604 315334
rect 494004 279654 494604 315098
rect 494004 279418 494186 279654
rect 494422 279418 494604 279654
rect 494004 279334 494604 279418
rect 494004 279098 494186 279334
rect 494422 279098 494604 279334
rect 494004 243654 494604 279098
rect 494004 243418 494186 243654
rect 494422 243418 494604 243654
rect 494004 243334 494604 243418
rect 494004 243098 494186 243334
rect 494422 243098 494604 243334
rect 494004 207654 494604 243098
rect 494004 207418 494186 207654
rect 494422 207418 494604 207654
rect 494004 207334 494604 207418
rect 494004 207098 494186 207334
rect 494422 207098 494604 207334
rect 494004 171654 494604 207098
rect 494004 171418 494186 171654
rect 494422 171418 494604 171654
rect 494004 171334 494604 171418
rect 494004 171098 494186 171334
rect 494422 171098 494604 171334
rect 494004 135654 494604 171098
rect 494004 135418 494186 135654
rect 494422 135418 494604 135654
rect 494004 135334 494604 135418
rect 494004 135098 494186 135334
rect 494422 135098 494604 135334
rect 494004 99654 494604 135098
rect 494004 99418 494186 99654
rect 494422 99418 494604 99654
rect 494004 99334 494604 99418
rect 494004 99098 494186 99334
rect 494422 99098 494604 99334
rect 492627 76124 492693 76125
rect 492627 76060 492628 76124
rect 492692 76060 492693 76124
rect 492627 76059 492693 76060
rect 492630 75853 492690 76059
rect 492627 75852 492693 75853
rect 492627 75788 492628 75852
rect 492692 75788 492693 75852
rect 492627 75787 492693 75788
rect 490404 59818 490586 60054
rect 490822 59818 491004 60054
rect 490404 59734 491004 59818
rect 490404 59498 490586 59734
rect 490822 59498 491004 59734
rect 490404 24054 491004 59498
rect 490404 23818 490586 24054
rect 490822 23818 491004 24054
rect 490404 23734 491004 23818
rect 490404 23498 490586 23734
rect 490822 23498 491004 23734
rect 490404 -3106 491004 23498
rect 490404 -3342 490586 -3106
rect 490822 -3342 491004 -3106
rect 490404 -3426 491004 -3342
rect 490404 -3662 490586 -3426
rect 490822 -3662 491004 -3426
rect 490404 -3684 491004 -3662
rect 494004 63654 494604 99098
rect 494004 63418 494186 63654
rect 494422 63418 494604 63654
rect 494004 63334 494604 63418
rect 494004 63098 494186 63334
rect 494422 63098 494604 63334
rect 494004 27654 494604 63098
rect 494004 27418 494186 27654
rect 494422 27418 494604 27654
rect 494004 27334 494604 27418
rect 494004 27098 494186 27334
rect 494422 27098 494604 27334
rect 494004 -4946 494604 27098
rect 494004 -5182 494186 -4946
rect 494422 -5182 494604 -4946
rect 494004 -5266 494604 -5182
rect 494004 -5502 494186 -5266
rect 494422 -5502 494604 -5266
rect 494004 -5524 494604 -5502
rect 497604 679254 498204 710722
rect 515604 710358 516204 711300
rect 515604 710122 515786 710358
rect 516022 710122 516204 710358
rect 515604 710038 516204 710122
rect 515604 709802 515786 710038
rect 516022 709802 516204 710038
rect 512004 708518 512604 709460
rect 512004 708282 512186 708518
rect 512422 708282 512604 708518
rect 512004 708198 512604 708282
rect 512004 707962 512186 708198
rect 512422 707962 512604 708198
rect 508404 706678 509004 707620
rect 508404 706442 508586 706678
rect 508822 706442 509004 706678
rect 508404 706358 509004 706442
rect 508404 706122 508586 706358
rect 508822 706122 509004 706358
rect 497604 679018 497786 679254
rect 498022 679018 498204 679254
rect 497604 678934 498204 679018
rect 497604 678698 497786 678934
rect 498022 678698 498204 678934
rect 497604 643254 498204 678698
rect 497604 643018 497786 643254
rect 498022 643018 498204 643254
rect 497604 642934 498204 643018
rect 497604 642698 497786 642934
rect 498022 642698 498204 642934
rect 497604 607254 498204 642698
rect 497604 607018 497786 607254
rect 498022 607018 498204 607254
rect 497604 606934 498204 607018
rect 497604 606698 497786 606934
rect 498022 606698 498204 606934
rect 497604 571254 498204 606698
rect 497604 571018 497786 571254
rect 498022 571018 498204 571254
rect 497604 570934 498204 571018
rect 497604 570698 497786 570934
rect 498022 570698 498204 570934
rect 497604 535254 498204 570698
rect 497604 535018 497786 535254
rect 498022 535018 498204 535254
rect 497604 534934 498204 535018
rect 497604 534698 497786 534934
rect 498022 534698 498204 534934
rect 497604 499254 498204 534698
rect 497604 499018 497786 499254
rect 498022 499018 498204 499254
rect 497604 498934 498204 499018
rect 497604 498698 497786 498934
rect 498022 498698 498204 498934
rect 497604 463254 498204 498698
rect 497604 463018 497786 463254
rect 498022 463018 498204 463254
rect 497604 462934 498204 463018
rect 497604 462698 497786 462934
rect 498022 462698 498204 462934
rect 497604 427254 498204 462698
rect 497604 427018 497786 427254
rect 498022 427018 498204 427254
rect 497604 426934 498204 427018
rect 497604 426698 497786 426934
rect 498022 426698 498204 426934
rect 497604 391254 498204 426698
rect 497604 391018 497786 391254
rect 498022 391018 498204 391254
rect 497604 390934 498204 391018
rect 497604 390698 497786 390934
rect 498022 390698 498204 390934
rect 497604 355254 498204 390698
rect 497604 355018 497786 355254
rect 498022 355018 498204 355254
rect 497604 354934 498204 355018
rect 497604 354698 497786 354934
rect 498022 354698 498204 354934
rect 497604 319254 498204 354698
rect 497604 319018 497786 319254
rect 498022 319018 498204 319254
rect 497604 318934 498204 319018
rect 497604 318698 497786 318934
rect 498022 318698 498204 318934
rect 497604 283254 498204 318698
rect 497604 283018 497786 283254
rect 498022 283018 498204 283254
rect 497604 282934 498204 283018
rect 497604 282698 497786 282934
rect 498022 282698 498204 282934
rect 497604 247254 498204 282698
rect 497604 247018 497786 247254
rect 498022 247018 498204 247254
rect 497604 246934 498204 247018
rect 497604 246698 497786 246934
rect 498022 246698 498204 246934
rect 497604 211254 498204 246698
rect 497604 211018 497786 211254
rect 498022 211018 498204 211254
rect 497604 210934 498204 211018
rect 497604 210698 497786 210934
rect 498022 210698 498204 210934
rect 497604 175254 498204 210698
rect 497604 175018 497786 175254
rect 498022 175018 498204 175254
rect 497604 174934 498204 175018
rect 497604 174698 497786 174934
rect 498022 174698 498204 174934
rect 497604 139254 498204 174698
rect 497604 139018 497786 139254
rect 498022 139018 498204 139254
rect 497604 138934 498204 139018
rect 497604 138698 497786 138934
rect 498022 138698 498204 138934
rect 497604 103254 498204 138698
rect 497604 103018 497786 103254
rect 498022 103018 498204 103254
rect 497604 102934 498204 103018
rect 497604 102698 497786 102934
rect 498022 102698 498204 102934
rect 497604 67254 498204 102698
rect 497604 67018 497786 67254
rect 498022 67018 498204 67254
rect 497604 66934 498204 67018
rect 497604 66698 497786 66934
rect 498022 66698 498204 66934
rect 497604 31254 498204 66698
rect 497604 31018 497786 31254
rect 498022 31018 498204 31254
rect 497604 30934 498204 31018
rect 497604 30698 497786 30934
rect 498022 30698 498204 30934
rect 479604 -6102 479786 -5866
rect 480022 -6102 480204 -5866
rect 479604 -6186 480204 -6102
rect 479604 -6422 479786 -6186
rect 480022 -6422 480204 -6186
rect 479604 -7364 480204 -6422
rect 497604 -6786 498204 30698
rect 504804 704838 505404 705780
rect 504804 704602 504986 704838
rect 505222 704602 505404 704838
rect 504804 704518 505404 704602
rect 504804 704282 504986 704518
rect 505222 704282 505404 704518
rect 504804 686454 505404 704282
rect 504804 686218 504986 686454
rect 505222 686218 505404 686454
rect 504804 686134 505404 686218
rect 504804 685898 504986 686134
rect 505222 685898 505404 686134
rect 504804 650454 505404 685898
rect 504804 650218 504986 650454
rect 505222 650218 505404 650454
rect 504804 650134 505404 650218
rect 504804 649898 504986 650134
rect 505222 649898 505404 650134
rect 504804 614454 505404 649898
rect 504804 614218 504986 614454
rect 505222 614218 505404 614454
rect 504804 614134 505404 614218
rect 504804 613898 504986 614134
rect 505222 613898 505404 614134
rect 504804 578454 505404 613898
rect 504804 578218 504986 578454
rect 505222 578218 505404 578454
rect 504804 578134 505404 578218
rect 504804 577898 504986 578134
rect 505222 577898 505404 578134
rect 504804 542454 505404 577898
rect 504804 542218 504986 542454
rect 505222 542218 505404 542454
rect 504804 542134 505404 542218
rect 504804 541898 504986 542134
rect 505222 541898 505404 542134
rect 504804 506454 505404 541898
rect 504804 506218 504986 506454
rect 505222 506218 505404 506454
rect 504804 506134 505404 506218
rect 504804 505898 504986 506134
rect 505222 505898 505404 506134
rect 504804 470454 505404 505898
rect 504804 470218 504986 470454
rect 505222 470218 505404 470454
rect 504804 470134 505404 470218
rect 504804 469898 504986 470134
rect 505222 469898 505404 470134
rect 504804 434454 505404 469898
rect 504804 434218 504986 434454
rect 505222 434218 505404 434454
rect 504804 434134 505404 434218
rect 504804 433898 504986 434134
rect 505222 433898 505404 434134
rect 504804 398454 505404 433898
rect 504804 398218 504986 398454
rect 505222 398218 505404 398454
rect 504804 398134 505404 398218
rect 504804 397898 504986 398134
rect 505222 397898 505404 398134
rect 504804 362454 505404 397898
rect 504804 362218 504986 362454
rect 505222 362218 505404 362454
rect 504804 362134 505404 362218
rect 504804 361898 504986 362134
rect 505222 361898 505404 362134
rect 504804 326454 505404 361898
rect 504804 326218 504986 326454
rect 505222 326218 505404 326454
rect 504804 326134 505404 326218
rect 504804 325898 504986 326134
rect 505222 325898 505404 326134
rect 504804 290454 505404 325898
rect 504804 290218 504986 290454
rect 505222 290218 505404 290454
rect 504804 290134 505404 290218
rect 504804 289898 504986 290134
rect 505222 289898 505404 290134
rect 504804 254454 505404 289898
rect 504804 254218 504986 254454
rect 505222 254218 505404 254454
rect 504804 254134 505404 254218
rect 504804 253898 504986 254134
rect 505222 253898 505404 254134
rect 504804 218454 505404 253898
rect 504804 218218 504986 218454
rect 505222 218218 505404 218454
rect 504804 218134 505404 218218
rect 504804 217898 504986 218134
rect 505222 217898 505404 218134
rect 504804 182454 505404 217898
rect 504804 182218 504986 182454
rect 505222 182218 505404 182454
rect 504804 182134 505404 182218
rect 504804 181898 504986 182134
rect 505222 181898 505404 182134
rect 504804 146454 505404 181898
rect 504804 146218 504986 146454
rect 505222 146218 505404 146454
rect 504804 146134 505404 146218
rect 504804 145898 504986 146134
rect 505222 145898 505404 146134
rect 504804 110454 505404 145898
rect 504804 110218 504986 110454
rect 505222 110218 505404 110454
rect 504804 110134 505404 110218
rect 504804 109898 504986 110134
rect 505222 109898 505404 110134
rect 504804 74454 505404 109898
rect 504804 74218 504986 74454
rect 505222 74218 505404 74454
rect 504804 74134 505404 74218
rect 504804 73898 504986 74134
rect 505222 73898 505404 74134
rect 504804 38454 505404 73898
rect 504804 38218 504986 38454
rect 505222 38218 505404 38454
rect 504804 38134 505404 38218
rect 504804 37898 504986 38134
rect 505222 37898 505404 38134
rect 504804 2454 505404 37898
rect 504804 2218 504986 2454
rect 505222 2218 505404 2454
rect 504804 2134 505404 2218
rect 504804 1898 504986 2134
rect 505222 1898 505404 2134
rect 504804 -346 505404 1898
rect 504804 -582 504986 -346
rect 505222 -582 505404 -346
rect 504804 -666 505404 -582
rect 504804 -902 504986 -666
rect 505222 -902 505404 -666
rect 504804 -1844 505404 -902
rect 508404 690054 509004 706122
rect 508404 689818 508586 690054
rect 508822 689818 509004 690054
rect 508404 689734 509004 689818
rect 508404 689498 508586 689734
rect 508822 689498 509004 689734
rect 508404 654054 509004 689498
rect 508404 653818 508586 654054
rect 508822 653818 509004 654054
rect 508404 653734 509004 653818
rect 508404 653498 508586 653734
rect 508822 653498 509004 653734
rect 508404 618054 509004 653498
rect 508404 617818 508586 618054
rect 508822 617818 509004 618054
rect 508404 617734 509004 617818
rect 508404 617498 508586 617734
rect 508822 617498 509004 617734
rect 508404 582054 509004 617498
rect 508404 581818 508586 582054
rect 508822 581818 509004 582054
rect 508404 581734 509004 581818
rect 508404 581498 508586 581734
rect 508822 581498 509004 581734
rect 508404 546054 509004 581498
rect 508404 545818 508586 546054
rect 508822 545818 509004 546054
rect 508404 545734 509004 545818
rect 508404 545498 508586 545734
rect 508822 545498 509004 545734
rect 508404 510054 509004 545498
rect 508404 509818 508586 510054
rect 508822 509818 509004 510054
rect 508404 509734 509004 509818
rect 508404 509498 508586 509734
rect 508822 509498 509004 509734
rect 508404 474054 509004 509498
rect 508404 473818 508586 474054
rect 508822 473818 509004 474054
rect 508404 473734 509004 473818
rect 508404 473498 508586 473734
rect 508822 473498 509004 473734
rect 508404 438054 509004 473498
rect 508404 437818 508586 438054
rect 508822 437818 509004 438054
rect 508404 437734 509004 437818
rect 508404 437498 508586 437734
rect 508822 437498 509004 437734
rect 508404 402054 509004 437498
rect 508404 401818 508586 402054
rect 508822 401818 509004 402054
rect 508404 401734 509004 401818
rect 508404 401498 508586 401734
rect 508822 401498 509004 401734
rect 508404 366054 509004 401498
rect 508404 365818 508586 366054
rect 508822 365818 509004 366054
rect 508404 365734 509004 365818
rect 508404 365498 508586 365734
rect 508822 365498 509004 365734
rect 508404 330054 509004 365498
rect 508404 329818 508586 330054
rect 508822 329818 509004 330054
rect 508404 329734 509004 329818
rect 508404 329498 508586 329734
rect 508822 329498 509004 329734
rect 508404 294054 509004 329498
rect 508404 293818 508586 294054
rect 508822 293818 509004 294054
rect 508404 293734 509004 293818
rect 508404 293498 508586 293734
rect 508822 293498 509004 293734
rect 508404 258054 509004 293498
rect 508404 257818 508586 258054
rect 508822 257818 509004 258054
rect 508404 257734 509004 257818
rect 508404 257498 508586 257734
rect 508822 257498 509004 257734
rect 508404 222054 509004 257498
rect 508404 221818 508586 222054
rect 508822 221818 509004 222054
rect 508404 221734 509004 221818
rect 508404 221498 508586 221734
rect 508822 221498 509004 221734
rect 508404 186054 509004 221498
rect 508404 185818 508586 186054
rect 508822 185818 509004 186054
rect 508404 185734 509004 185818
rect 508404 185498 508586 185734
rect 508822 185498 509004 185734
rect 508404 150054 509004 185498
rect 508404 149818 508586 150054
rect 508822 149818 509004 150054
rect 508404 149734 509004 149818
rect 508404 149498 508586 149734
rect 508822 149498 509004 149734
rect 508404 114054 509004 149498
rect 508404 113818 508586 114054
rect 508822 113818 509004 114054
rect 508404 113734 509004 113818
rect 508404 113498 508586 113734
rect 508822 113498 509004 113734
rect 508404 78054 509004 113498
rect 508404 77818 508586 78054
rect 508822 77818 509004 78054
rect 508404 77734 509004 77818
rect 508404 77498 508586 77734
rect 508822 77498 509004 77734
rect 508404 42054 509004 77498
rect 508404 41818 508586 42054
rect 508822 41818 509004 42054
rect 508404 41734 509004 41818
rect 508404 41498 508586 41734
rect 508822 41498 509004 41734
rect 508404 6054 509004 41498
rect 508404 5818 508586 6054
rect 508822 5818 509004 6054
rect 508404 5734 509004 5818
rect 508404 5498 508586 5734
rect 508822 5498 509004 5734
rect 508404 -2186 509004 5498
rect 508404 -2422 508586 -2186
rect 508822 -2422 509004 -2186
rect 508404 -2506 509004 -2422
rect 508404 -2742 508586 -2506
rect 508822 -2742 509004 -2506
rect 508404 -3684 509004 -2742
rect 512004 693654 512604 707962
rect 512004 693418 512186 693654
rect 512422 693418 512604 693654
rect 512004 693334 512604 693418
rect 512004 693098 512186 693334
rect 512422 693098 512604 693334
rect 512004 657654 512604 693098
rect 512004 657418 512186 657654
rect 512422 657418 512604 657654
rect 512004 657334 512604 657418
rect 512004 657098 512186 657334
rect 512422 657098 512604 657334
rect 512004 621654 512604 657098
rect 512004 621418 512186 621654
rect 512422 621418 512604 621654
rect 512004 621334 512604 621418
rect 512004 621098 512186 621334
rect 512422 621098 512604 621334
rect 512004 585654 512604 621098
rect 512004 585418 512186 585654
rect 512422 585418 512604 585654
rect 512004 585334 512604 585418
rect 512004 585098 512186 585334
rect 512422 585098 512604 585334
rect 512004 549654 512604 585098
rect 512004 549418 512186 549654
rect 512422 549418 512604 549654
rect 512004 549334 512604 549418
rect 512004 549098 512186 549334
rect 512422 549098 512604 549334
rect 512004 513654 512604 549098
rect 512004 513418 512186 513654
rect 512422 513418 512604 513654
rect 512004 513334 512604 513418
rect 512004 513098 512186 513334
rect 512422 513098 512604 513334
rect 512004 477654 512604 513098
rect 512004 477418 512186 477654
rect 512422 477418 512604 477654
rect 512004 477334 512604 477418
rect 512004 477098 512186 477334
rect 512422 477098 512604 477334
rect 512004 441654 512604 477098
rect 512004 441418 512186 441654
rect 512422 441418 512604 441654
rect 512004 441334 512604 441418
rect 512004 441098 512186 441334
rect 512422 441098 512604 441334
rect 512004 405654 512604 441098
rect 512004 405418 512186 405654
rect 512422 405418 512604 405654
rect 512004 405334 512604 405418
rect 512004 405098 512186 405334
rect 512422 405098 512604 405334
rect 512004 369654 512604 405098
rect 512004 369418 512186 369654
rect 512422 369418 512604 369654
rect 512004 369334 512604 369418
rect 512004 369098 512186 369334
rect 512422 369098 512604 369334
rect 512004 333654 512604 369098
rect 512004 333418 512186 333654
rect 512422 333418 512604 333654
rect 512004 333334 512604 333418
rect 512004 333098 512186 333334
rect 512422 333098 512604 333334
rect 512004 297654 512604 333098
rect 512004 297418 512186 297654
rect 512422 297418 512604 297654
rect 512004 297334 512604 297418
rect 512004 297098 512186 297334
rect 512422 297098 512604 297334
rect 512004 261654 512604 297098
rect 512004 261418 512186 261654
rect 512422 261418 512604 261654
rect 512004 261334 512604 261418
rect 512004 261098 512186 261334
rect 512422 261098 512604 261334
rect 512004 225654 512604 261098
rect 512004 225418 512186 225654
rect 512422 225418 512604 225654
rect 512004 225334 512604 225418
rect 512004 225098 512186 225334
rect 512422 225098 512604 225334
rect 512004 189654 512604 225098
rect 512004 189418 512186 189654
rect 512422 189418 512604 189654
rect 512004 189334 512604 189418
rect 512004 189098 512186 189334
rect 512422 189098 512604 189334
rect 512004 153654 512604 189098
rect 512004 153418 512186 153654
rect 512422 153418 512604 153654
rect 512004 153334 512604 153418
rect 512004 153098 512186 153334
rect 512422 153098 512604 153334
rect 512004 117654 512604 153098
rect 512004 117418 512186 117654
rect 512422 117418 512604 117654
rect 512004 117334 512604 117418
rect 512004 117098 512186 117334
rect 512422 117098 512604 117334
rect 512004 81654 512604 117098
rect 512004 81418 512186 81654
rect 512422 81418 512604 81654
rect 512004 81334 512604 81418
rect 512004 81098 512186 81334
rect 512422 81098 512604 81334
rect 512004 45654 512604 81098
rect 512004 45418 512186 45654
rect 512422 45418 512604 45654
rect 512004 45334 512604 45418
rect 512004 45098 512186 45334
rect 512422 45098 512604 45334
rect 512004 9654 512604 45098
rect 512004 9418 512186 9654
rect 512422 9418 512604 9654
rect 512004 9334 512604 9418
rect 512004 9098 512186 9334
rect 512422 9098 512604 9334
rect 512004 -4026 512604 9098
rect 512004 -4262 512186 -4026
rect 512422 -4262 512604 -4026
rect 512004 -4346 512604 -4262
rect 512004 -4582 512186 -4346
rect 512422 -4582 512604 -4346
rect 512004 -5524 512604 -4582
rect 515604 697254 516204 709802
rect 533604 711278 534204 711300
rect 533604 711042 533786 711278
rect 534022 711042 534204 711278
rect 533604 710958 534204 711042
rect 533604 710722 533786 710958
rect 534022 710722 534204 710958
rect 530004 709438 530604 709460
rect 530004 709202 530186 709438
rect 530422 709202 530604 709438
rect 530004 709118 530604 709202
rect 530004 708882 530186 709118
rect 530422 708882 530604 709118
rect 526404 707598 527004 707620
rect 526404 707362 526586 707598
rect 526822 707362 527004 707598
rect 526404 707278 527004 707362
rect 526404 707042 526586 707278
rect 526822 707042 527004 707278
rect 515604 697018 515786 697254
rect 516022 697018 516204 697254
rect 515604 696934 516204 697018
rect 515604 696698 515786 696934
rect 516022 696698 516204 696934
rect 515604 661254 516204 696698
rect 515604 661018 515786 661254
rect 516022 661018 516204 661254
rect 515604 660934 516204 661018
rect 515604 660698 515786 660934
rect 516022 660698 516204 660934
rect 515604 625254 516204 660698
rect 515604 625018 515786 625254
rect 516022 625018 516204 625254
rect 515604 624934 516204 625018
rect 515604 624698 515786 624934
rect 516022 624698 516204 624934
rect 515604 589254 516204 624698
rect 515604 589018 515786 589254
rect 516022 589018 516204 589254
rect 515604 588934 516204 589018
rect 515604 588698 515786 588934
rect 516022 588698 516204 588934
rect 515604 553254 516204 588698
rect 515604 553018 515786 553254
rect 516022 553018 516204 553254
rect 515604 552934 516204 553018
rect 515604 552698 515786 552934
rect 516022 552698 516204 552934
rect 515604 517254 516204 552698
rect 515604 517018 515786 517254
rect 516022 517018 516204 517254
rect 515604 516934 516204 517018
rect 515604 516698 515786 516934
rect 516022 516698 516204 516934
rect 515604 481254 516204 516698
rect 515604 481018 515786 481254
rect 516022 481018 516204 481254
rect 515604 480934 516204 481018
rect 515604 480698 515786 480934
rect 516022 480698 516204 480934
rect 515604 445254 516204 480698
rect 515604 445018 515786 445254
rect 516022 445018 516204 445254
rect 515604 444934 516204 445018
rect 515604 444698 515786 444934
rect 516022 444698 516204 444934
rect 515604 409254 516204 444698
rect 515604 409018 515786 409254
rect 516022 409018 516204 409254
rect 515604 408934 516204 409018
rect 515604 408698 515786 408934
rect 516022 408698 516204 408934
rect 515604 373254 516204 408698
rect 515604 373018 515786 373254
rect 516022 373018 516204 373254
rect 515604 372934 516204 373018
rect 515604 372698 515786 372934
rect 516022 372698 516204 372934
rect 515604 337254 516204 372698
rect 515604 337018 515786 337254
rect 516022 337018 516204 337254
rect 515604 336934 516204 337018
rect 515604 336698 515786 336934
rect 516022 336698 516204 336934
rect 515604 301254 516204 336698
rect 515604 301018 515786 301254
rect 516022 301018 516204 301254
rect 515604 300934 516204 301018
rect 515604 300698 515786 300934
rect 516022 300698 516204 300934
rect 515604 265254 516204 300698
rect 515604 265018 515786 265254
rect 516022 265018 516204 265254
rect 515604 264934 516204 265018
rect 515604 264698 515786 264934
rect 516022 264698 516204 264934
rect 515604 229254 516204 264698
rect 515604 229018 515786 229254
rect 516022 229018 516204 229254
rect 515604 228934 516204 229018
rect 515604 228698 515786 228934
rect 516022 228698 516204 228934
rect 515604 193254 516204 228698
rect 515604 193018 515786 193254
rect 516022 193018 516204 193254
rect 515604 192934 516204 193018
rect 515604 192698 515786 192934
rect 516022 192698 516204 192934
rect 515604 157254 516204 192698
rect 515604 157018 515786 157254
rect 516022 157018 516204 157254
rect 515604 156934 516204 157018
rect 515604 156698 515786 156934
rect 516022 156698 516204 156934
rect 515604 121254 516204 156698
rect 515604 121018 515786 121254
rect 516022 121018 516204 121254
rect 515604 120934 516204 121018
rect 515604 120698 515786 120934
rect 516022 120698 516204 120934
rect 515604 85254 516204 120698
rect 515604 85018 515786 85254
rect 516022 85018 516204 85254
rect 515604 84934 516204 85018
rect 515604 84698 515786 84934
rect 516022 84698 516204 84934
rect 515604 49254 516204 84698
rect 515604 49018 515786 49254
rect 516022 49018 516204 49254
rect 515604 48934 516204 49018
rect 515604 48698 515786 48934
rect 516022 48698 516204 48934
rect 515604 13254 516204 48698
rect 515604 13018 515786 13254
rect 516022 13018 516204 13254
rect 515604 12934 516204 13018
rect 515604 12698 515786 12934
rect 516022 12698 516204 12934
rect 497604 -7022 497786 -6786
rect 498022 -7022 498204 -6786
rect 497604 -7106 498204 -7022
rect 497604 -7342 497786 -7106
rect 498022 -7342 498204 -7106
rect 497604 -7364 498204 -7342
rect 515604 -5866 516204 12698
rect 522804 705758 523404 705780
rect 522804 705522 522986 705758
rect 523222 705522 523404 705758
rect 522804 705438 523404 705522
rect 522804 705202 522986 705438
rect 523222 705202 523404 705438
rect 522804 668454 523404 705202
rect 522804 668218 522986 668454
rect 523222 668218 523404 668454
rect 522804 668134 523404 668218
rect 522804 667898 522986 668134
rect 523222 667898 523404 668134
rect 522804 632454 523404 667898
rect 522804 632218 522986 632454
rect 523222 632218 523404 632454
rect 522804 632134 523404 632218
rect 522804 631898 522986 632134
rect 523222 631898 523404 632134
rect 522804 596454 523404 631898
rect 522804 596218 522986 596454
rect 523222 596218 523404 596454
rect 522804 596134 523404 596218
rect 522804 595898 522986 596134
rect 523222 595898 523404 596134
rect 522804 560454 523404 595898
rect 522804 560218 522986 560454
rect 523222 560218 523404 560454
rect 522804 560134 523404 560218
rect 522804 559898 522986 560134
rect 523222 559898 523404 560134
rect 522804 524454 523404 559898
rect 522804 524218 522986 524454
rect 523222 524218 523404 524454
rect 522804 524134 523404 524218
rect 522804 523898 522986 524134
rect 523222 523898 523404 524134
rect 522804 488454 523404 523898
rect 522804 488218 522986 488454
rect 523222 488218 523404 488454
rect 522804 488134 523404 488218
rect 522804 487898 522986 488134
rect 523222 487898 523404 488134
rect 522804 452454 523404 487898
rect 522804 452218 522986 452454
rect 523222 452218 523404 452454
rect 522804 452134 523404 452218
rect 522804 451898 522986 452134
rect 523222 451898 523404 452134
rect 522804 416454 523404 451898
rect 522804 416218 522986 416454
rect 523222 416218 523404 416454
rect 522804 416134 523404 416218
rect 522804 415898 522986 416134
rect 523222 415898 523404 416134
rect 522804 380454 523404 415898
rect 522804 380218 522986 380454
rect 523222 380218 523404 380454
rect 522804 380134 523404 380218
rect 522804 379898 522986 380134
rect 523222 379898 523404 380134
rect 522804 344454 523404 379898
rect 522804 344218 522986 344454
rect 523222 344218 523404 344454
rect 522804 344134 523404 344218
rect 522804 343898 522986 344134
rect 523222 343898 523404 344134
rect 522804 308454 523404 343898
rect 522804 308218 522986 308454
rect 523222 308218 523404 308454
rect 522804 308134 523404 308218
rect 522804 307898 522986 308134
rect 523222 307898 523404 308134
rect 522804 272454 523404 307898
rect 522804 272218 522986 272454
rect 523222 272218 523404 272454
rect 522804 272134 523404 272218
rect 522804 271898 522986 272134
rect 523222 271898 523404 272134
rect 522804 236454 523404 271898
rect 522804 236218 522986 236454
rect 523222 236218 523404 236454
rect 522804 236134 523404 236218
rect 522804 235898 522986 236134
rect 523222 235898 523404 236134
rect 522804 200454 523404 235898
rect 522804 200218 522986 200454
rect 523222 200218 523404 200454
rect 522804 200134 523404 200218
rect 522804 199898 522986 200134
rect 523222 199898 523404 200134
rect 522804 164454 523404 199898
rect 522804 164218 522986 164454
rect 523222 164218 523404 164454
rect 522804 164134 523404 164218
rect 522804 163898 522986 164134
rect 523222 163898 523404 164134
rect 522804 128454 523404 163898
rect 522804 128218 522986 128454
rect 523222 128218 523404 128454
rect 522804 128134 523404 128218
rect 522804 127898 522986 128134
rect 523222 127898 523404 128134
rect 522804 92454 523404 127898
rect 522804 92218 522986 92454
rect 523222 92218 523404 92454
rect 522804 92134 523404 92218
rect 522804 91898 522986 92134
rect 523222 91898 523404 92134
rect 522804 56454 523404 91898
rect 522804 56218 522986 56454
rect 523222 56218 523404 56454
rect 522804 56134 523404 56218
rect 522804 55898 522986 56134
rect 523222 55898 523404 56134
rect 522804 20454 523404 55898
rect 522804 20218 522986 20454
rect 523222 20218 523404 20454
rect 522804 20134 523404 20218
rect 522804 19898 522986 20134
rect 523222 19898 523404 20134
rect 522804 -1266 523404 19898
rect 522804 -1502 522986 -1266
rect 523222 -1502 523404 -1266
rect 522804 -1586 523404 -1502
rect 522804 -1822 522986 -1586
rect 523222 -1822 523404 -1586
rect 522804 -1844 523404 -1822
rect 526404 672054 527004 707042
rect 526404 671818 526586 672054
rect 526822 671818 527004 672054
rect 526404 671734 527004 671818
rect 526404 671498 526586 671734
rect 526822 671498 527004 671734
rect 526404 636054 527004 671498
rect 526404 635818 526586 636054
rect 526822 635818 527004 636054
rect 526404 635734 527004 635818
rect 526404 635498 526586 635734
rect 526822 635498 527004 635734
rect 526404 600054 527004 635498
rect 526404 599818 526586 600054
rect 526822 599818 527004 600054
rect 526404 599734 527004 599818
rect 526404 599498 526586 599734
rect 526822 599498 527004 599734
rect 526404 564054 527004 599498
rect 526404 563818 526586 564054
rect 526822 563818 527004 564054
rect 526404 563734 527004 563818
rect 526404 563498 526586 563734
rect 526822 563498 527004 563734
rect 526404 528054 527004 563498
rect 526404 527818 526586 528054
rect 526822 527818 527004 528054
rect 526404 527734 527004 527818
rect 526404 527498 526586 527734
rect 526822 527498 527004 527734
rect 526404 492054 527004 527498
rect 526404 491818 526586 492054
rect 526822 491818 527004 492054
rect 526404 491734 527004 491818
rect 526404 491498 526586 491734
rect 526822 491498 527004 491734
rect 526404 456054 527004 491498
rect 526404 455818 526586 456054
rect 526822 455818 527004 456054
rect 526404 455734 527004 455818
rect 526404 455498 526586 455734
rect 526822 455498 527004 455734
rect 526404 420054 527004 455498
rect 526404 419818 526586 420054
rect 526822 419818 527004 420054
rect 526404 419734 527004 419818
rect 526404 419498 526586 419734
rect 526822 419498 527004 419734
rect 526404 384054 527004 419498
rect 526404 383818 526586 384054
rect 526822 383818 527004 384054
rect 526404 383734 527004 383818
rect 526404 383498 526586 383734
rect 526822 383498 527004 383734
rect 526404 348054 527004 383498
rect 526404 347818 526586 348054
rect 526822 347818 527004 348054
rect 526404 347734 527004 347818
rect 526404 347498 526586 347734
rect 526822 347498 527004 347734
rect 526404 312054 527004 347498
rect 526404 311818 526586 312054
rect 526822 311818 527004 312054
rect 526404 311734 527004 311818
rect 526404 311498 526586 311734
rect 526822 311498 527004 311734
rect 526404 276054 527004 311498
rect 526404 275818 526586 276054
rect 526822 275818 527004 276054
rect 526404 275734 527004 275818
rect 526404 275498 526586 275734
rect 526822 275498 527004 275734
rect 526404 240054 527004 275498
rect 526404 239818 526586 240054
rect 526822 239818 527004 240054
rect 526404 239734 527004 239818
rect 526404 239498 526586 239734
rect 526822 239498 527004 239734
rect 526404 204054 527004 239498
rect 526404 203818 526586 204054
rect 526822 203818 527004 204054
rect 526404 203734 527004 203818
rect 526404 203498 526586 203734
rect 526822 203498 527004 203734
rect 526404 168054 527004 203498
rect 526404 167818 526586 168054
rect 526822 167818 527004 168054
rect 526404 167734 527004 167818
rect 526404 167498 526586 167734
rect 526822 167498 527004 167734
rect 526404 132054 527004 167498
rect 526404 131818 526586 132054
rect 526822 131818 527004 132054
rect 526404 131734 527004 131818
rect 526404 131498 526586 131734
rect 526822 131498 527004 131734
rect 526404 96054 527004 131498
rect 526404 95818 526586 96054
rect 526822 95818 527004 96054
rect 526404 95734 527004 95818
rect 526404 95498 526586 95734
rect 526822 95498 527004 95734
rect 526404 60054 527004 95498
rect 526404 59818 526586 60054
rect 526822 59818 527004 60054
rect 526404 59734 527004 59818
rect 526404 59498 526586 59734
rect 526822 59498 527004 59734
rect 526404 24054 527004 59498
rect 526404 23818 526586 24054
rect 526822 23818 527004 24054
rect 526404 23734 527004 23818
rect 526404 23498 526586 23734
rect 526822 23498 527004 23734
rect 526404 -3106 527004 23498
rect 526404 -3342 526586 -3106
rect 526822 -3342 527004 -3106
rect 526404 -3426 527004 -3342
rect 526404 -3662 526586 -3426
rect 526822 -3662 527004 -3426
rect 526404 -3684 527004 -3662
rect 530004 675654 530604 708882
rect 530004 675418 530186 675654
rect 530422 675418 530604 675654
rect 530004 675334 530604 675418
rect 530004 675098 530186 675334
rect 530422 675098 530604 675334
rect 530004 639654 530604 675098
rect 530004 639418 530186 639654
rect 530422 639418 530604 639654
rect 530004 639334 530604 639418
rect 530004 639098 530186 639334
rect 530422 639098 530604 639334
rect 530004 603654 530604 639098
rect 530004 603418 530186 603654
rect 530422 603418 530604 603654
rect 530004 603334 530604 603418
rect 530004 603098 530186 603334
rect 530422 603098 530604 603334
rect 530004 567654 530604 603098
rect 530004 567418 530186 567654
rect 530422 567418 530604 567654
rect 530004 567334 530604 567418
rect 530004 567098 530186 567334
rect 530422 567098 530604 567334
rect 530004 531654 530604 567098
rect 530004 531418 530186 531654
rect 530422 531418 530604 531654
rect 530004 531334 530604 531418
rect 530004 531098 530186 531334
rect 530422 531098 530604 531334
rect 530004 495654 530604 531098
rect 530004 495418 530186 495654
rect 530422 495418 530604 495654
rect 530004 495334 530604 495418
rect 530004 495098 530186 495334
rect 530422 495098 530604 495334
rect 530004 459654 530604 495098
rect 530004 459418 530186 459654
rect 530422 459418 530604 459654
rect 530004 459334 530604 459418
rect 530004 459098 530186 459334
rect 530422 459098 530604 459334
rect 530004 423654 530604 459098
rect 530004 423418 530186 423654
rect 530422 423418 530604 423654
rect 530004 423334 530604 423418
rect 530004 423098 530186 423334
rect 530422 423098 530604 423334
rect 530004 387654 530604 423098
rect 530004 387418 530186 387654
rect 530422 387418 530604 387654
rect 530004 387334 530604 387418
rect 530004 387098 530186 387334
rect 530422 387098 530604 387334
rect 530004 351654 530604 387098
rect 530004 351418 530186 351654
rect 530422 351418 530604 351654
rect 530004 351334 530604 351418
rect 530004 351098 530186 351334
rect 530422 351098 530604 351334
rect 530004 315654 530604 351098
rect 530004 315418 530186 315654
rect 530422 315418 530604 315654
rect 530004 315334 530604 315418
rect 530004 315098 530186 315334
rect 530422 315098 530604 315334
rect 530004 279654 530604 315098
rect 530004 279418 530186 279654
rect 530422 279418 530604 279654
rect 530004 279334 530604 279418
rect 530004 279098 530186 279334
rect 530422 279098 530604 279334
rect 530004 243654 530604 279098
rect 530004 243418 530186 243654
rect 530422 243418 530604 243654
rect 530004 243334 530604 243418
rect 530004 243098 530186 243334
rect 530422 243098 530604 243334
rect 530004 207654 530604 243098
rect 530004 207418 530186 207654
rect 530422 207418 530604 207654
rect 530004 207334 530604 207418
rect 530004 207098 530186 207334
rect 530422 207098 530604 207334
rect 530004 171654 530604 207098
rect 530004 171418 530186 171654
rect 530422 171418 530604 171654
rect 530004 171334 530604 171418
rect 530004 171098 530186 171334
rect 530422 171098 530604 171334
rect 530004 135654 530604 171098
rect 530004 135418 530186 135654
rect 530422 135418 530604 135654
rect 530004 135334 530604 135418
rect 530004 135098 530186 135334
rect 530422 135098 530604 135334
rect 530004 99654 530604 135098
rect 530004 99418 530186 99654
rect 530422 99418 530604 99654
rect 530004 99334 530604 99418
rect 530004 99098 530186 99334
rect 530422 99098 530604 99334
rect 530004 63654 530604 99098
rect 530004 63418 530186 63654
rect 530422 63418 530604 63654
rect 530004 63334 530604 63418
rect 530004 63098 530186 63334
rect 530422 63098 530604 63334
rect 530004 27654 530604 63098
rect 530004 27418 530186 27654
rect 530422 27418 530604 27654
rect 530004 27334 530604 27418
rect 530004 27098 530186 27334
rect 530422 27098 530604 27334
rect 530004 -4946 530604 27098
rect 530004 -5182 530186 -4946
rect 530422 -5182 530604 -4946
rect 530004 -5266 530604 -5182
rect 530004 -5502 530186 -5266
rect 530422 -5502 530604 -5266
rect 530004 -5524 530604 -5502
rect 533604 679254 534204 710722
rect 551604 710358 552204 711300
rect 551604 710122 551786 710358
rect 552022 710122 552204 710358
rect 551604 710038 552204 710122
rect 551604 709802 551786 710038
rect 552022 709802 552204 710038
rect 548004 708518 548604 709460
rect 548004 708282 548186 708518
rect 548422 708282 548604 708518
rect 548004 708198 548604 708282
rect 548004 707962 548186 708198
rect 548422 707962 548604 708198
rect 544404 706678 545004 707620
rect 544404 706442 544586 706678
rect 544822 706442 545004 706678
rect 544404 706358 545004 706442
rect 544404 706122 544586 706358
rect 544822 706122 545004 706358
rect 533604 679018 533786 679254
rect 534022 679018 534204 679254
rect 533604 678934 534204 679018
rect 533604 678698 533786 678934
rect 534022 678698 534204 678934
rect 533604 643254 534204 678698
rect 533604 643018 533786 643254
rect 534022 643018 534204 643254
rect 533604 642934 534204 643018
rect 533604 642698 533786 642934
rect 534022 642698 534204 642934
rect 533604 607254 534204 642698
rect 533604 607018 533786 607254
rect 534022 607018 534204 607254
rect 533604 606934 534204 607018
rect 533604 606698 533786 606934
rect 534022 606698 534204 606934
rect 533604 571254 534204 606698
rect 533604 571018 533786 571254
rect 534022 571018 534204 571254
rect 533604 570934 534204 571018
rect 533604 570698 533786 570934
rect 534022 570698 534204 570934
rect 533604 535254 534204 570698
rect 533604 535018 533786 535254
rect 534022 535018 534204 535254
rect 533604 534934 534204 535018
rect 533604 534698 533786 534934
rect 534022 534698 534204 534934
rect 533604 499254 534204 534698
rect 533604 499018 533786 499254
rect 534022 499018 534204 499254
rect 533604 498934 534204 499018
rect 533604 498698 533786 498934
rect 534022 498698 534204 498934
rect 533604 463254 534204 498698
rect 533604 463018 533786 463254
rect 534022 463018 534204 463254
rect 533604 462934 534204 463018
rect 533604 462698 533786 462934
rect 534022 462698 534204 462934
rect 533604 427254 534204 462698
rect 533604 427018 533786 427254
rect 534022 427018 534204 427254
rect 533604 426934 534204 427018
rect 533604 426698 533786 426934
rect 534022 426698 534204 426934
rect 533604 391254 534204 426698
rect 533604 391018 533786 391254
rect 534022 391018 534204 391254
rect 533604 390934 534204 391018
rect 533604 390698 533786 390934
rect 534022 390698 534204 390934
rect 533604 355254 534204 390698
rect 533604 355018 533786 355254
rect 534022 355018 534204 355254
rect 533604 354934 534204 355018
rect 533604 354698 533786 354934
rect 534022 354698 534204 354934
rect 533604 319254 534204 354698
rect 533604 319018 533786 319254
rect 534022 319018 534204 319254
rect 533604 318934 534204 319018
rect 533604 318698 533786 318934
rect 534022 318698 534204 318934
rect 533604 283254 534204 318698
rect 533604 283018 533786 283254
rect 534022 283018 534204 283254
rect 533604 282934 534204 283018
rect 533604 282698 533786 282934
rect 534022 282698 534204 282934
rect 533604 247254 534204 282698
rect 533604 247018 533786 247254
rect 534022 247018 534204 247254
rect 533604 246934 534204 247018
rect 533604 246698 533786 246934
rect 534022 246698 534204 246934
rect 533604 211254 534204 246698
rect 533604 211018 533786 211254
rect 534022 211018 534204 211254
rect 533604 210934 534204 211018
rect 533604 210698 533786 210934
rect 534022 210698 534204 210934
rect 533604 175254 534204 210698
rect 533604 175018 533786 175254
rect 534022 175018 534204 175254
rect 533604 174934 534204 175018
rect 533604 174698 533786 174934
rect 534022 174698 534204 174934
rect 533604 139254 534204 174698
rect 533604 139018 533786 139254
rect 534022 139018 534204 139254
rect 533604 138934 534204 139018
rect 533604 138698 533786 138934
rect 534022 138698 534204 138934
rect 533604 103254 534204 138698
rect 533604 103018 533786 103254
rect 534022 103018 534204 103254
rect 533604 102934 534204 103018
rect 533604 102698 533786 102934
rect 534022 102698 534204 102934
rect 533604 67254 534204 102698
rect 533604 67018 533786 67254
rect 534022 67018 534204 67254
rect 533604 66934 534204 67018
rect 533604 66698 533786 66934
rect 534022 66698 534204 66934
rect 533604 31254 534204 66698
rect 533604 31018 533786 31254
rect 534022 31018 534204 31254
rect 533604 30934 534204 31018
rect 533604 30698 533786 30934
rect 534022 30698 534204 30934
rect 515604 -6102 515786 -5866
rect 516022 -6102 516204 -5866
rect 515604 -6186 516204 -6102
rect 515604 -6422 515786 -6186
rect 516022 -6422 516204 -6186
rect 515604 -7364 516204 -6422
rect 533604 -6786 534204 30698
rect 540804 704838 541404 705780
rect 540804 704602 540986 704838
rect 541222 704602 541404 704838
rect 540804 704518 541404 704602
rect 540804 704282 540986 704518
rect 541222 704282 541404 704518
rect 540804 686454 541404 704282
rect 540804 686218 540986 686454
rect 541222 686218 541404 686454
rect 540804 686134 541404 686218
rect 540804 685898 540986 686134
rect 541222 685898 541404 686134
rect 540804 650454 541404 685898
rect 540804 650218 540986 650454
rect 541222 650218 541404 650454
rect 540804 650134 541404 650218
rect 540804 649898 540986 650134
rect 541222 649898 541404 650134
rect 540804 614454 541404 649898
rect 540804 614218 540986 614454
rect 541222 614218 541404 614454
rect 540804 614134 541404 614218
rect 540804 613898 540986 614134
rect 541222 613898 541404 614134
rect 540804 578454 541404 613898
rect 540804 578218 540986 578454
rect 541222 578218 541404 578454
rect 540804 578134 541404 578218
rect 540804 577898 540986 578134
rect 541222 577898 541404 578134
rect 540804 542454 541404 577898
rect 540804 542218 540986 542454
rect 541222 542218 541404 542454
rect 540804 542134 541404 542218
rect 540804 541898 540986 542134
rect 541222 541898 541404 542134
rect 540804 506454 541404 541898
rect 540804 506218 540986 506454
rect 541222 506218 541404 506454
rect 540804 506134 541404 506218
rect 540804 505898 540986 506134
rect 541222 505898 541404 506134
rect 540804 470454 541404 505898
rect 540804 470218 540986 470454
rect 541222 470218 541404 470454
rect 540804 470134 541404 470218
rect 540804 469898 540986 470134
rect 541222 469898 541404 470134
rect 540804 434454 541404 469898
rect 540804 434218 540986 434454
rect 541222 434218 541404 434454
rect 540804 434134 541404 434218
rect 540804 433898 540986 434134
rect 541222 433898 541404 434134
rect 540804 398454 541404 433898
rect 540804 398218 540986 398454
rect 541222 398218 541404 398454
rect 540804 398134 541404 398218
rect 540804 397898 540986 398134
rect 541222 397898 541404 398134
rect 540804 362454 541404 397898
rect 540804 362218 540986 362454
rect 541222 362218 541404 362454
rect 540804 362134 541404 362218
rect 540804 361898 540986 362134
rect 541222 361898 541404 362134
rect 540804 326454 541404 361898
rect 540804 326218 540986 326454
rect 541222 326218 541404 326454
rect 540804 326134 541404 326218
rect 540804 325898 540986 326134
rect 541222 325898 541404 326134
rect 540804 290454 541404 325898
rect 540804 290218 540986 290454
rect 541222 290218 541404 290454
rect 540804 290134 541404 290218
rect 540804 289898 540986 290134
rect 541222 289898 541404 290134
rect 540804 254454 541404 289898
rect 540804 254218 540986 254454
rect 541222 254218 541404 254454
rect 540804 254134 541404 254218
rect 540804 253898 540986 254134
rect 541222 253898 541404 254134
rect 540804 218454 541404 253898
rect 540804 218218 540986 218454
rect 541222 218218 541404 218454
rect 540804 218134 541404 218218
rect 540804 217898 540986 218134
rect 541222 217898 541404 218134
rect 540804 182454 541404 217898
rect 540804 182218 540986 182454
rect 541222 182218 541404 182454
rect 540804 182134 541404 182218
rect 540804 181898 540986 182134
rect 541222 181898 541404 182134
rect 540804 146454 541404 181898
rect 540804 146218 540986 146454
rect 541222 146218 541404 146454
rect 540804 146134 541404 146218
rect 540804 145898 540986 146134
rect 541222 145898 541404 146134
rect 540804 110454 541404 145898
rect 540804 110218 540986 110454
rect 541222 110218 541404 110454
rect 540804 110134 541404 110218
rect 540804 109898 540986 110134
rect 541222 109898 541404 110134
rect 540804 74454 541404 109898
rect 540804 74218 540986 74454
rect 541222 74218 541404 74454
rect 540804 74134 541404 74218
rect 540804 73898 540986 74134
rect 541222 73898 541404 74134
rect 540804 38454 541404 73898
rect 540804 38218 540986 38454
rect 541222 38218 541404 38454
rect 540804 38134 541404 38218
rect 540804 37898 540986 38134
rect 541222 37898 541404 38134
rect 540804 2454 541404 37898
rect 540804 2218 540986 2454
rect 541222 2218 541404 2454
rect 540804 2134 541404 2218
rect 540804 1898 540986 2134
rect 541222 1898 541404 2134
rect 540804 -346 541404 1898
rect 540804 -582 540986 -346
rect 541222 -582 541404 -346
rect 540804 -666 541404 -582
rect 540804 -902 540986 -666
rect 541222 -902 541404 -666
rect 540804 -1844 541404 -902
rect 544404 690054 545004 706122
rect 544404 689818 544586 690054
rect 544822 689818 545004 690054
rect 544404 689734 545004 689818
rect 544404 689498 544586 689734
rect 544822 689498 545004 689734
rect 544404 654054 545004 689498
rect 544404 653818 544586 654054
rect 544822 653818 545004 654054
rect 544404 653734 545004 653818
rect 544404 653498 544586 653734
rect 544822 653498 545004 653734
rect 544404 618054 545004 653498
rect 544404 617818 544586 618054
rect 544822 617818 545004 618054
rect 544404 617734 545004 617818
rect 544404 617498 544586 617734
rect 544822 617498 545004 617734
rect 544404 582054 545004 617498
rect 544404 581818 544586 582054
rect 544822 581818 545004 582054
rect 544404 581734 545004 581818
rect 544404 581498 544586 581734
rect 544822 581498 545004 581734
rect 544404 546054 545004 581498
rect 544404 545818 544586 546054
rect 544822 545818 545004 546054
rect 544404 545734 545004 545818
rect 544404 545498 544586 545734
rect 544822 545498 545004 545734
rect 544404 510054 545004 545498
rect 544404 509818 544586 510054
rect 544822 509818 545004 510054
rect 544404 509734 545004 509818
rect 544404 509498 544586 509734
rect 544822 509498 545004 509734
rect 544404 474054 545004 509498
rect 544404 473818 544586 474054
rect 544822 473818 545004 474054
rect 544404 473734 545004 473818
rect 544404 473498 544586 473734
rect 544822 473498 545004 473734
rect 544404 438054 545004 473498
rect 544404 437818 544586 438054
rect 544822 437818 545004 438054
rect 544404 437734 545004 437818
rect 544404 437498 544586 437734
rect 544822 437498 545004 437734
rect 544404 402054 545004 437498
rect 544404 401818 544586 402054
rect 544822 401818 545004 402054
rect 544404 401734 545004 401818
rect 544404 401498 544586 401734
rect 544822 401498 545004 401734
rect 544404 366054 545004 401498
rect 544404 365818 544586 366054
rect 544822 365818 545004 366054
rect 544404 365734 545004 365818
rect 544404 365498 544586 365734
rect 544822 365498 545004 365734
rect 544404 330054 545004 365498
rect 544404 329818 544586 330054
rect 544822 329818 545004 330054
rect 544404 329734 545004 329818
rect 544404 329498 544586 329734
rect 544822 329498 545004 329734
rect 544404 294054 545004 329498
rect 544404 293818 544586 294054
rect 544822 293818 545004 294054
rect 544404 293734 545004 293818
rect 544404 293498 544586 293734
rect 544822 293498 545004 293734
rect 544404 258054 545004 293498
rect 544404 257818 544586 258054
rect 544822 257818 545004 258054
rect 544404 257734 545004 257818
rect 544404 257498 544586 257734
rect 544822 257498 545004 257734
rect 544404 222054 545004 257498
rect 544404 221818 544586 222054
rect 544822 221818 545004 222054
rect 544404 221734 545004 221818
rect 544404 221498 544586 221734
rect 544822 221498 545004 221734
rect 544404 186054 545004 221498
rect 544404 185818 544586 186054
rect 544822 185818 545004 186054
rect 544404 185734 545004 185818
rect 544404 185498 544586 185734
rect 544822 185498 545004 185734
rect 544404 150054 545004 185498
rect 544404 149818 544586 150054
rect 544822 149818 545004 150054
rect 544404 149734 545004 149818
rect 544404 149498 544586 149734
rect 544822 149498 545004 149734
rect 544404 114054 545004 149498
rect 544404 113818 544586 114054
rect 544822 113818 545004 114054
rect 544404 113734 545004 113818
rect 544404 113498 544586 113734
rect 544822 113498 545004 113734
rect 544404 78054 545004 113498
rect 544404 77818 544586 78054
rect 544822 77818 545004 78054
rect 544404 77734 545004 77818
rect 544404 77498 544586 77734
rect 544822 77498 545004 77734
rect 544404 42054 545004 77498
rect 544404 41818 544586 42054
rect 544822 41818 545004 42054
rect 544404 41734 545004 41818
rect 544404 41498 544586 41734
rect 544822 41498 545004 41734
rect 544404 6054 545004 41498
rect 544404 5818 544586 6054
rect 544822 5818 545004 6054
rect 544404 5734 545004 5818
rect 544404 5498 544586 5734
rect 544822 5498 545004 5734
rect 544404 -2186 545004 5498
rect 544404 -2422 544586 -2186
rect 544822 -2422 545004 -2186
rect 544404 -2506 545004 -2422
rect 544404 -2742 544586 -2506
rect 544822 -2742 545004 -2506
rect 544404 -3684 545004 -2742
rect 548004 693654 548604 707962
rect 548004 693418 548186 693654
rect 548422 693418 548604 693654
rect 548004 693334 548604 693418
rect 548004 693098 548186 693334
rect 548422 693098 548604 693334
rect 548004 657654 548604 693098
rect 548004 657418 548186 657654
rect 548422 657418 548604 657654
rect 548004 657334 548604 657418
rect 548004 657098 548186 657334
rect 548422 657098 548604 657334
rect 548004 621654 548604 657098
rect 548004 621418 548186 621654
rect 548422 621418 548604 621654
rect 548004 621334 548604 621418
rect 548004 621098 548186 621334
rect 548422 621098 548604 621334
rect 548004 585654 548604 621098
rect 548004 585418 548186 585654
rect 548422 585418 548604 585654
rect 548004 585334 548604 585418
rect 548004 585098 548186 585334
rect 548422 585098 548604 585334
rect 548004 549654 548604 585098
rect 548004 549418 548186 549654
rect 548422 549418 548604 549654
rect 548004 549334 548604 549418
rect 548004 549098 548186 549334
rect 548422 549098 548604 549334
rect 548004 513654 548604 549098
rect 548004 513418 548186 513654
rect 548422 513418 548604 513654
rect 548004 513334 548604 513418
rect 548004 513098 548186 513334
rect 548422 513098 548604 513334
rect 548004 477654 548604 513098
rect 548004 477418 548186 477654
rect 548422 477418 548604 477654
rect 548004 477334 548604 477418
rect 548004 477098 548186 477334
rect 548422 477098 548604 477334
rect 548004 441654 548604 477098
rect 548004 441418 548186 441654
rect 548422 441418 548604 441654
rect 548004 441334 548604 441418
rect 548004 441098 548186 441334
rect 548422 441098 548604 441334
rect 548004 405654 548604 441098
rect 548004 405418 548186 405654
rect 548422 405418 548604 405654
rect 548004 405334 548604 405418
rect 548004 405098 548186 405334
rect 548422 405098 548604 405334
rect 548004 369654 548604 405098
rect 548004 369418 548186 369654
rect 548422 369418 548604 369654
rect 548004 369334 548604 369418
rect 548004 369098 548186 369334
rect 548422 369098 548604 369334
rect 548004 333654 548604 369098
rect 548004 333418 548186 333654
rect 548422 333418 548604 333654
rect 548004 333334 548604 333418
rect 548004 333098 548186 333334
rect 548422 333098 548604 333334
rect 548004 297654 548604 333098
rect 551604 697254 552204 709802
rect 569604 711278 570204 711300
rect 569604 711042 569786 711278
rect 570022 711042 570204 711278
rect 569604 710958 570204 711042
rect 569604 710722 569786 710958
rect 570022 710722 570204 710958
rect 566004 709438 566604 709460
rect 566004 709202 566186 709438
rect 566422 709202 566604 709438
rect 566004 709118 566604 709202
rect 566004 708882 566186 709118
rect 566422 708882 566604 709118
rect 562404 707598 563004 707620
rect 562404 707362 562586 707598
rect 562822 707362 563004 707598
rect 562404 707278 563004 707362
rect 562404 707042 562586 707278
rect 562822 707042 563004 707278
rect 551604 697018 551786 697254
rect 552022 697018 552204 697254
rect 551604 696934 552204 697018
rect 551604 696698 551786 696934
rect 552022 696698 552204 696934
rect 551604 661254 552204 696698
rect 551604 661018 551786 661254
rect 552022 661018 552204 661254
rect 551604 660934 552204 661018
rect 551604 660698 551786 660934
rect 552022 660698 552204 660934
rect 551604 625254 552204 660698
rect 551604 625018 551786 625254
rect 552022 625018 552204 625254
rect 551604 624934 552204 625018
rect 551604 624698 551786 624934
rect 552022 624698 552204 624934
rect 551604 589254 552204 624698
rect 551604 589018 551786 589254
rect 552022 589018 552204 589254
rect 551604 588934 552204 589018
rect 551604 588698 551786 588934
rect 552022 588698 552204 588934
rect 551604 553254 552204 588698
rect 551604 553018 551786 553254
rect 552022 553018 552204 553254
rect 551604 552934 552204 553018
rect 551604 552698 551786 552934
rect 552022 552698 552204 552934
rect 551604 517254 552204 552698
rect 551604 517018 551786 517254
rect 552022 517018 552204 517254
rect 551604 516934 552204 517018
rect 551604 516698 551786 516934
rect 552022 516698 552204 516934
rect 551604 481254 552204 516698
rect 551604 481018 551786 481254
rect 552022 481018 552204 481254
rect 551604 480934 552204 481018
rect 551604 480698 551786 480934
rect 552022 480698 552204 480934
rect 551604 445254 552204 480698
rect 551604 445018 551786 445254
rect 552022 445018 552204 445254
rect 551604 444934 552204 445018
rect 551604 444698 551786 444934
rect 552022 444698 552204 444934
rect 551604 409254 552204 444698
rect 551604 409018 551786 409254
rect 552022 409018 552204 409254
rect 551604 408934 552204 409018
rect 551604 408698 551786 408934
rect 552022 408698 552204 408934
rect 551604 373254 552204 408698
rect 551604 373018 551786 373254
rect 552022 373018 552204 373254
rect 551604 372934 552204 373018
rect 551604 372698 551786 372934
rect 552022 372698 552204 372934
rect 551604 337254 552204 372698
rect 551604 337018 551786 337254
rect 552022 337018 552204 337254
rect 551604 336934 552204 337018
rect 551604 336698 551786 336934
rect 552022 336698 552204 336934
rect 550587 310588 550653 310589
rect 550587 310524 550588 310588
rect 550652 310524 550653 310588
rect 550587 310523 550653 310524
rect 550590 310317 550650 310523
rect 550587 310316 550653 310317
rect 550587 310252 550588 310316
rect 550652 310252 550653 310316
rect 550587 310251 550653 310252
rect 548004 297418 548186 297654
rect 548422 297418 548604 297654
rect 548004 297334 548604 297418
rect 548004 297098 548186 297334
rect 548422 297098 548604 297334
rect 548004 261654 548604 297098
rect 548004 261418 548186 261654
rect 548422 261418 548604 261654
rect 548004 261334 548604 261418
rect 548004 261098 548186 261334
rect 548422 261098 548604 261334
rect 548004 225654 548604 261098
rect 548004 225418 548186 225654
rect 548422 225418 548604 225654
rect 548004 225334 548604 225418
rect 548004 225098 548186 225334
rect 548422 225098 548604 225334
rect 548004 189654 548604 225098
rect 548004 189418 548186 189654
rect 548422 189418 548604 189654
rect 548004 189334 548604 189418
rect 548004 189098 548186 189334
rect 548422 189098 548604 189334
rect 548004 153654 548604 189098
rect 548004 153418 548186 153654
rect 548422 153418 548604 153654
rect 548004 153334 548604 153418
rect 548004 153098 548186 153334
rect 548422 153098 548604 153334
rect 548004 117654 548604 153098
rect 548004 117418 548186 117654
rect 548422 117418 548604 117654
rect 548004 117334 548604 117418
rect 548004 117098 548186 117334
rect 548422 117098 548604 117334
rect 548004 81654 548604 117098
rect 548004 81418 548186 81654
rect 548422 81418 548604 81654
rect 548004 81334 548604 81418
rect 548004 81098 548186 81334
rect 548422 81098 548604 81334
rect 548004 45654 548604 81098
rect 548004 45418 548186 45654
rect 548422 45418 548604 45654
rect 548004 45334 548604 45418
rect 548004 45098 548186 45334
rect 548422 45098 548604 45334
rect 548004 9654 548604 45098
rect 548004 9418 548186 9654
rect 548422 9418 548604 9654
rect 548004 9334 548604 9418
rect 548004 9098 548186 9334
rect 548422 9098 548604 9334
rect 548004 -4026 548604 9098
rect 548004 -4262 548186 -4026
rect 548422 -4262 548604 -4026
rect 548004 -4346 548604 -4262
rect 548004 -4582 548186 -4346
rect 548422 -4582 548604 -4346
rect 548004 -5524 548604 -4582
rect 551604 301254 552204 336698
rect 551604 301018 551786 301254
rect 552022 301018 552204 301254
rect 551604 300934 552204 301018
rect 551604 300698 551786 300934
rect 552022 300698 552204 300934
rect 551604 265254 552204 300698
rect 551604 265018 551786 265254
rect 552022 265018 552204 265254
rect 551604 264934 552204 265018
rect 551604 264698 551786 264934
rect 552022 264698 552204 264934
rect 551604 229254 552204 264698
rect 551604 229018 551786 229254
rect 552022 229018 552204 229254
rect 551604 228934 552204 229018
rect 551604 228698 551786 228934
rect 552022 228698 552204 228934
rect 551604 193254 552204 228698
rect 551604 193018 551786 193254
rect 552022 193018 552204 193254
rect 551604 192934 552204 193018
rect 551604 192698 551786 192934
rect 552022 192698 552204 192934
rect 551604 157254 552204 192698
rect 551604 157018 551786 157254
rect 552022 157018 552204 157254
rect 551604 156934 552204 157018
rect 551604 156698 551786 156934
rect 552022 156698 552204 156934
rect 551604 121254 552204 156698
rect 551604 121018 551786 121254
rect 552022 121018 552204 121254
rect 551604 120934 552204 121018
rect 551604 120698 551786 120934
rect 552022 120698 552204 120934
rect 551604 85254 552204 120698
rect 551604 85018 551786 85254
rect 552022 85018 552204 85254
rect 551604 84934 552204 85018
rect 551604 84698 551786 84934
rect 552022 84698 552204 84934
rect 551604 49254 552204 84698
rect 551604 49018 551786 49254
rect 552022 49018 552204 49254
rect 551604 48934 552204 49018
rect 551604 48698 551786 48934
rect 552022 48698 552204 48934
rect 551604 13254 552204 48698
rect 551604 13018 551786 13254
rect 552022 13018 552204 13254
rect 551604 12934 552204 13018
rect 551604 12698 551786 12934
rect 552022 12698 552204 12934
rect 533604 -7022 533786 -6786
rect 534022 -7022 534204 -6786
rect 533604 -7106 534204 -7022
rect 533604 -7342 533786 -7106
rect 534022 -7342 534204 -7106
rect 533604 -7364 534204 -7342
rect 551604 -5866 552204 12698
rect 558804 705758 559404 705780
rect 558804 705522 558986 705758
rect 559222 705522 559404 705758
rect 558804 705438 559404 705522
rect 558804 705202 558986 705438
rect 559222 705202 559404 705438
rect 558804 668454 559404 705202
rect 558804 668218 558986 668454
rect 559222 668218 559404 668454
rect 558804 668134 559404 668218
rect 558804 667898 558986 668134
rect 559222 667898 559404 668134
rect 558804 632454 559404 667898
rect 558804 632218 558986 632454
rect 559222 632218 559404 632454
rect 558804 632134 559404 632218
rect 558804 631898 558986 632134
rect 559222 631898 559404 632134
rect 558804 596454 559404 631898
rect 558804 596218 558986 596454
rect 559222 596218 559404 596454
rect 558804 596134 559404 596218
rect 558804 595898 558986 596134
rect 559222 595898 559404 596134
rect 558804 560454 559404 595898
rect 558804 560218 558986 560454
rect 559222 560218 559404 560454
rect 558804 560134 559404 560218
rect 558804 559898 558986 560134
rect 559222 559898 559404 560134
rect 558804 524454 559404 559898
rect 558804 524218 558986 524454
rect 559222 524218 559404 524454
rect 558804 524134 559404 524218
rect 558804 523898 558986 524134
rect 559222 523898 559404 524134
rect 558804 488454 559404 523898
rect 558804 488218 558986 488454
rect 559222 488218 559404 488454
rect 558804 488134 559404 488218
rect 558804 487898 558986 488134
rect 559222 487898 559404 488134
rect 558804 452454 559404 487898
rect 558804 452218 558986 452454
rect 559222 452218 559404 452454
rect 558804 452134 559404 452218
rect 558804 451898 558986 452134
rect 559222 451898 559404 452134
rect 558804 416454 559404 451898
rect 558804 416218 558986 416454
rect 559222 416218 559404 416454
rect 558804 416134 559404 416218
rect 558804 415898 558986 416134
rect 559222 415898 559404 416134
rect 558804 380454 559404 415898
rect 558804 380218 558986 380454
rect 559222 380218 559404 380454
rect 558804 380134 559404 380218
rect 558804 379898 558986 380134
rect 559222 379898 559404 380134
rect 558804 344454 559404 379898
rect 558804 344218 558986 344454
rect 559222 344218 559404 344454
rect 558804 344134 559404 344218
rect 558804 343898 558986 344134
rect 559222 343898 559404 344134
rect 558804 308454 559404 343898
rect 562404 672054 563004 707042
rect 562404 671818 562586 672054
rect 562822 671818 563004 672054
rect 562404 671734 563004 671818
rect 562404 671498 562586 671734
rect 562822 671498 563004 671734
rect 562404 636054 563004 671498
rect 562404 635818 562586 636054
rect 562822 635818 563004 636054
rect 562404 635734 563004 635818
rect 562404 635498 562586 635734
rect 562822 635498 563004 635734
rect 562404 600054 563004 635498
rect 562404 599818 562586 600054
rect 562822 599818 563004 600054
rect 562404 599734 563004 599818
rect 562404 599498 562586 599734
rect 562822 599498 563004 599734
rect 562404 564054 563004 599498
rect 562404 563818 562586 564054
rect 562822 563818 563004 564054
rect 562404 563734 563004 563818
rect 562404 563498 562586 563734
rect 562822 563498 563004 563734
rect 562404 528054 563004 563498
rect 562404 527818 562586 528054
rect 562822 527818 563004 528054
rect 562404 527734 563004 527818
rect 562404 527498 562586 527734
rect 562822 527498 563004 527734
rect 562404 492054 563004 527498
rect 562404 491818 562586 492054
rect 562822 491818 563004 492054
rect 562404 491734 563004 491818
rect 562404 491498 562586 491734
rect 562822 491498 563004 491734
rect 562404 456054 563004 491498
rect 562404 455818 562586 456054
rect 562822 455818 563004 456054
rect 562404 455734 563004 455818
rect 562404 455498 562586 455734
rect 562822 455498 563004 455734
rect 562404 420054 563004 455498
rect 562404 419818 562586 420054
rect 562822 419818 563004 420054
rect 562404 419734 563004 419818
rect 562404 419498 562586 419734
rect 562822 419498 563004 419734
rect 562404 384054 563004 419498
rect 562404 383818 562586 384054
rect 562822 383818 563004 384054
rect 562404 383734 563004 383818
rect 562404 383498 562586 383734
rect 562822 383498 563004 383734
rect 562404 348054 563004 383498
rect 562404 347818 562586 348054
rect 562822 347818 563004 348054
rect 562404 347734 563004 347818
rect 562404 347498 562586 347734
rect 562822 347498 563004 347734
rect 562404 312054 563004 347498
rect 562404 311818 562586 312054
rect 562822 311818 563004 312054
rect 562404 311734 563004 311818
rect 562404 311498 562586 311734
rect 562822 311498 563004 311734
rect 560342 311070 560586 311130
rect 560342 310861 560402 311070
rect 560339 310860 560405 310861
rect 560339 310796 560340 310860
rect 560404 310796 560405 310860
rect 560339 310795 560405 310796
rect 560526 310725 560586 311070
rect 560523 310724 560589 310725
rect 560523 310660 560524 310724
rect 560588 310660 560589 310724
rect 560523 310659 560589 310660
rect 558804 308218 558986 308454
rect 559222 308218 559404 308454
rect 558804 308134 559404 308218
rect 558804 307898 558986 308134
rect 559222 307898 559404 308134
rect 558804 272454 559404 307898
rect 558804 272218 558986 272454
rect 559222 272218 559404 272454
rect 558804 272134 559404 272218
rect 558804 271898 558986 272134
rect 559222 271898 559404 272134
rect 558804 236454 559404 271898
rect 558804 236218 558986 236454
rect 559222 236218 559404 236454
rect 558804 236134 559404 236218
rect 558804 235898 558986 236134
rect 559222 235898 559404 236134
rect 558804 200454 559404 235898
rect 558804 200218 558986 200454
rect 559222 200218 559404 200454
rect 558804 200134 559404 200218
rect 558804 199898 558986 200134
rect 559222 199898 559404 200134
rect 558804 164454 559404 199898
rect 558804 164218 558986 164454
rect 559222 164218 559404 164454
rect 558804 164134 559404 164218
rect 558804 163898 558986 164134
rect 559222 163898 559404 164134
rect 558804 128454 559404 163898
rect 558804 128218 558986 128454
rect 559222 128218 559404 128454
rect 558804 128134 559404 128218
rect 558804 127898 558986 128134
rect 559222 127898 559404 128134
rect 558804 92454 559404 127898
rect 558804 92218 558986 92454
rect 559222 92218 559404 92454
rect 558804 92134 559404 92218
rect 558804 91898 558986 92134
rect 559222 91898 559404 92134
rect 558804 56454 559404 91898
rect 558804 56218 558986 56454
rect 559222 56218 559404 56454
rect 558804 56134 559404 56218
rect 558804 55898 558986 56134
rect 559222 55898 559404 56134
rect 558804 20454 559404 55898
rect 558804 20218 558986 20454
rect 559222 20218 559404 20454
rect 558804 20134 559404 20218
rect 558804 19898 558986 20134
rect 559222 19898 559404 20134
rect 558804 -1266 559404 19898
rect 558804 -1502 558986 -1266
rect 559222 -1502 559404 -1266
rect 558804 -1586 559404 -1502
rect 558804 -1822 558986 -1586
rect 559222 -1822 559404 -1586
rect 558804 -1844 559404 -1822
rect 562404 276054 563004 311498
rect 562404 275818 562586 276054
rect 562822 275818 563004 276054
rect 562404 275734 563004 275818
rect 562404 275498 562586 275734
rect 562822 275498 563004 275734
rect 562404 240054 563004 275498
rect 562404 239818 562586 240054
rect 562822 239818 563004 240054
rect 562404 239734 563004 239818
rect 562404 239498 562586 239734
rect 562822 239498 563004 239734
rect 562404 204054 563004 239498
rect 562404 203818 562586 204054
rect 562822 203818 563004 204054
rect 562404 203734 563004 203818
rect 562404 203498 562586 203734
rect 562822 203498 563004 203734
rect 562404 168054 563004 203498
rect 562404 167818 562586 168054
rect 562822 167818 563004 168054
rect 562404 167734 563004 167818
rect 562404 167498 562586 167734
rect 562822 167498 563004 167734
rect 562404 132054 563004 167498
rect 562404 131818 562586 132054
rect 562822 131818 563004 132054
rect 562404 131734 563004 131818
rect 562404 131498 562586 131734
rect 562822 131498 563004 131734
rect 562404 96054 563004 131498
rect 562404 95818 562586 96054
rect 562822 95818 563004 96054
rect 562404 95734 563004 95818
rect 562404 95498 562586 95734
rect 562822 95498 563004 95734
rect 562404 60054 563004 95498
rect 562404 59818 562586 60054
rect 562822 59818 563004 60054
rect 562404 59734 563004 59818
rect 562404 59498 562586 59734
rect 562822 59498 563004 59734
rect 562404 24054 563004 59498
rect 562404 23818 562586 24054
rect 562822 23818 563004 24054
rect 562404 23734 563004 23818
rect 562404 23498 562586 23734
rect 562822 23498 563004 23734
rect 562404 -3106 563004 23498
rect 562404 -3342 562586 -3106
rect 562822 -3342 563004 -3106
rect 562404 -3426 563004 -3342
rect 562404 -3662 562586 -3426
rect 562822 -3662 563004 -3426
rect 562404 -3684 563004 -3662
rect 566004 675654 566604 708882
rect 566004 675418 566186 675654
rect 566422 675418 566604 675654
rect 566004 675334 566604 675418
rect 566004 675098 566186 675334
rect 566422 675098 566604 675334
rect 566004 639654 566604 675098
rect 566004 639418 566186 639654
rect 566422 639418 566604 639654
rect 566004 639334 566604 639418
rect 566004 639098 566186 639334
rect 566422 639098 566604 639334
rect 566004 603654 566604 639098
rect 566004 603418 566186 603654
rect 566422 603418 566604 603654
rect 566004 603334 566604 603418
rect 566004 603098 566186 603334
rect 566422 603098 566604 603334
rect 566004 567654 566604 603098
rect 566004 567418 566186 567654
rect 566422 567418 566604 567654
rect 566004 567334 566604 567418
rect 566004 567098 566186 567334
rect 566422 567098 566604 567334
rect 566004 531654 566604 567098
rect 566004 531418 566186 531654
rect 566422 531418 566604 531654
rect 566004 531334 566604 531418
rect 566004 531098 566186 531334
rect 566422 531098 566604 531334
rect 566004 495654 566604 531098
rect 566004 495418 566186 495654
rect 566422 495418 566604 495654
rect 566004 495334 566604 495418
rect 566004 495098 566186 495334
rect 566422 495098 566604 495334
rect 566004 459654 566604 495098
rect 566004 459418 566186 459654
rect 566422 459418 566604 459654
rect 566004 459334 566604 459418
rect 566004 459098 566186 459334
rect 566422 459098 566604 459334
rect 566004 423654 566604 459098
rect 566004 423418 566186 423654
rect 566422 423418 566604 423654
rect 566004 423334 566604 423418
rect 566004 423098 566186 423334
rect 566422 423098 566604 423334
rect 566004 387654 566604 423098
rect 566004 387418 566186 387654
rect 566422 387418 566604 387654
rect 566004 387334 566604 387418
rect 566004 387098 566186 387334
rect 566422 387098 566604 387334
rect 566004 351654 566604 387098
rect 566004 351418 566186 351654
rect 566422 351418 566604 351654
rect 566004 351334 566604 351418
rect 566004 351098 566186 351334
rect 566422 351098 566604 351334
rect 566004 315654 566604 351098
rect 566004 315418 566186 315654
rect 566422 315418 566604 315654
rect 566004 315334 566604 315418
rect 566004 315098 566186 315334
rect 566422 315098 566604 315334
rect 566004 279654 566604 315098
rect 566004 279418 566186 279654
rect 566422 279418 566604 279654
rect 566004 279334 566604 279418
rect 566004 279098 566186 279334
rect 566422 279098 566604 279334
rect 566004 243654 566604 279098
rect 566004 243418 566186 243654
rect 566422 243418 566604 243654
rect 566004 243334 566604 243418
rect 566004 243098 566186 243334
rect 566422 243098 566604 243334
rect 566004 207654 566604 243098
rect 566004 207418 566186 207654
rect 566422 207418 566604 207654
rect 566004 207334 566604 207418
rect 566004 207098 566186 207334
rect 566422 207098 566604 207334
rect 566004 171654 566604 207098
rect 566004 171418 566186 171654
rect 566422 171418 566604 171654
rect 566004 171334 566604 171418
rect 566004 171098 566186 171334
rect 566422 171098 566604 171334
rect 566004 135654 566604 171098
rect 566004 135418 566186 135654
rect 566422 135418 566604 135654
rect 566004 135334 566604 135418
rect 566004 135098 566186 135334
rect 566422 135098 566604 135334
rect 566004 99654 566604 135098
rect 566004 99418 566186 99654
rect 566422 99418 566604 99654
rect 566004 99334 566604 99418
rect 566004 99098 566186 99334
rect 566422 99098 566604 99334
rect 566004 63654 566604 99098
rect 566004 63418 566186 63654
rect 566422 63418 566604 63654
rect 566004 63334 566604 63418
rect 566004 63098 566186 63334
rect 566422 63098 566604 63334
rect 566004 27654 566604 63098
rect 566004 27418 566186 27654
rect 566422 27418 566604 27654
rect 566004 27334 566604 27418
rect 566004 27098 566186 27334
rect 566422 27098 566604 27334
rect 566004 -4946 566604 27098
rect 566004 -5182 566186 -4946
rect 566422 -5182 566604 -4946
rect 566004 -5266 566604 -5182
rect 566004 -5502 566186 -5266
rect 566422 -5502 566604 -5266
rect 566004 -5524 566604 -5502
rect 569604 679254 570204 710722
rect 591760 711278 592360 711300
rect 591760 711042 591942 711278
rect 592178 711042 592360 711278
rect 591760 710958 592360 711042
rect 591760 710722 591942 710958
rect 592178 710722 592360 710958
rect 590840 710358 591440 710380
rect 590840 710122 591022 710358
rect 591258 710122 591440 710358
rect 590840 710038 591440 710122
rect 590840 709802 591022 710038
rect 591258 709802 591440 710038
rect 589920 709438 590520 709460
rect 589920 709202 590102 709438
rect 590338 709202 590520 709438
rect 589920 709118 590520 709202
rect 589920 708882 590102 709118
rect 590338 708882 590520 709118
rect 589000 708518 589600 708540
rect 589000 708282 589182 708518
rect 589418 708282 589600 708518
rect 589000 708198 589600 708282
rect 589000 707962 589182 708198
rect 589418 707962 589600 708198
rect 580404 706678 581004 707620
rect 588080 707598 588680 707620
rect 588080 707362 588262 707598
rect 588498 707362 588680 707598
rect 588080 707278 588680 707362
rect 588080 707042 588262 707278
rect 588498 707042 588680 707278
rect 580404 706442 580586 706678
rect 580822 706442 581004 706678
rect 580404 706358 581004 706442
rect 580404 706122 580586 706358
rect 580822 706122 581004 706358
rect 569604 679018 569786 679254
rect 570022 679018 570204 679254
rect 569604 678934 570204 679018
rect 569604 678698 569786 678934
rect 570022 678698 570204 678934
rect 569604 643254 570204 678698
rect 569604 643018 569786 643254
rect 570022 643018 570204 643254
rect 569604 642934 570204 643018
rect 569604 642698 569786 642934
rect 570022 642698 570204 642934
rect 569604 607254 570204 642698
rect 569604 607018 569786 607254
rect 570022 607018 570204 607254
rect 569604 606934 570204 607018
rect 569604 606698 569786 606934
rect 570022 606698 570204 606934
rect 569604 571254 570204 606698
rect 569604 571018 569786 571254
rect 570022 571018 570204 571254
rect 569604 570934 570204 571018
rect 569604 570698 569786 570934
rect 570022 570698 570204 570934
rect 569604 535254 570204 570698
rect 569604 535018 569786 535254
rect 570022 535018 570204 535254
rect 569604 534934 570204 535018
rect 569604 534698 569786 534934
rect 570022 534698 570204 534934
rect 569604 499254 570204 534698
rect 569604 499018 569786 499254
rect 570022 499018 570204 499254
rect 569604 498934 570204 499018
rect 569604 498698 569786 498934
rect 570022 498698 570204 498934
rect 569604 463254 570204 498698
rect 569604 463018 569786 463254
rect 570022 463018 570204 463254
rect 569604 462934 570204 463018
rect 569604 462698 569786 462934
rect 570022 462698 570204 462934
rect 569604 427254 570204 462698
rect 569604 427018 569786 427254
rect 570022 427018 570204 427254
rect 569604 426934 570204 427018
rect 569604 426698 569786 426934
rect 570022 426698 570204 426934
rect 569604 391254 570204 426698
rect 569604 391018 569786 391254
rect 570022 391018 570204 391254
rect 569604 390934 570204 391018
rect 569604 390698 569786 390934
rect 570022 390698 570204 390934
rect 569604 355254 570204 390698
rect 569604 355018 569786 355254
rect 570022 355018 570204 355254
rect 569604 354934 570204 355018
rect 569604 354698 569786 354934
rect 570022 354698 570204 354934
rect 569604 319254 570204 354698
rect 569604 319018 569786 319254
rect 570022 319018 570204 319254
rect 569604 318934 570204 319018
rect 569604 318698 569786 318934
rect 570022 318698 570204 318934
rect 569604 283254 570204 318698
rect 569604 283018 569786 283254
rect 570022 283018 570204 283254
rect 569604 282934 570204 283018
rect 569604 282698 569786 282934
rect 570022 282698 570204 282934
rect 569604 247254 570204 282698
rect 569604 247018 569786 247254
rect 570022 247018 570204 247254
rect 569604 246934 570204 247018
rect 569604 246698 569786 246934
rect 570022 246698 570204 246934
rect 569604 211254 570204 246698
rect 569604 211018 569786 211254
rect 570022 211018 570204 211254
rect 569604 210934 570204 211018
rect 569604 210698 569786 210934
rect 570022 210698 570204 210934
rect 569604 175254 570204 210698
rect 569604 175018 569786 175254
rect 570022 175018 570204 175254
rect 569604 174934 570204 175018
rect 569604 174698 569786 174934
rect 570022 174698 570204 174934
rect 569604 139254 570204 174698
rect 569604 139018 569786 139254
rect 570022 139018 570204 139254
rect 569604 138934 570204 139018
rect 569604 138698 569786 138934
rect 570022 138698 570204 138934
rect 569604 103254 570204 138698
rect 569604 103018 569786 103254
rect 570022 103018 570204 103254
rect 569604 102934 570204 103018
rect 569604 102698 569786 102934
rect 570022 102698 570204 102934
rect 569604 67254 570204 102698
rect 569604 67018 569786 67254
rect 570022 67018 570204 67254
rect 569604 66934 570204 67018
rect 569604 66698 569786 66934
rect 570022 66698 570204 66934
rect 569604 31254 570204 66698
rect 569604 31018 569786 31254
rect 570022 31018 570204 31254
rect 569604 30934 570204 31018
rect 569604 30698 569786 30934
rect 570022 30698 570204 30934
rect 551604 -6102 551786 -5866
rect 552022 -6102 552204 -5866
rect 551604 -6186 552204 -6102
rect 551604 -6422 551786 -6186
rect 552022 -6422 552204 -6186
rect 551604 -7364 552204 -6422
rect 569604 -6786 570204 30698
rect 576804 704838 577404 705780
rect 576804 704602 576986 704838
rect 577222 704602 577404 704838
rect 576804 704518 577404 704602
rect 576804 704282 576986 704518
rect 577222 704282 577404 704518
rect 576804 686454 577404 704282
rect 576804 686218 576986 686454
rect 577222 686218 577404 686454
rect 576804 686134 577404 686218
rect 576804 685898 576986 686134
rect 577222 685898 577404 686134
rect 576804 650454 577404 685898
rect 576804 650218 576986 650454
rect 577222 650218 577404 650454
rect 576804 650134 577404 650218
rect 576804 649898 576986 650134
rect 577222 649898 577404 650134
rect 576804 614454 577404 649898
rect 576804 614218 576986 614454
rect 577222 614218 577404 614454
rect 576804 614134 577404 614218
rect 576804 613898 576986 614134
rect 577222 613898 577404 614134
rect 576804 578454 577404 613898
rect 576804 578218 576986 578454
rect 577222 578218 577404 578454
rect 576804 578134 577404 578218
rect 576804 577898 576986 578134
rect 577222 577898 577404 578134
rect 576804 542454 577404 577898
rect 576804 542218 576986 542454
rect 577222 542218 577404 542454
rect 576804 542134 577404 542218
rect 576804 541898 576986 542134
rect 577222 541898 577404 542134
rect 576804 506454 577404 541898
rect 576804 506218 576986 506454
rect 577222 506218 577404 506454
rect 576804 506134 577404 506218
rect 576804 505898 576986 506134
rect 577222 505898 577404 506134
rect 576804 470454 577404 505898
rect 576804 470218 576986 470454
rect 577222 470218 577404 470454
rect 576804 470134 577404 470218
rect 576804 469898 576986 470134
rect 577222 469898 577404 470134
rect 576804 434454 577404 469898
rect 576804 434218 576986 434454
rect 577222 434218 577404 434454
rect 576804 434134 577404 434218
rect 576804 433898 576986 434134
rect 577222 433898 577404 434134
rect 576804 398454 577404 433898
rect 576804 398218 576986 398454
rect 577222 398218 577404 398454
rect 576804 398134 577404 398218
rect 576804 397898 576986 398134
rect 577222 397898 577404 398134
rect 576804 362454 577404 397898
rect 576804 362218 576986 362454
rect 577222 362218 577404 362454
rect 576804 362134 577404 362218
rect 576804 361898 576986 362134
rect 577222 361898 577404 362134
rect 576804 326454 577404 361898
rect 576804 326218 576986 326454
rect 577222 326218 577404 326454
rect 576804 326134 577404 326218
rect 576804 325898 576986 326134
rect 577222 325898 577404 326134
rect 576804 290454 577404 325898
rect 576804 290218 576986 290454
rect 577222 290218 577404 290454
rect 576804 290134 577404 290218
rect 576804 289898 576986 290134
rect 577222 289898 577404 290134
rect 576804 254454 577404 289898
rect 576804 254218 576986 254454
rect 577222 254218 577404 254454
rect 576804 254134 577404 254218
rect 576804 253898 576986 254134
rect 577222 253898 577404 254134
rect 576804 218454 577404 253898
rect 576804 218218 576986 218454
rect 577222 218218 577404 218454
rect 576804 218134 577404 218218
rect 576804 217898 576986 218134
rect 577222 217898 577404 218134
rect 576804 182454 577404 217898
rect 576804 182218 576986 182454
rect 577222 182218 577404 182454
rect 576804 182134 577404 182218
rect 576804 181898 576986 182134
rect 577222 181898 577404 182134
rect 576804 146454 577404 181898
rect 576804 146218 576986 146454
rect 577222 146218 577404 146454
rect 576804 146134 577404 146218
rect 576804 145898 576986 146134
rect 577222 145898 577404 146134
rect 576804 110454 577404 145898
rect 576804 110218 576986 110454
rect 577222 110218 577404 110454
rect 576804 110134 577404 110218
rect 576804 109898 576986 110134
rect 577222 109898 577404 110134
rect 576804 74454 577404 109898
rect 576804 74218 576986 74454
rect 577222 74218 577404 74454
rect 576804 74134 577404 74218
rect 576804 73898 576986 74134
rect 577222 73898 577404 74134
rect 576804 38454 577404 73898
rect 576804 38218 576986 38454
rect 577222 38218 577404 38454
rect 576804 38134 577404 38218
rect 576804 37898 576986 38134
rect 577222 37898 577404 38134
rect 576804 2454 577404 37898
rect 576804 2218 576986 2454
rect 577222 2218 577404 2454
rect 576804 2134 577404 2218
rect 576804 1898 576986 2134
rect 577222 1898 577404 2134
rect 576804 -346 577404 1898
rect 576804 -582 576986 -346
rect 577222 -582 577404 -346
rect 576804 -666 577404 -582
rect 576804 -902 576986 -666
rect 577222 -902 577404 -666
rect 576804 -1844 577404 -902
rect 580404 690054 581004 706122
rect 587160 706678 587760 706700
rect 587160 706442 587342 706678
rect 587578 706442 587760 706678
rect 587160 706358 587760 706442
rect 587160 706122 587342 706358
rect 587578 706122 587760 706358
rect 586240 705758 586840 705780
rect 586240 705522 586422 705758
rect 586658 705522 586840 705758
rect 586240 705438 586840 705522
rect 586240 705202 586422 705438
rect 586658 705202 586840 705438
rect 580404 689818 580586 690054
rect 580822 689818 581004 690054
rect 580404 689734 581004 689818
rect 580404 689498 580586 689734
rect 580822 689498 581004 689734
rect 580404 654054 581004 689498
rect 580404 653818 580586 654054
rect 580822 653818 581004 654054
rect 580404 653734 581004 653818
rect 580404 653498 580586 653734
rect 580822 653498 581004 653734
rect 580404 618054 581004 653498
rect 580404 617818 580586 618054
rect 580822 617818 581004 618054
rect 580404 617734 581004 617818
rect 580404 617498 580586 617734
rect 580822 617498 581004 617734
rect 580404 582054 581004 617498
rect 580404 581818 580586 582054
rect 580822 581818 581004 582054
rect 580404 581734 581004 581818
rect 580404 581498 580586 581734
rect 580822 581498 581004 581734
rect 580404 546054 581004 581498
rect 580404 545818 580586 546054
rect 580822 545818 581004 546054
rect 580404 545734 581004 545818
rect 580404 545498 580586 545734
rect 580822 545498 581004 545734
rect 580404 510054 581004 545498
rect 580404 509818 580586 510054
rect 580822 509818 581004 510054
rect 580404 509734 581004 509818
rect 580404 509498 580586 509734
rect 580822 509498 581004 509734
rect 580404 474054 581004 509498
rect 580404 473818 580586 474054
rect 580822 473818 581004 474054
rect 580404 473734 581004 473818
rect 580404 473498 580586 473734
rect 580822 473498 581004 473734
rect 580404 438054 581004 473498
rect 580404 437818 580586 438054
rect 580822 437818 581004 438054
rect 580404 437734 581004 437818
rect 580404 437498 580586 437734
rect 580822 437498 581004 437734
rect 580404 402054 581004 437498
rect 580404 401818 580586 402054
rect 580822 401818 581004 402054
rect 580404 401734 581004 401818
rect 580404 401498 580586 401734
rect 580822 401498 581004 401734
rect 580404 366054 581004 401498
rect 580404 365818 580586 366054
rect 580822 365818 581004 366054
rect 580404 365734 581004 365818
rect 580404 365498 580586 365734
rect 580822 365498 581004 365734
rect 580404 330054 581004 365498
rect 580404 329818 580586 330054
rect 580822 329818 581004 330054
rect 580404 329734 581004 329818
rect 580404 329498 580586 329734
rect 580822 329498 581004 329734
rect 580404 294054 581004 329498
rect 580404 293818 580586 294054
rect 580822 293818 581004 294054
rect 580404 293734 581004 293818
rect 580404 293498 580586 293734
rect 580822 293498 581004 293734
rect 580404 258054 581004 293498
rect 580404 257818 580586 258054
rect 580822 257818 581004 258054
rect 580404 257734 581004 257818
rect 580404 257498 580586 257734
rect 580822 257498 581004 257734
rect 580404 222054 581004 257498
rect 580404 221818 580586 222054
rect 580822 221818 581004 222054
rect 580404 221734 581004 221818
rect 580404 221498 580586 221734
rect 580822 221498 581004 221734
rect 580404 186054 581004 221498
rect 580404 185818 580586 186054
rect 580822 185818 581004 186054
rect 580404 185734 581004 185818
rect 580404 185498 580586 185734
rect 580822 185498 581004 185734
rect 580404 150054 581004 185498
rect 580404 149818 580586 150054
rect 580822 149818 581004 150054
rect 580404 149734 581004 149818
rect 580404 149498 580586 149734
rect 580822 149498 581004 149734
rect 580404 114054 581004 149498
rect 580404 113818 580586 114054
rect 580822 113818 581004 114054
rect 580404 113734 581004 113818
rect 580404 113498 580586 113734
rect 580822 113498 581004 113734
rect 580404 78054 581004 113498
rect 580404 77818 580586 78054
rect 580822 77818 581004 78054
rect 580404 77734 581004 77818
rect 580404 77498 580586 77734
rect 580822 77498 581004 77734
rect 580404 42054 581004 77498
rect 580404 41818 580586 42054
rect 580822 41818 581004 42054
rect 580404 41734 581004 41818
rect 580404 41498 580586 41734
rect 580822 41498 581004 41734
rect 580404 6054 581004 41498
rect 580404 5818 580586 6054
rect 580822 5818 581004 6054
rect 580404 5734 581004 5818
rect 580404 5498 580586 5734
rect 580822 5498 581004 5734
rect 580404 -2186 581004 5498
rect 585320 704838 585920 704860
rect 585320 704602 585502 704838
rect 585738 704602 585920 704838
rect 585320 704518 585920 704602
rect 585320 704282 585502 704518
rect 585738 704282 585920 704518
rect 585320 686454 585920 704282
rect 585320 686218 585502 686454
rect 585738 686218 585920 686454
rect 585320 686134 585920 686218
rect 585320 685898 585502 686134
rect 585738 685898 585920 686134
rect 585320 650454 585920 685898
rect 585320 650218 585502 650454
rect 585738 650218 585920 650454
rect 585320 650134 585920 650218
rect 585320 649898 585502 650134
rect 585738 649898 585920 650134
rect 585320 614454 585920 649898
rect 585320 614218 585502 614454
rect 585738 614218 585920 614454
rect 585320 614134 585920 614218
rect 585320 613898 585502 614134
rect 585738 613898 585920 614134
rect 585320 578454 585920 613898
rect 585320 578218 585502 578454
rect 585738 578218 585920 578454
rect 585320 578134 585920 578218
rect 585320 577898 585502 578134
rect 585738 577898 585920 578134
rect 585320 542454 585920 577898
rect 585320 542218 585502 542454
rect 585738 542218 585920 542454
rect 585320 542134 585920 542218
rect 585320 541898 585502 542134
rect 585738 541898 585920 542134
rect 585320 506454 585920 541898
rect 585320 506218 585502 506454
rect 585738 506218 585920 506454
rect 585320 506134 585920 506218
rect 585320 505898 585502 506134
rect 585738 505898 585920 506134
rect 585320 470454 585920 505898
rect 585320 470218 585502 470454
rect 585738 470218 585920 470454
rect 585320 470134 585920 470218
rect 585320 469898 585502 470134
rect 585738 469898 585920 470134
rect 585320 434454 585920 469898
rect 585320 434218 585502 434454
rect 585738 434218 585920 434454
rect 585320 434134 585920 434218
rect 585320 433898 585502 434134
rect 585738 433898 585920 434134
rect 585320 398454 585920 433898
rect 585320 398218 585502 398454
rect 585738 398218 585920 398454
rect 585320 398134 585920 398218
rect 585320 397898 585502 398134
rect 585738 397898 585920 398134
rect 585320 362454 585920 397898
rect 585320 362218 585502 362454
rect 585738 362218 585920 362454
rect 585320 362134 585920 362218
rect 585320 361898 585502 362134
rect 585738 361898 585920 362134
rect 585320 326454 585920 361898
rect 585320 326218 585502 326454
rect 585738 326218 585920 326454
rect 585320 326134 585920 326218
rect 585320 325898 585502 326134
rect 585738 325898 585920 326134
rect 585320 290454 585920 325898
rect 585320 290218 585502 290454
rect 585738 290218 585920 290454
rect 585320 290134 585920 290218
rect 585320 289898 585502 290134
rect 585738 289898 585920 290134
rect 585320 254454 585920 289898
rect 585320 254218 585502 254454
rect 585738 254218 585920 254454
rect 585320 254134 585920 254218
rect 585320 253898 585502 254134
rect 585738 253898 585920 254134
rect 585320 218454 585920 253898
rect 585320 218218 585502 218454
rect 585738 218218 585920 218454
rect 585320 218134 585920 218218
rect 585320 217898 585502 218134
rect 585738 217898 585920 218134
rect 585320 182454 585920 217898
rect 585320 182218 585502 182454
rect 585738 182218 585920 182454
rect 585320 182134 585920 182218
rect 585320 181898 585502 182134
rect 585738 181898 585920 182134
rect 585320 146454 585920 181898
rect 585320 146218 585502 146454
rect 585738 146218 585920 146454
rect 585320 146134 585920 146218
rect 585320 145898 585502 146134
rect 585738 145898 585920 146134
rect 585320 110454 585920 145898
rect 585320 110218 585502 110454
rect 585738 110218 585920 110454
rect 585320 110134 585920 110218
rect 585320 109898 585502 110134
rect 585738 109898 585920 110134
rect 585320 74454 585920 109898
rect 585320 74218 585502 74454
rect 585738 74218 585920 74454
rect 585320 74134 585920 74218
rect 585320 73898 585502 74134
rect 585738 73898 585920 74134
rect 585320 38454 585920 73898
rect 585320 38218 585502 38454
rect 585738 38218 585920 38454
rect 585320 38134 585920 38218
rect 585320 37898 585502 38134
rect 585738 37898 585920 38134
rect 585320 2454 585920 37898
rect 585320 2218 585502 2454
rect 585738 2218 585920 2454
rect 585320 2134 585920 2218
rect 585320 1898 585502 2134
rect 585738 1898 585920 2134
rect 585320 -346 585920 1898
rect 585320 -582 585502 -346
rect 585738 -582 585920 -346
rect 585320 -666 585920 -582
rect 585320 -902 585502 -666
rect 585738 -902 585920 -666
rect 585320 -924 585920 -902
rect 586240 668454 586840 705202
rect 586240 668218 586422 668454
rect 586658 668218 586840 668454
rect 586240 668134 586840 668218
rect 586240 667898 586422 668134
rect 586658 667898 586840 668134
rect 586240 632454 586840 667898
rect 586240 632218 586422 632454
rect 586658 632218 586840 632454
rect 586240 632134 586840 632218
rect 586240 631898 586422 632134
rect 586658 631898 586840 632134
rect 586240 596454 586840 631898
rect 586240 596218 586422 596454
rect 586658 596218 586840 596454
rect 586240 596134 586840 596218
rect 586240 595898 586422 596134
rect 586658 595898 586840 596134
rect 586240 560454 586840 595898
rect 586240 560218 586422 560454
rect 586658 560218 586840 560454
rect 586240 560134 586840 560218
rect 586240 559898 586422 560134
rect 586658 559898 586840 560134
rect 586240 524454 586840 559898
rect 586240 524218 586422 524454
rect 586658 524218 586840 524454
rect 586240 524134 586840 524218
rect 586240 523898 586422 524134
rect 586658 523898 586840 524134
rect 586240 488454 586840 523898
rect 586240 488218 586422 488454
rect 586658 488218 586840 488454
rect 586240 488134 586840 488218
rect 586240 487898 586422 488134
rect 586658 487898 586840 488134
rect 586240 452454 586840 487898
rect 586240 452218 586422 452454
rect 586658 452218 586840 452454
rect 586240 452134 586840 452218
rect 586240 451898 586422 452134
rect 586658 451898 586840 452134
rect 586240 416454 586840 451898
rect 586240 416218 586422 416454
rect 586658 416218 586840 416454
rect 586240 416134 586840 416218
rect 586240 415898 586422 416134
rect 586658 415898 586840 416134
rect 586240 380454 586840 415898
rect 586240 380218 586422 380454
rect 586658 380218 586840 380454
rect 586240 380134 586840 380218
rect 586240 379898 586422 380134
rect 586658 379898 586840 380134
rect 586240 344454 586840 379898
rect 586240 344218 586422 344454
rect 586658 344218 586840 344454
rect 586240 344134 586840 344218
rect 586240 343898 586422 344134
rect 586658 343898 586840 344134
rect 586240 308454 586840 343898
rect 586240 308218 586422 308454
rect 586658 308218 586840 308454
rect 586240 308134 586840 308218
rect 586240 307898 586422 308134
rect 586658 307898 586840 308134
rect 586240 272454 586840 307898
rect 586240 272218 586422 272454
rect 586658 272218 586840 272454
rect 586240 272134 586840 272218
rect 586240 271898 586422 272134
rect 586658 271898 586840 272134
rect 586240 236454 586840 271898
rect 586240 236218 586422 236454
rect 586658 236218 586840 236454
rect 586240 236134 586840 236218
rect 586240 235898 586422 236134
rect 586658 235898 586840 236134
rect 586240 200454 586840 235898
rect 586240 200218 586422 200454
rect 586658 200218 586840 200454
rect 586240 200134 586840 200218
rect 586240 199898 586422 200134
rect 586658 199898 586840 200134
rect 586240 164454 586840 199898
rect 586240 164218 586422 164454
rect 586658 164218 586840 164454
rect 586240 164134 586840 164218
rect 586240 163898 586422 164134
rect 586658 163898 586840 164134
rect 586240 128454 586840 163898
rect 586240 128218 586422 128454
rect 586658 128218 586840 128454
rect 586240 128134 586840 128218
rect 586240 127898 586422 128134
rect 586658 127898 586840 128134
rect 586240 92454 586840 127898
rect 586240 92218 586422 92454
rect 586658 92218 586840 92454
rect 586240 92134 586840 92218
rect 586240 91898 586422 92134
rect 586658 91898 586840 92134
rect 586240 56454 586840 91898
rect 586240 56218 586422 56454
rect 586658 56218 586840 56454
rect 586240 56134 586840 56218
rect 586240 55898 586422 56134
rect 586658 55898 586840 56134
rect 586240 20454 586840 55898
rect 586240 20218 586422 20454
rect 586658 20218 586840 20454
rect 586240 20134 586840 20218
rect 586240 19898 586422 20134
rect 586658 19898 586840 20134
rect 586240 -1266 586840 19898
rect 586240 -1502 586422 -1266
rect 586658 -1502 586840 -1266
rect 586240 -1586 586840 -1502
rect 586240 -1822 586422 -1586
rect 586658 -1822 586840 -1586
rect 586240 -1844 586840 -1822
rect 587160 690054 587760 706122
rect 587160 689818 587342 690054
rect 587578 689818 587760 690054
rect 587160 689734 587760 689818
rect 587160 689498 587342 689734
rect 587578 689498 587760 689734
rect 587160 654054 587760 689498
rect 587160 653818 587342 654054
rect 587578 653818 587760 654054
rect 587160 653734 587760 653818
rect 587160 653498 587342 653734
rect 587578 653498 587760 653734
rect 587160 618054 587760 653498
rect 587160 617818 587342 618054
rect 587578 617818 587760 618054
rect 587160 617734 587760 617818
rect 587160 617498 587342 617734
rect 587578 617498 587760 617734
rect 587160 582054 587760 617498
rect 587160 581818 587342 582054
rect 587578 581818 587760 582054
rect 587160 581734 587760 581818
rect 587160 581498 587342 581734
rect 587578 581498 587760 581734
rect 587160 546054 587760 581498
rect 587160 545818 587342 546054
rect 587578 545818 587760 546054
rect 587160 545734 587760 545818
rect 587160 545498 587342 545734
rect 587578 545498 587760 545734
rect 587160 510054 587760 545498
rect 587160 509818 587342 510054
rect 587578 509818 587760 510054
rect 587160 509734 587760 509818
rect 587160 509498 587342 509734
rect 587578 509498 587760 509734
rect 587160 474054 587760 509498
rect 587160 473818 587342 474054
rect 587578 473818 587760 474054
rect 587160 473734 587760 473818
rect 587160 473498 587342 473734
rect 587578 473498 587760 473734
rect 587160 438054 587760 473498
rect 587160 437818 587342 438054
rect 587578 437818 587760 438054
rect 587160 437734 587760 437818
rect 587160 437498 587342 437734
rect 587578 437498 587760 437734
rect 587160 402054 587760 437498
rect 587160 401818 587342 402054
rect 587578 401818 587760 402054
rect 587160 401734 587760 401818
rect 587160 401498 587342 401734
rect 587578 401498 587760 401734
rect 587160 366054 587760 401498
rect 587160 365818 587342 366054
rect 587578 365818 587760 366054
rect 587160 365734 587760 365818
rect 587160 365498 587342 365734
rect 587578 365498 587760 365734
rect 587160 330054 587760 365498
rect 587160 329818 587342 330054
rect 587578 329818 587760 330054
rect 587160 329734 587760 329818
rect 587160 329498 587342 329734
rect 587578 329498 587760 329734
rect 587160 294054 587760 329498
rect 587160 293818 587342 294054
rect 587578 293818 587760 294054
rect 587160 293734 587760 293818
rect 587160 293498 587342 293734
rect 587578 293498 587760 293734
rect 587160 258054 587760 293498
rect 587160 257818 587342 258054
rect 587578 257818 587760 258054
rect 587160 257734 587760 257818
rect 587160 257498 587342 257734
rect 587578 257498 587760 257734
rect 587160 222054 587760 257498
rect 587160 221818 587342 222054
rect 587578 221818 587760 222054
rect 587160 221734 587760 221818
rect 587160 221498 587342 221734
rect 587578 221498 587760 221734
rect 587160 186054 587760 221498
rect 587160 185818 587342 186054
rect 587578 185818 587760 186054
rect 587160 185734 587760 185818
rect 587160 185498 587342 185734
rect 587578 185498 587760 185734
rect 587160 150054 587760 185498
rect 587160 149818 587342 150054
rect 587578 149818 587760 150054
rect 587160 149734 587760 149818
rect 587160 149498 587342 149734
rect 587578 149498 587760 149734
rect 587160 114054 587760 149498
rect 587160 113818 587342 114054
rect 587578 113818 587760 114054
rect 587160 113734 587760 113818
rect 587160 113498 587342 113734
rect 587578 113498 587760 113734
rect 587160 78054 587760 113498
rect 587160 77818 587342 78054
rect 587578 77818 587760 78054
rect 587160 77734 587760 77818
rect 587160 77498 587342 77734
rect 587578 77498 587760 77734
rect 587160 42054 587760 77498
rect 587160 41818 587342 42054
rect 587578 41818 587760 42054
rect 587160 41734 587760 41818
rect 587160 41498 587342 41734
rect 587578 41498 587760 41734
rect 587160 6054 587760 41498
rect 587160 5818 587342 6054
rect 587578 5818 587760 6054
rect 587160 5734 587760 5818
rect 587160 5498 587342 5734
rect 587578 5498 587760 5734
rect 580404 -2422 580586 -2186
rect 580822 -2422 581004 -2186
rect 580404 -2506 581004 -2422
rect 580404 -2742 580586 -2506
rect 580822 -2742 581004 -2506
rect 580404 -3684 581004 -2742
rect 587160 -2186 587760 5498
rect 587160 -2422 587342 -2186
rect 587578 -2422 587760 -2186
rect 587160 -2506 587760 -2422
rect 587160 -2742 587342 -2506
rect 587578 -2742 587760 -2506
rect 587160 -2764 587760 -2742
rect 588080 672054 588680 707042
rect 588080 671818 588262 672054
rect 588498 671818 588680 672054
rect 588080 671734 588680 671818
rect 588080 671498 588262 671734
rect 588498 671498 588680 671734
rect 588080 636054 588680 671498
rect 588080 635818 588262 636054
rect 588498 635818 588680 636054
rect 588080 635734 588680 635818
rect 588080 635498 588262 635734
rect 588498 635498 588680 635734
rect 588080 600054 588680 635498
rect 588080 599818 588262 600054
rect 588498 599818 588680 600054
rect 588080 599734 588680 599818
rect 588080 599498 588262 599734
rect 588498 599498 588680 599734
rect 588080 564054 588680 599498
rect 588080 563818 588262 564054
rect 588498 563818 588680 564054
rect 588080 563734 588680 563818
rect 588080 563498 588262 563734
rect 588498 563498 588680 563734
rect 588080 528054 588680 563498
rect 588080 527818 588262 528054
rect 588498 527818 588680 528054
rect 588080 527734 588680 527818
rect 588080 527498 588262 527734
rect 588498 527498 588680 527734
rect 588080 492054 588680 527498
rect 588080 491818 588262 492054
rect 588498 491818 588680 492054
rect 588080 491734 588680 491818
rect 588080 491498 588262 491734
rect 588498 491498 588680 491734
rect 588080 456054 588680 491498
rect 588080 455818 588262 456054
rect 588498 455818 588680 456054
rect 588080 455734 588680 455818
rect 588080 455498 588262 455734
rect 588498 455498 588680 455734
rect 588080 420054 588680 455498
rect 588080 419818 588262 420054
rect 588498 419818 588680 420054
rect 588080 419734 588680 419818
rect 588080 419498 588262 419734
rect 588498 419498 588680 419734
rect 588080 384054 588680 419498
rect 588080 383818 588262 384054
rect 588498 383818 588680 384054
rect 588080 383734 588680 383818
rect 588080 383498 588262 383734
rect 588498 383498 588680 383734
rect 588080 348054 588680 383498
rect 588080 347818 588262 348054
rect 588498 347818 588680 348054
rect 588080 347734 588680 347818
rect 588080 347498 588262 347734
rect 588498 347498 588680 347734
rect 588080 312054 588680 347498
rect 588080 311818 588262 312054
rect 588498 311818 588680 312054
rect 588080 311734 588680 311818
rect 588080 311498 588262 311734
rect 588498 311498 588680 311734
rect 588080 276054 588680 311498
rect 588080 275818 588262 276054
rect 588498 275818 588680 276054
rect 588080 275734 588680 275818
rect 588080 275498 588262 275734
rect 588498 275498 588680 275734
rect 588080 240054 588680 275498
rect 588080 239818 588262 240054
rect 588498 239818 588680 240054
rect 588080 239734 588680 239818
rect 588080 239498 588262 239734
rect 588498 239498 588680 239734
rect 588080 204054 588680 239498
rect 588080 203818 588262 204054
rect 588498 203818 588680 204054
rect 588080 203734 588680 203818
rect 588080 203498 588262 203734
rect 588498 203498 588680 203734
rect 588080 168054 588680 203498
rect 588080 167818 588262 168054
rect 588498 167818 588680 168054
rect 588080 167734 588680 167818
rect 588080 167498 588262 167734
rect 588498 167498 588680 167734
rect 588080 132054 588680 167498
rect 588080 131818 588262 132054
rect 588498 131818 588680 132054
rect 588080 131734 588680 131818
rect 588080 131498 588262 131734
rect 588498 131498 588680 131734
rect 588080 96054 588680 131498
rect 588080 95818 588262 96054
rect 588498 95818 588680 96054
rect 588080 95734 588680 95818
rect 588080 95498 588262 95734
rect 588498 95498 588680 95734
rect 588080 60054 588680 95498
rect 588080 59818 588262 60054
rect 588498 59818 588680 60054
rect 588080 59734 588680 59818
rect 588080 59498 588262 59734
rect 588498 59498 588680 59734
rect 588080 24054 588680 59498
rect 588080 23818 588262 24054
rect 588498 23818 588680 24054
rect 588080 23734 588680 23818
rect 588080 23498 588262 23734
rect 588498 23498 588680 23734
rect 588080 -3106 588680 23498
rect 588080 -3342 588262 -3106
rect 588498 -3342 588680 -3106
rect 588080 -3426 588680 -3342
rect 588080 -3662 588262 -3426
rect 588498 -3662 588680 -3426
rect 588080 -3684 588680 -3662
rect 589000 693654 589600 707962
rect 589000 693418 589182 693654
rect 589418 693418 589600 693654
rect 589000 693334 589600 693418
rect 589000 693098 589182 693334
rect 589418 693098 589600 693334
rect 589000 657654 589600 693098
rect 589000 657418 589182 657654
rect 589418 657418 589600 657654
rect 589000 657334 589600 657418
rect 589000 657098 589182 657334
rect 589418 657098 589600 657334
rect 589000 621654 589600 657098
rect 589000 621418 589182 621654
rect 589418 621418 589600 621654
rect 589000 621334 589600 621418
rect 589000 621098 589182 621334
rect 589418 621098 589600 621334
rect 589000 585654 589600 621098
rect 589000 585418 589182 585654
rect 589418 585418 589600 585654
rect 589000 585334 589600 585418
rect 589000 585098 589182 585334
rect 589418 585098 589600 585334
rect 589000 549654 589600 585098
rect 589000 549418 589182 549654
rect 589418 549418 589600 549654
rect 589000 549334 589600 549418
rect 589000 549098 589182 549334
rect 589418 549098 589600 549334
rect 589000 513654 589600 549098
rect 589000 513418 589182 513654
rect 589418 513418 589600 513654
rect 589000 513334 589600 513418
rect 589000 513098 589182 513334
rect 589418 513098 589600 513334
rect 589000 477654 589600 513098
rect 589000 477418 589182 477654
rect 589418 477418 589600 477654
rect 589000 477334 589600 477418
rect 589000 477098 589182 477334
rect 589418 477098 589600 477334
rect 589000 441654 589600 477098
rect 589000 441418 589182 441654
rect 589418 441418 589600 441654
rect 589000 441334 589600 441418
rect 589000 441098 589182 441334
rect 589418 441098 589600 441334
rect 589000 405654 589600 441098
rect 589000 405418 589182 405654
rect 589418 405418 589600 405654
rect 589000 405334 589600 405418
rect 589000 405098 589182 405334
rect 589418 405098 589600 405334
rect 589000 369654 589600 405098
rect 589000 369418 589182 369654
rect 589418 369418 589600 369654
rect 589000 369334 589600 369418
rect 589000 369098 589182 369334
rect 589418 369098 589600 369334
rect 589000 333654 589600 369098
rect 589000 333418 589182 333654
rect 589418 333418 589600 333654
rect 589000 333334 589600 333418
rect 589000 333098 589182 333334
rect 589418 333098 589600 333334
rect 589000 297654 589600 333098
rect 589000 297418 589182 297654
rect 589418 297418 589600 297654
rect 589000 297334 589600 297418
rect 589000 297098 589182 297334
rect 589418 297098 589600 297334
rect 589000 261654 589600 297098
rect 589000 261418 589182 261654
rect 589418 261418 589600 261654
rect 589000 261334 589600 261418
rect 589000 261098 589182 261334
rect 589418 261098 589600 261334
rect 589000 225654 589600 261098
rect 589000 225418 589182 225654
rect 589418 225418 589600 225654
rect 589000 225334 589600 225418
rect 589000 225098 589182 225334
rect 589418 225098 589600 225334
rect 589000 189654 589600 225098
rect 589000 189418 589182 189654
rect 589418 189418 589600 189654
rect 589000 189334 589600 189418
rect 589000 189098 589182 189334
rect 589418 189098 589600 189334
rect 589000 153654 589600 189098
rect 589000 153418 589182 153654
rect 589418 153418 589600 153654
rect 589000 153334 589600 153418
rect 589000 153098 589182 153334
rect 589418 153098 589600 153334
rect 589000 117654 589600 153098
rect 589000 117418 589182 117654
rect 589418 117418 589600 117654
rect 589000 117334 589600 117418
rect 589000 117098 589182 117334
rect 589418 117098 589600 117334
rect 589000 81654 589600 117098
rect 589000 81418 589182 81654
rect 589418 81418 589600 81654
rect 589000 81334 589600 81418
rect 589000 81098 589182 81334
rect 589418 81098 589600 81334
rect 589000 45654 589600 81098
rect 589000 45418 589182 45654
rect 589418 45418 589600 45654
rect 589000 45334 589600 45418
rect 589000 45098 589182 45334
rect 589418 45098 589600 45334
rect 589000 9654 589600 45098
rect 589000 9418 589182 9654
rect 589418 9418 589600 9654
rect 589000 9334 589600 9418
rect 589000 9098 589182 9334
rect 589418 9098 589600 9334
rect 589000 -4026 589600 9098
rect 589000 -4262 589182 -4026
rect 589418 -4262 589600 -4026
rect 589000 -4346 589600 -4262
rect 589000 -4582 589182 -4346
rect 589418 -4582 589600 -4346
rect 589000 -4604 589600 -4582
rect 589920 675654 590520 708882
rect 589920 675418 590102 675654
rect 590338 675418 590520 675654
rect 589920 675334 590520 675418
rect 589920 675098 590102 675334
rect 590338 675098 590520 675334
rect 589920 639654 590520 675098
rect 589920 639418 590102 639654
rect 590338 639418 590520 639654
rect 589920 639334 590520 639418
rect 589920 639098 590102 639334
rect 590338 639098 590520 639334
rect 589920 603654 590520 639098
rect 589920 603418 590102 603654
rect 590338 603418 590520 603654
rect 589920 603334 590520 603418
rect 589920 603098 590102 603334
rect 590338 603098 590520 603334
rect 589920 567654 590520 603098
rect 589920 567418 590102 567654
rect 590338 567418 590520 567654
rect 589920 567334 590520 567418
rect 589920 567098 590102 567334
rect 590338 567098 590520 567334
rect 589920 531654 590520 567098
rect 589920 531418 590102 531654
rect 590338 531418 590520 531654
rect 589920 531334 590520 531418
rect 589920 531098 590102 531334
rect 590338 531098 590520 531334
rect 589920 495654 590520 531098
rect 589920 495418 590102 495654
rect 590338 495418 590520 495654
rect 589920 495334 590520 495418
rect 589920 495098 590102 495334
rect 590338 495098 590520 495334
rect 589920 459654 590520 495098
rect 589920 459418 590102 459654
rect 590338 459418 590520 459654
rect 589920 459334 590520 459418
rect 589920 459098 590102 459334
rect 590338 459098 590520 459334
rect 589920 423654 590520 459098
rect 589920 423418 590102 423654
rect 590338 423418 590520 423654
rect 589920 423334 590520 423418
rect 589920 423098 590102 423334
rect 590338 423098 590520 423334
rect 589920 387654 590520 423098
rect 589920 387418 590102 387654
rect 590338 387418 590520 387654
rect 589920 387334 590520 387418
rect 589920 387098 590102 387334
rect 590338 387098 590520 387334
rect 589920 351654 590520 387098
rect 589920 351418 590102 351654
rect 590338 351418 590520 351654
rect 589920 351334 590520 351418
rect 589920 351098 590102 351334
rect 590338 351098 590520 351334
rect 589920 315654 590520 351098
rect 589920 315418 590102 315654
rect 590338 315418 590520 315654
rect 589920 315334 590520 315418
rect 589920 315098 590102 315334
rect 590338 315098 590520 315334
rect 589920 279654 590520 315098
rect 589920 279418 590102 279654
rect 590338 279418 590520 279654
rect 589920 279334 590520 279418
rect 589920 279098 590102 279334
rect 590338 279098 590520 279334
rect 589920 243654 590520 279098
rect 589920 243418 590102 243654
rect 590338 243418 590520 243654
rect 589920 243334 590520 243418
rect 589920 243098 590102 243334
rect 590338 243098 590520 243334
rect 589920 207654 590520 243098
rect 589920 207418 590102 207654
rect 590338 207418 590520 207654
rect 589920 207334 590520 207418
rect 589920 207098 590102 207334
rect 590338 207098 590520 207334
rect 589920 171654 590520 207098
rect 589920 171418 590102 171654
rect 590338 171418 590520 171654
rect 589920 171334 590520 171418
rect 589920 171098 590102 171334
rect 590338 171098 590520 171334
rect 589920 135654 590520 171098
rect 589920 135418 590102 135654
rect 590338 135418 590520 135654
rect 589920 135334 590520 135418
rect 589920 135098 590102 135334
rect 590338 135098 590520 135334
rect 589920 99654 590520 135098
rect 589920 99418 590102 99654
rect 590338 99418 590520 99654
rect 589920 99334 590520 99418
rect 589920 99098 590102 99334
rect 590338 99098 590520 99334
rect 589920 63654 590520 99098
rect 589920 63418 590102 63654
rect 590338 63418 590520 63654
rect 589920 63334 590520 63418
rect 589920 63098 590102 63334
rect 590338 63098 590520 63334
rect 589920 27654 590520 63098
rect 589920 27418 590102 27654
rect 590338 27418 590520 27654
rect 589920 27334 590520 27418
rect 589920 27098 590102 27334
rect 590338 27098 590520 27334
rect 589920 -4946 590520 27098
rect 589920 -5182 590102 -4946
rect 590338 -5182 590520 -4946
rect 589920 -5266 590520 -5182
rect 589920 -5502 590102 -5266
rect 590338 -5502 590520 -5266
rect 589920 -5524 590520 -5502
rect 590840 697254 591440 709802
rect 590840 697018 591022 697254
rect 591258 697018 591440 697254
rect 590840 696934 591440 697018
rect 590840 696698 591022 696934
rect 591258 696698 591440 696934
rect 590840 661254 591440 696698
rect 590840 661018 591022 661254
rect 591258 661018 591440 661254
rect 590840 660934 591440 661018
rect 590840 660698 591022 660934
rect 591258 660698 591440 660934
rect 590840 625254 591440 660698
rect 590840 625018 591022 625254
rect 591258 625018 591440 625254
rect 590840 624934 591440 625018
rect 590840 624698 591022 624934
rect 591258 624698 591440 624934
rect 590840 589254 591440 624698
rect 590840 589018 591022 589254
rect 591258 589018 591440 589254
rect 590840 588934 591440 589018
rect 590840 588698 591022 588934
rect 591258 588698 591440 588934
rect 590840 553254 591440 588698
rect 590840 553018 591022 553254
rect 591258 553018 591440 553254
rect 590840 552934 591440 553018
rect 590840 552698 591022 552934
rect 591258 552698 591440 552934
rect 590840 517254 591440 552698
rect 590840 517018 591022 517254
rect 591258 517018 591440 517254
rect 590840 516934 591440 517018
rect 590840 516698 591022 516934
rect 591258 516698 591440 516934
rect 590840 481254 591440 516698
rect 590840 481018 591022 481254
rect 591258 481018 591440 481254
rect 590840 480934 591440 481018
rect 590840 480698 591022 480934
rect 591258 480698 591440 480934
rect 590840 445254 591440 480698
rect 590840 445018 591022 445254
rect 591258 445018 591440 445254
rect 590840 444934 591440 445018
rect 590840 444698 591022 444934
rect 591258 444698 591440 444934
rect 590840 409254 591440 444698
rect 590840 409018 591022 409254
rect 591258 409018 591440 409254
rect 590840 408934 591440 409018
rect 590840 408698 591022 408934
rect 591258 408698 591440 408934
rect 590840 373254 591440 408698
rect 590840 373018 591022 373254
rect 591258 373018 591440 373254
rect 590840 372934 591440 373018
rect 590840 372698 591022 372934
rect 591258 372698 591440 372934
rect 590840 337254 591440 372698
rect 590840 337018 591022 337254
rect 591258 337018 591440 337254
rect 590840 336934 591440 337018
rect 590840 336698 591022 336934
rect 591258 336698 591440 336934
rect 590840 301254 591440 336698
rect 590840 301018 591022 301254
rect 591258 301018 591440 301254
rect 590840 300934 591440 301018
rect 590840 300698 591022 300934
rect 591258 300698 591440 300934
rect 590840 265254 591440 300698
rect 590840 265018 591022 265254
rect 591258 265018 591440 265254
rect 590840 264934 591440 265018
rect 590840 264698 591022 264934
rect 591258 264698 591440 264934
rect 590840 229254 591440 264698
rect 590840 229018 591022 229254
rect 591258 229018 591440 229254
rect 590840 228934 591440 229018
rect 590840 228698 591022 228934
rect 591258 228698 591440 228934
rect 590840 193254 591440 228698
rect 590840 193018 591022 193254
rect 591258 193018 591440 193254
rect 590840 192934 591440 193018
rect 590840 192698 591022 192934
rect 591258 192698 591440 192934
rect 590840 157254 591440 192698
rect 590840 157018 591022 157254
rect 591258 157018 591440 157254
rect 590840 156934 591440 157018
rect 590840 156698 591022 156934
rect 591258 156698 591440 156934
rect 590840 121254 591440 156698
rect 590840 121018 591022 121254
rect 591258 121018 591440 121254
rect 590840 120934 591440 121018
rect 590840 120698 591022 120934
rect 591258 120698 591440 120934
rect 590840 85254 591440 120698
rect 590840 85018 591022 85254
rect 591258 85018 591440 85254
rect 590840 84934 591440 85018
rect 590840 84698 591022 84934
rect 591258 84698 591440 84934
rect 590840 49254 591440 84698
rect 590840 49018 591022 49254
rect 591258 49018 591440 49254
rect 590840 48934 591440 49018
rect 590840 48698 591022 48934
rect 591258 48698 591440 48934
rect 590840 13254 591440 48698
rect 590840 13018 591022 13254
rect 591258 13018 591440 13254
rect 590840 12934 591440 13018
rect 590840 12698 591022 12934
rect 591258 12698 591440 12934
rect 590840 -5866 591440 12698
rect 590840 -6102 591022 -5866
rect 591258 -6102 591440 -5866
rect 590840 -6186 591440 -6102
rect 590840 -6422 591022 -6186
rect 591258 -6422 591440 -6186
rect 590840 -6444 591440 -6422
rect 591760 679254 592360 710722
rect 591760 679018 591942 679254
rect 592178 679018 592360 679254
rect 591760 678934 592360 679018
rect 591760 678698 591942 678934
rect 592178 678698 592360 678934
rect 591760 643254 592360 678698
rect 591760 643018 591942 643254
rect 592178 643018 592360 643254
rect 591760 642934 592360 643018
rect 591760 642698 591942 642934
rect 592178 642698 592360 642934
rect 591760 607254 592360 642698
rect 591760 607018 591942 607254
rect 592178 607018 592360 607254
rect 591760 606934 592360 607018
rect 591760 606698 591942 606934
rect 592178 606698 592360 606934
rect 591760 571254 592360 606698
rect 591760 571018 591942 571254
rect 592178 571018 592360 571254
rect 591760 570934 592360 571018
rect 591760 570698 591942 570934
rect 592178 570698 592360 570934
rect 591760 535254 592360 570698
rect 591760 535018 591942 535254
rect 592178 535018 592360 535254
rect 591760 534934 592360 535018
rect 591760 534698 591942 534934
rect 592178 534698 592360 534934
rect 591760 499254 592360 534698
rect 591760 499018 591942 499254
rect 592178 499018 592360 499254
rect 591760 498934 592360 499018
rect 591760 498698 591942 498934
rect 592178 498698 592360 498934
rect 591760 463254 592360 498698
rect 591760 463018 591942 463254
rect 592178 463018 592360 463254
rect 591760 462934 592360 463018
rect 591760 462698 591942 462934
rect 592178 462698 592360 462934
rect 591760 427254 592360 462698
rect 591760 427018 591942 427254
rect 592178 427018 592360 427254
rect 591760 426934 592360 427018
rect 591760 426698 591942 426934
rect 592178 426698 592360 426934
rect 591760 391254 592360 426698
rect 591760 391018 591942 391254
rect 592178 391018 592360 391254
rect 591760 390934 592360 391018
rect 591760 390698 591942 390934
rect 592178 390698 592360 390934
rect 591760 355254 592360 390698
rect 591760 355018 591942 355254
rect 592178 355018 592360 355254
rect 591760 354934 592360 355018
rect 591760 354698 591942 354934
rect 592178 354698 592360 354934
rect 591760 319254 592360 354698
rect 591760 319018 591942 319254
rect 592178 319018 592360 319254
rect 591760 318934 592360 319018
rect 591760 318698 591942 318934
rect 592178 318698 592360 318934
rect 591760 283254 592360 318698
rect 591760 283018 591942 283254
rect 592178 283018 592360 283254
rect 591760 282934 592360 283018
rect 591760 282698 591942 282934
rect 592178 282698 592360 282934
rect 591760 247254 592360 282698
rect 591760 247018 591942 247254
rect 592178 247018 592360 247254
rect 591760 246934 592360 247018
rect 591760 246698 591942 246934
rect 592178 246698 592360 246934
rect 591760 211254 592360 246698
rect 591760 211018 591942 211254
rect 592178 211018 592360 211254
rect 591760 210934 592360 211018
rect 591760 210698 591942 210934
rect 592178 210698 592360 210934
rect 591760 175254 592360 210698
rect 591760 175018 591942 175254
rect 592178 175018 592360 175254
rect 591760 174934 592360 175018
rect 591760 174698 591942 174934
rect 592178 174698 592360 174934
rect 591760 139254 592360 174698
rect 591760 139018 591942 139254
rect 592178 139018 592360 139254
rect 591760 138934 592360 139018
rect 591760 138698 591942 138934
rect 592178 138698 592360 138934
rect 591760 103254 592360 138698
rect 591760 103018 591942 103254
rect 592178 103018 592360 103254
rect 591760 102934 592360 103018
rect 591760 102698 591942 102934
rect 592178 102698 592360 102934
rect 591760 67254 592360 102698
rect 591760 67018 591942 67254
rect 592178 67018 592360 67254
rect 591760 66934 592360 67018
rect 591760 66698 591942 66934
rect 592178 66698 592360 66934
rect 591760 31254 592360 66698
rect 591760 31018 591942 31254
rect 592178 31018 592360 31254
rect 591760 30934 592360 31018
rect 591760 30698 591942 30934
rect 592178 30698 592360 30934
rect 569604 -7022 569786 -6786
rect 570022 -7022 570204 -6786
rect 569604 -7106 570204 -7022
rect 569604 -7342 569786 -7106
rect 570022 -7342 570204 -7106
rect 569604 -7364 570204 -7342
rect 591760 -6786 592360 30698
rect 591760 -7022 591942 -6786
rect 592178 -7022 592360 -6786
rect 591760 -7106 592360 -7022
rect 591760 -7342 591942 -7106
rect 592178 -7342 592360 -7106
rect 591760 -7364 592360 -7342
<< via4 >>
rect -8254 711042 -8018 711278
rect -8254 710722 -8018 710958
rect -8254 679018 -8018 679254
rect -8254 678698 -8018 678934
rect -8254 643018 -8018 643254
rect -8254 642698 -8018 642934
rect -8254 607018 -8018 607254
rect -8254 606698 -8018 606934
rect -8254 571018 -8018 571254
rect -8254 570698 -8018 570934
rect -8254 535018 -8018 535254
rect -8254 534698 -8018 534934
rect -8254 499018 -8018 499254
rect -8254 498698 -8018 498934
rect -8254 463018 -8018 463254
rect -8254 462698 -8018 462934
rect -8254 427018 -8018 427254
rect -8254 426698 -8018 426934
rect -8254 391018 -8018 391254
rect -8254 390698 -8018 390934
rect -8254 355018 -8018 355254
rect -8254 354698 -8018 354934
rect -8254 319018 -8018 319254
rect -8254 318698 -8018 318934
rect -8254 283018 -8018 283254
rect -8254 282698 -8018 282934
rect -8254 247018 -8018 247254
rect -8254 246698 -8018 246934
rect -8254 211018 -8018 211254
rect -8254 210698 -8018 210934
rect -8254 175018 -8018 175254
rect -8254 174698 -8018 174934
rect -8254 139018 -8018 139254
rect -8254 138698 -8018 138934
rect -8254 103018 -8018 103254
rect -8254 102698 -8018 102934
rect -8254 67018 -8018 67254
rect -8254 66698 -8018 66934
rect -8254 31018 -8018 31254
rect -8254 30698 -8018 30934
rect -7334 710122 -7098 710358
rect -7334 709802 -7098 710038
rect 11786 710122 12022 710358
rect 11786 709802 12022 710038
rect -7334 697018 -7098 697254
rect -7334 696698 -7098 696934
rect -7334 661018 -7098 661254
rect -7334 660698 -7098 660934
rect -7334 625018 -7098 625254
rect -7334 624698 -7098 624934
rect -7334 589018 -7098 589254
rect -7334 588698 -7098 588934
rect -7334 553018 -7098 553254
rect -7334 552698 -7098 552934
rect -7334 517018 -7098 517254
rect -7334 516698 -7098 516934
rect -7334 481018 -7098 481254
rect -7334 480698 -7098 480934
rect -7334 445018 -7098 445254
rect -7334 444698 -7098 444934
rect -7334 409018 -7098 409254
rect -7334 408698 -7098 408934
rect -7334 373018 -7098 373254
rect -7334 372698 -7098 372934
rect -7334 337018 -7098 337254
rect -7334 336698 -7098 336934
rect -7334 301018 -7098 301254
rect -7334 300698 -7098 300934
rect -7334 265018 -7098 265254
rect -7334 264698 -7098 264934
rect -7334 229018 -7098 229254
rect -7334 228698 -7098 228934
rect -7334 193018 -7098 193254
rect -7334 192698 -7098 192934
rect -7334 157018 -7098 157254
rect -7334 156698 -7098 156934
rect -7334 121018 -7098 121254
rect -7334 120698 -7098 120934
rect -7334 85018 -7098 85254
rect -7334 84698 -7098 84934
rect -7334 49018 -7098 49254
rect -7334 48698 -7098 48934
rect -7334 13018 -7098 13254
rect -7334 12698 -7098 12934
rect -6414 709202 -6178 709438
rect -6414 708882 -6178 709118
rect -6414 675418 -6178 675654
rect -6414 675098 -6178 675334
rect -6414 639418 -6178 639654
rect -6414 639098 -6178 639334
rect -6414 603418 -6178 603654
rect -6414 603098 -6178 603334
rect -6414 567418 -6178 567654
rect -6414 567098 -6178 567334
rect -6414 531418 -6178 531654
rect -6414 531098 -6178 531334
rect -6414 495418 -6178 495654
rect -6414 495098 -6178 495334
rect -6414 459418 -6178 459654
rect -6414 459098 -6178 459334
rect -6414 423418 -6178 423654
rect -6414 423098 -6178 423334
rect -6414 387418 -6178 387654
rect -6414 387098 -6178 387334
rect -6414 351418 -6178 351654
rect -6414 351098 -6178 351334
rect -6414 315418 -6178 315654
rect -6414 315098 -6178 315334
rect -6414 279418 -6178 279654
rect -6414 279098 -6178 279334
rect -6414 243418 -6178 243654
rect -6414 243098 -6178 243334
rect -6414 207418 -6178 207654
rect -6414 207098 -6178 207334
rect -6414 171418 -6178 171654
rect -6414 171098 -6178 171334
rect -6414 135418 -6178 135654
rect -6414 135098 -6178 135334
rect -6414 99418 -6178 99654
rect -6414 99098 -6178 99334
rect -6414 63418 -6178 63654
rect -6414 63098 -6178 63334
rect -6414 27418 -6178 27654
rect -6414 27098 -6178 27334
rect -5494 708282 -5258 708518
rect -5494 707962 -5258 708198
rect 8186 708282 8422 708518
rect 8186 707962 8422 708198
rect -5494 693418 -5258 693654
rect -5494 693098 -5258 693334
rect -5494 657418 -5258 657654
rect -5494 657098 -5258 657334
rect -5494 621418 -5258 621654
rect -5494 621098 -5258 621334
rect -5494 585418 -5258 585654
rect -5494 585098 -5258 585334
rect -5494 549418 -5258 549654
rect -5494 549098 -5258 549334
rect -5494 513418 -5258 513654
rect -5494 513098 -5258 513334
rect -5494 477418 -5258 477654
rect -5494 477098 -5258 477334
rect -5494 441418 -5258 441654
rect -5494 441098 -5258 441334
rect -5494 405418 -5258 405654
rect -5494 405098 -5258 405334
rect -5494 369418 -5258 369654
rect -5494 369098 -5258 369334
rect -5494 333418 -5258 333654
rect -5494 333098 -5258 333334
rect -5494 297418 -5258 297654
rect -5494 297098 -5258 297334
rect -5494 261418 -5258 261654
rect -5494 261098 -5258 261334
rect -5494 225418 -5258 225654
rect -5494 225098 -5258 225334
rect -5494 189418 -5258 189654
rect -5494 189098 -5258 189334
rect -5494 153418 -5258 153654
rect -5494 153098 -5258 153334
rect -5494 117418 -5258 117654
rect -5494 117098 -5258 117334
rect -5494 81418 -5258 81654
rect -5494 81098 -5258 81334
rect -5494 45418 -5258 45654
rect -5494 45098 -5258 45334
rect -5494 9418 -5258 9654
rect -5494 9098 -5258 9334
rect -4574 707362 -4338 707598
rect -4574 707042 -4338 707278
rect -4574 671818 -4338 672054
rect -4574 671498 -4338 671734
rect -4574 635818 -4338 636054
rect -4574 635498 -4338 635734
rect -4574 599818 -4338 600054
rect -4574 599498 -4338 599734
rect -4574 563818 -4338 564054
rect -4574 563498 -4338 563734
rect -4574 527818 -4338 528054
rect -4574 527498 -4338 527734
rect -4574 491818 -4338 492054
rect -4574 491498 -4338 491734
rect -4574 455818 -4338 456054
rect -4574 455498 -4338 455734
rect -4574 419818 -4338 420054
rect -4574 419498 -4338 419734
rect -4574 383818 -4338 384054
rect -4574 383498 -4338 383734
rect -4574 347818 -4338 348054
rect -4574 347498 -4338 347734
rect -4574 311818 -4338 312054
rect -4574 311498 -4338 311734
rect -4574 275818 -4338 276054
rect -4574 275498 -4338 275734
rect -4574 239818 -4338 240054
rect -4574 239498 -4338 239734
rect -4574 203818 -4338 204054
rect -4574 203498 -4338 203734
rect -4574 167818 -4338 168054
rect -4574 167498 -4338 167734
rect -4574 131818 -4338 132054
rect -4574 131498 -4338 131734
rect -4574 95818 -4338 96054
rect -4574 95498 -4338 95734
rect -4574 59818 -4338 60054
rect -4574 59498 -4338 59734
rect -4574 23818 -4338 24054
rect -4574 23498 -4338 23734
rect -3654 706442 -3418 706678
rect -3654 706122 -3418 706358
rect 4586 706442 4822 706678
rect 4586 706122 4822 706358
rect -3654 689818 -3418 690054
rect -3654 689498 -3418 689734
rect -3654 653818 -3418 654054
rect -3654 653498 -3418 653734
rect -3654 617818 -3418 618054
rect -3654 617498 -3418 617734
rect -3654 581818 -3418 582054
rect -3654 581498 -3418 581734
rect -3654 545818 -3418 546054
rect -3654 545498 -3418 545734
rect -3654 509818 -3418 510054
rect -3654 509498 -3418 509734
rect -3654 473818 -3418 474054
rect -3654 473498 -3418 473734
rect -3654 437818 -3418 438054
rect -3654 437498 -3418 437734
rect -3654 401818 -3418 402054
rect -3654 401498 -3418 401734
rect -3654 365818 -3418 366054
rect -3654 365498 -3418 365734
rect -3654 329818 -3418 330054
rect -3654 329498 -3418 329734
rect -3654 293818 -3418 294054
rect -3654 293498 -3418 293734
rect -3654 257818 -3418 258054
rect -3654 257498 -3418 257734
rect -3654 221818 -3418 222054
rect -3654 221498 -3418 221734
rect -3654 185818 -3418 186054
rect -3654 185498 -3418 185734
rect -3654 149818 -3418 150054
rect -3654 149498 -3418 149734
rect -3654 113818 -3418 114054
rect -3654 113498 -3418 113734
rect -3654 77818 -3418 78054
rect -3654 77498 -3418 77734
rect -3654 41818 -3418 42054
rect -3654 41498 -3418 41734
rect -3654 5818 -3418 6054
rect -3654 5498 -3418 5734
rect -2734 705522 -2498 705758
rect -2734 705202 -2498 705438
rect -2734 668218 -2498 668454
rect -2734 667898 -2498 668134
rect -2734 632218 -2498 632454
rect -2734 631898 -2498 632134
rect -2734 596218 -2498 596454
rect -2734 595898 -2498 596134
rect -2734 560218 -2498 560454
rect -2734 559898 -2498 560134
rect -2734 524218 -2498 524454
rect -2734 523898 -2498 524134
rect -2734 488218 -2498 488454
rect -2734 487898 -2498 488134
rect -2734 452218 -2498 452454
rect -2734 451898 -2498 452134
rect -2734 416218 -2498 416454
rect -2734 415898 -2498 416134
rect -2734 380218 -2498 380454
rect -2734 379898 -2498 380134
rect -2734 344218 -2498 344454
rect -2734 343898 -2498 344134
rect -2734 308218 -2498 308454
rect -2734 307898 -2498 308134
rect -2734 272218 -2498 272454
rect -2734 271898 -2498 272134
rect -2734 236218 -2498 236454
rect -2734 235898 -2498 236134
rect -2734 200218 -2498 200454
rect -2734 199898 -2498 200134
rect -2734 164218 -2498 164454
rect -2734 163898 -2498 164134
rect -2734 128218 -2498 128454
rect -2734 127898 -2498 128134
rect -2734 92218 -2498 92454
rect -2734 91898 -2498 92134
rect -2734 56218 -2498 56454
rect -2734 55898 -2498 56134
rect -2734 20218 -2498 20454
rect -2734 19898 -2498 20134
rect -1814 704602 -1578 704838
rect -1814 704282 -1578 704518
rect -1814 686218 -1578 686454
rect -1814 685898 -1578 686134
rect -1814 650218 -1578 650454
rect -1814 649898 -1578 650134
rect -1814 614218 -1578 614454
rect -1814 613898 -1578 614134
rect -1814 578218 -1578 578454
rect -1814 577898 -1578 578134
rect -1814 542218 -1578 542454
rect -1814 541898 -1578 542134
rect -1814 506218 -1578 506454
rect -1814 505898 -1578 506134
rect -1814 470218 -1578 470454
rect -1814 469898 -1578 470134
rect -1814 434218 -1578 434454
rect -1814 433898 -1578 434134
rect -1814 398218 -1578 398454
rect -1814 397898 -1578 398134
rect -1814 362218 -1578 362454
rect -1814 361898 -1578 362134
rect -1814 326218 -1578 326454
rect -1814 325898 -1578 326134
rect -1814 290218 -1578 290454
rect -1814 289898 -1578 290134
rect -1814 254218 -1578 254454
rect -1814 253898 -1578 254134
rect -1814 218218 -1578 218454
rect -1814 217898 -1578 218134
rect -1814 182218 -1578 182454
rect -1814 181898 -1578 182134
rect -1814 146218 -1578 146454
rect -1814 145898 -1578 146134
rect -1814 110218 -1578 110454
rect -1814 109898 -1578 110134
rect -1814 74218 -1578 74454
rect -1814 73898 -1578 74134
rect -1814 38218 -1578 38454
rect -1814 37898 -1578 38134
rect -1814 2218 -1578 2454
rect -1814 1898 -1578 2134
rect -1814 -582 -1578 -346
rect -1814 -902 -1578 -666
rect 986 704602 1222 704838
rect 986 704282 1222 704518
rect 986 686218 1222 686454
rect 986 685898 1222 686134
rect 986 650218 1222 650454
rect 986 649898 1222 650134
rect 986 614218 1222 614454
rect 986 613898 1222 614134
rect 986 578218 1222 578454
rect 986 577898 1222 578134
rect 986 542218 1222 542454
rect 986 541898 1222 542134
rect 986 506218 1222 506454
rect 986 505898 1222 506134
rect 986 470218 1222 470454
rect 986 469898 1222 470134
rect 986 434218 1222 434454
rect 986 433898 1222 434134
rect 986 398218 1222 398454
rect 986 397898 1222 398134
rect 986 362218 1222 362454
rect 986 361898 1222 362134
rect 986 326218 1222 326454
rect 986 325898 1222 326134
rect 986 290218 1222 290454
rect 986 289898 1222 290134
rect 986 254218 1222 254454
rect 986 253898 1222 254134
rect 986 218218 1222 218454
rect 986 217898 1222 218134
rect 986 182218 1222 182454
rect 986 181898 1222 182134
rect 986 146218 1222 146454
rect 986 145898 1222 146134
rect 986 110218 1222 110454
rect 986 109898 1222 110134
rect 986 74218 1222 74454
rect 986 73898 1222 74134
rect 986 38218 1222 38454
rect 986 37898 1222 38134
rect 986 2218 1222 2454
rect 986 1898 1222 2134
rect 986 -582 1222 -346
rect 986 -902 1222 -666
rect -2734 -1502 -2498 -1266
rect -2734 -1822 -2498 -1586
rect 4586 689818 4822 690054
rect 4586 689498 4822 689734
rect 4586 653818 4822 654054
rect 4586 653498 4822 653734
rect 4586 617818 4822 618054
rect 4586 617498 4822 617734
rect 4586 581818 4822 582054
rect 4586 581498 4822 581734
rect 4586 545818 4822 546054
rect 4586 545498 4822 545734
rect 4586 509818 4822 510054
rect 4586 509498 4822 509734
rect 4586 473818 4822 474054
rect 4586 473498 4822 473734
rect 4586 437818 4822 438054
rect 4586 437498 4822 437734
rect 4586 401818 4822 402054
rect 4586 401498 4822 401734
rect 4586 365818 4822 366054
rect 4586 365498 4822 365734
rect 4586 329818 4822 330054
rect 4586 329498 4822 329734
rect 4586 293818 4822 294054
rect 4586 293498 4822 293734
rect 4586 257818 4822 258054
rect 4586 257498 4822 257734
rect 4586 221818 4822 222054
rect 4586 221498 4822 221734
rect 4586 185818 4822 186054
rect 4586 185498 4822 185734
rect 4586 149818 4822 150054
rect 4586 149498 4822 149734
rect 4586 113818 4822 114054
rect 4586 113498 4822 113734
rect 4586 77818 4822 78054
rect 4586 77498 4822 77734
rect 4586 41818 4822 42054
rect 4586 41498 4822 41734
rect 4586 5818 4822 6054
rect 4586 5498 4822 5734
rect -3654 -2422 -3418 -2186
rect -3654 -2742 -3418 -2506
rect 4586 -2422 4822 -2186
rect 4586 -2742 4822 -2506
rect -4574 -3342 -4338 -3106
rect -4574 -3662 -4338 -3426
rect 8186 693418 8422 693654
rect 8186 693098 8422 693334
rect 8186 657418 8422 657654
rect 8186 657098 8422 657334
rect 8186 621418 8422 621654
rect 8186 621098 8422 621334
rect 8186 585418 8422 585654
rect 8186 585098 8422 585334
rect 8186 549418 8422 549654
rect 8186 549098 8422 549334
rect 8186 513418 8422 513654
rect 8186 513098 8422 513334
rect 8186 477418 8422 477654
rect 8186 477098 8422 477334
rect 8186 441418 8422 441654
rect 8186 441098 8422 441334
rect 8186 405418 8422 405654
rect 8186 405098 8422 405334
rect 8186 369418 8422 369654
rect 8186 369098 8422 369334
rect 8186 333418 8422 333654
rect 8186 333098 8422 333334
rect 8186 297418 8422 297654
rect 8186 297098 8422 297334
rect 8186 261418 8422 261654
rect 8186 261098 8422 261334
rect 8186 225418 8422 225654
rect 8186 225098 8422 225334
rect 8186 189418 8422 189654
rect 8186 189098 8422 189334
rect 8186 153418 8422 153654
rect 8186 153098 8422 153334
rect 8186 117418 8422 117654
rect 8186 117098 8422 117334
rect 8186 81418 8422 81654
rect 8186 81098 8422 81334
rect 8186 45418 8422 45654
rect 8186 45098 8422 45334
rect 8186 9418 8422 9654
rect 8186 9098 8422 9334
rect -5494 -4262 -5258 -4026
rect -5494 -4582 -5258 -4346
rect 8186 -4262 8422 -4026
rect 8186 -4582 8422 -4346
rect -6414 -5182 -6178 -4946
rect -6414 -5502 -6178 -5266
rect 29786 711042 30022 711278
rect 29786 710722 30022 710958
rect 26186 709202 26422 709438
rect 26186 708882 26422 709118
rect 22586 707362 22822 707598
rect 22586 707042 22822 707278
rect 11786 697018 12022 697254
rect 11786 696698 12022 696934
rect 11786 661018 12022 661254
rect 11786 660698 12022 660934
rect 11786 625018 12022 625254
rect 11786 624698 12022 624934
rect 11786 589018 12022 589254
rect 11786 588698 12022 588934
rect 11786 553018 12022 553254
rect 11786 552698 12022 552934
rect 11786 517018 12022 517254
rect 11786 516698 12022 516934
rect 11786 481018 12022 481254
rect 11786 480698 12022 480934
rect 11786 445018 12022 445254
rect 11786 444698 12022 444934
rect 11786 409018 12022 409254
rect 11786 408698 12022 408934
rect 11786 373018 12022 373254
rect 11786 372698 12022 372934
rect 11786 337018 12022 337254
rect 11786 336698 12022 336934
rect 11786 301018 12022 301254
rect 11786 300698 12022 300934
rect 11786 265018 12022 265254
rect 11786 264698 12022 264934
rect 11786 229018 12022 229254
rect 11786 228698 12022 228934
rect 11786 193018 12022 193254
rect 11786 192698 12022 192934
rect 11786 157018 12022 157254
rect 11786 156698 12022 156934
rect 11786 121018 12022 121254
rect 11786 120698 12022 120934
rect 11786 85018 12022 85254
rect 11786 84698 12022 84934
rect 11786 49018 12022 49254
rect 11786 48698 12022 48934
rect 11786 13018 12022 13254
rect 11786 12698 12022 12934
rect -7334 -6102 -7098 -5866
rect -7334 -6422 -7098 -6186
rect 18986 705522 19222 705758
rect 18986 705202 19222 705438
rect 18986 668218 19222 668454
rect 18986 667898 19222 668134
rect 18986 632218 19222 632454
rect 18986 631898 19222 632134
rect 18986 596218 19222 596454
rect 18986 595898 19222 596134
rect 18986 560218 19222 560454
rect 18986 559898 19222 560134
rect 18986 524218 19222 524454
rect 18986 523898 19222 524134
rect 18986 488218 19222 488454
rect 18986 487898 19222 488134
rect 18986 452218 19222 452454
rect 18986 451898 19222 452134
rect 18986 416218 19222 416454
rect 18986 415898 19222 416134
rect 18986 380218 19222 380454
rect 18986 379898 19222 380134
rect 18986 344218 19222 344454
rect 18986 343898 19222 344134
rect 18986 308218 19222 308454
rect 18986 307898 19222 308134
rect 18986 272218 19222 272454
rect 18986 271898 19222 272134
rect 18986 236218 19222 236454
rect 18986 235898 19222 236134
rect 18986 200218 19222 200454
rect 18986 199898 19222 200134
rect 18986 164218 19222 164454
rect 18986 163898 19222 164134
rect 18986 128218 19222 128454
rect 18986 127898 19222 128134
rect 18986 92218 19222 92454
rect 18986 91898 19222 92134
rect 18986 56218 19222 56454
rect 18986 55898 19222 56134
rect 18986 20218 19222 20454
rect 18986 19898 19222 20134
rect 18986 -1502 19222 -1266
rect 18986 -1822 19222 -1586
rect 22586 671818 22822 672054
rect 22586 671498 22822 671734
rect 22586 635818 22822 636054
rect 22586 635498 22822 635734
rect 22586 599818 22822 600054
rect 22586 599498 22822 599734
rect 22586 563818 22822 564054
rect 22586 563498 22822 563734
rect 22586 527818 22822 528054
rect 22586 527498 22822 527734
rect 22586 491818 22822 492054
rect 22586 491498 22822 491734
rect 22586 455818 22822 456054
rect 22586 455498 22822 455734
rect 22586 419818 22822 420054
rect 22586 419498 22822 419734
rect 22586 383818 22822 384054
rect 22586 383498 22822 383734
rect 22586 347818 22822 348054
rect 22586 347498 22822 347734
rect 22586 311818 22822 312054
rect 22586 311498 22822 311734
rect 22586 275818 22822 276054
rect 22586 275498 22822 275734
rect 22586 239818 22822 240054
rect 22586 239498 22822 239734
rect 22586 203818 22822 204054
rect 22586 203498 22822 203734
rect 22586 167818 22822 168054
rect 22586 167498 22822 167734
rect 22586 131818 22822 132054
rect 22586 131498 22822 131734
rect 22586 95818 22822 96054
rect 22586 95498 22822 95734
rect 22586 59818 22822 60054
rect 22586 59498 22822 59734
rect 22586 23818 22822 24054
rect 22586 23498 22822 23734
rect 22586 -3342 22822 -3106
rect 22586 -3662 22822 -3426
rect 26186 675418 26422 675654
rect 26186 675098 26422 675334
rect 26186 639418 26422 639654
rect 26186 639098 26422 639334
rect 26186 603418 26422 603654
rect 26186 603098 26422 603334
rect 26186 567418 26422 567654
rect 26186 567098 26422 567334
rect 26186 531418 26422 531654
rect 26186 531098 26422 531334
rect 26186 495418 26422 495654
rect 26186 495098 26422 495334
rect 26186 459418 26422 459654
rect 26186 459098 26422 459334
rect 26186 423418 26422 423654
rect 26186 423098 26422 423334
rect 26186 387418 26422 387654
rect 26186 387098 26422 387334
rect 26186 351418 26422 351654
rect 26186 351098 26422 351334
rect 26186 315418 26422 315654
rect 26186 315098 26422 315334
rect 26186 279418 26422 279654
rect 26186 279098 26422 279334
rect 26186 243418 26422 243654
rect 26186 243098 26422 243334
rect 26186 207418 26422 207654
rect 26186 207098 26422 207334
rect 26186 171418 26422 171654
rect 26186 171098 26422 171334
rect 26186 135418 26422 135654
rect 26186 135098 26422 135334
rect 26186 99418 26422 99654
rect 26186 99098 26422 99334
rect 26186 63418 26422 63654
rect 26186 63098 26422 63334
rect 26186 27418 26422 27654
rect 26186 27098 26422 27334
rect 26186 -5182 26422 -4946
rect 26186 -5502 26422 -5266
rect 47786 710122 48022 710358
rect 47786 709802 48022 710038
rect 44186 708282 44422 708518
rect 44186 707962 44422 708198
rect 40586 706442 40822 706678
rect 40586 706122 40822 706358
rect 29786 679018 30022 679254
rect 29786 678698 30022 678934
rect 29786 643018 30022 643254
rect 29786 642698 30022 642934
rect 29786 607018 30022 607254
rect 29786 606698 30022 606934
rect 29786 571018 30022 571254
rect 29786 570698 30022 570934
rect 29786 535018 30022 535254
rect 29786 534698 30022 534934
rect 29786 499018 30022 499254
rect 29786 498698 30022 498934
rect 29786 463018 30022 463254
rect 29786 462698 30022 462934
rect 29786 427018 30022 427254
rect 29786 426698 30022 426934
rect 29786 391018 30022 391254
rect 29786 390698 30022 390934
rect 29786 355018 30022 355254
rect 29786 354698 30022 354934
rect 29786 319018 30022 319254
rect 29786 318698 30022 318934
rect 29786 283018 30022 283254
rect 29786 282698 30022 282934
rect 29786 247018 30022 247254
rect 29786 246698 30022 246934
rect 29786 211018 30022 211254
rect 29786 210698 30022 210934
rect 29786 175018 30022 175254
rect 29786 174698 30022 174934
rect 29786 139018 30022 139254
rect 29786 138698 30022 138934
rect 29786 103018 30022 103254
rect 29786 102698 30022 102934
rect 29786 67018 30022 67254
rect 29786 66698 30022 66934
rect 29786 31018 30022 31254
rect 29786 30698 30022 30934
rect 11786 -6102 12022 -5866
rect 11786 -6422 12022 -6186
rect -8254 -7022 -8018 -6786
rect -8254 -7342 -8018 -7106
rect 36986 704602 37222 704838
rect 36986 704282 37222 704518
rect 36986 686218 37222 686454
rect 36986 685898 37222 686134
rect 36986 650218 37222 650454
rect 36986 649898 37222 650134
rect 36986 614218 37222 614454
rect 36986 613898 37222 614134
rect 36986 578218 37222 578454
rect 36986 577898 37222 578134
rect 36986 542218 37222 542454
rect 36986 541898 37222 542134
rect 36986 506218 37222 506454
rect 36986 505898 37222 506134
rect 36986 470218 37222 470454
rect 36986 469898 37222 470134
rect 36986 434218 37222 434454
rect 36986 433898 37222 434134
rect 36986 398218 37222 398454
rect 36986 397898 37222 398134
rect 36986 362218 37222 362454
rect 36986 361898 37222 362134
rect 36986 326218 37222 326454
rect 36986 325898 37222 326134
rect 36986 290218 37222 290454
rect 36986 289898 37222 290134
rect 36986 254218 37222 254454
rect 36986 253898 37222 254134
rect 36986 218218 37222 218454
rect 36986 217898 37222 218134
rect 36986 182218 37222 182454
rect 36986 181898 37222 182134
rect 36986 146218 37222 146454
rect 36986 145898 37222 146134
rect 36986 110218 37222 110454
rect 36986 109898 37222 110134
rect 36986 74218 37222 74454
rect 36986 73898 37222 74134
rect 36986 38218 37222 38454
rect 36986 37898 37222 38134
rect 36986 2218 37222 2454
rect 36986 1898 37222 2134
rect 36986 -582 37222 -346
rect 36986 -902 37222 -666
rect 40586 689818 40822 690054
rect 40586 689498 40822 689734
rect 40586 653818 40822 654054
rect 40586 653498 40822 653734
rect 40586 617818 40822 618054
rect 40586 617498 40822 617734
rect 40586 581818 40822 582054
rect 40586 581498 40822 581734
rect 40586 545818 40822 546054
rect 40586 545498 40822 545734
rect 40586 509818 40822 510054
rect 40586 509498 40822 509734
rect 40586 473818 40822 474054
rect 40586 473498 40822 473734
rect 40586 437818 40822 438054
rect 40586 437498 40822 437734
rect 40586 401818 40822 402054
rect 40586 401498 40822 401734
rect 40586 365818 40822 366054
rect 40586 365498 40822 365734
rect 40586 329818 40822 330054
rect 40586 329498 40822 329734
rect 40586 293818 40822 294054
rect 40586 293498 40822 293734
rect 40586 257818 40822 258054
rect 40586 257498 40822 257734
rect 40586 221818 40822 222054
rect 40586 221498 40822 221734
rect 40586 185818 40822 186054
rect 40586 185498 40822 185734
rect 40586 149818 40822 150054
rect 40586 149498 40822 149734
rect 40586 113818 40822 114054
rect 40586 113498 40822 113734
rect 40586 77818 40822 78054
rect 40586 77498 40822 77734
rect 40586 41818 40822 42054
rect 40586 41498 40822 41734
rect 40586 5818 40822 6054
rect 40586 5498 40822 5734
rect 40586 -2422 40822 -2186
rect 40586 -2742 40822 -2506
rect 44186 693418 44422 693654
rect 44186 693098 44422 693334
rect 44186 657418 44422 657654
rect 44186 657098 44422 657334
rect 44186 621418 44422 621654
rect 44186 621098 44422 621334
rect 44186 585418 44422 585654
rect 44186 585098 44422 585334
rect 44186 549418 44422 549654
rect 44186 549098 44422 549334
rect 44186 513418 44422 513654
rect 44186 513098 44422 513334
rect 44186 477418 44422 477654
rect 44186 477098 44422 477334
rect 44186 441418 44422 441654
rect 44186 441098 44422 441334
rect 44186 405418 44422 405654
rect 44186 405098 44422 405334
rect 44186 369418 44422 369654
rect 44186 369098 44422 369334
rect 44186 333418 44422 333654
rect 44186 333098 44422 333334
rect 44186 297418 44422 297654
rect 44186 297098 44422 297334
rect 44186 261418 44422 261654
rect 44186 261098 44422 261334
rect 44186 225418 44422 225654
rect 44186 225098 44422 225334
rect 44186 189418 44422 189654
rect 44186 189098 44422 189334
rect 44186 153418 44422 153654
rect 44186 153098 44422 153334
rect 44186 117418 44422 117654
rect 44186 117098 44422 117334
rect 44186 81418 44422 81654
rect 44186 81098 44422 81334
rect 44186 45418 44422 45654
rect 44186 45098 44422 45334
rect 44186 9418 44422 9654
rect 44186 9098 44422 9334
rect 44186 -4262 44422 -4026
rect 44186 -4582 44422 -4346
rect 65786 711042 66022 711278
rect 65786 710722 66022 710958
rect 62186 709202 62422 709438
rect 62186 708882 62422 709118
rect 58586 707362 58822 707598
rect 58586 707042 58822 707278
rect 47786 697018 48022 697254
rect 47786 696698 48022 696934
rect 47786 661018 48022 661254
rect 47786 660698 48022 660934
rect 47786 625018 48022 625254
rect 47786 624698 48022 624934
rect 47786 589018 48022 589254
rect 47786 588698 48022 588934
rect 47786 553018 48022 553254
rect 47786 552698 48022 552934
rect 47786 517018 48022 517254
rect 47786 516698 48022 516934
rect 47786 481018 48022 481254
rect 47786 480698 48022 480934
rect 47786 445018 48022 445254
rect 47786 444698 48022 444934
rect 47786 409018 48022 409254
rect 47786 408698 48022 408934
rect 47786 373018 48022 373254
rect 47786 372698 48022 372934
rect 47786 337018 48022 337254
rect 47786 336698 48022 336934
rect 47786 301018 48022 301254
rect 47786 300698 48022 300934
rect 47786 265018 48022 265254
rect 47786 264698 48022 264934
rect 47786 229018 48022 229254
rect 47786 228698 48022 228934
rect 47786 193018 48022 193254
rect 47786 192698 48022 192934
rect 47786 157018 48022 157254
rect 47786 156698 48022 156934
rect 47786 121018 48022 121254
rect 47786 120698 48022 120934
rect 47786 85018 48022 85254
rect 47786 84698 48022 84934
rect 47786 49018 48022 49254
rect 47786 48698 48022 48934
rect 47786 13018 48022 13254
rect 47786 12698 48022 12934
rect 29786 -7022 30022 -6786
rect 29786 -7342 30022 -7106
rect 54986 705522 55222 705758
rect 54986 705202 55222 705438
rect 54986 668218 55222 668454
rect 54986 667898 55222 668134
rect 54986 632218 55222 632454
rect 54986 631898 55222 632134
rect 54986 596218 55222 596454
rect 54986 595898 55222 596134
rect 54986 560218 55222 560454
rect 54986 559898 55222 560134
rect 54986 524218 55222 524454
rect 54986 523898 55222 524134
rect 54986 488218 55222 488454
rect 54986 487898 55222 488134
rect 54986 452218 55222 452454
rect 54986 451898 55222 452134
rect 54986 416218 55222 416454
rect 54986 415898 55222 416134
rect 54986 380218 55222 380454
rect 54986 379898 55222 380134
rect 54986 344218 55222 344454
rect 54986 343898 55222 344134
rect 54986 308218 55222 308454
rect 54986 307898 55222 308134
rect 54986 272218 55222 272454
rect 54986 271898 55222 272134
rect 54986 236218 55222 236454
rect 54986 235898 55222 236134
rect 54986 200218 55222 200454
rect 54986 199898 55222 200134
rect 54986 164218 55222 164454
rect 54986 163898 55222 164134
rect 54986 128218 55222 128454
rect 54986 127898 55222 128134
rect 54986 92218 55222 92454
rect 54986 91898 55222 92134
rect 54986 56218 55222 56454
rect 54986 55898 55222 56134
rect 54986 20218 55222 20454
rect 54986 19898 55222 20134
rect 54986 -1502 55222 -1266
rect 54986 -1822 55222 -1586
rect 58586 671818 58822 672054
rect 58586 671498 58822 671734
rect 58586 635818 58822 636054
rect 58586 635498 58822 635734
rect 58586 599818 58822 600054
rect 58586 599498 58822 599734
rect 58586 563818 58822 564054
rect 58586 563498 58822 563734
rect 58586 527818 58822 528054
rect 58586 527498 58822 527734
rect 58586 491818 58822 492054
rect 58586 491498 58822 491734
rect 58586 455818 58822 456054
rect 58586 455498 58822 455734
rect 58586 419818 58822 420054
rect 58586 419498 58822 419734
rect 58586 383818 58822 384054
rect 58586 383498 58822 383734
rect 58586 347818 58822 348054
rect 58586 347498 58822 347734
rect 58586 311818 58822 312054
rect 58586 311498 58822 311734
rect 58586 275818 58822 276054
rect 58586 275498 58822 275734
rect 58586 239818 58822 240054
rect 58586 239498 58822 239734
rect 58586 203818 58822 204054
rect 58586 203498 58822 203734
rect 58586 167818 58822 168054
rect 58586 167498 58822 167734
rect 58586 131818 58822 132054
rect 58586 131498 58822 131734
rect 58586 95818 58822 96054
rect 58586 95498 58822 95734
rect 58586 59818 58822 60054
rect 58586 59498 58822 59734
rect 58586 23818 58822 24054
rect 58586 23498 58822 23734
rect 58586 -3342 58822 -3106
rect 58586 -3662 58822 -3426
rect 62186 675418 62422 675654
rect 62186 675098 62422 675334
rect 62186 639418 62422 639654
rect 62186 639098 62422 639334
rect 62186 603418 62422 603654
rect 62186 603098 62422 603334
rect 62186 567418 62422 567654
rect 62186 567098 62422 567334
rect 62186 531418 62422 531654
rect 62186 531098 62422 531334
rect 62186 495418 62422 495654
rect 62186 495098 62422 495334
rect 62186 459418 62422 459654
rect 62186 459098 62422 459334
rect 62186 423418 62422 423654
rect 62186 423098 62422 423334
rect 62186 387418 62422 387654
rect 62186 387098 62422 387334
rect 62186 351418 62422 351654
rect 62186 351098 62422 351334
rect 62186 315418 62422 315654
rect 62186 315098 62422 315334
rect 62186 279418 62422 279654
rect 62186 279098 62422 279334
rect 62186 243418 62422 243654
rect 62186 243098 62422 243334
rect 62186 207418 62422 207654
rect 62186 207098 62422 207334
rect 62186 171418 62422 171654
rect 62186 171098 62422 171334
rect 62186 135418 62422 135654
rect 62186 135098 62422 135334
rect 62186 99418 62422 99654
rect 62186 99098 62422 99334
rect 62186 63418 62422 63654
rect 62186 63098 62422 63334
rect 62186 27418 62422 27654
rect 62186 27098 62422 27334
rect 62186 -5182 62422 -4946
rect 62186 -5502 62422 -5266
rect 83786 710122 84022 710358
rect 83786 709802 84022 710038
rect 80186 708282 80422 708518
rect 80186 707962 80422 708198
rect 76586 706442 76822 706678
rect 76586 706122 76822 706358
rect 65786 679018 66022 679254
rect 65786 678698 66022 678934
rect 65786 643018 66022 643254
rect 65786 642698 66022 642934
rect 65786 607018 66022 607254
rect 65786 606698 66022 606934
rect 65786 571018 66022 571254
rect 65786 570698 66022 570934
rect 65786 535018 66022 535254
rect 65786 534698 66022 534934
rect 65786 499018 66022 499254
rect 65786 498698 66022 498934
rect 65786 463018 66022 463254
rect 65786 462698 66022 462934
rect 65786 427018 66022 427254
rect 65786 426698 66022 426934
rect 65786 391018 66022 391254
rect 65786 390698 66022 390934
rect 65786 355018 66022 355254
rect 65786 354698 66022 354934
rect 65786 319018 66022 319254
rect 65786 318698 66022 318934
rect 65786 283018 66022 283254
rect 65786 282698 66022 282934
rect 65786 247018 66022 247254
rect 65786 246698 66022 246934
rect 65786 211018 66022 211254
rect 65786 210698 66022 210934
rect 65786 175018 66022 175254
rect 65786 174698 66022 174934
rect 65786 139018 66022 139254
rect 65786 138698 66022 138934
rect 65786 103018 66022 103254
rect 65786 102698 66022 102934
rect 65786 67018 66022 67254
rect 65786 66698 66022 66934
rect 65786 31018 66022 31254
rect 65786 30698 66022 30934
rect 47786 -6102 48022 -5866
rect 47786 -6422 48022 -6186
rect 72986 704602 73222 704838
rect 72986 704282 73222 704518
rect 72986 686218 73222 686454
rect 72986 685898 73222 686134
rect 72986 650218 73222 650454
rect 72986 649898 73222 650134
rect 72986 614218 73222 614454
rect 72986 613898 73222 614134
rect 72986 578218 73222 578454
rect 72986 577898 73222 578134
rect 72986 542218 73222 542454
rect 72986 541898 73222 542134
rect 72986 506218 73222 506454
rect 72986 505898 73222 506134
rect 72986 470218 73222 470454
rect 72986 469898 73222 470134
rect 72986 434218 73222 434454
rect 72986 433898 73222 434134
rect 72986 398218 73222 398454
rect 72986 397898 73222 398134
rect 72986 362218 73222 362454
rect 72986 361898 73222 362134
rect 72986 326218 73222 326454
rect 72986 325898 73222 326134
rect 72986 290218 73222 290454
rect 72986 289898 73222 290134
rect 72986 254218 73222 254454
rect 72986 253898 73222 254134
rect 72986 218218 73222 218454
rect 72986 217898 73222 218134
rect 72986 182218 73222 182454
rect 72986 181898 73222 182134
rect 72986 146218 73222 146454
rect 72986 145898 73222 146134
rect 72986 110218 73222 110454
rect 72986 109898 73222 110134
rect 72986 74218 73222 74454
rect 72986 73898 73222 74134
rect 72986 38218 73222 38454
rect 72986 37898 73222 38134
rect 72986 2218 73222 2454
rect 72986 1898 73222 2134
rect 72986 -582 73222 -346
rect 72986 -902 73222 -666
rect 76586 689818 76822 690054
rect 76586 689498 76822 689734
rect 76586 653818 76822 654054
rect 76586 653498 76822 653734
rect 76586 617818 76822 618054
rect 76586 617498 76822 617734
rect 76586 581818 76822 582054
rect 76586 581498 76822 581734
rect 76586 545818 76822 546054
rect 76586 545498 76822 545734
rect 76586 509818 76822 510054
rect 76586 509498 76822 509734
rect 76586 473818 76822 474054
rect 76586 473498 76822 473734
rect 76586 437818 76822 438054
rect 76586 437498 76822 437734
rect 76586 401818 76822 402054
rect 76586 401498 76822 401734
rect 76586 365818 76822 366054
rect 76586 365498 76822 365734
rect 76586 329818 76822 330054
rect 76586 329498 76822 329734
rect 76586 293818 76822 294054
rect 76586 293498 76822 293734
rect 76586 257818 76822 258054
rect 76586 257498 76822 257734
rect 76586 221818 76822 222054
rect 76586 221498 76822 221734
rect 76586 185818 76822 186054
rect 76586 185498 76822 185734
rect 76586 149818 76822 150054
rect 76586 149498 76822 149734
rect 76586 113818 76822 114054
rect 76586 113498 76822 113734
rect 76586 77818 76822 78054
rect 76586 77498 76822 77734
rect 76586 41818 76822 42054
rect 76586 41498 76822 41734
rect 76586 5818 76822 6054
rect 76586 5498 76822 5734
rect 76586 -2422 76822 -2186
rect 76586 -2742 76822 -2506
rect 80186 693418 80422 693654
rect 80186 693098 80422 693334
rect 80186 657418 80422 657654
rect 80186 657098 80422 657334
rect 80186 621418 80422 621654
rect 80186 621098 80422 621334
rect 80186 585418 80422 585654
rect 80186 585098 80422 585334
rect 80186 549418 80422 549654
rect 80186 549098 80422 549334
rect 80186 513418 80422 513654
rect 80186 513098 80422 513334
rect 80186 477418 80422 477654
rect 80186 477098 80422 477334
rect 80186 441418 80422 441654
rect 80186 441098 80422 441334
rect 80186 405418 80422 405654
rect 80186 405098 80422 405334
rect 80186 369418 80422 369654
rect 80186 369098 80422 369334
rect 80186 333418 80422 333654
rect 80186 333098 80422 333334
rect 80186 297418 80422 297654
rect 80186 297098 80422 297334
rect 80186 261418 80422 261654
rect 80186 261098 80422 261334
rect 80186 225418 80422 225654
rect 80186 225098 80422 225334
rect 80186 189418 80422 189654
rect 80186 189098 80422 189334
rect 80186 153418 80422 153654
rect 80186 153098 80422 153334
rect 80186 117418 80422 117654
rect 80186 117098 80422 117334
rect 80186 81418 80422 81654
rect 80186 81098 80422 81334
rect 80186 45418 80422 45654
rect 80186 45098 80422 45334
rect 80186 9418 80422 9654
rect 80186 9098 80422 9334
rect 80186 -4262 80422 -4026
rect 80186 -4582 80422 -4346
rect 101786 711042 102022 711278
rect 101786 710722 102022 710958
rect 98186 709202 98422 709438
rect 98186 708882 98422 709118
rect 94586 707362 94822 707598
rect 94586 707042 94822 707278
rect 83786 697018 84022 697254
rect 83786 696698 84022 696934
rect 83786 661018 84022 661254
rect 83786 660698 84022 660934
rect 83786 625018 84022 625254
rect 83786 624698 84022 624934
rect 83786 589018 84022 589254
rect 83786 588698 84022 588934
rect 83786 553018 84022 553254
rect 83786 552698 84022 552934
rect 83786 517018 84022 517254
rect 83786 516698 84022 516934
rect 83786 481018 84022 481254
rect 83786 480698 84022 480934
rect 83786 445018 84022 445254
rect 83786 444698 84022 444934
rect 83786 409018 84022 409254
rect 83786 408698 84022 408934
rect 83786 373018 84022 373254
rect 83786 372698 84022 372934
rect 83786 337018 84022 337254
rect 83786 336698 84022 336934
rect 83786 301018 84022 301254
rect 83786 300698 84022 300934
rect 83786 265018 84022 265254
rect 83786 264698 84022 264934
rect 83786 229018 84022 229254
rect 83786 228698 84022 228934
rect 83786 193018 84022 193254
rect 83786 192698 84022 192934
rect 83786 157018 84022 157254
rect 83786 156698 84022 156934
rect 83786 121018 84022 121254
rect 83786 120698 84022 120934
rect 83786 85018 84022 85254
rect 83786 84698 84022 84934
rect 83786 49018 84022 49254
rect 83786 48698 84022 48934
rect 83786 13018 84022 13254
rect 83786 12698 84022 12934
rect 65786 -7022 66022 -6786
rect 65786 -7342 66022 -7106
rect 90986 705522 91222 705758
rect 90986 705202 91222 705438
rect 90986 668218 91222 668454
rect 90986 667898 91222 668134
rect 90986 632218 91222 632454
rect 90986 631898 91222 632134
rect 90986 596218 91222 596454
rect 90986 595898 91222 596134
rect 90986 560218 91222 560454
rect 90986 559898 91222 560134
rect 90986 524218 91222 524454
rect 90986 523898 91222 524134
rect 90986 488218 91222 488454
rect 90986 487898 91222 488134
rect 90986 452218 91222 452454
rect 90986 451898 91222 452134
rect 90986 416218 91222 416454
rect 90986 415898 91222 416134
rect 90986 380218 91222 380454
rect 90986 379898 91222 380134
rect 90986 344218 91222 344454
rect 90986 343898 91222 344134
rect 90986 308218 91222 308454
rect 90986 307898 91222 308134
rect 90986 272218 91222 272454
rect 90986 271898 91222 272134
rect 90986 236218 91222 236454
rect 90986 235898 91222 236134
rect 90986 200218 91222 200454
rect 90986 199898 91222 200134
rect 90986 164218 91222 164454
rect 90986 163898 91222 164134
rect 90986 128218 91222 128454
rect 90986 127898 91222 128134
rect 90986 92218 91222 92454
rect 90986 91898 91222 92134
rect 90986 56218 91222 56454
rect 90986 55898 91222 56134
rect 90986 20218 91222 20454
rect 90986 19898 91222 20134
rect 90986 -1502 91222 -1266
rect 90986 -1822 91222 -1586
rect 94586 671818 94822 672054
rect 94586 671498 94822 671734
rect 94586 635818 94822 636054
rect 94586 635498 94822 635734
rect 94586 599818 94822 600054
rect 94586 599498 94822 599734
rect 94586 563818 94822 564054
rect 94586 563498 94822 563734
rect 94586 527818 94822 528054
rect 94586 527498 94822 527734
rect 94586 491818 94822 492054
rect 94586 491498 94822 491734
rect 94586 455818 94822 456054
rect 94586 455498 94822 455734
rect 94586 419818 94822 420054
rect 94586 419498 94822 419734
rect 94586 383818 94822 384054
rect 94586 383498 94822 383734
rect 94586 347818 94822 348054
rect 94586 347498 94822 347734
rect 94586 311818 94822 312054
rect 94586 311498 94822 311734
rect 94586 275818 94822 276054
rect 94586 275498 94822 275734
rect 94586 239818 94822 240054
rect 94586 239498 94822 239734
rect 94586 203818 94822 204054
rect 94586 203498 94822 203734
rect 94586 167818 94822 168054
rect 94586 167498 94822 167734
rect 94586 131818 94822 132054
rect 94586 131498 94822 131734
rect 94586 95818 94822 96054
rect 94586 95498 94822 95734
rect 94586 59818 94822 60054
rect 94586 59498 94822 59734
rect 94586 23818 94822 24054
rect 94586 23498 94822 23734
rect 94586 -3342 94822 -3106
rect 94586 -3662 94822 -3426
rect 98186 675418 98422 675654
rect 98186 675098 98422 675334
rect 98186 639418 98422 639654
rect 98186 639098 98422 639334
rect 98186 603418 98422 603654
rect 98186 603098 98422 603334
rect 98186 567418 98422 567654
rect 98186 567098 98422 567334
rect 98186 531418 98422 531654
rect 98186 531098 98422 531334
rect 98186 495418 98422 495654
rect 98186 495098 98422 495334
rect 98186 459418 98422 459654
rect 98186 459098 98422 459334
rect 98186 423418 98422 423654
rect 98186 423098 98422 423334
rect 98186 387418 98422 387654
rect 98186 387098 98422 387334
rect 98186 351418 98422 351654
rect 98186 351098 98422 351334
rect 98186 315418 98422 315654
rect 98186 315098 98422 315334
rect 98186 279418 98422 279654
rect 98186 279098 98422 279334
rect 98186 243418 98422 243654
rect 98186 243098 98422 243334
rect 98186 207418 98422 207654
rect 98186 207098 98422 207334
rect 98186 171418 98422 171654
rect 98186 171098 98422 171334
rect 98186 135418 98422 135654
rect 98186 135098 98422 135334
rect 98186 99418 98422 99654
rect 98186 99098 98422 99334
rect 98186 63418 98422 63654
rect 98186 63098 98422 63334
rect 98186 27418 98422 27654
rect 98186 27098 98422 27334
rect 98186 -5182 98422 -4946
rect 98186 -5502 98422 -5266
rect 119786 710122 120022 710358
rect 119786 709802 120022 710038
rect 116186 708282 116422 708518
rect 116186 707962 116422 708198
rect 112586 706442 112822 706678
rect 112586 706122 112822 706358
rect 101786 679018 102022 679254
rect 101786 678698 102022 678934
rect 101786 643018 102022 643254
rect 101786 642698 102022 642934
rect 101786 607018 102022 607254
rect 101786 606698 102022 606934
rect 101786 571018 102022 571254
rect 101786 570698 102022 570934
rect 101786 535018 102022 535254
rect 101786 534698 102022 534934
rect 101786 499018 102022 499254
rect 101786 498698 102022 498934
rect 101786 463018 102022 463254
rect 101786 462698 102022 462934
rect 101786 427018 102022 427254
rect 101786 426698 102022 426934
rect 101786 391018 102022 391254
rect 101786 390698 102022 390934
rect 101786 355018 102022 355254
rect 101786 354698 102022 354934
rect 101786 319018 102022 319254
rect 101786 318698 102022 318934
rect 101786 283018 102022 283254
rect 101786 282698 102022 282934
rect 101786 247018 102022 247254
rect 101786 246698 102022 246934
rect 101786 211018 102022 211254
rect 101786 210698 102022 210934
rect 101786 175018 102022 175254
rect 101786 174698 102022 174934
rect 101786 139018 102022 139254
rect 101786 138698 102022 138934
rect 101786 103018 102022 103254
rect 101786 102698 102022 102934
rect 101786 67018 102022 67254
rect 101786 66698 102022 66934
rect 101786 31018 102022 31254
rect 101786 30698 102022 30934
rect 83786 -6102 84022 -5866
rect 83786 -6422 84022 -6186
rect 108986 704602 109222 704838
rect 108986 704282 109222 704518
rect 108986 686218 109222 686454
rect 108986 685898 109222 686134
rect 108986 650218 109222 650454
rect 108986 649898 109222 650134
rect 108986 614218 109222 614454
rect 108986 613898 109222 614134
rect 108986 578218 109222 578454
rect 108986 577898 109222 578134
rect 108986 542218 109222 542454
rect 108986 541898 109222 542134
rect 108986 506218 109222 506454
rect 108986 505898 109222 506134
rect 108986 470218 109222 470454
rect 108986 469898 109222 470134
rect 108986 434218 109222 434454
rect 108986 433898 109222 434134
rect 108986 398218 109222 398454
rect 108986 397898 109222 398134
rect 108986 362218 109222 362454
rect 108986 361898 109222 362134
rect 108986 326218 109222 326454
rect 108986 325898 109222 326134
rect 108986 290218 109222 290454
rect 108986 289898 109222 290134
rect 108986 254218 109222 254454
rect 108986 253898 109222 254134
rect 108986 218218 109222 218454
rect 108986 217898 109222 218134
rect 108986 182218 109222 182454
rect 108986 181898 109222 182134
rect 108986 146218 109222 146454
rect 108986 145898 109222 146134
rect 108986 110218 109222 110454
rect 108986 109898 109222 110134
rect 108986 74218 109222 74454
rect 108986 73898 109222 74134
rect 108986 38218 109222 38454
rect 108986 37898 109222 38134
rect 108986 2218 109222 2454
rect 108986 1898 109222 2134
rect 108986 -582 109222 -346
rect 108986 -902 109222 -666
rect 112586 689818 112822 690054
rect 112586 689498 112822 689734
rect 112586 653818 112822 654054
rect 112586 653498 112822 653734
rect 112586 617818 112822 618054
rect 112586 617498 112822 617734
rect 112586 581818 112822 582054
rect 112586 581498 112822 581734
rect 112586 545818 112822 546054
rect 112586 545498 112822 545734
rect 112586 509818 112822 510054
rect 112586 509498 112822 509734
rect 112586 473818 112822 474054
rect 112586 473498 112822 473734
rect 112586 437818 112822 438054
rect 112586 437498 112822 437734
rect 112586 401818 112822 402054
rect 112586 401498 112822 401734
rect 112586 365818 112822 366054
rect 112586 365498 112822 365734
rect 112586 329818 112822 330054
rect 112586 329498 112822 329734
rect 112586 293818 112822 294054
rect 112586 293498 112822 293734
rect 112586 257818 112822 258054
rect 112586 257498 112822 257734
rect 112586 221818 112822 222054
rect 112586 221498 112822 221734
rect 112586 185818 112822 186054
rect 112586 185498 112822 185734
rect 112586 149818 112822 150054
rect 112586 149498 112822 149734
rect 112586 113818 112822 114054
rect 112586 113498 112822 113734
rect 112586 77818 112822 78054
rect 112586 77498 112822 77734
rect 112586 41818 112822 42054
rect 112586 41498 112822 41734
rect 112586 5818 112822 6054
rect 112586 5498 112822 5734
rect 112586 -2422 112822 -2186
rect 112586 -2742 112822 -2506
rect 116186 693418 116422 693654
rect 116186 693098 116422 693334
rect 116186 657418 116422 657654
rect 116186 657098 116422 657334
rect 116186 621418 116422 621654
rect 116186 621098 116422 621334
rect 116186 585418 116422 585654
rect 116186 585098 116422 585334
rect 116186 549418 116422 549654
rect 116186 549098 116422 549334
rect 116186 513418 116422 513654
rect 116186 513098 116422 513334
rect 116186 477418 116422 477654
rect 116186 477098 116422 477334
rect 116186 441418 116422 441654
rect 116186 441098 116422 441334
rect 116186 405418 116422 405654
rect 116186 405098 116422 405334
rect 116186 369418 116422 369654
rect 116186 369098 116422 369334
rect 116186 333418 116422 333654
rect 116186 333098 116422 333334
rect 116186 297418 116422 297654
rect 116186 297098 116422 297334
rect 116186 261418 116422 261654
rect 116186 261098 116422 261334
rect 116186 225418 116422 225654
rect 116186 225098 116422 225334
rect 116186 189418 116422 189654
rect 116186 189098 116422 189334
rect 116186 153418 116422 153654
rect 116186 153098 116422 153334
rect 116186 117418 116422 117654
rect 116186 117098 116422 117334
rect 116186 81418 116422 81654
rect 116186 81098 116422 81334
rect 116186 45418 116422 45654
rect 116186 45098 116422 45334
rect 116186 9418 116422 9654
rect 116186 9098 116422 9334
rect 116186 -4262 116422 -4026
rect 116186 -4582 116422 -4346
rect 137786 711042 138022 711278
rect 137786 710722 138022 710958
rect 134186 709202 134422 709438
rect 134186 708882 134422 709118
rect 130586 707362 130822 707598
rect 130586 707042 130822 707278
rect 119786 697018 120022 697254
rect 119786 696698 120022 696934
rect 119786 661018 120022 661254
rect 119786 660698 120022 660934
rect 119786 625018 120022 625254
rect 119786 624698 120022 624934
rect 119786 589018 120022 589254
rect 119786 588698 120022 588934
rect 119786 553018 120022 553254
rect 119786 552698 120022 552934
rect 119786 517018 120022 517254
rect 119786 516698 120022 516934
rect 119786 481018 120022 481254
rect 119786 480698 120022 480934
rect 119786 445018 120022 445254
rect 119786 444698 120022 444934
rect 119786 409018 120022 409254
rect 119786 408698 120022 408934
rect 119786 373018 120022 373254
rect 119786 372698 120022 372934
rect 119786 337018 120022 337254
rect 119786 336698 120022 336934
rect 119786 301018 120022 301254
rect 119786 300698 120022 300934
rect 119786 265018 120022 265254
rect 119786 264698 120022 264934
rect 119786 229018 120022 229254
rect 119786 228698 120022 228934
rect 119786 193018 120022 193254
rect 119786 192698 120022 192934
rect 119786 157018 120022 157254
rect 119786 156698 120022 156934
rect 119786 121018 120022 121254
rect 119786 120698 120022 120934
rect 119786 85018 120022 85254
rect 119786 84698 120022 84934
rect 119786 49018 120022 49254
rect 119786 48698 120022 48934
rect 119786 13018 120022 13254
rect 119786 12698 120022 12934
rect 101786 -7022 102022 -6786
rect 101786 -7342 102022 -7106
rect 126986 705522 127222 705758
rect 126986 705202 127222 705438
rect 126986 668218 127222 668454
rect 126986 667898 127222 668134
rect 126986 632218 127222 632454
rect 126986 631898 127222 632134
rect 126986 596218 127222 596454
rect 126986 595898 127222 596134
rect 126986 560218 127222 560454
rect 126986 559898 127222 560134
rect 126986 524218 127222 524454
rect 126986 523898 127222 524134
rect 126986 488218 127222 488454
rect 126986 487898 127222 488134
rect 126986 452218 127222 452454
rect 126986 451898 127222 452134
rect 126986 416218 127222 416454
rect 126986 415898 127222 416134
rect 126986 380218 127222 380454
rect 126986 379898 127222 380134
rect 126986 344218 127222 344454
rect 126986 343898 127222 344134
rect 126986 308218 127222 308454
rect 126986 307898 127222 308134
rect 126986 272218 127222 272454
rect 126986 271898 127222 272134
rect 126986 236218 127222 236454
rect 126986 235898 127222 236134
rect 126986 200218 127222 200454
rect 126986 199898 127222 200134
rect 126986 164218 127222 164454
rect 126986 163898 127222 164134
rect 126986 128218 127222 128454
rect 126986 127898 127222 128134
rect 126986 92218 127222 92454
rect 126986 91898 127222 92134
rect 126986 56218 127222 56454
rect 126986 55898 127222 56134
rect 126986 20218 127222 20454
rect 126986 19898 127222 20134
rect 126986 -1502 127222 -1266
rect 126986 -1822 127222 -1586
rect 130586 671818 130822 672054
rect 130586 671498 130822 671734
rect 130586 635818 130822 636054
rect 130586 635498 130822 635734
rect 130586 599818 130822 600054
rect 130586 599498 130822 599734
rect 130586 563818 130822 564054
rect 130586 563498 130822 563734
rect 130586 527818 130822 528054
rect 130586 527498 130822 527734
rect 130586 491818 130822 492054
rect 130586 491498 130822 491734
rect 130586 455818 130822 456054
rect 130586 455498 130822 455734
rect 130586 419818 130822 420054
rect 130586 419498 130822 419734
rect 130586 383818 130822 384054
rect 130586 383498 130822 383734
rect 130586 347818 130822 348054
rect 130586 347498 130822 347734
rect 130586 311818 130822 312054
rect 130586 311498 130822 311734
rect 130586 275818 130822 276054
rect 130586 275498 130822 275734
rect 130586 239818 130822 240054
rect 130586 239498 130822 239734
rect 130586 203818 130822 204054
rect 130586 203498 130822 203734
rect 130586 167818 130822 168054
rect 130586 167498 130822 167734
rect 130586 131818 130822 132054
rect 130586 131498 130822 131734
rect 130586 95818 130822 96054
rect 130586 95498 130822 95734
rect 130586 59818 130822 60054
rect 130586 59498 130822 59734
rect 130586 23818 130822 24054
rect 130586 23498 130822 23734
rect 130586 -3342 130822 -3106
rect 130586 -3662 130822 -3426
rect 134186 675418 134422 675654
rect 134186 675098 134422 675334
rect 134186 639418 134422 639654
rect 134186 639098 134422 639334
rect 134186 603418 134422 603654
rect 134186 603098 134422 603334
rect 134186 567418 134422 567654
rect 134186 567098 134422 567334
rect 134186 531418 134422 531654
rect 134186 531098 134422 531334
rect 134186 495418 134422 495654
rect 134186 495098 134422 495334
rect 134186 459418 134422 459654
rect 134186 459098 134422 459334
rect 134186 423418 134422 423654
rect 134186 423098 134422 423334
rect 134186 387418 134422 387654
rect 134186 387098 134422 387334
rect 134186 351418 134422 351654
rect 134186 351098 134422 351334
rect 134186 315418 134422 315654
rect 134186 315098 134422 315334
rect 134186 279418 134422 279654
rect 134186 279098 134422 279334
rect 134186 243418 134422 243654
rect 134186 243098 134422 243334
rect 134186 207418 134422 207654
rect 134186 207098 134422 207334
rect 134186 171418 134422 171654
rect 134186 171098 134422 171334
rect 134186 135418 134422 135654
rect 134186 135098 134422 135334
rect 134186 99418 134422 99654
rect 134186 99098 134422 99334
rect 134186 63418 134422 63654
rect 134186 63098 134422 63334
rect 134186 27418 134422 27654
rect 134186 27098 134422 27334
rect 134186 -5182 134422 -4946
rect 134186 -5502 134422 -5266
rect 155786 710122 156022 710358
rect 155786 709802 156022 710038
rect 152186 708282 152422 708518
rect 152186 707962 152422 708198
rect 148586 706442 148822 706678
rect 148586 706122 148822 706358
rect 137786 679018 138022 679254
rect 137786 678698 138022 678934
rect 137786 643018 138022 643254
rect 137786 642698 138022 642934
rect 137786 607018 138022 607254
rect 137786 606698 138022 606934
rect 137786 571018 138022 571254
rect 137786 570698 138022 570934
rect 137786 535018 138022 535254
rect 137786 534698 138022 534934
rect 137786 499018 138022 499254
rect 137786 498698 138022 498934
rect 137786 463018 138022 463254
rect 137786 462698 138022 462934
rect 137786 427018 138022 427254
rect 137786 426698 138022 426934
rect 137786 391018 138022 391254
rect 137786 390698 138022 390934
rect 137786 355018 138022 355254
rect 137786 354698 138022 354934
rect 137786 319018 138022 319254
rect 137786 318698 138022 318934
rect 137786 283018 138022 283254
rect 137786 282698 138022 282934
rect 137786 247018 138022 247254
rect 137786 246698 138022 246934
rect 137786 211018 138022 211254
rect 137786 210698 138022 210934
rect 137786 175018 138022 175254
rect 137786 174698 138022 174934
rect 137786 139018 138022 139254
rect 137786 138698 138022 138934
rect 137786 103018 138022 103254
rect 137786 102698 138022 102934
rect 137786 67018 138022 67254
rect 137786 66698 138022 66934
rect 137786 31018 138022 31254
rect 137786 30698 138022 30934
rect 119786 -6102 120022 -5866
rect 119786 -6422 120022 -6186
rect 144986 704602 145222 704838
rect 144986 704282 145222 704518
rect 144986 686218 145222 686454
rect 144986 685898 145222 686134
rect 144986 650218 145222 650454
rect 144986 649898 145222 650134
rect 144986 614218 145222 614454
rect 144986 613898 145222 614134
rect 144986 578218 145222 578454
rect 144986 577898 145222 578134
rect 144986 542218 145222 542454
rect 144986 541898 145222 542134
rect 144986 506218 145222 506454
rect 144986 505898 145222 506134
rect 144986 470218 145222 470454
rect 144986 469898 145222 470134
rect 144986 434218 145222 434454
rect 144986 433898 145222 434134
rect 144986 398218 145222 398454
rect 144986 397898 145222 398134
rect 144986 362218 145222 362454
rect 144986 361898 145222 362134
rect 144986 326218 145222 326454
rect 144986 325898 145222 326134
rect 144986 290218 145222 290454
rect 144986 289898 145222 290134
rect 144986 254218 145222 254454
rect 144986 253898 145222 254134
rect 144986 218218 145222 218454
rect 144986 217898 145222 218134
rect 144986 182218 145222 182454
rect 144986 181898 145222 182134
rect 144986 146218 145222 146454
rect 144986 145898 145222 146134
rect 144986 110218 145222 110454
rect 144986 109898 145222 110134
rect 144986 74218 145222 74454
rect 144986 73898 145222 74134
rect 144986 38218 145222 38454
rect 144986 37898 145222 38134
rect 144986 2218 145222 2454
rect 144986 1898 145222 2134
rect 144986 -582 145222 -346
rect 144986 -902 145222 -666
rect 148586 689818 148822 690054
rect 148586 689498 148822 689734
rect 148586 653818 148822 654054
rect 148586 653498 148822 653734
rect 148586 617818 148822 618054
rect 148586 617498 148822 617734
rect 148586 581818 148822 582054
rect 148586 581498 148822 581734
rect 148586 545818 148822 546054
rect 148586 545498 148822 545734
rect 148586 509818 148822 510054
rect 148586 509498 148822 509734
rect 148586 473818 148822 474054
rect 148586 473498 148822 473734
rect 148586 437818 148822 438054
rect 148586 437498 148822 437734
rect 148586 401818 148822 402054
rect 148586 401498 148822 401734
rect 148586 365818 148822 366054
rect 148586 365498 148822 365734
rect 148586 329818 148822 330054
rect 148586 329498 148822 329734
rect 148586 293818 148822 294054
rect 148586 293498 148822 293734
rect 148586 257818 148822 258054
rect 148586 257498 148822 257734
rect 148586 221818 148822 222054
rect 148586 221498 148822 221734
rect 148586 185818 148822 186054
rect 148586 185498 148822 185734
rect 148586 149818 148822 150054
rect 148586 149498 148822 149734
rect 148586 113818 148822 114054
rect 148586 113498 148822 113734
rect 148586 77818 148822 78054
rect 148586 77498 148822 77734
rect 148586 41818 148822 42054
rect 148586 41498 148822 41734
rect 148586 5818 148822 6054
rect 148586 5498 148822 5734
rect 148586 -2422 148822 -2186
rect 148586 -2742 148822 -2506
rect 152186 693418 152422 693654
rect 152186 693098 152422 693334
rect 152186 657418 152422 657654
rect 152186 657098 152422 657334
rect 152186 621418 152422 621654
rect 152186 621098 152422 621334
rect 152186 585418 152422 585654
rect 152186 585098 152422 585334
rect 152186 549418 152422 549654
rect 152186 549098 152422 549334
rect 152186 513418 152422 513654
rect 152186 513098 152422 513334
rect 152186 477418 152422 477654
rect 152186 477098 152422 477334
rect 152186 441418 152422 441654
rect 152186 441098 152422 441334
rect 152186 405418 152422 405654
rect 152186 405098 152422 405334
rect 152186 369418 152422 369654
rect 152186 369098 152422 369334
rect 152186 333418 152422 333654
rect 152186 333098 152422 333334
rect 152186 297418 152422 297654
rect 152186 297098 152422 297334
rect 152186 261418 152422 261654
rect 152186 261098 152422 261334
rect 152186 225418 152422 225654
rect 152186 225098 152422 225334
rect 152186 189418 152422 189654
rect 152186 189098 152422 189334
rect 152186 153418 152422 153654
rect 152186 153098 152422 153334
rect 152186 117418 152422 117654
rect 152186 117098 152422 117334
rect 152186 81418 152422 81654
rect 152186 81098 152422 81334
rect 152186 45418 152422 45654
rect 152186 45098 152422 45334
rect 152186 9418 152422 9654
rect 152186 9098 152422 9334
rect 152186 -4262 152422 -4026
rect 152186 -4582 152422 -4346
rect 173786 711042 174022 711278
rect 173786 710722 174022 710958
rect 170186 709202 170422 709438
rect 170186 708882 170422 709118
rect 166586 707362 166822 707598
rect 166586 707042 166822 707278
rect 155786 697018 156022 697254
rect 155786 696698 156022 696934
rect 155786 661018 156022 661254
rect 155786 660698 156022 660934
rect 155786 625018 156022 625254
rect 155786 624698 156022 624934
rect 155786 589018 156022 589254
rect 155786 588698 156022 588934
rect 155786 553018 156022 553254
rect 155786 552698 156022 552934
rect 155786 517018 156022 517254
rect 155786 516698 156022 516934
rect 155786 481018 156022 481254
rect 155786 480698 156022 480934
rect 155786 445018 156022 445254
rect 155786 444698 156022 444934
rect 155786 409018 156022 409254
rect 155786 408698 156022 408934
rect 155786 373018 156022 373254
rect 155786 372698 156022 372934
rect 155786 337018 156022 337254
rect 155786 336698 156022 336934
rect 155786 301018 156022 301254
rect 155786 300698 156022 300934
rect 155786 265018 156022 265254
rect 155786 264698 156022 264934
rect 155786 229018 156022 229254
rect 155786 228698 156022 228934
rect 155786 193018 156022 193254
rect 155786 192698 156022 192934
rect 155786 157018 156022 157254
rect 155786 156698 156022 156934
rect 155786 121018 156022 121254
rect 155786 120698 156022 120934
rect 155786 85018 156022 85254
rect 155786 84698 156022 84934
rect 155786 49018 156022 49254
rect 155786 48698 156022 48934
rect 155786 13018 156022 13254
rect 155786 12698 156022 12934
rect 137786 -7022 138022 -6786
rect 137786 -7342 138022 -7106
rect 162986 705522 163222 705758
rect 162986 705202 163222 705438
rect 162986 668218 163222 668454
rect 162986 667898 163222 668134
rect 162986 632218 163222 632454
rect 162986 631898 163222 632134
rect 162986 596218 163222 596454
rect 162986 595898 163222 596134
rect 162986 560218 163222 560454
rect 162986 559898 163222 560134
rect 162986 524218 163222 524454
rect 162986 523898 163222 524134
rect 162986 488218 163222 488454
rect 162986 487898 163222 488134
rect 162986 452218 163222 452454
rect 162986 451898 163222 452134
rect 162986 416218 163222 416454
rect 162986 415898 163222 416134
rect 162986 380218 163222 380454
rect 162986 379898 163222 380134
rect 162986 344218 163222 344454
rect 162986 343898 163222 344134
rect 162986 308218 163222 308454
rect 162986 307898 163222 308134
rect 162986 272218 163222 272454
rect 162986 271898 163222 272134
rect 162986 236218 163222 236454
rect 162986 235898 163222 236134
rect 162986 200218 163222 200454
rect 162986 199898 163222 200134
rect 162986 164218 163222 164454
rect 162986 163898 163222 164134
rect 162986 128218 163222 128454
rect 162986 127898 163222 128134
rect 162986 92218 163222 92454
rect 162986 91898 163222 92134
rect 162986 56218 163222 56454
rect 162986 55898 163222 56134
rect 162986 20218 163222 20454
rect 162986 19898 163222 20134
rect 162986 -1502 163222 -1266
rect 162986 -1822 163222 -1586
rect 166586 671818 166822 672054
rect 166586 671498 166822 671734
rect 166586 635818 166822 636054
rect 166586 635498 166822 635734
rect 166586 599818 166822 600054
rect 166586 599498 166822 599734
rect 166586 563818 166822 564054
rect 166586 563498 166822 563734
rect 166586 527818 166822 528054
rect 166586 527498 166822 527734
rect 166586 491818 166822 492054
rect 166586 491498 166822 491734
rect 166586 455818 166822 456054
rect 166586 455498 166822 455734
rect 166586 419818 166822 420054
rect 166586 419498 166822 419734
rect 166586 383818 166822 384054
rect 166586 383498 166822 383734
rect 166586 347818 166822 348054
rect 166586 347498 166822 347734
rect 166586 311818 166822 312054
rect 166586 311498 166822 311734
rect 166586 275818 166822 276054
rect 166586 275498 166822 275734
rect 166586 239818 166822 240054
rect 166586 239498 166822 239734
rect 166586 203818 166822 204054
rect 166586 203498 166822 203734
rect 166586 167818 166822 168054
rect 166586 167498 166822 167734
rect 166586 131818 166822 132054
rect 166586 131498 166822 131734
rect 166586 95818 166822 96054
rect 166586 95498 166822 95734
rect 166586 59818 166822 60054
rect 166586 59498 166822 59734
rect 166586 23818 166822 24054
rect 166586 23498 166822 23734
rect 166586 -3342 166822 -3106
rect 166586 -3662 166822 -3426
rect 170186 675418 170422 675654
rect 170186 675098 170422 675334
rect 170186 639418 170422 639654
rect 170186 639098 170422 639334
rect 170186 603418 170422 603654
rect 170186 603098 170422 603334
rect 170186 567418 170422 567654
rect 170186 567098 170422 567334
rect 170186 531418 170422 531654
rect 170186 531098 170422 531334
rect 170186 495418 170422 495654
rect 170186 495098 170422 495334
rect 170186 459418 170422 459654
rect 170186 459098 170422 459334
rect 170186 423418 170422 423654
rect 170186 423098 170422 423334
rect 170186 387418 170422 387654
rect 170186 387098 170422 387334
rect 170186 351418 170422 351654
rect 170186 351098 170422 351334
rect 170186 315418 170422 315654
rect 170186 315098 170422 315334
rect 170186 279418 170422 279654
rect 170186 279098 170422 279334
rect 170186 243418 170422 243654
rect 170186 243098 170422 243334
rect 170186 207418 170422 207654
rect 170186 207098 170422 207334
rect 170186 171418 170422 171654
rect 170186 171098 170422 171334
rect 170186 135418 170422 135654
rect 170186 135098 170422 135334
rect 170186 99418 170422 99654
rect 170186 99098 170422 99334
rect 170186 63418 170422 63654
rect 170186 63098 170422 63334
rect 170186 27418 170422 27654
rect 170186 27098 170422 27334
rect 170186 -5182 170422 -4946
rect 170186 -5502 170422 -5266
rect 191786 710122 192022 710358
rect 191786 709802 192022 710038
rect 188186 708282 188422 708518
rect 188186 707962 188422 708198
rect 184586 706442 184822 706678
rect 184586 706122 184822 706358
rect 173786 679018 174022 679254
rect 173786 678698 174022 678934
rect 173786 643018 174022 643254
rect 173786 642698 174022 642934
rect 173786 607018 174022 607254
rect 173786 606698 174022 606934
rect 173786 571018 174022 571254
rect 173786 570698 174022 570934
rect 173786 535018 174022 535254
rect 173786 534698 174022 534934
rect 173786 499018 174022 499254
rect 173786 498698 174022 498934
rect 173786 463018 174022 463254
rect 173786 462698 174022 462934
rect 173786 427018 174022 427254
rect 173786 426698 174022 426934
rect 173786 391018 174022 391254
rect 173786 390698 174022 390934
rect 173786 355018 174022 355254
rect 173786 354698 174022 354934
rect 173786 319018 174022 319254
rect 173786 318698 174022 318934
rect 173786 283018 174022 283254
rect 173786 282698 174022 282934
rect 173786 247018 174022 247254
rect 173786 246698 174022 246934
rect 173786 211018 174022 211254
rect 173786 210698 174022 210934
rect 173786 175018 174022 175254
rect 173786 174698 174022 174934
rect 173786 139018 174022 139254
rect 173786 138698 174022 138934
rect 173786 103018 174022 103254
rect 173786 102698 174022 102934
rect 173786 67018 174022 67254
rect 173786 66698 174022 66934
rect 173786 31018 174022 31254
rect 173786 30698 174022 30934
rect 155786 -6102 156022 -5866
rect 155786 -6422 156022 -6186
rect 180986 704602 181222 704838
rect 180986 704282 181222 704518
rect 180986 686218 181222 686454
rect 180986 685898 181222 686134
rect 180986 650218 181222 650454
rect 180986 649898 181222 650134
rect 180986 614218 181222 614454
rect 180986 613898 181222 614134
rect 180986 578218 181222 578454
rect 180986 577898 181222 578134
rect 180986 542218 181222 542454
rect 180986 541898 181222 542134
rect 180986 506218 181222 506454
rect 180986 505898 181222 506134
rect 180986 470218 181222 470454
rect 180986 469898 181222 470134
rect 180986 434218 181222 434454
rect 180986 433898 181222 434134
rect 180986 398218 181222 398454
rect 180986 397898 181222 398134
rect 180986 362218 181222 362454
rect 180986 361898 181222 362134
rect 180986 326218 181222 326454
rect 180986 325898 181222 326134
rect 180986 290218 181222 290454
rect 180986 289898 181222 290134
rect 180986 254218 181222 254454
rect 180986 253898 181222 254134
rect 180986 218218 181222 218454
rect 180986 217898 181222 218134
rect 180986 182218 181222 182454
rect 180986 181898 181222 182134
rect 180986 146218 181222 146454
rect 180986 145898 181222 146134
rect 180986 110218 181222 110454
rect 180986 109898 181222 110134
rect 180986 74218 181222 74454
rect 180986 73898 181222 74134
rect 180986 38218 181222 38454
rect 180986 37898 181222 38134
rect 180986 2218 181222 2454
rect 180986 1898 181222 2134
rect 180986 -582 181222 -346
rect 180986 -902 181222 -666
rect 184586 689818 184822 690054
rect 184586 689498 184822 689734
rect 184586 653818 184822 654054
rect 184586 653498 184822 653734
rect 184586 617818 184822 618054
rect 184586 617498 184822 617734
rect 184586 581818 184822 582054
rect 184586 581498 184822 581734
rect 184586 545818 184822 546054
rect 184586 545498 184822 545734
rect 184586 509818 184822 510054
rect 184586 509498 184822 509734
rect 184586 473818 184822 474054
rect 184586 473498 184822 473734
rect 184586 437818 184822 438054
rect 184586 437498 184822 437734
rect 184586 401818 184822 402054
rect 184586 401498 184822 401734
rect 184586 365818 184822 366054
rect 184586 365498 184822 365734
rect 184586 329818 184822 330054
rect 184586 329498 184822 329734
rect 184586 293818 184822 294054
rect 184586 293498 184822 293734
rect 184586 257818 184822 258054
rect 184586 257498 184822 257734
rect 184586 221818 184822 222054
rect 184586 221498 184822 221734
rect 184586 185818 184822 186054
rect 184586 185498 184822 185734
rect 184586 149818 184822 150054
rect 184586 149498 184822 149734
rect 184586 113818 184822 114054
rect 184586 113498 184822 113734
rect 184586 77818 184822 78054
rect 184586 77498 184822 77734
rect 184586 41818 184822 42054
rect 184586 41498 184822 41734
rect 184586 5818 184822 6054
rect 184586 5498 184822 5734
rect 184586 -2422 184822 -2186
rect 184586 -2742 184822 -2506
rect 188186 693418 188422 693654
rect 188186 693098 188422 693334
rect 188186 657418 188422 657654
rect 188186 657098 188422 657334
rect 188186 621418 188422 621654
rect 188186 621098 188422 621334
rect 188186 585418 188422 585654
rect 188186 585098 188422 585334
rect 188186 549418 188422 549654
rect 188186 549098 188422 549334
rect 188186 513418 188422 513654
rect 188186 513098 188422 513334
rect 188186 477418 188422 477654
rect 188186 477098 188422 477334
rect 188186 441418 188422 441654
rect 188186 441098 188422 441334
rect 188186 405418 188422 405654
rect 188186 405098 188422 405334
rect 188186 369418 188422 369654
rect 188186 369098 188422 369334
rect 188186 333418 188422 333654
rect 188186 333098 188422 333334
rect 188186 297418 188422 297654
rect 188186 297098 188422 297334
rect 188186 261418 188422 261654
rect 188186 261098 188422 261334
rect 188186 225418 188422 225654
rect 188186 225098 188422 225334
rect 188186 189418 188422 189654
rect 188186 189098 188422 189334
rect 188186 153418 188422 153654
rect 188186 153098 188422 153334
rect 188186 117418 188422 117654
rect 188186 117098 188422 117334
rect 188186 81418 188422 81654
rect 188186 81098 188422 81334
rect 188186 45418 188422 45654
rect 188186 45098 188422 45334
rect 188186 9418 188422 9654
rect 188186 9098 188422 9334
rect 188186 -4262 188422 -4026
rect 188186 -4582 188422 -4346
rect 209786 711042 210022 711278
rect 209786 710722 210022 710958
rect 206186 709202 206422 709438
rect 206186 708882 206422 709118
rect 202586 707362 202822 707598
rect 202586 707042 202822 707278
rect 191786 697018 192022 697254
rect 191786 696698 192022 696934
rect 191786 661018 192022 661254
rect 191786 660698 192022 660934
rect 191786 625018 192022 625254
rect 191786 624698 192022 624934
rect 191786 589018 192022 589254
rect 191786 588698 192022 588934
rect 191786 553018 192022 553254
rect 191786 552698 192022 552934
rect 191786 517018 192022 517254
rect 191786 516698 192022 516934
rect 191786 481018 192022 481254
rect 191786 480698 192022 480934
rect 191786 445018 192022 445254
rect 191786 444698 192022 444934
rect 191786 409018 192022 409254
rect 191786 408698 192022 408934
rect 191786 373018 192022 373254
rect 191786 372698 192022 372934
rect 191786 337018 192022 337254
rect 191786 336698 192022 336934
rect 191786 301018 192022 301254
rect 191786 300698 192022 300934
rect 191786 265018 192022 265254
rect 191786 264698 192022 264934
rect 191786 229018 192022 229254
rect 191786 228698 192022 228934
rect 191786 193018 192022 193254
rect 191786 192698 192022 192934
rect 191786 157018 192022 157254
rect 191786 156698 192022 156934
rect 191786 121018 192022 121254
rect 191786 120698 192022 120934
rect 191786 85018 192022 85254
rect 191786 84698 192022 84934
rect 191786 49018 192022 49254
rect 191786 48698 192022 48934
rect 191786 13018 192022 13254
rect 191786 12698 192022 12934
rect 173786 -7022 174022 -6786
rect 173786 -7342 174022 -7106
rect 198986 705522 199222 705758
rect 198986 705202 199222 705438
rect 198986 668218 199222 668454
rect 198986 667898 199222 668134
rect 198986 632218 199222 632454
rect 198986 631898 199222 632134
rect 198986 596218 199222 596454
rect 198986 595898 199222 596134
rect 198986 560218 199222 560454
rect 198986 559898 199222 560134
rect 198986 524218 199222 524454
rect 198986 523898 199222 524134
rect 198986 488218 199222 488454
rect 198986 487898 199222 488134
rect 198986 452218 199222 452454
rect 198986 451898 199222 452134
rect 198986 416218 199222 416454
rect 198986 415898 199222 416134
rect 198986 380218 199222 380454
rect 198986 379898 199222 380134
rect 198986 344218 199222 344454
rect 198986 343898 199222 344134
rect 198986 308218 199222 308454
rect 198986 307898 199222 308134
rect 198986 272218 199222 272454
rect 198986 271898 199222 272134
rect 198986 236218 199222 236454
rect 198986 235898 199222 236134
rect 198986 200218 199222 200454
rect 198986 199898 199222 200134
rect 198986 164218 199222 164454
rect 198986 163898 199222 164134
rect 198986 128218 199222 128454
rect 198986 127898 199222 128134
rect 198986 92218 199222 92454
rect 198986 91898 199222 92134
rect 198986 56218 199222 56454
rect 198986 55898 199222 56134
rect 198986 20218 199222 20454
rect 198986 19898 199222 20134
rect 198986 -1502 199222 -1266
rect 198986 -1822 199222 -1586
rect 202586 671818 202822 672054
rect 202586 671498 202822 671734
rect 202586 635818 202822 636054
rect 202586 635498 202822 635734
rect 202586 599818 202822 600054
rect 202586 599498 202822 599734
rect 202586 563818 202822 564054
rect 202586 563498 202822 563734
rect 202586 527818 202822 528054
rect 202586 527498 202822 527734
rect 202586 491818 202822 492054
rect 202586 491498 202822 491734
rect 202586 455818 202822 456054
rect 202586 455498 202822 455734
rect 202586 419818 202822 420054
rect 202586 419498 202822 419734
rect 202586 383818 202822 384054
rect 202586 383498 202822 383734
rect 202586 347818 202822 348054
rect 202586 347498 202822 347734
rect 202586 311818 202822 312054
rect 202586 311498 202822 311734
rect 202586 275818 202822 276054
rect 202586 275498 202822 275734
rect 202586 239818 202822 240054
rect 202586 239498 202822 239734
rect 202586 203818 202822 204054
rect 202586 203498 202822 203734
rect 202586 167818 202822 168054
rect 202586 167498 202822 167734
rect 202586 131818 202822 132054
rect 202586 131498 202822 131734
rect 202586 95818 202822 96054
rect 202586 95498 202822 95734
rect 202586 59818 202822 60054
rect 202586 59498 202822 59734
rect 202586 23818 202822 24054
rect 202586 23498 202822 23734
rect 202586 -3342 202822 -3106
rect 202586 -3662 202822 -3426
rect 206186 675418 206422 675654
rect 206186 675098 206422 675334
rect 206186 639418 206422 639654
rect 206186 639098 206422 639334
rect 206186 603418 206422 603654
rect 206186 603098 206422 603334
rect 206186 567418 206422 567654
rect 206186 567098 206422 567334
rect 206186 531418 206422 531654
rect 206186 531098 206422 531334
rect 206186 495418 206422 495654
rect 206186 495098 206422 495334
rect 206186 459418 206422 459654
rect 206186 459098 206422 459334
rect 206186 423418 206422 423654
rect 206186 423098 206422 423334
rect 206186 387418 206422 387654
rect 206186 387098 206422 387334
rect 206186 351418 206422 351654
rect 206186 351098 206422 351334
rect 206186 315418 206422 315654
rect 206186 315098 206422 315334
rect 206186 279418 206422 279654
rect 206186 279098 206422 279334
rect 206186 243418 206422 243654
rect 206186 243098 206422 243334
rect 206186 207418 206422 207654
rect 206186 207098 206422 207334
rect 206186 171418 206422 171654
rect 206186 171098 206422 171334
rect 206186 135418 206422 135654
rect 206186 135098 206422 135334
rect 206186 99418 206422 99654
rect 206186 99098 206422 99334
rect 206186 63418 206422 63654
rect 206186 63098 206422 63334
rect 206186 27418 206422 27654
rect 206186 27098 206422 27334
rect 206186 -5182 206422 -4946
rect 206186 -5502 206422 -5266
rect 227786 710122 228022 710358
rect 227786 709802 228022 710038
rect 224186 708282 224422 708518
rect 224186 707962 224422 708198
rect 220586 706442 220822 706678
rect 220586 706122 220822 706358
rect 209786 679018 210022 679254
rect 209786 678698 210022 678934
rect 209786 643018 210022 643254
rect 209786 642698 210022 642934
rect 209786 607018 210022 607254
rect 209786 606698 210022 606934
rect 209786 571018 210022 571254
rect 209786 570698 210022 570934
rect 209786 535018 210022 535254
rect 209786 534698 210022 534934
rect 209786 499018 210022 499254
rect 209786 498698 210022 498934
rect 209786 463018 210022 463254
rect 209786 462698 210022 462934
rect 209786 427018 210022 427254
rect 209786 426698 210022 426934
rect 209786 391018 210022 391254
rect 209786 390698 210022 390934
rect 209786 355018 210022 355254
rect 209786 354698 210022 354934
rect 209786 319018 210022 319254
rect 209786 318698 210022 318934
rect 209786 283018 210022 283254
rect 209786 282698 210022 282934
rect 209786 247018 210022 247254
rect 209786 246698 210022 246934
rect 209786 211018 210022 211254
rect 209786 210698 210022 210934
rect 209786 175018 210022 175254
rect 209786 174698 210022 174934
rect 209786 139018 210022 139254
rect 209786 138698 210022 138934
rect 209786 103018 210022 103254
rect 209786 102698 210022 102934
rect 209786 67018 210022 67254
rect 209786 66698 210022 66934
rect 209786 31018 210022 31254
rect 209786 30698 210022 30934
rect 191786 -6102 192022 -5866
rect 191786 -6422 192022 -6186
rect 216986 704602 217222 704838
rect 216986 704282 217222 704518
rect 216986 686218 217222 686454
rect 216986 685898 217222 686134
rect 216986 650218 217222 650454
rect 216986 649898 217222 650134
rect 216986 614218 217222 614454
rect 216986 613898 217222 614134
rect 216986 578218 217222 578454
rect 216986 577898 217222 578134
rect 216986 542218 217222 542454
rect 216986 541898 217222 542134
rect 216986 506218 217222 506454
rect 216986 505898 217222 506134
rect 216986 470218 217222 470454
rect 216986 469898 217222 470134
rect 216986 434218 217222 434454
rect 216986 433898 217222 434134
rect 216986 398218 217222 398454
rect 216986 397898 217222 398134
rect 216986 362218 217222 362454
rect 216986 361898 217222 362134
rect 216986 326218 217222 326454
rect 216986 325898 217222 326134
rect 216986 290218 217222 290454
rect 216986 289898 217222 290134
rect 216986 254218 217222 254454
rect 216986 253898 217222 254134
rect 216986 218218 217222 218454
rect 216986 217898 217222 218134
rect 216986 182218 217222 182454
rect 216986 181898 217222 182134
rect 216986 146218 217222 146454
rect 216986 145898 217222 146134
rect 216986 110218 217222 110454
rect 216986 109898 217222 110134
rect 216986 74218 217222 74454
rect 216986 73898 217222 74134
rect 216986 38218 217222 38454
rect 216986 37898 217222 38134
rect 216986 2218 217222 2454
rect 216986 1898 217222 2134
rect 216986 -582 217222 -346
rect 216986 -902 217222 -666
rect 220586 689818 220822 690054
rect 220586 689498 220822 689734
rect 220586 653818 220822 654054
rect 220586 653498 220822 653734
rect 220586 617818 220822 618054
rect 220586 617498 220822 617734
rect 220586 581818 220822 582054
rect 220586 581498 220822 581734
rect 220586 545818 220822 546054
rect 220586 545498 220822 545734
rect 220586 509818 220822 510054
rect 220586 509498 220822 509734
rect 220586 473818 220822 474054
rect 220586 473498 220822 473734
rect 220586 437818 220822 438054
rect 220586 437498 220822 437734
rect 220586 401818 220822 402054
rect 220586 401498 220822 401734
rect 220586 365818 220822 366054
rect 220586 365498 220822 365734
rect 220586 329818 220822 330054
rect 220586 329498 220822 329734
rect 220586 293818 220822 294054
rect 220586 293498 220822 293734
rect 220586 257818 220822 258054
rect 220586 257498 220822 257734
rect 220586 221818 220822 222054
rect 220586 221498 220822 221734
rect 220586 185818 220822 186054
rect 220586 185498 220822 185734
rect 220586 149818 220822 150054
rect 220586 149498 220822 149734
rect 220586 113818 220822 114054
rect 220586 113498 220822 113734
rect 220586 77818 220822 78054
rect 220586 77498 220822 77734
rect 220586 41818 220822 42054
rect 220586 41498 220822 41734
rect 220586 5818 220822 6054
rect 220586 5498 220822 5734
rect 220586 -2422 220822 -2186
rect 220586 -2742 220822 -2506
rect 224186 693418 224422 693654
rect 224186 693098 224422 693334
rect 224186 657418 224422 657654
rect 224186 657098 224422 657334
rect 224186 621418 224422 621654
rect 224186 621098 224422 621334
rect 224186 585418 224422 585654
rect 224186 585098 224422 585334
rect 224186 549418 224422 549654
rect 224186 549098 224422 549334
rect 224186 513418 224422 513654
rect 224186 513098 224422 513334
rect 224186 477418 224422 477654
rect 224186 477098 224422 477334
rect 224186 441418 224422 441654
rect 224186 441098 224422 441334
rect 224186 405418 224422 405654
rect 224186 405098 224422 405334
rect 224186 369418 224422 369654
rect 224186 369098 224422 369334
rect 224186 333418 224422 333654
rect 224186 333098 224422 333334
rect 224186 297418 224422 297654
rect 224186 297098 224422 297334
rect 224186 261418 224422 261654
rect 224186 261098 224422 261334
rect 224186 225418 224422 225654
rect 224186 225098 224422 225334
rect 224186 189418 224422 189654
rect 224186 189098 224422 189334
rect 224186 153418 224422 153654
rect 224186 153098 224422 153334
rect 224186 117418 224422 117654
rect 224186 117098 224422 117334
rect 224186 81418 224422 81654
rect 224186 81098 224422 81334
rect 224186 45418 224422 45654
rect 224186 45098 224422 45334
rect 224186 9418 224422 9654
rect 224186 9098 224422 9334
rect 224186 -4262 224422 -4026
rect 224186 -4582 224422 -4346
rect 245786 711042 246022 711278
rect 245786 710722 246022 710958
rect 242186 709202 242422 709438
rect 242186 708882 242422 709118
rect 238586 707362 238822 707598
rect 238586 707042 238822 707278
rect 227786 697018 228022 697254
rect 227786 696698 228022 696934
rect 227786 661018 228022 661254
rect 227786 660698 228022 660934
rect 227786 625018 228022 625254
rect 227786 624698 228022 624934
rect 227786 589018 228022 589254
rect 227786 588698 228022 588934
rect 227786 553018 228022 553254
rect 227786 552698 228022 552934
rect 227786 517018 228022 517254
rect 227786 516698 228022 516934
rect 227786 481018 228022 481254
rect 227786 480698 228022 480934
rect 227786 445018 228022 445254
rect 227786 444698 228022 444934
rect 227786 409018 228022 409254
rect 227786 408698 228022 408934
rect 234986 705522 235222 705758
rect 234986 705202 235222 705438
rect 234986 668218 235222 668454
rect 234986 667898 235222 668134
rect 234986 632218 235222 632454
rect 234986 631898 235222 632134
rect 234986 596218 235222 596454
rect 234986 595898 235222 596134
rect 234986 560218 235222 560454
rect 234986 559898 235222 560134
rect 234986 524218 235222 524454
rect 234986 523898 235222 524134
rect 234986 488218 235222 488454
rect 234986 487898 235222 488134
rect 234986 452218 235222 452454
rect 234986 451898 235222 452134
rect 234986 416218 235222 416454
rect 234986 415898 235222 416134
rect 227786 373018 228022 373254
rect 227786 372698 228022 372934
rect 227786 337018 228022 337254
rect 227786 336698 228022 336934
rect 227786 301018 228022 301254
rect 227786 300698 228022 300934
rect 227786 265018 228022 265254
rect 227786 264698 228022 264934
rect 227786 229018 228022 229254
rect 227786 228698 228022 228934
rect 227786 193018 228022 193254
rect 227786 192698 228022 192934
rect 227786 157018 228022 157254
rect 227786 156698 228022 156934
rect 227786 121018 228022 121254
rect 227786 120698 228022 120934
rect 227786 85018 228022 85254
rect 227786 84698 228022 84934
rect 227786 49018 228022 49254
rect 227786 48698 228022 48934
rect 238586 671818 238822 672054
rect 238586 671498 238822 671734
rect 238586 635818 238822 636054
rect 238586 635498 238822 635734
rect 238586 599818 238822 600054
rect 238586 599498 238822 599734
rect 238586 563818 238822 564054
rect 238586 563498 238822 563734
rect 238586 527818 238822 528054
rect 238586 527498 238822 527734
rect 238586 491818 238822 492054
rect 238586 491498 238822 491734
rect 238586 455818 238822 456054
rect 238586 455498 238822 455734
rect 238586 419818 238822 420054
rect 238586 419498 238822 419734
rect 234986 380218 235222 380454
rect 234986 379898 235222 380134
rect 234986 344218 235222 344454
rect 234986 343898 235222 344134
rect 234986 308218 235222 308454
rect 234986 307898 235222 308134
rect 234986 272218 235222 272454
rect 234986 271898 235222 272134
rect 234986 236218 235222 236454
rect 234986 235898 235222 236134
rect 242186 675418 242422 675654
rect 242186 675098 242422 675334
rect 242186 639418 242422 639654
rect 242186 639098 242422 639334
rect 242186 603418 242422 603654
rect 242186 603098 242422 603334
rect 242186 567418 242422 567654
rect 242186 567098 242422 567334
rect 242186 531418 242422 531654
rect 242186 531098 242422 531334
rect 242186 495418 242422 495654
rect 242186 495098 242422 495334
rect 242186 459418 242422 459654
rect 242186 459098 242422 459334
rect 242186 423418 242422 423654
rect 242186 423098 242422 423334
rect 238586 383818 238822 384054
rect 238586 383498 238822 383734
rect 238586 347818 238822 348054
rect 238586 347498 238822 347734
rect 238586 311818 238822 312054
rect 238586 311498 238822 311734
rect 263786 710122 264022 710358
rect 263786 709802 264022 710038
rect 260186 708282 260422 708518
rect 260186 707962 260422 708198
rect 256586 706442 256822 706678
rect 256586 706122 256822 706358
rect 245786 679018 246022 679254
rect 245786 678698 246022 678934
rect 245786 643018 246022 643254
rect 245786 642698 246022 642934
rect 245786 607018 246022 607254
rect 245786 606698 246022 606934
rect 245786 571018 246022 571254
rect 245786 570698 246022 570934
rect 245786 535018 246022 535254
rect 245786 534698 246022 534934
rect 245786 499018 246022 499254
rect 245786 498698 246022 498934
rect 245786 463018 246022 463254
rect 245786 462698 246022 462934
rect 245786 427018 246022 427254
rect 245786 426698 246022 426934
rect 242186 387418 242422 387654
rect 242186 387098 242422 387334
rect 242186 351418 242422 351654
rect 242186 351098 242422 351334
rect 245786 391018 246022 391254
rect 245786 390698 246022 390934
rect 245786 355018 246022 355254
rect 245786 354698 246022 354934
rect 242186 315418 242422 315654
rect 242186 315098 242422 315334
rect 238586 275818 238822 276054
rect 238586 275498 238822 275734
rect 238586 239818 238822 240054
rect 238586 239498 238822 239734
rect 234986 200218 235222 200454
rect 234986 199898 235222 200134
rect 234986 164218 235222 164454
rect 234986 163898 235222 164134
rect 234986 128218 235222 128454
rect 234986 127898 235222 128134
rect 234986 92218 235222 92454
rect 234986 91898 235222 92134
rect 234986 56218 235222 56454
rect 234986 55898 235222 56134
rect 227786 13018 228022 13254
rect 227786 12698 228022 12934
rect 209786 -7022 210022 -6786
rect 209786 -7342 210022 -7106
rect 234986 20218 235222 20454
rect 234986 19898 235222 20134
rect 234986 -1502 235222 -1266
rect 234986 -1822 235222 -1586
rect 238586 203818 238822 204054
rect 238586 203498 238822 203734
rect 238586 167818 238822 168054
rect 238586 167498 238822 167734
rect 238586 131818 238822 132054
rect 238586 131498 238822 131734
rect 238586 95818 238822 96054
rect 238586 95498 238822 95734
rect 242186 279418 242422 279654
rect 242186 279098 242422 279334
rect 242186 243418 242422 243654
rect 242186 243098 242422 243334
rect 242186 207418 242422 207654
rect 242186 207098 242422 207334
rect 242186 171418 242422 171654
rect 242186 171098 242422 171334
rect 242186 135418 242422 135654
rect 242186 135098 242422 135334
rect 242186 99418 242422 99654
rect 242186 99098 242422 99334
rect 238586 59818 238822 60054
rect 238586 59498 238822 59734
rect 238586 23818 238822 24054
rect 238586 23498 238822 23734
rect 238586 -3342 238822 -3106
rect 238586 -3662 238822 -3426
rect 242186 63418 242422 63654
rect 242186 63098 242422 63334
rect 242186 27418 242422 27654
rect 242186 27098 242422 27334
rect 242186 -5182 242422 -4946
rect 242186 -5502 242422 -5266
rect 245786 319018 246022 319254
rect 245786 318698 246022 318934
rect 245786 283018 246022 283254
rect 245786 282698 246022 282934
rect 245786 247018 246022 247254
rect 245786 246698 246022 246934
rect 245786 211018 246022 211254
rect 245786 210698 246022 210934
rect 245786 175018 246022 175254
rect 245786 174698 246022 174934
rect 245786 139018 246022 139254
rect 245786 138698 246022 138934
rect 245786 103018 246022 103254
rect 245786 102698 246022 102934
rect 245786 67018 246022 67254
rect 245786 66698 246022 66934
rect 245786 31018 246022 31254
rect 245786 30698 246022 30934
rect 227786 -6102 228022 -5866
rect 227786 -6422 228022 -6186
rect 252986 704602 253222 704838
rect 252986 704282 253222 704518
rect 252986 686218 253222 686454
rect 252986 685898 253222 686134
rect 252986 650218 253222 650454
rect 252986 649898 253222 650134
rect 252986 614218 253222 614454
rect 252986 613898 253222 614134
rect 252986 578218 253222 578454
rect 252986 577898 253222 578134
rect 252986 542218 253222 542454
rect 252986 541898 253222 542134
rect 252986 506218 253222 506454
rect 252986 505898 253222 506134
rect 252986 470218 253222 470454
rect 252986 469898 253222 470134
rect 252986 434218 253222 434454
rect 252986 433898 253222 434134
rect 252986 398218 253222 398454
rect 252986 397898 253222 398134
rect 252986 362218 253222 362454
rect 252986 361898 253222 362134
rect 252986 326218 253222 326454
rect 252986 325898 253222 326134
rect 252986 290218 253222 290454
rect 252986 289898 253222 290134
rect 252986 254218 253222 254454
rect 252986 253898 253222 254134
rect 252986 218218 253222 218454
rect 252986 217898 253222 218134
rect 252986 182218 253222 182454
rect 252986 181898 253222 182134
rect 252986 146218 253222 146454
rect 252986 145898 253222 146134
rect 252986 110218 253222 110454
rect 252986 109898 253222 110134
rect 252986 74218 253222 74454
rect 252986 73898 253222 74134
rect 252986 38218 253222 38454
rect 252986 37898 253222 38134
rect 252986 2218 253222 2454
rect 252986 1898 253222 2134
rect 252986 -582 253222 -346
rect 252986 -902 253222 -666
rect 256586 689818 256822 690054
rect 256586 689498 256822 689734
rect 256586 653818 256822 654054
rect 256586 653498 256822 653734
rect 256586 617818 256822 618054
rect 256586 617498 256822 617734
rect 256586 581818 256822 582054
rect 256586 581498 256822 581734
rect 256586 545818 256822 546054
rect 256586 545498 256822 545734
rect 256586 509818 256822 510054
rect 256586 509498 256822 509734
rect 256586 473818 256822 474054
rect 256586 473498 256822 473734
rect 256586 437818 256822 438054
rect 256586 437498 256822 437734
rect 256586 401818 256822 402054
rect 256586 401498 256822 401734
rect 256586 365818 256822 366054
rect 256586 365498 256822 365734
rect 256586 329818 256822 330054
rect 256586 329498 256822 329734
rect 260186 693418 260422 693654
rect 260186 693098 260422 693334
rect 260186 657418 260422 657654
rect 260186 657098 260422 657334
rect 260186 621418 260422 621654
rect 260186 621098 260422 621334
rect 260186 585418 260422 585654
rect 260186 585098 260422 585334
rect 260186 549418 260422 549654
rect 260186 549098 260422 549334
rect 260186 513418 260422 513654
rect 260186 513098 260422 513334
rect 260186 477418 260422 477654
rect 260186 477098 260422 477334
rect 260186 441418 260422 441654
rect 260186 441098 260422 441334
rect 260186 405418 260422 405654
rect 260186 405098 260422 405334
rect 281786 711042 282022 711278
rect 281786 710722 282022 710958
rect 278186 709202 278422 709438
rect 278186 708882 278422 709118
rect 274586 707362 274822 707598
rect 274586 707042 274822 707278
rect 263786 697018 264022 697254
rect 263786 696698 264022 696934
rect 263786 661018 264022 661254
rect 263786 660698 264022 660934
rect 263786 625018 264022 625254
rect 263786 624698 264022 624934
rect 263786 589018 264022 589254
rect 263786 588698 264022 588934
rect 263786 553018 264022 553254
rect 263786 552698 264022 552934
rect 263786 517018 264022 517254
rect 263786 516698 264022 516934
rect 263786 481018 264022 481254
rect 263786 480698 264022 480934
rect 263786 445018 264022 445254
rect 263786 444698 264022 444934
rect 263786 409018 264022 409254
rect 263786 408698 264022 408934
rect 260186 369418 260422 369654
rect 260186 369098 260422 369334
rect 263786 373018 264022 373254
rect 263786 372698 264022 372934
rect 263786 337018 264022 337254
rect 263786 336698 264022 336934
rect 260186 333418 260422 333654
rect 260186 333098 260422 333334
rect 256586 293818 256822 294054
rect 256586 293498 256822 293734
rect 256586 257818 256822 258054
rect 256586 257498 256822 257734
rect 260186 297418 260422 297654
rect 260186 297098 260422 297334
rect 260186 261418 260422 261654
rect 260186 261098 260422 261334
rect 256586 221818 256822 222054
rect 256586 221498 256822 221734
rect 256586 185818 256822 186054
rect 256586 185498 256822 185734
rect 256586 149818 256822 150054
rect 256586 149498 256822 149734
rect 256586 113818 256822 114054
rect 256586 113498 256822 113734
rect 256586 77818 256822 78054
rect 256586 77498 256822 77734
rect 256586 41818 256822 42054
rect 256586 41498 256822 41734
rect 256586 5818 256822 6054
rect 256586 5498 256822 5734
rect 256586 -2422 256822 -2186
rect 256586 -2742 256822 -2506
rect 260186 225418 260422 225654
rect 260186 225098 260422 225334
rect 260186 189418 260422 189654
rect 260186 189098 260422 189334
rect 260186 153418 260422 153654
rect 260186 153098 260422 153334
rect 260186 117418 260422 117654
rect 260186 117098 260422 117334
rect 260186 81418 260422 81654
rect 260186 81098 260422 81334
rect 263786 301018 264022 301254
rect 263786 300698 264022 300934
rect 263786 265018 264022 265254
rect 263786 264698 264022 264934
rect 263786 229018 264022 229254
rect 263786 228698 264022 228934
rect 263786 193018 264022 193254
rect 263786 192698 264022 192934
rect 263786 157018 264022 157254
rect 263786 156698 264022 156934
rect 263786 121018 264022 121254
rect 263786 120698 264022 120934
rect 263786 85018 264022 85254
rect 263786 84698 264022 84934
rect 260186 45418 260422 45654
rect 260186 45098 260422 45334
rect 260186 9418 260422 9654
rect 260186 9098 260422 9334
rect 260186 -4262 260422 -4026
rect 260186 -4582 260422 -4346
rect 263786 49018 264022 49254
rect 263786 48698 264022 48934
rect 270986 705522 271222 705758
rect 270986 705202 271222 705438
rect 270986 668218 271222 668454
rect 270986 667898 271222 668134
rect 270986 632218 271222 632454
rect 270986 631898 271222 632134
rect 270986 596218 271222 596454
rect 270986 595898 271222 596134
rect 270986 560218 271222 560454
rect 270986 559898 271222 560134
rect 270986 524218 271222 524454
rect 270986 523898 271222 524134
rect 270986 488218 271222 488454
rect 270986 487898 271222 488134
rect 270986 452218 271222 452454
rect 270986 451898 271222 452134
rect 270986 416218 271222 416454
rect 270986 415898 271222 416134
rect 270986 380218 271222 380454
rect 270986 379898 271222 380134
rect 270986 344218 271222 344454
rect 270986 343898 271222 344134
rect 270986 308218 271222 308454
rect 270986 307898 271222 308134
rect 270986 272218 271222 272454
rect 270986 271898 271222 272134
rect 270986 236218 271222 236454
rect 270986 235898 271222 236134
rect 270986 200218 271222 200454
rect 270986 199898 271222 200134
rect 270986 164218 271222 164454
rect 270986 163898 271222 164134
rect 270986 128218 271222 128454
rect 270986 127898 271222 128134
rect 270986 92218 271222 92454
rect 270986 91898 271222 92134
rect 270986 56218 271222 56454
rect 270986 55898 271222 56134
rect 263786 13018 264022 13254
rect 263786 12698 264022 12934
rect 245786 -7022 246022 -6786
rect 245786 -7342 246022 -7106
rect 270986 20218 271222 20454
rect 270986 19898 271222 20134
rect 270986 -1502 271222 -1266
rect 270986 -1822 271222 -1586
rect 274586 671818 274822 672054
rect 274586 671498 274822 671734
rect 274586 635818 274822 636054
rect 274586 635498 274822 635734
rect 274586 599818 274822 600054
rect 274586 599498 274822 599734
rect 274586 563818 274822 564054
rect 274586 563498 274822 563734
rect 274586 527818 274822 528054
rect 274586 527498 274822 527734
rect 274586 491818 274822 492054
rect 274586 491498 274822 491734
rect 274586 455818 274822 456054
rect 274586 455498 274822 455734
rect 274586 419818 274822 420054
rect 274586 419498 274822 419734
rect 274586 383818 274822 384054
rect 274586 383498 274822 383734
rect 274586 347818 274822 348054
rect 274586 347498 274822 347734
rect 278186 675418 278422 675654
rect 278186 675098 278422 675334
rect 278186 639418 278422 639654
rect 278186 639098 278422 639334
rect 278186 603418 278422 603654
rect 278186 603098 278422 603334
rect 278186 567418 278422 567654
rect 278186 567098 278422 567334
rect 278186 531418 278422 531654
rect 278186 531098 278422 531334
rect 278186 495418 278422 495654
rect 278186 495098 278422 495334
rect 278186 459418 278422 459654
rect 278186 459098 278422 459334
rect 278186 423418 278422 423654
rect 278186 423098 278422 423334
rect 278186 387418 278422 387654
rect 278186 387098 278422 387334
rect 278186 351418 278422 351654
rect 278186 351098 278422 351334
rect 278186 315418 278422 315654
rect 278186 315098 278422 315334
rect 274586 311818 274822 312054
rect 274586 311498 274822 311734
rect 274586 275818 274822 276054
rect 274586 275498 274822 275734
rect 274586 239818 274822 240054
rect 274586 239498 274822 239734
rect 274586 203818 274822 204054
rect 274586 203498 274822 203734
rect 274586 167818 274822 168054
rect 274586 167498 274822 167734
rect 274586 131818 274822 132054
rect 274586 131498 274822 131734
rect 274586 95818 274822 96054
rect 274586 95498 274822 95734
rect 274586 59818 274822 60054
rect 274586 59498 274822 59734
rect 274586 23818 274822 24054
rect 274586 23498 274822 23734
rect 274586 -3342 274822 -3106
rect 274586 -3662 274822 -3426
rect 278186 279418 278422 279654
rect 278186 279098 278422 279334
rect 278186 243418 278422 243654
rect 278186 243098 278422 243334
rect 278186 207418 278422 207654
rect 278186 207098 278422 207334
rect 278186 171418 278422 171654
rect 278186 171098 278422 171334
rect 278186 135418 278422 135654
rect 278186 135098 278422 135334
rect 278186 99418 278422 99654
rect 278186 99098 278422 99334
rect 278186 63418 278422 63654
rect 278186 63098 278422 63334
rect 278186 27418 278422 27654
rect 278186 27098 278422 27334
rect 278186 -5182 278422 -4946
rect 278186 -5502 278422 -5266
rect 299786 710122 300022 710358
rect 299786 709802 300022 710038
rect 296186 708282 296422 708518
rect 296186 707962 296422 708198
rect 292586 706442 292822 706678
rect 292586 706122 292822 706358
rect 281786 679018 282022 679254
rect 281786 678698 282022 678934
rect 281786 643018 282022 643254
rect 281786 642698 282022 642934
rect 281786 607018 282022 607254
rect 281786 606698 282022 606934
rect 281786 571018 282022 571254
rect 281786 570698 282022 570934
rect 281786 535018 282022 535254
rect 281786 534698 282022 534934
rect 281786 499018 282022 499254
rect 281786 498698 282022 498934
rect 281786 463018 282022 463254
rect 281786 462698 282022 462934
rect 281786 427018 282022 427254
rect 281786 426698 282022 426934
rect 288986 704602 289222 704838
rect 288986 704282 289222 704518
rect 288986 686218 289222 686454
rect 288986 685898 289222 686134
rect 288986 650218 289222 650454
rect 288986 649898 289222 650134
rect 288986 614218 289222 614454
rect 288986 613898 289222 614134
rect 288986 578218 289222 578454
rect 288986 577898 289222 578134
rect 288986 542218 289222 542454
rect 288986 541898 289222 542134
rect 288986 506218 289222 506454
rect 288986 505898 289222 506134
rect 288986 470218 289222 470454
rect 288986 469898 289222 470134
rect 288986 434218 289222 434454
rect 288986 433898 289222 434134
rect 281786 391018 282022 391254
rect 281786 390698 282022 390934
rect 281786 355018 282022 355254
rect 281786 354698 282022 354934
rect 281786 319018 282022 319254
rect 281786 318698 282022 318934
rect 281786 283018 282022 283254
rect 281786 282698 282022 282934
rect 281786 247018 282022 247254
rect 281786 246698 282022 246934
rect 281786 211018 282022 211254
rect 281786 210698 282022 210934
rect 281786 175018 282022 175254
rect 281786 174698 282022 174934
rect 281786 139018 282022 139254
rect 281786 138698 282022 138934
rect 281786 103018 282022 103254
rect 281786 102698 282022 102934
rect 281786 67018 282022 67254
rect 281786 66698 282022 66934
rect 288986 398218 289222 398454
rect 288986 397898 289222 398134
rect 288986 362218 289222 362454
rect 288986 361898 289222 362134
rect 288986 326218 289222 326454
rect 288986 325898 289222 326134
rect 288986 290218 289222 290454
rect 288986 289898 289222 290134
rect 288986 254218 289222 254454
rect 288986 253898 289222 254134
rect 288986 218218 289222 218454
rect 288986 217898 289222 218134
rect 288986 182218 289222 182454
rect 288986 181898 289222 182134
rect 288986 146218 289222 146454
rect 288986 145898 289222 146134
rect 288986 110218 289222 110454
rect 288986 109898 289222 110134
rect 288986 74218 289222 74454
rect 288986 73898 289222 74134
rect 281786 31018 282022 31254
rect 281786 30698 282022 30934
rect 263786 -6102 264022 -5866
rect 263786 -6422 264022 -6186
rect 288986 38218 289222 38454
rect 288986 37898 289222 38134
rect 288986 2218 289222 2454
rect 288986 1898 289222 2134
rect 288986 -582 289222 -346
rect 288986 -902 289222 -666
rect 292586 689818 292822 690054
rect 292586 689498 292822 689734
rect 292586 653818 292822 654054
rect 292586 653498 292822 653734
rect 292586 617818 292822 618054
rect 292586 617498 292822 617734
rect 292586 581818 292822 582054
rect 292586 581498 292822 581734
rect 292586 545818 292822 546054
rect 292586 545498 292822 545734
rect 292586 509818 292822 510054
rect 292586 509498 292822 509734
rect 292586 473818 292822 474054
rect 292586 473498 292822 473734
rect 292586 437818 292822 438054
rect 292586 437498 292822 437734
rect 292586 401818 292822 402054
rect 292586 401498 292822 401734
rect 292586 365818 292822 366054
rect 292586 365498 292822 365734
rect 292586 329818 292822 330054
rect 292586 329498 292822 329734
rect 292586 293818 292822 294054
rect 292586 293498 292822 293734
rect 292586 257818 292822 258054
rect 292586 257498 292822 257734
rect 292586 221818 292822 222054
rect 292586 221498 292822 221734
rect 292586 185818 292822 186054
rect 292586 185498 292822 185734
rect 292586 149818 292822 150054
rect 292586 149498 292822 149734
rect 292586 113818 292822 114054
rect 292586 113498 292822 113734
rect 292586 77818 292822 78054
rect 292586 77498 292822 77734
rect 292586 41818 292822 42054
rect 292586 41498 292822 41734
rect 292586 5818 292822 6054
rect 292586 5498 292822 5734
rect 292586 -2422 292822 -2186
rect 292586 -2742 292822 -2506
rect 296186 693418 296422 693654
rect 296186 693098 296422 693334
rect 296186 657418 296422 657654
rect 296186 657098 296422 657334
rect 296186 621418 296422 621654
rect 296186 621098 296422 621334
rect 296186 585418 296422 585654
rect 296186 585098 296422 585334
rect 296186 549418 296422 549654
rect 296186 549098 296422 549334
rect 296186 513418 296422 513654
rect 296186 513098 296422 513334
rect 296186 477418 296422 477654
rect 296186 477098 296422 477334
rect 296186 441418 296422 441654
rect 296186 441098 296422 441334
rect 296186 405418 296422 405654
rect 296186 405098 296422 405334
rect 296186 369418 296422 369654
rect 296186 369098 296422 369334
rect 296186 333418 296422 333654
rect 296186 333098 296422 333334
rect 317786 711042 318022 711278
rect 317786 710722 318022 710958
rect 314186 709202 314422 709438
rect 314186 708882 314422 709118
rect 310586 707362 310822 707598
rect 310586 707042 310822 707278
rect 299786 697018 300022 697254
rect 299786 696698 300022 696934
rect 299786 661018 300022 661254
rect 299786 660698 300022 660934
rect 299786 625018 300022 625254
rect 299786 624698 300022 624934
rect 299786 589018 300022 589254
rect 299786 588698 300022 588934
rect 299786 553018 300022 553254
rect 299786 552698 300022 552934
rect 299786 517018 300022 517254
rect 299786 516698 300022 516934
rect 299786 481018 300022 481254
rect 299786 480698 300022 480934
rect 299786 445018 300022 445254
rect 299786 444698 300022 444934
rect 299786 409018 300022 409254
rect 299786 408698 300022 408934
rect 299786 373018 300022 373254
rect 299786 372698 300022 372934
rect 299786 337018 300022 337254
rect 299786 336698 300022 336934
rect 296186 297418 296422 297654
rect 296186 297098 296422 297334
rect 296186 261418 296422 261654
rect 296186 261098 296422 261334
rect 296186 225418 296422 225654
rect 296186 225098 296422 225334
rect 296186 189418 296422 189654
rect 296186 189098 296422 189334
rect 296186 153418 296422 153654
rect 296186 153098 296422 153334
rect 296186 117418 296422 117654
rect 296186 117098 296422 117334
rect 296186 81418 296422 81654
rect 296186 81098 296422 81334
rect 296186 45418 296422 45654
rect 296186 45098 296422 45334
rect 296186 9418 296422 9654
rect 296186 9098 296422 9334
rect 296186 -4262 296422 -4026
rect 296186 -4582 296422 -4346
rect 299786 301018 300022 301254
rect 299786 300698 300022 300934
rect 299786 265018 300022 265254
rect 299786 264698 300022 264934
rect 299786 229018 300022 229254
rect 299786 228698 300022 228934
rect 299786 193018 300022 193254
rect 299786 192698 300022 192934
rect 299786 157018 300022 157254
rect 299786 156698 300022 156934
rect 299786 121018 300022 121254
rect 299786 120698 300022 120934
rect 299786 85018 300022 85254
rect 299786 84698 300022 84934
rect 299786 49018 300022 49254
rect 299786 48698 300022 48934
rect 299786 13018 300022 13254
rect 299786 12698 300022 12934
rect 281786 -7022 282022 -6786
rect 281786 -7342 282022 -7106
rect 306986 705522 307222 705758
rect 306986 705202 307222 705438
rect 306986 668218 307222 668454
rect 306986 667898 307222 668134
rect 306986 632218 307222 632454
rect 306986 631898 307222 632134
rect 306986 596218 307222 596454
rect 306986 595898 307222 596134
rect 306986 560218 307222 560454
rect 306986 559898 307222 560134
rect 306986 524218 307222 524454
rect 306986 523898 307222 524134
rect 306986 488218 307222 488454
rect 306986 487898 307222 488134
rect 306986 452218 307222 452454
rect 306986 451898 307222 452134
rect 306986 416218 307222 416454
rect 306986 415898 307222 416134
rect 306986 380218 307222 380454
rect 306986 379898 307222 380134
rect 306986 344218 307222 344454
rect 306986 343898 307222 344134
rect 306986 308218 307222 308454
rect 306986 307898 307222 308134
rect 306986 272218 307222 272454
rect 306986 271898 307222 272134
rect 306986 236218 307222 236454
rect 306986 235898 307222 236134
rect 306986 200218 307222 200454
rect 306986 199898 307222 200134
rect 306986 164218 307222 164454
rect 306986 163898 307222 164134
rect 306986 128218 307222 128454
rect 306986 127898 307222 128134
rect 306986 92218 307222 92454
rect 306986 91898 307222 92134
rect 306986 56218 307222 56454
rect 306986 55898 307222 56134
rect 306986 20218 307222 20454
rect 306986 19898 307222 20134
rect 306986 -1502 307222 -1266
rect 306986 -1822 307222 -1586
rect 310586 671818 310822 672054
rect 310586 671498 310822 671734
rect 310586 635818 310822 636054
rect 310586 635498 310822 635734
rect 310586 599818 310822 600054
rect 310586 599498 310822 599734
rect 310586 563818 310822 564054
rect 310586 563498 310822 563734
rect 310586 527818 310822 528054
rect 310586 527498 310822 527734
rect 310586 491818 310822 492054
rect 310586 491498 310822 491734
rect 310586 455818 310822 456054
rect 310586 455498 310822 455734
rect 310586 419818 310822 420054
rect 310586 419498 310822 419734
rect 310586 383818 310822 384054
rect 310586 383498 310822 383734
rect 310586 347818 310822 348054
rect 310586 347498 310822 347734
rect 310586 311818 310822 312054
rect 310586 311498 310822 311734
rect 310586 275818 310822 276054
rect 310586 275498 310822 275734
rect 310586 239818 310822 240054
rect 310586 239498 310822 239734
rect 310586 203818 310822 204054
rect 310586 203498 310822 203734
rect 310586 167818 310822 168054
rect 310586 167498 310822 167734
rect 310586 131818 310822 132054
rect 310586 131498 310822 131734
rect 310586 95818 310822 96054
rect 310586 95498 310822 95734
rect 310586 59818 310822 60054
rect 310586 59498 310822 59734
rect 310586 23818 310822 24054
rect 310586 23498 310822 23734
rect 310586 -3342 310822 -3106
rect 310586 -3662 310822 -3426
rect 314186 675418 314422 675654
rect 314186 675098 314422 675334
rect 314186 639418 314422 639654
rect 314186 639098 314422 639334
rect 314186 603418 314422 603654
rect 314186 603098 314422 603334
rect 314186 567418 314422 567654
rect 314186 567098 314422 567334
rect 314186 531418 314422 531654
rect 314186 531098 314422 531334
rect 314186 495418 314422 495654
rect 314186 495098 314422 495334
rect 314186 459418 314422 459654
rect 314186 459098 314422 459334
rect 314186 423418 314422 423654
rect 314186 423098 314422 423334
rect 314186 387418 314422 387654
rect 314186 387098 314422 387334
rect 314186 351418 314422 351654
rect 314186 351098 314422 351334
rect 314186 315418 314422 315654
rect 314186 315098 314422 315334
rect 314186 279418 314422 279654
rect 314186 279098 314422 279334
rect 314186 243418 314422 243654
rect 314186 243098 314422 243334
rect 314186 207418 314422 207654
rect 314186 207098 314422 207334
rect 314186 171418 314422 171654
rect 314186 171098 314422 171334
rect 314186 135418 314422 135654
rect 314186 135098 314422 135334
rect 314186 99418 314422 99654
rect 314186 99098 314422 99334
rect 314186 63418 314422 63654
rect 314186 63098 314422 63334
rect 314186 27418 314422 27654
rect 314186 27098 314422 27334
rect 314186 -5182 314422 -4946
rect 314186 -5502 314422 -5266
rect 335786 710122 336022 710358
rect 335786 709802 336022 710038
rect 332186 708282 332422 708518
rect 332186 707962 332422 708198
rect 328586 706442 328822 706678
rect 328586 706122 328822 706358
rect 317786 679018 318022 679254
rect 317786 678698 318022 678934
rect 317786 643018 318022 643254
rect 317786 642698 318022 642934
rect 317786 607018 318022 607254
rect 317786 606698 318022 606934
rect 317786 571018 318022 571254
rect 317786 570698 318022 570934
rect 317786 535018 318022 535254
rect 317786 534698 318022 534934
rect 317786 499018 318022 499254
rect 317786 498698 318022 498934
rect 317786 463018 318022 463254
rect 317786 462698 318022 462934
rect 317786 427018 318022 427254
rect 317786 426698 318022 426934
rect 317786 391018 318022 391254
rect 317786 390698 318022 390934
rect 317786 355018 318022 355254
rect 317786 354698 318022 354934
rect 317786 319018 318022 319254
rect 317786 318698 318022 318934
rect 317786 283018 318022 283254
rect 317786 282698 318022 282934
rect 317786 247018 318022 247254
rect 317786 246698 318022 246934
rect 317786 211018 318022 211254
rect 317786 210698 318022 210934
rect 317786 175018 318022 175254
rect 317786 174698 318022 174934
rect 317786 139018 318022 139254
rect 317786 138698 318022 138934
rect 317786 103018 318022 103254
rect 317786 102698 318022 102934
rect 317786 67018 318022 67254
rect 317786 66698 318022 66934
rect 317786 31018 318022 31254
rect 317786 30698 318022 30934
rect 299786 -6102 300022 -5866
rect 299786 -6422 300022 -6186
rect 324986 704602 325222 704838
rect 324986 704282 325222 704518
rect 324986 686218 325222 686454
rect 324986 685898 325222 686134
rect 324986 650218 325222 650454
rect 324986 649898 325222 650134
rect 324986 614218 325222 614454
rect 324986 613898 325222 614134
rect 324986 578218 325222 578454
rect 324986 577898 325222 578134
rect 324986 542218 325222 542454
rect 324986 541898 325222 542134
rect 324986 506218 325222 506454
rect 324986 505898 325222 506134
rect 324986 470218 325222 470454
rect 324986 469898 325222 470134
rect 324986 434218 325222 434454
rect 324986 433898 325222 434134
rect 324986 398218 325222 398454
rect 324986 397898 325222 398134
rect 324986 362218 325222 362454
rect 324986 361898 325222 362134
rect 324986 326218 325222 326454
rect 324986 325898 325222 326134
rect 324986 290218 325222 290454
rect 324986 289898 325222 290134
rect 324986 254218 325222 254454
rect 324986 253898 325222 254134
rect 324986 218218 325222 218454
rect 324986 217898 325222 218134
rect 324986 182218 325222 182454
rect 324986 181898 325222 182134
rect 324986 146218 325222 146454
rect 324986 145898 325222 146134
rect 324986 110218 325222 110454
rect 324986 109898 325222 110134
rect 324986 74218 325222 74454
rect 324986 73898 325222 74134
rect 324986 38218 325222 38454
rect 324986 37898 325222 38134
rect 324986 2218 325222 2454
rect 324986 1898 325222 2134
rect 324986 -582 325222 -346
rect 324986 -902 325222 -666
rect 328586 689818 328822 690054
rect 328586 689498 328822 689734
rect 328586 653818 328822 654054
rect 328586 653498 328822 653734
rect 328586 617818 328822 618054
rect 328586 617498 328822 617734
rect 328586 581818 328822 582054
rect 328586 581498 328822 581734
rect 328586 545818 328822 546054
rect 328586 545498 328822 545734
rect 328586 509818 328822 510054
rect 328586 509498 328822 509734
rect 328586 473818 328822 474054
rect 328586 473498 328822 473734
rect 328586 437818 328822 438054
rect 328586 437498 328822 437734
rect 328586 401818 328822 402054
rect 328586 401498 328822 401734
rect 328586 365818 328822 366054
rect 328586 365498 328822 365734
rect 328586 329818 328822 330054
rect 328586 329498 328822 329734
rect 328586 293818 328822 294054
rect 328586 293498 328822 293734
rect 328586 257818 328822 258054
rect 328586 257498 328822 257734
rect 328586 221818 328822 222054
rect 328586 221498 328822 221734
rect 328586 185818 328822 186054
rect 328586 185498 328822 185734
rect 328586 149818 328822 150054
rect 328586 149498 328822 149734
rect 328586 113818 328822 114054
rect 328586 113498 328822 113734
rect 328586 77818 328822 78054
rect 328586 77498 328822 77734
rect 328586 41818 328822 42054
rect 328586 41498 328822 41734
rect 328586 5818 328822 6054
rect 328586 5498 328822 5734
rect 328586 -2422 328822 -2186
rect 328586 -2742 328822 -2506
rect 332186 693418 332422 693654
rect 332186 693098 332422 693334
rect 332186 657418 332422 657654
rect 332186 657098 332422 657334
rect 332186 621418 332422 621654
rect 332186 621098 332422 621334
rect 332186 585418 332422 585654
rect 332186 585098 332422 585334
rect 332186 549418 332422 549654
rect 332186 549098 332422 549334
rect 332186 513418 332422 513654
rect 332186 513098 332422 513334
rect 332186 477418 332422 477654
rect 332186 477098 332422 477334
rect 332186 441418 332422 441654
rect 332186 441098 332422 441334
rect 332186 405418 332422 405654
rect 332186 405098 332422 405334
rect 332186 369418 332422 369654
rect 332186 369098 332422 369334
rect 332186 333418 332422 333654
rect 332186 333098 332422 333334
rect 332186 297418 332422 297654
rect 332186 297098 332422 297334
rect 332186 261418 332422 261654
rect 332186 261098 332422 261334
rect 332186 225418 332422 225654
rect 332186 225098 332422 225334
rect 332186 189418 332422 189654
rect 332186 189098 332422 189334
rect 332186 153418 332422 153654
rect 332186 153098 332422 153334
rect 332186 117418 332422 117654
rect 332186 117098 332422 117334
rect 332186 81418 332422 81654
rect 332186 81098 332422 81334
rect 332186 45418 332422 45654
rect 332186 45098 332422 45334
rect 332186 9418 332422 9654
rect 332186 9098 332422 9334
rect 332186 -4262 332422 -4026
rect 332186 -4582 332422 -4346
rect 353786 711042 354022 711278
rect 353786 710722 354022 710958
rect 350186 709202 350422 709438
rect 350186 708882 350422 709118
rect 346586 707362 346822 707598
rect 346586 707042 346822 707278
rect 335786 697018 336022 697254
rect 335786 696698 336022 696934
rect 335786 661018 336022 661254
rect 335786 660698 336022 660934
rect 335786 625018 336022 625254
rect 335786 624698 336022 624934
rect 335786 589018 336022 589254
rect 335786 588698 336022 588934
rect 335786 553018 336022 553254
rect 335786 552698 336022 552934
rect 335786 517018 336022 517254
rect 335786 516698 336022 516934
rect 335786 481018 336022 481254
rect 335786 480698 336022 480934
rect 335786 445018 336022 445254
rect 335786 444698 336022 444934
rect 335786 409018 336022 409254
rect 335786 408698 336022 408934
rect 335786 373018 336022 373254
rect 335786 372698 336022 372934
rect 335786 337018 336022 337254
rect 335786 336698 336022 336934
rect 335786 301018 336022 301254
rect 335786 300698 336022 300934
rect 335786 265018 336022 265254
rect 335786 264698 336022 264934
rect 335786 229018 336022 229254
rect 335786 228698 336022 228934
rect 335786 193018 336022 193254
rect 335786 192698 336022 192934
rect 335786 157018 336022 157254
rect 335786 156698 336022 156934
rect 335786 121018 336022 121254
rect 335786 120698 336022 120934
rect 335786 85018 336022 85254
rect 335786 84698 336022 84934
rect 335786 49018 336022 49254
rect 335786 48698 336022 48934
rect 335786 13018 336022 13254
rect 335786 12698 336022 12934
rect 317786 -7022 318022 -6786
rect 317786 -7342 318022 -7106
rect 342986 705522 343222 705758
rect 342986 705202 343222 705438
rect 342986 668218 343222 668454
rect 342986 667898 343222 668134
rect 342986 632218 343222 632454
rect 342986 631898 343222 632134
rect 342986 596218 343222 596454
rect 342986 595898 343222 596134
rect 342986 560218 343222 560454
rect 342986 559898 343222 560134
rect 342986 524218 343222 524454
rect 342986 523898 343222 524134
rect 342986 488218 343222 488454
rect 342986 487898 343222 488134
rect 342986 452218 343222 452454
rect 342986 451898 343222 452134
rect 342986 416218 343222 416454
rect 342986 415898 343222 416134
rect 342986 380218 343222 380454
rect 342986 379898 343222 380134
rect 342986 344218 343222 344454
rect 342986 343898 343222 344134
rect 342986 308218 343222 308454
rect 342986 307898 343222 308134
rect 342986 272218 343222 272454
rect 342986 271898 343222 272134
rect 342986 236218 343222 236454
rect 342986 235898 343222 236134
rect 342986 200218 343222 200454
rect 342986 199898 343222 200134
rect 342986 164218 343222 164454
rect 342986 163898 343222 164134
rect 342986 128218 343222 128454
rect 342986 127898 343222 128134
rect 342986 92218 343222 92454
rect 342986 91898 343222 92134
rect 342986 56218 343222 56454
rect 342986 55898 343222 56134
rect 342986 20218 343222 20454
rect 342986 19898 343222 20134
rect 342986 -1502 343222 -1266
rect 342986 -1822 343222 -1586
rect 346586 671818 346822 672054
rect 346586 671498 346822 671734
rect 346586 635818 346822 636054
rect 346586 635498 346822 635734
rect 346586 599818 346822 600054
rect 346586 599498 346822 599734
rect 346586 563818 346822 564054
rect 346586 563498 346822 563734
rect 346586 527818 346822 528054
rect 346586 527498 346822 527734
rect 346586 491818 346822 492054
rect 346586 491498 346822 491734
rect 346586 455818 346822 456054
rect 346586 455498 346822 455734
rect 346586 419818 346822 420054
rect 346586 419498 346822 419734
rect 346586 383818 346822 384054
rect 346586 383498 346822 383734
rect 346586 347818 346822 348054
rect 346586 347498 346822 347734
rect 346586 311818 346822 312054
rect 346586 311498 346822 311734
rect 346586 275818 346822 276054
rect 346586 275498 346822 275734
rect 346586 239818 346822 240054
rect 346586 239498 346822 239734
rect 346586 203818 346822 204054
rect 346586 203498 346822 203734
rect 346586 167818 346822 168054
rect 346586 167498 346822 167734
rect 346586 131818 346822 132054
rect 346586 131498 346822 131734
rect 346586 95818 346822 96054
rect 346586 95498 346822 95734
rect 346586 59818 346822 60054
rect 346586 59498 346822 59734
rect 346586 23818 346822 24054
rect 346586 23498 346822 23734
rect 346586 -3342 346822 -3106
rect 346586 -3662 346822 -3426
rect 350186 675418 350422 675654
rect 350186 675098 350422 675334
rect 350186 639418 350422 639654
rect 350186 639098 350422 639334
rect 350186 603418 350422 603654
rect 350186 603098 350422 603334
rect 350186 567418 350422 567654
rect 350186 567098 350422 567334
rect 350186 531418 350422 531654
rect 350186 531098 350422 531334
rect 350186 495418 350422 495654
rect 350186 495098 350422 495334
rect 350186 459418 350422 459654
rect 350186 459098 350422 459334
rect 350186 423418 350422 423654
rect 350186 423098 350422 423334
rect 350186 387418 350422 387654
rect 350186 387098 350422 387334
rect 350186 351418 350422 351654
rect 350186 351098 350422 351334
rect 350186 315418 350422 315654
rect 350186 315098 350422 315334
rect 350186 279418 350422 279654
rect 350186 279098 350422 279334
rect 350186 243418 350422 243654
rect 350186 243098 350422 243334
rect 350186 207418 350422 207654
rect 350186 207098 350422 207334
rect 350186 171418 350422 171654
rect 350186 171098 350422 171334
rect 350186 135418 350422 135654
rect 350186 135098 350422 135334
rect 350186 99418 350422 99654
rect 350186 99098 350422 99334
rect 350186 63418 350422 63654
rect 350186 63098 350422 63334
rect 350186 27418 350422 27654
rect 350186 27098 350422 27334
rect 350186 -5182 350422 -4946
rect 350186 -5502 350422 -5266
rect 371786 710122 372022 710358
rect 371786 709802 372022 710038
rect 368186 708282 368422 708518
rect 368186 707962 368422 708198
rect 364586 706442 364822 706678
rect 364586 706122 364822 706358
rect 353786 679018 354022 679254
rect 353786 678698 354022 678934
rect 353786 643018 354022 643254
rect 353786 642698 354022 642934
rect 353786 607018 354022 607254
rect 353786 606698 354022 606934
rect 353786 571018 354022 571254
rect 353786 570698 354022 570934
rect 353786 535018 354022 535254
rect 353786 534698 354022 534934
rect 353786 499018 354022 499254
rect 353786 498698 354022 498934
rect 353786 463018 354022 463254
rect 353786 462698 354022 462934
rect 353786 427018 354022 427254
rect 353786 426698 354022 426934
rect 353786 391018 354022 391254
rect 353786 390698 354022 390934
rect 353786 355018 354022 355254
rect 353786 354698 354022 354934
rect 360986 704602 361222 704838
rect 360986 704282 361222 704518
rect 360986 686218 361222 686454
rect 360986 685898 361222 686134
rect 360986 650218 361222 650454
rect 360986 649898 361222 650134
rect 360986 614218 361222 614454
rect 360986 613898 361222 614134
rect 360986 578218 361222 578454
rect 360986 577898 361222 578134
rect 360986 542218 361222 542454
rect 360986 541898 361222 542134
rect 360986 506218 361222 506454
rect 360986 505898 361222 506134
rect 360986 470218 361222 470454
rect 360986 469898 361222 470134
rect 360986 434218 361222 434454
rect 360986 433898 361222 434134
rect 360986 398218 361222 398454
rect 360986 397898 361222 398134
rect 360986 362218 361222 362454
rect 360986 361898 361222 362134
rect 360986 326218 361222 326454
rect 360986 325898 361222 326134
rect 353786 319018 354022 319254
rect 353786 318698 354022 318934
rect 353786 283018 354022 283254
rect 353786 282698 354022 282934
rect 353786 247018 354022 247254
rect 353786 246698 354022 246934
rect 353786 211018 354022 211254
rect 353786 210698 354022 210934
rect 353786 175018 354022 175254
rect 353786 174698 354022 174934
rect 353786 139018 354022 139254
rect 353786 138698 354022 138934
rect 353786 103018 354022 103254
rect 353786 102698 354022 102934
rect 353786 67018 354022 67254
rect 353786 66698 354022 66934
rect 353786 31018 354022 31254
rect 353786 30698 354022 30934
rect 335786 -6102 336022 -5866
rect 335786 -6422 336022 -6186
rect 360986 290218 361222 290454
rect 360986 289898 361222 290134
rect 360986 254218 361222 254454
rect 360986 253898 361222 254134
rect 360986 218218 361222 218454
rect 360986 217898 361222 218134
rect 360986 182218 361222 182454
rect 360986 181898 361222 182134
rect 360986 146218 361222 146454
rect 360986 145898 361222 146134
rect 360986 110218 361222 110454
rect 360986 109898 361222 110134
rect 360986 74218 361222 74454
rect 360986 73898 361222 74134
rect 360986 38218 361222 38454
rect 360986 37898 361222 38134
rect 360986 2218 361222 2454
rect 360986 1898 361222 2134
rect 360986 -582 361222 -346
rect 360986 -902 361222 -666
rect 364586 689818 364822 690054
rect 364586 689498 364822 689734
rect 364586 653818 364822 654054
rect 364586 653498 364822 653734
rect 364586 617818 364822 618054
rect 364586 617498 364822 617734
rect 364586 581818 364822 582054
rect 364586 581498 364822 581734
rect 364586 545818 364822 546054
rect 364586 545498 364822 545734
rect 364586 509818 364822 510054
rect 364586 509498 364822 509734
rect 364586 473818 364822 474054
rect 364586 473498 364822 473734
rect 364586 437818 364822 438054
rect 364586 437498 364822 437734
rect 364586 401818 364822 402054
rect 364586 401498 364822 401734
rect 364586 365818 364822 366054
rect 364586 365498 364822 365734
rect 364586 329818 364822 330054
rect 364586 329498 364822 329734
rect 364586 293818 364822 294054
rect 364586 293498 364822 293734
rect 364586 257818 364822 258054
rect 364586 257498 364822 257734
rect 364586 221818 364822 222054
rect 364586 221498 364822 221734
rect 364586 185818 364822 186054
rect 364586 185498 364822 185734
rect 364586 149818 364822 150054
rect 364586 149498 364822 149734
rect 364586 113818 364822 114054
rect 364586 113498 364822 113734
rect 364586 77818 364822 78054
rect 364586 77498 364822 77734
rect 364586 41818 364822 42054
rect 364586 41498 364822 41734
rect 364586 5818 364822 6054
rect 364586 5498 364822 5734
rect 364586 -2422 364822 -2186
rect 364586 -2742 364822 -2506
rect 368186 693418 368422 693654
rect 368186 693098 368422 693334
rect 368186 657418 368422 657654
rect 368186 657098 368422 657334
rect 368186 621418 368422 621654
rect 368186 621098 368422 621334
rect 368186 585418 368422 585654
rect 368186 585098 368422 585334
rect 368186 549418 368422 549654
rect 368186 549098 368422 549334
rect 368186 513418 368422 513654
rect 368186 513098 368422 513334
rect 368186 477418 368422 477654
rect 368186 477098 368422 477334
rect 368186 441418 368422 441654
rect 368186 441098 368422 441334
rect 368186 405418 368422 405654
rect 368186 405098 368422 405334
rect 368186 369418 368422 369654
rect 368186 369098 368422 369334
rect 368186 333418 368422 333654
rect 368186 333098 368422 333334
rect 368186 297418 368422 297654
rect 368186 297098 368422 297334
rect 368186 261418 368422 261654
rect 368186 261098 368422 261334
rect 368186 225418 368422 225654
rect 368186 225098 368422 225334
rect 368186 189418 368422 189654
rect 368186 189098 368422 189334
rect 368186 153418 368422 153654
rect 368186 153098 368422 153334
rect 368186 117418 368422 117654
rect 368186 117098 368422 117334
rect 368186 81418 368422 81654
rect 368186 81098 368422 81334
rect 368186 45418 368422 45654
rect 368186 45098 368422 45334
rect 368186 9418 368422 9654
rect 368186 9098 368422 9334
rect 368186 -4262 368422 -4026
rect 368186 -4582 368422 -4346
rect 389786 711042 390022 711278
rect 389786 710722 390022 710958
rect 386186 709202 386422 709438
rect 386186 708882 386422 709118
rect 382586 707362 382822 707598
rect 382586 707042 382822 707278
rect 371786 697018 372022 697254
rect 371786 696698 372022 696934
rect 371786 661018 372022 661254
rect 371786 660698 372022 660934
rect 371786 625018 372022 625254
rect 371786 624698 372022 624934
rect 371786 589018 372022 589254
rect 371786 588698 372022 588934
rect 371786 553018 372022 553254
rect 371786 552698 372022 552934
rect 371786 517018 372022 517254
rect 371786 516698 372022 516934
rect 371786 481018 372022 481254
rect 371786 480698 372022 480934
rect 371786 445018 372022 445254
rect 371786 444698 372022 444934
rect 371786 409018 372022 409254
rect 371786 408698 372022 408934
rect 371786 373018 372022 373254
rect 371786 372698 372022 372934
rect 371786 337018 372022 337254
rect 371786 336698 372022 336934
rect 371786 301018 372022 301254
rect 371786 300698 372022 300934
rect 371786 265018 372022 265254
rect 371786 264698 372022 264934
rect 371786 229018 372022 229254
rect 371786 228698 372022 228934
rect 371786 193018 372022 193254
rect 371786 192698 372022 192934
rect 371786 157018 372022 157254
rect 371786 156698 372022 156934
rect 371786 121018 372022 121254
rect 371786 120698 372022 120934
rect 371786 85018 372022 85254
rect 371786 84698 372022 84934
rect 371786 49018 372022 49254
rect 371786 48698 372022 48934
rect 371786 13018 372022 13254
rect 371786 12698 372022 12934
rect 353786 -7022 354022 -6786
rect 353786 -7342 354022 -7106
rect 378986 705522 379222 705758
rect 378986 705202 379222 705438
rect 378986 668218 379222 668454
rect 378986 667898 379222 668134
rect 378986 632218 379222 632454
rect 378986 631898 379222 632134
rect 378986 596218 379222 596454
rect 378986 595898 379222 596134
rect 378986 560218 379222 560454
rect 378986 559898 379222 560134
rect 378986 524218 379222 524454
rect 378986 523898 379222 524134
rect 378986 488218 379222 488454
rect 378986 487898 379222 488134
rect 378986 452218 379222 452454
rect 378986 451898 379222 452134
rect 378986 416218 379222 416454
rect 378986 415898 379222 416134
rect 378986 380218 379222 380454
rect 378986 379898 379222 380134
rect 378986 344218 379222 344454
rect 378986 343898 379222 344134
rect 378986 308218 379222 308454
rect 378986 307898 379222 308134
rect 378986 272218 379222 272454
rect 378986 271898 379222 272134
rect 378986 236218 379222 236454
rect 378986 235898 379222 236134
rect 378986 200218 379222 200454
rect 378986 199898 379222 200134
rect 378986 164218 379222 164454
rect 378986 163898 379222 164134
rect 378986 128218 379222 128454
rect 378986 127898 379222 128134
rect 378986 92218 379222 92454
rect 378986 91898 379222 92134
rect 378986 56218 379222 56454
rect 378986 55898 379222 56134
rect 378986 20218 379222 20454
rect 378986 19898 379222 20134
rect 378986 -1502 379222 -1266
rect 378986 -1822 379222 -1586
rect 382586 671818 382822 672054
rect 382586 671498 382822 671734
rect 382586 635818 382822 636054
rect 382586 635498 382822 635734
rect 382586 599818 382822 600054
rect 382586 599498 382822 599734
rect 382586 563818 382822 564054
rect 382586 563498 382822 563734
rect 382586 527818 382822 528054
rect 382586 527498 382822 527734
rect 382586 491818 382822 492054
rect 382586 491498 382822 491734
rect 382586 455818 382822 456054
rect 382586 455498 382822 455734
rect 382586 419818 382822 420054
rect 382586 419498 382822 419734
rect 382586 383818 382822 384054
rect 382586 383498 382822 383734
rect 382586 347818 382822 348054
rect 382586 347498 382822 347734
rect 382586 311818 382822 312054
rect 382586 311498 382822 311734
rect 382586 275818 382822 276054
rect 382586 275498 382822 275734
rect 382586 239818 382822 240054
rect 382586 239498 382822 239734
rect 382586 203818 382822 204054
rect 382586 203498 382822 203734
rect 382586 167818 382822 168054
rect 382586 167498 382822 167734
rect 382586 131818 382822 132054
rect 382586 131498 382822 131734
rect 382586 95818 382822 96054
rect 382586 95498 382822 95734
rect 382586 59818 382822 60054
rect 382586 59498 382822 59734
rect 382586 23818 382822 24054
rect 382586 23498 382822 23734
rect 382586 -3342 382822 -3106
rect 382586 -3662 382822 -3426
rect 386186 675418 386422 675654
rect 386186 675098 386422 675334
rect 386186 639418 386422 639654
rect 386186 639098 386422 639334
rect 386186 603418 386422 603654
rect 386186 603098 386422 603334
rect 386186 567418 386422 567654
rect 386186 567098 386422 567334
rect 386186 531418 386422 531654
rect 386186 531098 386422 531334
rect 386186 495418 386422 495654
rect 386186 495098 386422 495334
rect 386186 459418 386422 459654
rect 386186 459098 386422 459334
rect 386186 423418 386422 423654
rect 386186 423098 386422 423334
rect 386186 387418 386422 387654
rect 386186 387098 386422 387334
rect 386186 351418 386422 351654
rect 386186 351098 386422 351334
rect 386186 315418 386422 315654
rect 386186 315098 386422 315334
rect 386186 279418 386422 279654
rect 386186 279098 386422 279334
rect 386186 243418 386422 243654
rect 386186 243098 386422 243334
rect 386186 207418 386422 207654
rect 386186 207098 386422 207334
rect 386186 171418 386422 171654
rect 386186 171098 386422 171334
rect 386186 135418 386422 135654
rect 386186 135098 386422 135334
rect 386186 99418 386422 99654
rect 386186 99098 386422 99334
rect 386186 63418 386422 63654
rect 386186 63098 386422 63334
rect 386186 27418 386422 27654
rect 386186 27098 386422 27334
rect 386186 -5182 386422 -4946
rect 386186 -5502 386422 -5266
rect 407786 710122 408022 710358
rect 407786 709802 408022 710038
rect 404186 708282 404422 708518
rect 404186 707962 404422 708198
rect 400586 706442 400822 706678
rect 400586 706122 400822 706358
rect 389786 679018 390022 679254
rect 389786 678698 390022 678934
rect 389786 643018 390022 643254
rect 389786 642698 390022 642934
rect 389786 607018 390022 607254
rect 389786 606698 390022 606934
rect 389786 571018 390022 571254
rect 389786 570698 390022 570934
rect 389786 535018 390022 535254
rect 389786 534698 390022 534934
rect 389786 499018 390022 499254
rect 389786 498698 390022 498934
rect 389786 463018 390022 463254
rect 389786 462698 390022 462934
rect 389786 427018 390022 427254
rect 389786 426698 390022 426934
rect 389786 391018 390022 391254
rect 389786 390698 390022 390934
rect 389786 355018 390022 355254
rect 389786 354698 390022 354934
rect 396986 704602 397222 704838
rect 396986 704282 397222 704518
rect 396986 686218 397222 686454
rect 396986 685898 397222 686134
rect 396986 650218 397222 650454
rect 396986 649898 397222 650134
rect 396986 614218 397222 614454
rect 396986 613898 397222 614134
rect 396986 578218 397222 578454
rect 396986 577898 397222 578134
rect 396986 542218 397222 542454
rect 396986 541898 397222 542134
rect 396986 506218 397222 506454
rect 396986 505898 397222 506134
rect 396986 470218 397222 470454
rect 396986 469898 397222 470134
rect 396986 434218 397222 434454
rect 396986 433898 397222 434134
rect 396986 398218 397222 398454
rect 396986 397898 397222 398134
rect 396986 362218 397222 362454
rect 396986 361898 397222 362134
rect 396986 326218 397222 326454
rect 396986 325898 397222 326134
rect 389786 319018 390022 319254
rect 389786 318698 390022 318934
rect 389786 283018 390022 283254
rect 389786 282698 390022 282934
rect 389786 247018 390022 247254
rect 389786 246698 390022 246934
rect 389786 211018 390022 211254
rect 389786 210698 390022 210934
rect 389786 175018 390022 175254
rect 389786 174698 390022 174934
rect 389786 139018 390022 139254
rect 389786 138698 390022 138934
rect 389786 103018 390022 103254
rect 389786 102698 390022 102934
rect 389786 67018 390022 67254
rect 389786 66698 390022 66934
rect 389786 31018 390022 31254
rect 389786 30698 390022 30934
rect 371786 -6102 372022 -5866
rect 371786 -6422 372022 -6186
rect 396986 290218 397222 290454
rect 396986 289898 397222 290134
rect 396986 254218 397222 254454
rect 396986 253898 397222 254134
rect 396986 218218 397222 218454
rect 396986 217898 397222 218134
rect 396986 182218 397222 182454
rect 396986 181898 397222 182134
rect 396986 146218 397222 146454
rect 396986 145898 397222 146134
rect 396986 110218 397222 110454
rect 396986 109898 397222 110134
rect 396986 74218 397222 74454
rect 396986 73898 397222 74134
rect 396986 38218 397222 38454
rect 396986 37898 397222 38134
rect 396986 2218 397222 2454
rect 396986 1898 397222 2134
rect 396986 -582 397222 -346
rect 396986 -902 397222 -666
rect 400586 689818 400822 690054
rect 400586 689498 400822 689734
rect 400586 653818 400822 654054
rect 400586 653498 400822 653734
rect 400586 617818 400822 618054
rect 400586 617498 400822 617734
rect 400586 581818 400822 582054
rect 400586 581498 400822 581734
rect 400586 545818 400822 546054
rect 400586 545498 400822 545734
rect 400586 509818 400822 510054
rect 400586 509498 400822 509734
rect 400586 473818 400822 474054
rect 400586 473498 400822 473734
rect 400586 437818 400822 438054
rect 400586 437498 400822 437734
rect 400586 401818 400822 402054
rect 400586 401498 400822 401734
rect 400586 365818 400822 366054
rect 400586 365498 400822 365734
rect 400586 329818 400822 330054
rect 400586 329498 400822 329734
rect 400586 293818 400822 294054
rect 400586 293498 400822 293734
rect 400586 257818 400822 258054
rect 400586 257498 400822 257734
rect 400586 221818 400822 222054
rect 400586 221498 400822 221734
rect 400586 185818 400822 186054
rect 400586 185498 400822 185734
rect 400586 149818 400822 150054
rect 400586 149498 400822 149734
rect 400586 113818 400822 114054
rect 400586 113498 400822 113734
rect 400586 77818 400822 78054
rect 400586 77498 400822 77734
rect 400586 41818 400822 42054
rect 400586 41498 400822 41734
rect 400586 5818 400822 6054
rect 400586 5498 400822 5734
rect 400586 -2422 400822 -2186
rect 400586 -2742 400822 -2506
rect 404186 693418 404422 693654
rect 404186 693098 404422 693334
rect 404186 657418 404422 657654
rect 404186 657098 404422 657334
rect 404186 621418 404422 621654
rect 404186 621098 404422 621334
rect 404186 585418 404422 585654
rect 404186 585098 404422 585334
rect 404186 549418 404422 549654
rect 404186 549098 404422 549334
rect 404186 513418 404422 513654
rect 404186 513098 404422 513334
rect 404186 477418 404422 477654
rect 404186 477098 404422 477334
rect 404186 441418 404422 441654
rect 404186 441098 404422 441334
rect 404186 405418 404422 405654
rect 404186 405098 404422 405334
rect 404186 369418 404422 369654
rect 404186 369098 404422 369334
rect 404186 333418 404422 333654
rect 404186 333098 404422 333334
rect 404186 297418 404422 297654
rect 404186 297098 404422 297334
rect 404186 261418 404422 261654
rect 404186 261098 404422 261334
rect 404186 225418 404422 225654
rect 404186 225098 404422 225334
rect 404186 189418 404422 189654
rect 404186 189098 404422 189334
rect 404186 153418 404422 153654
rect 404186 153098 404422 153334
rect 404186 117418 404422 117654
rect 404186 117098 404422 117334
rect 404186 81418 404422 81654
rect 404186 81098 404422 81334
rect 404186 45418 404422 45654
rect 404186 45098 404422 45334
rect 404186 9418 404422 9654
rect 404186 9098 404422 9334
rect 404186 -4262 404422 -4026
rect 404186 -4582 404422 -4346
rect 425786 711042 426022 711278
rect 425786 710722 426022 710958
rect 422186 709202 422422 709438
rect 422186 708882 422422 709118
rect 418586 707362 418822 707598
rect 418586 707042 418822 707278
rect 407786 697018 408022 697254
rect 407786 696698 408022 696934
rect 407786 661018 408022 661254
rect 407786 660698 408022 660934
rect 407786 625018 408022 625254
rect 407786 624698 408022 624934
rect 407786 589018 408022 589254
rect 407786 588698 408022 588934
rect 407786 553018 408022 553254
rect 407786 552698 408022 552934
rect 407786 517018 408022 517254
rect 407786 516698 408022 516934
rect 407786 481018 408022 481254
rect 407786 480698 408022 480934
rect 407786 445018 408022 445254
rect 407786 444698 408022 444934
rect 407786 409018 408022 409254
rect 407786 408698 408022 408934
rect 407786 373018 408022 373254
rect 407786 372698 408022 372934
rect 407786 337018 408022 337254
rect 407786 336698 408022 336934
rect 407786 301018 408022 301254
rect 407786 300698 408022 300934
rect 407786 265018 408022 265254
rect 407786 264698 408022 264934
rect 407786 229018 408022 229254
rect 407786 228698 408022 228934
rect 407786 193018 408022 193254
rect 407786 192698 408022 192934
rect 407786 157018 408022 157254
rect 407786 156698 408022 156934
rect 407786 121018 408022 121254
rect 407786 120698 408022 120934
rect 407786 85018 408022 85254
rect 407786 84698 408022 84934
rect 407786 49018 408022 49254
rect 407786 48698 408022 48934
rect 407786 13018 408022 13254
rect 407786 12698 408022 12934
rect 389786 -7022 390022 -6786
rect 389786 -7342 390022 -7106
rect 414986 705522 415222 705758
rect 414986 705202 415222 705438
rect 414986 668218 415222 668454
rect 414986 667898 415222 668134
rect 414986 632218 415222 632454
rect 414986 631898 415222 632134
rect 414986 596218 415222 596454
rect 414986 595898 415222 596134
rect 414986 560218 415222 560454
rect 414986 559898 415222 560134
rect 414986 524218 415222 524454
rect 414986 523898 415222 524134
rect 414986 488218 415222 488454
rect 414986 487898 415222 488134
rect 414986 452218 415222 452454
rect 414986 451898 415222 452134
rect 414986 416218 415222 416454
rect 414986 415898 415222 416134
rect 414986 380218 415222 380454
rect 414986 379898 415222 380134
rect 414986 344218 415222 344454
rect 414986 343898 415222 344134
rect 414986 308218 415222 308454
rect 414986 307898 415222 308134
rect 414986 272218 415222 272454
rect 414986 271898 415222 272134
rect 414986 236218 415222 236454
rect 414986 235898 415222 236134
rect 414986 200218 415222 200454
rect 414986 199898 415222 200134
rect 414986 164218 415222 164454
rect 414986 163898 415222 164134
rect 414986 128218 415222 128454
rect 414986 127898 415222 128134
rect 414986 92218 415222 92454
rect 414986 91898 415222 92134
rect 414986 56218 415222 56454
rect 414986 55898 415222 56134
rect 414986 20218 415222 20454
rect 414986 19898 415222 20134
rect 414986 -1502 415222 -1266
rect 414986 -1822 415222 -1586
rect 418586 671818 418822 672054
rect 418586 671498 418822 671734
rect 418586 635818 418822 636054
rect 418586 635498 418822 635734
rect 418586 599818 418822 600054
rect 418586 599498 418822 599734
rect 418586 563818 418822 564054
rect 418586 563498 418822 563734
rect 418586 527818 418822 528054
rect 418586 527498 418822 527734
rect 418586 491818 418822 492054
rect 418586 491498 418822 491734
rect 418586 455818 418822 456054
rect 418586 455498 418822 455734
rect 418586 419818 418822 420054
rect 418586 419498 418822 419734
rect 418586 383818 418822 384054
rect 418586 383498 418822 383734
rect 418586 347818 418822 348054
rect 418586 347498 418822 347734
rect 418586 311818 418822 312054
rect 418586 311498 418822 311734
rect 418586 275818 418822 276054
rect 418586 275498 418822 275734
rect 418586 239818 418822 240054
rect 418586 239498 418822 239734
rect 418586 203818 418822 204054
rect 418586 203498 418822 203734
rect 418586 167818 418822 168054
rect 418586 167498 418822 167734
rect 418586 131818 418822 132054
rect 418586 131498 418822 131734
rect 418586 95818 418822 96054
rect 418586 95498 418822 95734
rect 418586 59818 418822 60054
rect 418586 59498 418822 59734
rect 418586 23818 418822 24054
rect 418586 23498 418822 23734
rect 418586 -3342 418822 -3106
rect 418586 -3662 418822 -3426
rect 422186 675418 422422 675654
rect 422186 675098 422422 675334
rect 422186 639418 422422 639654
rect 422186 639098 422422 639334
rect 422186 603418 422422 603654
rect 422186 603098 422422 603334
rect 422186 567418 422422 567654
rect 422186 567098 422422 567334
rect 422186 531418 422422 531654
rect 422186 531098 422422 531334
rect 422186 495418 422422 495654
rect 422186 495098 422422 495334
rect 422186 459418 422422 459654
rect 422186 459098 422422 459334
rect 422186 423418 422422 423654
rect 422186 423098 422422 423334
rect 422186 387418 422422 387654
rect 422186 387098 422422 387334
rect 422186 351418 422422 351654
rect 422186 351098 422422 351334
rect 422186 315418 422422 315654
rect 422186 315098 422422 315334
rect 422186 279418 422422 279654
rect 422186 279098 422422 279334
rect 422186 243418 422422 243654
rect 422186 243098 422422 243334
rect 422186 207418 422422 207654
rect 422186 207098 422422 207334
rect 422186 171418 422422 171654
rect 422186 171098 422422 171334
rect 422186 135418 422422 135654
rect 422186 135098 422422 135334
rect 422186 99418 422422 99654
rect 422186 99098 422422 99334
rect 422186 63418 422422 63654
rect 422186 63098 422422 63334
rect 422186 27418 422422 27654
rect 422186 27098 422422 27334
rect 422186 -5182 422422 -4946
rect 422186 -5502 422422 -5266
rect 443786 710122 444022 710358
rect 443786 709802 444022 710038
rect 440186 708282 440422 708518
rect 440186 707962 440422 708198
rect 436586 706442 436822 706678
rect 436586 706122 436822 706358
rect 425786 679018 426022 679254
rect 425786 678698 426022 678934
rect 425786 643018 426022 643254
rect 425786 642698 426022 642934
rect 425786 607018 426022 607254
rect 425786 606698 426022 606934
rect 425786 571018 426022 571254
rect 425786 570698 426022 570934
rect 425786 535018 426022 535254
rect 425786 534698 426022 534934
rect 425786 499018 426022 499254
rect 425786 498698 426022 498934
rect 425786 463018 426022 463254
rect 425786 462698 426022 462934
rect 425786 427018 426022 427254
rect 425786 426698 426022 426934
rect 425786 391018 426022 391254
rect 425786 390698 426022 390934
rect 425786 355018 426022 355254
rect 425786 354698 426022 354934
rect 425786 319018 426022 319254
rect 425786 318698 426022 318934
rect 425786 283018 426022 283254
rect 425786 282698 426022 282934
rect 425786 247018 426022 247254
rect 425786 246698 426022 246934
rect 425786 211018 426022 211254
rect 425786 210698 426022 210934
rect 425786 175018 426022 175254
rect 425786 174698 426022 174934
rect 425786 139018 426022 139254
rect 425786 138698 426022 138934
rect 425786 103018 426022 103254
rect 425786 102698 426022 102934
rect 425786 67018 426022 67254
rect 425786 66698 426022 66934
rect 425786 31018 426022 31254
rect 425786 30698 426022 30934
rect 407786 -6102 408022 -5866
rect 407786 -6422 408022 -6186
rect 432986 704602 433222 704838
rect 432986 704282 433222 704518
rect 432986 686218 433222 686454
rect 432986 685898 433222 686134
rect 432986 650218 433222 650454
rect 432986 649898 433222 650134
rect 432986 614218 433222 614454
rect 432986 613898 433222 614134
rect 432986 578218 433222 578454
rect 432986 577898 433222 578134
rect 432986 542218 433222 542454
rect 432986 541898 433222 542134
rect 432986 506218 433222 506454
rect 432986 505898 433222 506134
rect 432986 470218 433222 470454
rect 432986 469898 433222 470134
rect 432986 434218 433222 434454
rect 432986 433898 433222 434134
rect 432986 398218 433222 398454
rect 432986 397898 433222 398134
rect 432986 362218 433222 362454
rect 432986 361898 433222 362134
rect 432986 326218 433222 326454
rect 432986 325898 433222 326134
rect 432986 290218 433222 290454
rect 432986 289898 433222 290134
rect 432986 254218 433222 254454
rect 432986 253898 433222 254134
rect 432986 218218 433222 218454
rect 432986 217898 433222 218134
rect 432986 182218 433222 182454
rect 432986 181898 433222 182134
rect 432986 146218 433222 146454
rect 432986 145898 433222 146134
rect 432986 110218 433222 110454
rect 432986 109898 433222 110134
rect 432986 74218 433222 74454
rect 432986 73898 433222 74134
rect 432986 38218 433222 38454
rect 432986 37898 433222 38134
rect 432986 2218 433222 2454
rect 432986 1898 433222 2134
rect 432986 -582 433222 -346
rect 432986 -902 433222 -666
rect 436586 689818 436822 690054
rect 436586 689498 436822 689734
rect 436586 653818 436822 654054
rect 436586 653498 436822 653734
rect 436586 617818 436822 618054
rect 436586 617498 436822 617734
rect 436586 581818 436822 582054
rect 436586 581498 436822 581734
rect 436586 545818 436822 546054
rect 436586 545498 436822 545734
rect 436586 509818 436822 510054
rect 436586 509498 436822 509734
rect 436586 473818 436822 474054
rect 436586 473498 436822 473734
rect 436586 437818 436822 438054
rect 436586 437498 436822 437734
rect 436586 401818 436822 402054
rect 436586 401498 436822 401734
rect 436586 365818 436822 366054
rect 436586 365498 436822 365734
rect 436586 329818 436822 330054
rect 436586 329498 436822 329734
rect 436586 293818 436822 294054
rect 436586 293498 436822 293734
rect 436586 257818 436822 258054
rect 436586 257498 436822 257734
rect 436586 221818 436822 222054
rect 436586 221498 436822 221734
rect 436586 185818 436822 186054
rect 436586 185498 436822 185734
rect 436586 149818 436822 150054
rect 436586 149498 436822 149734
rect 436586 113818 436822 114054
rect 436586 113498 436822 113734
rect 436586 77818 436822 78054
rect 436586 77498 436822 77734
rect 436586 41818 436822 42054
rect 436586 41498 436822 41734
rect 436586 5818 436822 6054
rect 436586 5498 436822 5734
rect 436586 -2422 436822 -2186
rect 436586 -2742 436822 -2506
rect 440186 693418 440422 693654
rect 440186 693098 440422 693334
rect 440186 657418 440422 657654
rect 440186 657098 440422 657334
rect 440186 621418 440422 621654
rect 440186 621098 440422 621334
rect 440186 585418 440422 585654
rect 440186 585098 440422 585334
rect 440186 549418 440422 549654
rect 440186 549098 440422 549334
rect 440186 513418 440422 513654
rect 440186 513098 440422 513334
rect 440186 477418 440422 477654
rect 440186 477098 440422 477334
rect 440186 441418 440422 441654
rect 440186 441098 440422 441334
rect 440186 405418 440422 405654
rect 440186 405098 440422 405334
rect 440186 369418 440422 369654
rect 440186 369098 440422 369334
rect 440186 333418 440422 333654
rect 440186 333098 440422 333334
rect 440186 297418 440422 297654
rect 440186 297098 440422 297334
rect 440186 261418 440422 261654
rect 440186 261098 440422 261334
rect 440186 225418 440422 225654
rect 440186 225098 440422 225334
rect 440186 189418 440422 189654
rect 440186 189098 440422 189334
rect 440186 153418 440422 153654
rect 440186 153098 440422 153334
rect 440186 117418 440422 117654
rect 440186 117098 440422 117334
rect 440186 81418 440422 81654
rect 440186 81098 440422 81334
rect 440186 45418 440422 45654
rect 440186 45098 440422 45334
rect 440186 9418 440422 9654
rect 440186 9098 440422 9334
rect 440186 -4262 440422 -4026
rect 440186 -4582 440422 -4346
rect 461786 711042 462022 711278
rect 461786 710722 462022 710958
rect 458186 709202 458422 709438
rect 458186 708882 458422 709118
rect 454586 707362 454822 707598
rect 454586 707042 454822 707278
rect 443786 697018 444022 697254
rect 443786 696698 444022 696934
rect 443786 661018 444022 661254
rect 443786 660698 444022 660934
rect 443786 625018 444022 625254
rect 443786 624698 444022 624934
rect 443786 589018 444022 589254
rect 443786 588698 444022 588934
rect 443786 553018 444022 553254
rect 443786 552698 444022 552934
rect 443786 517018 444022 517254
rect 443786 516698 444022 516934
rect 443786 481018 444022 481254
rect 443786 480698 444022 480934
rect 443786 445018 444022 445254
rect 443786 444698 444022 444934
rect 443786 409018 444022 409254
rect 443786 408698 444022 408934
rect 443786 373018 444022 373254
rect 443786 372698 444022 372934
rect 443786 337018 444022 337254
rect 443786 336698 444022 336934
rect 443786 301018 444022 301254
rect 443786 300698 444022 300934
rect 443786 265018 444022 265254
rect 443786 264698 444022 264934
rect 443786 229018 444022 229254
rect 443786 228698 444022 228934
rect 443786 193018 444022 193254
rect 443786 192698 444022 192934
rect 443786 157018 444022 157254
rect 443786 156698 444022 156934
rect 443786 121018 444022 121254
rect 443786 120698 444022 120934
rect 443786 85018 444022 85254
rect 443786 84698 444022 84934
rect 443786 49018 444022 49254
rect 443786 48698 444022 48934
rect 443786 13018 444022 13254
rect 443786 12698 444022 12934
rect 425786 -7022 426022 -6786
rect 425786 -7342 426022 -7106
rect 450986 705522 451222 705758
rect 450986 705202 451222 705438
rect 450986 668218 451222 668454
rect 450986 667898 451222 668134
rect 450986 632218 451222 632454
rect 450986 631898 451222 632134
rect 450986 596218 451222 596454
rect 450986 595898 451222 596134
rect 450986 560218 451222 560454
rect 450986 559898 451222 560134
rect 450986 524218 451222 524454
rect 450986 523898 451222 524134
rect 450986 488218 451222 488454
rect 450986 487898 451222 488134
rect 450986 452218 451222 452454
rect 450986 451898 451222 452134
rect 450986 416218 451222 416454
rect 450986 415898 451222 416134
rect 450986 380218 451222 380454
rect 450986 379898 451222 380134
rect 450986 344218 451222 344454
rect 450986 343898 451222 344134
rect 450986 308218 451222 308454
rect 450986 307898 451222 308134
rect 450986 272218 451222 272454
rect 450986 271898 451222 272134
rect 450986 236218 451222 236454
rect 450986 235898 451222 236134
rect 450986 200218 451222 200454
rect 450986 199898 451222 200134
rect 450986 164218 451222 164454
rect 450986 163898 451222 164134
rect 450986 128218 451222 128454
rect 450986 127898 451222 128134
rect 450986 92218 451222 92454
rect 450986 91898 451222 92134
rect 450986 56218 451222 56454
rect 450986 55898 451222 56134
rect 450986 20218 451222 20454
rect 450986 19898 451222 20134
rect 450986 -1502 451222 -1266
rect 450986 -1822 451222 -1586
rect 454586 671818 454822 672054
rect 454586 671498 454822 671734
rect 454586 635818 454822 636054
rect 454586 635498 454822 635734
rect 454586 599818 454822 600054
rect 454586 599498 454822 599734
rect 454586 563818 454822 564054
rect 454586 563498 454822 563734
rect 454586 527818 454822 528054
rect 454586 527498 454822 527734
rect 454586 491818 454822 492054
rect 454586 491498 454822 491734
rect 454586 455818 454822 456054
rect 454586 455498 454822 455734
rect 454586 419818 454822 420054
rect 454586 419498 454822 419734
rect 454586 383818 454822 384054
rect 454586 383498 454822 383734
rect 454586 347818 454822 348054
rect 454586 347498 454822 347734
rect 454586 311818 454822 312054
rect 454586 311498 454822 311734
rect 454586 275818 454822 276054
rect 454586 275498 454822 275734
rect 454586 239818 454822 240054
rect 454586 239498 454822 239734
rect 454586 203818 454822 204054
rect 454586 203498 454822 203734
rect 454586 167818 454822 168054
rect 454586 167498 454822 167734
rect 454586 131818 454822 132054
rect 454586 131498 454822 131734
rect 454586 95818 454822 96054
rect 454586 95498 454822 95734
rect 454586 59818 454822 60054
rect 454586 59498 454822 59734
rect 454586 23818 454822 24054
rect 454586 23498 454822 23734
rect 454586 -3342 454822 -3106
rect 454586 -3662 454822 -3426
rect 458186 675418 458422 675654
rect 458186 675098 458422 675334
rect 458186 639418 458422 639654
rect 458186 639098 458422 639334
rect 458186 603418 458422 603654
rect 458186 603098 458422 603334
rect 458186 567418 458422 567654
rect 458186 567098 458422 567334
rect 458186 531418 458422 531654
rect 458186 531098 458422 531334
rect 458186 495418 458422 495654
rect 458186 495098 458422 495334
rect 458186 459418 458422 459654
rect 458186 459098 458422 459334
rect 458186 423418 458422 423654
rect 458186 423098 458422 423334
rect 458186 387418 458422 387654
rect 458186 387098 458422 387334
rect 458186 351418 458422 351654
rect 458186 351098 458422 351334
rect 458186 315418 458422 315654
rect 458186 315098 458422 315334
rect 458186 279418 458422 279654
rect 458186 279098 458422 279334
rect 458186 243418 458422 243654
rect 458186 243098 458422 243334
rect 458186 207418 458422 207654
rect 458186 207098 458422 207334
rect 458186 171418 458422 171654
rect 458186 171098 458422 171334
rect 458186 135418 458422 135654
rect 458186 135098 458422 135334
rect 458186 99418 458422 99654
rect 458186 99098 458422 99334
rect 458186 63418 458422 63654
rect 458186 63098 458422 63334
rect 458186 27418 458422 27654
rect 458186 27098 458422 27334
rect 458186 -5182 458422 -4946
rect 458186 -5502 458422 -5266
rect 479786 710122 480022 710358
rect 479786 709802 480022 710038
rect 476186 708282 476422 708518
rect 476186 707962 476422 708198
rect 472586 706442 472822 706678
rect 472586 706122 472822 706358
rect 461786 679018 462022 679254
rect 461786 678698 462022 678934
rect 461786 643018 462022 643254
rect 461786 642698 462022 642934
rect 461786 607018 462022 607254
rect 461786 606698 462022 606934
rect 461786 571018 462022 571254
rect 461786 570698 462022 570934
rect 461786 535018 462022 535254
rect 461786 534698 462022 534934
rect 461786 499018 462022 499254
rect 461786 498698 462022 498934
rect 461786 463018 462022 463254
rect 461786 462698 462022 462934
rect 461786 427018 462022 427254
rect 461786 426698 462022 426934
rect 461786 391018 462022 391254
rect 461786 390698 462022 390934
rect 461786 355018 462022 355254
rect 461786 354698 462022 354934
rect 461786 319018 462022 319254
rect 461786 318698 462022 318934
rect 461786 283018 462022 283254
rect 461786 282698 462022 282934
rect 461786 247018 462022 247254
rect 461786 246698 462022 246934
rect 461786 211018 462022 211254
rect 461786 210698 462022 210934
rect 461786 175018 462022 175254
rect 461786 174698 462022 174934
rect 461786 139018 462022 139254
rect 461786 138698 462022 138934
rect 461786 103018 462022 103254
rect 461786 102698 462022 102934
rect 461786 67018 462022 67254
rect 461786 66698 462022 66934
rect 461786 31018 462022 31254
rect 461786 30698 462022 30934
rect 443786 -6102 444022 -5866
rect 443786 -6422 444022 -6186
rect 468986 704602 469222 704838
rect 468986 704282 469222 704518
rect 468986 686218 469222 686454
rect 468986 685898 469222 686134
rect 468986 650218 469222 650454
rect 468986 649898 469222 650134
rect 468986 614218 469222 614454
rect 468986 613898 469222 614134
rect 468986 578218 469222 578454
rect 468986 577898 469222 578134
rect 468986 542218 469222 542454
rect 468986 541898 469222 542134
rect 468986 506218 469222 506454
rect 468986 505898 469222 506134
rect 468986 470218 469222 470454
rect 468986 469898 469222 470134
rect 468986 434218 469222 434454
rect 468986 433898 469222 434134
rect 468986 398218 469222 398454
rect 468986 397898 469222 398134
rect 468986 362218 469222 362454
rect 468986 361898 469222 362134
rect 468986 326218 469222 326454
rect 468986 325898 469222 326134
rect 468986 290218 469222 290454
rect 468986 289898 469222 290134
rect 468986 254218 469222 254454
rect 468986 253898 469222 254134
rect 468986 218218 469222 218454
rect 468986 217898 469222 218134
rect 468986 182218 469222 182454
rect 468986 181898 469222 182134
rect 468986 146218 469222 146454
rect 468986 145898 469222 146134
rect 468986 110218 469222 110454
rect 468986 109898 469222 110134
rect 468986 74218 469222 74454
rect 468986 73898 469222 74134
rect 468986 38218 469222 38454
rect 468986 37898 469222 38134
rect 468986 2218 469222 2454
rect 468986 1898 469222 2134
rect 468986 -582 469222 -346
rect 468986 -902 469222 -666
rect 472586 689818 472822 690054
rect 472586 689498 472822 689734
rect 472586 653818 472822 654054
rect 472586 653498 472822 653734
rect 472586 617818 472822 618054
rect 472586 617498 472822 617734
rect 472586 581818 472822 582054
rect 472586 581498 472822 581734
rect 472586 545818 472822 546054
rect 472586 545498 472822 545734
rect 472586 509818 472822 510054
rect 472586 509498 472822 509734
rect 472586 473818 472822 474054
rect 472586 473498 472822 473734
rect 472586 437818 472822 438054
rect 472586 437498 472822 437734
rect 472586 401818 472822 402054
rect 472586 401498 472822 401734
rect 472586 365818 472822 366054
rect 472586 365498 472822 365734
rect 472586 329818 472822 330054
rect 472586 329498 472822 329734
rect 472586 293818 472822 294054
rect 472586 293498 472822 293734
rect 472586 257818 472822 258054
rect 472586 257498 472822 257734
rect 472586 221818 472822 222054
rect 472586 221498 472822 221734
rect 472586 185818 472822 186054
rect 472586 185498 472822 185734
rect 472586 149818 472822 150054
rect 472586 149498 472822 149734
rect 472586 113818 472822 114054
rect 472586 113498 472822 113734
rect 472586 77818 472822 78054
rect 472586 77498 472822 77734
rect 472586 41818 472822 42054
rect 472586 41498 472822 41734
rect 472586 5818 472822 6054
rect 472586 5498 472822 5734
rect 472586 -2422 472822 -2186
rect 472586 -2742 472822 -2506
rect 476186 693418 476422 693654
rect 476186 693098 476422 693334
rect 476186 657418 476422 657654
rect 476186 657098 476422 657334
rect 476186 621418 476422 621654
rect 476186 621098 476422 621334
rect 476186 585418 476422 585654
rect 476186 585098 476422 585334
rect 476186 549418 476422 549654
rect 476186 549098 476422 549334
rect 476186 513418 476422 513654
rect 476186 513098 476422 513334
rect 476186 477418 476422 477654
rect 476186 477098 476422 477334
rect 476186 441418 476422 441654
rect 476186 441098 476422 441334
rect 476186 405418 476422 405654
rect 476186 405098 476422 405334
rect 476186 369418 476422 369654
rect 476186 369098 476422 369334
rect 476186 333418 476422 333654
rect 476186 333098 476422 333334
rect 476186 297418 476422 297654
rect 476186 297098 476422 297334
rect 476186 261418 476422 261654
rect 476186 261098 476422 261334
rect 476186 225418 476422 225654
rect 476186 225098 476422 225334
rect 476186 189418 476422 189654
rect 476186 189098 476422 189334
rect 476186 153418 476422 153654
rect 476186 153098 476422 153334
rect 476186 117418 476422 117654
rect 476186 117098 476422 117334
rect 476186 81418 476422 81654
rect 476186 81098 476422 81334
rect 476186 45418 476422 45654
rect 476186 45098 476422 45334
rect 476186 9418 476422 9654
rect 476186 9098 476422 9334
rect 476186 -4262 476422 -4026
rect 476186 -4582 476422 -4346
rect 497786 711042 498022 711278
rect 497786 710722 498022 710958
rect 494186 709202 494422 709438
rect 494186 708882 494422 709118
rect 490586 707362 490822 707598
rect 490586 707042 490822 707278
rect 479786 697018 480022 697254
rect 479786 696698 480022 696934
rect 479786 661018 480022 661254
rect 479786 660698 480022 660934
rect 479786 625018 480022 625254
rect 479786 624698 480022 624934
rect 479786 589018 480022 589254
rect 479786 588698 480022 588934
rect 479786 553018 480022 553254
rect 479786 552698 480022 552934
rect 479786 517018 480022 517254
rect 479786 516698 480022 516934
rect 479786 481018 480022 481254
rect 479786 480698 480022 480934
rect 479786 445018 480022 445254
rect 479786 444698 480022 444934
rect 479786 409018 480022 409254
rect 479786 408698 480022 408934
rect 479786 373018 480022 373254
rect 479786 372698 480022 372934
rect 479786 337018 480022 337254
rect 479786 336698 480022 336934
rect 479786 301018 480022 301254
rect 479786 300698 480022 300934
rect 479786 265018 480022 265254
rect 479786 264698 480022 264934
rect 479786 229018 480022 229254
rect 479786 228698 480022 228934
rect 479786 193018 480022 193254
rect 479786 192698 480022 192934
rect 479786 157018 480022 157254
rect 479786 156698 480022 156934
rect 479786 121018 480022 121254
rect 479786 120698 480022 120934
rect 479786 85018 480022 85254
rect 479786 84698 480022 84934
rect 479786 49018 480022 49254
rect 479786 48698 480022 48934
rect 486986 705522 487222 705758
rect 486986 705202 487222 705438
rect 486986 668218 487222 668454
rect 486986 667898 487222 668134
rect 486986 632218 487222 632454
rect 486986 631898 487222 632134
rect 486986 596218 487222 596454
rect 486986 595898 487222 596134
rect 486986 560218 487222 560454
rect 486986 559898 487222 560134
rect 486986 524218 487222 524454
rect 486986 523898 487222 524134
rect 486986 488218 487222 488454
rect 486986 487898 487222 488134
rect 486986 452218 487222 452454
rect 486986 451898 487222 452134
rect 486986 416218 487222 416454
rect 486986 415898 487222 416134
rect 486986 380218 487222 380454
rect 486986 379898 487222 380134
rect 486986 344218 487222 344454
rect 486986 343898 487222 344134
rect 486986 308218 487222 308454
rect 486986 307898 487222 308134
rect 486986 272218 487222 272454
rect 486986 271898 487222 272134
rect 486986 236218 487222 236454
rect 486986 235898 487222 236134
rect 486986 200218 487222 200454
rect 486986 199898 487222 200134
rect 486986 164218 487222 164454
rect 486986 163898 487222 164134
rect 486986 128218 487222 128454
rect 486986 127898 487222 128134
rect 486986 92218 487222 92454
rect 486986 91898 487222 92134
rect 486986 56218 487222 56454
rect 486986 55898 487222 56134
rect 479786 13018 480022 13254
rect 479786 12698 480022 12934
rect 461786 -7022 462022 -6786
rect 461786 -7342 462022 -7106
rect 486986 20218 487222 20454
rect 486986 19898 487222 20134
rect 486986 -1502 487222 -1266
rect 486986 -1822 487222 -1586
rect 490586 671818 490822 672054
rect 490586 671498 490822 671734
rect 490586 635818 490822 636054
rect 490586 635498 490822 635734
rect 490586 599818 490822 600054
rect 490586 599498 490822 599734
rect 490586 563818 490822 564054
rect 490586 563498 490822 563734
rect 490586 527818 490822 528054
rect 490586 527498 490822 527734
rect 490586 491818 490822 492054
rect 490586 491498 490822 491734
rect 490586 455818 490822 456054
rect 490586 455498 490822 455734
rect 490586 419818 490822 420054
rect 490586 419498 490822 419734
rect 490586 383818 490822 384054
rect 490586 383498 490822 383734
rect 490586 347818 490822 348054
rect 490586 347498 490822 347734
rect 490586 311818 490822 312054
rect 490586 311498 490822 311734
rect 490586 275818 490822 276054
rect 490586 275498 490822 275734
rect 490586 239818 490822 240054
rect 490586 239498 490822 239734
rect 490586 203818 490822 204054
rect 490586 203498 490822 203734
rect 490586 167818 490822 168054
rect 490586 167498 490822 167734
rect 490586 131818 490822 132054
rect 490586 131498 490822 131734
rect 490586 95818 490822 96054
rect 490586 95498 490822 95734
rect 494186 675418 494422 675654
rect 494186 675098 494422 675334
rect 494186 639418 494422 639654
rect 494186 639098 494422 639334
rect 494186 603418 494422 603654
rect 494186 603098 494422 603334
rect 494186 567418 494422 567654
rect 494186 567098 494422 567334
rect 494186 531418 494422 531654
rect 494186 531098 494422 531334
rect 494186 495418 494422 495654
rect 494186 495098 494422 495334
rect 494186 459418 494422 459654
rect 494186 459098 494422 459334
rect 494186 423418 494422 423654
rect 494186 423098 494422 423334
rect 494186 387418 494422 387654
rect 494186 387098 494422 387334
rect 494186 351418 494422 351654
rect 494186 351098 494422 351334
rect 494186 315418 494422 315654
rect 494186 315098 494422 315334
rect 494186 279418 494422 279654
rect 494186 279098 494422 279334
rect 494186 243418 494422 243654
rect 494186 243098 494422 243334
rect 494186 207418 494422 207654
rect 494186 207098 494422 207334
rect 494186 171418 494422 171654
rect 494186 171098 494422 171334
rect 494186 135418 494422 135654
rect 494186 135098 494422 135334
rect 494186 99418 494422 99654
rect 494186 99098 494422 99334
rect 490586 59818 490822 60054
rect 490586 59498 490822 59734
rect 490586 23818 490822 24054
rect 490586 23498 490822 23734
rect 490586 -3342 490822 -3106
rect 490586 -3662 490822 -3426
rect 494186 63418 494422 63654
rect 494186 63098 494422 63334
rect 494186 27418 494422 27654
rect 494186 27098 494422 27334
rect 494186 -5182 494422 -4946
rect 494186 -5502 494422 -5266
rect 515786 710122 516022 710358
rect 515786 709802 516022 710038
rect 512186 708282 512422 708518
rect 512186 707962 512422 708198
rect 508586 706442 508822 706678
rect 508586 706122 508822 706358
rect 497786 679018 498022 679254
rect 497786 678698 498022 678934
rect 497786 643018 498022 643254
rect 497786 642698 498022 642934
rect 497786 607018 498022 607254
rect 497786 606698 498022 606934
rect 497786 571018 498022 571254
rect 497786 570698 498022 570934
rect 497786 535018 498022 535254
rect 497786 534698 498022 534934
rect 497786 499018 498022 499254
rect 497786 498698 498022 498934
rect 497786 463018 498022 463254
rect 497786 462698 498022 462934
rect 497786 427018 498022 427254
rect 497786 426698 498022 426934
rect 497786 391018 498022 391254
rect 497786 390698 498022 390934
rect 497786 355018 498022 355254
rect 497786 354698 498022 354934
rect 497786 319018 498022 319254
rect 497786 318698 498022 318934
rect 497786 283018 498022 283254
rect 497786 282698 498022 282934
rect 497786 247018 498022 247254
rect 497786 246698 498022 246934
rect 497786 211018 498022 211254
rect 497786 210698 498022 210934
rect 497786 175018 498022 175254
rect 497786 174698 498022 174934
rect 497786 139018 498022 139254
rect 497786 138698 498022 138934
rect 497786 103018 498022 103254
rect 497786 102698 498022 102934
rect 497786 67018 498022 67254
rect 497786 66698 498022 66934
rect 497786 31018 498022 31254
rect 497786 30698 498022 30934
rect 479786 -6102 480022 -5866
rect 479786 -6422 480022 -6186
rect 504986 704602 505222 704838
rect 504986 704282 505222 704518
rect 504986 686218 505222 686454
rect 504986 685898 505222 686134
rect 504986 650218 505222 650454
rect 504986 649898 505222 650134
rect 504986 614218 505222 614454
rect 504986 613898 505222 614134
rect 504986 578218 505222 578454
rect 504986 577898 505222 578134
rect 504986 542218 505222 542454
rect 504986 541898 505222 542134
rect 504986 506218 505222 506454
rect 504986 505898 505222 506134
rect 504986 470218 505222 470454
rect 504986 469898 505222 470134
rect 504986 434218 505222 434454
rect 504986 433898 505222 434134
rect 504986 398218 505222 398454
rect 504986 397898 505222 398134
rect 504986 362218 505222 362454
rect 504986 361898 505222 362134
rect 504986 326218 505222 326454
rect 504986 325898 505222 326134
rect 504986 290218 505222 290454
rect 504986 289898 505222 290134
rect 504986 254218 505222 254454
rect 504986 253898 505222 254134
rect 504986 218218 505222 218454
rect 504986 217898 505222 218134
rect 504986 182218 505222 182454
rect 504986 181898 505222 182134
rect 504986 146218 505222 146454
rect 504986 145898 505222 146134
rect 504986 110218 505222 110454
rect 504986 109898 505222 110134
rect 504986 74218 505222 74454
rect 504986 73898 505222 74134
rect 504986 38218 505222 38454
rect 504986 37898 505222 38134
rect 504986 2218 505222 2454
rect 504986 1898 505222 2134
rect 504986 -582 505222 -346
rect 504986 -902 505222 -666
rect 508586 689818 508822 690054
rect 508586 689498 508822 689734
rect 508586 653818 508822 654054
rect 508586 653498 508822 653734
rect 508586 617818 508822 618054
rect 508586 617498 508822 617734
rect 508586 581818 508822 582054
rect 508586 581498 508822 581734
rect 508586 545818 508822 546054
rect 508586 545498 508822 545734
rect 508586 509818 508822 510054
rect 508586 509498 508822 509734
rect 508586 473818 508822 474054
rect 508586 473498 508822 473734
rect 508586 437818 508822 438054
rect 508586 437498 508822 437734
rect 508586 401818 508822 402054
rect 508586 401498 508822 401734
rect 508586 365818 508822 366054
rect 508586 365498 508822 365734
rect 508586 329818 508822 330054
rect 508586 329498 508822 329734
rect 508586 293818 508822 294054
rect 508586 293498 508822 293734
rect 508586 257818 508822 258054
rect 508586 257498 508822 257734
rect 508586 221818 508822 222054
rect 508586 221498 508822 221734
rect 508586 185818 508822 186054
rect 508586 185498 508822 185734
rect 508586 149818 508822 150054
rect 508586 149498 508822 149734
rect 508586 113818 508822 114054
rect 508586 113498 508822 113734
rect 508586 77818 508822 78054
rect 508586 77498 508822 77734
rect 508586 41818 508822 42054
rect 508586 41498 508822 41734
rect 508586 5818 508822 6054
rect 508586 5498 508822 5734
rect 508586 -2422 508822 -2186
rect 508586 -2742 508822 -2506
rect 512186 693418 512422 693654
rect 512186 693098 512422 693334
rect 512186 657418 512422 657654
rect 512186 657098 512422 657334
rect 512186 621418 512422 621654
rect 512186 621098 512422 621334
rect 512186 585418 512422 585654
rect 512186 585098 512422 585334
rect 512186 549418 512422 549654
rect 512186 549098 512422 549334
rect 512186 513418 512422 513654
rect 512186 513098 512422 513334
rect 512186 477418 512422 477654
rect 512186 477098 512422 477334
rect 512186 441418 512422 441654
rect 512186 441098 512422 441334
rect 512186 405418 512422 405654
rect 512186 405098 512422 405334
rect 512186 369418 512422 369654
rect 512186 369098 512422 369334
rect 512186 333418 512422 333654
rect 512186 333098 512422 333334
rect 512186 297418 512422 297654
rect 512186 297098 512422 297334
rect 512186 261418 512422 261654
rect 512186 261098 512422 261334
rect 512186 225418 512422 225654
rect 512186 225098 512422 225334
rect 512186 189418 512422 189654
rect 512186 189098 512422 189334
rect 512186 153418 512422 153654
rect 512186 153098 512422 153334
rect 512186 117418 512422 117654
rect 512186 117098 512422 117334
rect 512186 81418 512422 81654
rect 512186 81098 512422 81334
rect 512186 45418 512422 45654
rect 512186 45098 512422 45334
rect 512186 9418 512422 9654
rect 512186 9098 512422 9334
rect 512186 -4262 512422 -4026
rect 512186 -4582 512422 -4346
rect 533786 711042 534022 711278
rect 533786 710722 534022 710958
rect 530186 709202 530422 709438
rect 530186 708882 530422 709118
rect 526586 707362 526822 707598
rect 526586 707042 526822 707278
rect 515786 697018 516022 697254
rect 515786 696698 516022 696934
rect 515786 661018 516022 661254
rect 515786 660698 516022 660934
rect 515786 625018 516022 625254
rect 515786 624698 516022 624934
rect 515786 589018 516022 589254
rect 515786 588698 516022 588934
rect 515786 553018 516022 553254
rect 515786 552698 516022 552934
rect 515786 517018 516022 517254
rect 515786 516698 516022 516934
rect 515786 481018 516022 481254
rect 515786 480698 516022 480934
rect 515786 445018 516022 445254
rect 515786 444698 516022 444934
rect 515786 409018 516022 409254
rect 515786 408698 516022 408934
rect 515786 373018 516022 373254
rect 515786 372698 516022 372934
rect 515786 337018 516022 337254
rect 515786 336698 516022 336934
rect 515786 301018 516022 301254
rect 515786 300698 516022 300934
rect 515786 265018 516022 265254
rect 515786 264698 516022 264934
rect 515786 229018 516022 229254
rect 515786 228698 516022 228934
rect 515786 193018 516022 193254
rect 515786 192698 516022 192934
rect 515786 157018 516022 157254
rect 515786 156698 516022 156934
rect 515786 121018 516022 121254
rect 515786 120698 516022 120934
rect 515786 85018 516022 85254
rect 515786 84698 516022 84934
rect 515786 49018 516022 49254
rect 515786 48698 516022 48934
rect 515786 13018 516022 13254
rect 515786 12698 516022 12934
rect 497786 -7022 498022 -6786
rect 497786 -7342 498022 -7106
rect 522986 705522 523222 705758
rect 522986 705202 523222 705438
rect 522986 668218 523222 668454
rect 522986 667898 523222 668134
rect 522986 632218 523222 632454
rect 522986 631898 523222 632134
rect 522986 596218 523222 596454
rect 522986 595898 523222 596134
rect 522986 560218 523222 560454
rect 522986 559898 523222 560134
rect 522986 524218 523222 524454
rect 522986 523898 523222 524134
rect 522986 488218 523222 488454
rect 522986 487898 523222 488134
rect 522986 452218 523222 452454
rect 522986 451898 523222 452134
rect 522986 416218 523222 416454
rect 522986 415898 523222 416134
rect 522986 380218 523222 380454
rect 522986 379898 523222 380134
rect 522986 344218 523222 344454
rect 522986 343898 523222 344134
rect 522986 308218 523222 308454
rect 522986 307898 523222 308134
rect 522986 272218 523222 272454
rect 522986 271898 523222 272134
rect 522986 236218 523222 236454
rect 522986 235898 523222 236134
rect 522986 200218 523222 200454
rect 522986 199898 523222 200134
rect 522986 164218 523222 164454
rect 522986 163898 523222 164134
rect 522986 128218 523222 128454
rect 522986 127898 523222 128134
rect 522986 92218 523222 92454
rect 522986 91898 523222 92134
rect 522986 56218 523222 56454
rect 522986 55898 523222 56134
rect 522986 20218 523222 20454
rect 522986 19898 523222 20134
rect 522986 -1502 523222 -1266
rect 522986 -1822 523222 -1586
rect 526586 671818 526822 672054
rect 526586 671498 526822 671734
rect 526586 635818 526822 636054
rect 526586 635498 526822 635734
rect 526586 599818 526822 600054
rect 526586 599498 526822 599734
rect 526586 563818 526822 564054
rect 526586 563498 526822 563734
rect 526586 527818 526822 528054
rect 526586 527498 526822 527734
rect 526586 491818 526822 492054
rect 526586 491498 526822 491734
rect 526586 455818 526822 456054
rect 526586 455498 526822 455734
rect 526586 419818 526822 420054
rect 526586 419498 526822 419734
rect 526586 383818 526822 384054
rect 526586 383498 526822 383734
rect 526586 347818 526822 348054
rect 526586 347498 526822 347734
rect 526586 311818 526822 312054
rect 526586 311498 526822 311734
rect 526586 275818 526822 276054
rect 526586 275498 526822 275734
rect 526586 239818 526822 240054
rect 526586 239498 526822 239734
rect 526586 203818 526822 204054
rect 526586 203498 526822 203734
rect 526586 167818 526822 168054
rect 526586 167498 526822 167734
rect 526586 131818 526822 132054
rect 526586 131498 526822 131734
rect 526586 95818 526822 96054
rect 526586 95498 526822 95734
rect 526586 59818 526822 60054
rect 526586 59498 526822 59734
rect 526586 23818 526822 24054
rect 526586 23498 526822 23734
rect 526586 -3342 526822 -3106
rect 526586 -3662 526822 -3426
rect 530186 675418 530422 675654
rect 530186 675098 530422 675334
rect 530186 639418 530422 639654
rect 530186 639098 530422 639334
rect 530186 603418 530422 603654
rect 530186 603098 530422 603334
rect 530186 567418 530422 567654
rect 530186 567098 530422 567334
rect 530186 531418 530422 531654
rect 530186 531098 530422 531334
rect 530186 495418 530422 495654
rect 530186 495098 530422 495334
rect 530186 459418 530422 459654
rect 530186 459098 530422 459334
rect 530186 423418 530422 423654
rect 530186 423098 530422 423334
rect 530186 387418 530422 387654
rect 530186 387098 530422 387334
rect 530186 351418 530422 351654
rect 530186 351098 530422 351334
rect 530186 315418 530422 315654
rect 530186 315098 530422 315334
rect 530186 279418 530422 279654
rect 530186 279098 530422 279334
rect 530186 243418 530422 243654
rect 530186 243098 530422 243334
rect 530186 207418 530422 207654
rect 530186 207098 530422 207334
rect 530186 171418 530422 171654
rect 530186 171098 530422 171334
rect 530186 135418 530422 135654
rect 530186 135098 530422 135334
rect 530186 99418 530422 99654
rect 530186 99098 530422 99334
rect 530186 63418 530422 63654
rect 530186 63098 530422 63334
rect 530186 27418 530422 27654
rect 530186 27098 530422 27334
rect 530186 -5182 530422 -4946
rect 530186 -5502 530422 -5266
rect 551786 710122 552022 710358
rect 551786 709802 552022 710038
rect 548186 708282 548422 708518
rect 548186 707962 548422 708198
rect 544586 706442 544822 706678
rect 544586 706122 544822 706358
rect 533786 679018 534022 679254
rect 533786 678698 534022 678934
rect 533786 643018 534022 643254
rect 533786 642698 534022 642934
rect 533786 607018 534022 607254
rect 533786 606698 534022 606934
rect 533786 571018 534022 571254
rect 533786 570698 534022 570934
rect 533786 535018 534022 535254
rect 533786 534698 534022 534934
rect 533786 499018 534022 499254
rect 533786 498698 534022 498934
rect 533786 463018 534022 463254
rect 533786 462698 534022 462934
rect 533786 427018 534022 427254
rect 533786 426698 534022 426934
rect 533786 391018 534022 391254
rect 533786 390698 534022 390934
rect 533786 355018 534022 355254
rect 533786 354698 534022 354934
rect 533786 319018 534022 319254
rect 533786 318698 534022 318934
rect 533786 283018 534022 283254
rect 533786 282698 534022 282934
rect 533786 247018 534022 247254
rect 533786 246698 534022 246934
rect 533786 211018 534022 211254
rect 533786 210698 534022 210934
rect 533786 175018 534022 175254
rect 533786 174698 534022 174934
rect 533786 139018 534022 139254
rect 533786 138698 534022 138934
rect 533786 103018 534022 103254
rect 533786 102698 534022 102934
rect 533786 67018 534022 67254
rect 533786 66698 534022 66934
rect 533786 31018 534022 31254
rect 533786 30698 534022 30934
rect 515786 -6102 516022 -5866
rect 515786 -6422 516022 -6186
rect 540986 704602 541222 704838
rect 540986 704282 541222 704518
rect 540986 686218 541222 686454
rect 540986 685898 541222 686134
rect 540986 650218 541222 650454
rect 540986 649898 541222 650134
rect 540986 614218 541222 614454
rect 540986 613898 541222 614134
rect 540986 578218 541222 578454
rect 540986 577898 541222 578134
rect 540986 542218 541222 542454
rect 540986 541898 541222 542134
rect 540986 506218 541222 506454
rect 540986 505898 541222 506134
rect 540986 470218 541222 470454
rect 540986 469898 541222 470134
rect 540986 434218 541222 434454
rect 540986 433898 541222 434134
rect 540986 398218 541222 398454
rect 540986 397898 541222 398134
rect 540986 362218 541222 362454
rect 540986 361898 541222 362134
rect 540986 326218 541222 326454
rect 540986 325898 541222 326134
rect 540986 290218 541222 290454
rect 540986 289898 541222 290134
rect 540986 254218 541222 254454
rect 540986 253898 541222 254134
rect 540986 218218 541222 218454
rect 540986 217898 541222 218134
rect 540986 182218 541222 182454
rect 540986 181898 541222 182134
rect 540986 146218 541222 146454
rect 540986 145898 541222 146134
rect 540986 110218 541222 110454
rect 540986 109898 541222 110134
rect 540986 74218 541222 74454
rect 540986 73898 541222 74134
rect 540986 38218 541222 38454
rect 540986 37898 541222 38134
rect 540986 2218 541222 2454
rect 540986 1898 541222 2134
rect 540986 -582 541222 -346
rect 540986 -902 541222 -666
rect 544586 689818 544822 690054
rect 544586 689498 544822 689734
rect 544586 653818 544822 654054
rect 544586 653498 544822 653734
rect 544586 617818 544822 618054
rect 544586 617498 544822 617734
rect 544586 581818 544822 582054
rect 544586 581498 544822 581734
rect 544586 545818 544822 546054
rect 544586 545498 544822 545734
rect 544586 509818 544822 510054
rect 544586 509498 544822 509734
rect 544586 473818 544822 474054
rect 544586 473498 544822 473734
rect 544586 437818 544822 438054
rect 544586 437498 544822 437734
rect 544586 401818 544822 402054
rect 544586 401498 544822 401734
rect 544586 365818 544822 366054
rect 544586 365498 544822 365734
rect 544586 329818 544822 330054
rect 544586 329498 544822 329734
rect 544586 293818 544822 294054
rect 544586 293498 544822 293734
rect 544586 257818 544822 258054
rect 544586 257498 544822 257734
rect 544586 221818 544822 222054
rect 544586 221498 544822 221734
rect 544586 185818 544822 186054
rect 544586 185498 544822 185734
rect 544586 149818 544822 150054
rect 544586 149498 544822 149734
rect 544586 113818 544822 114054
rect 544586 113498 544822 113734
rect 544586 77818 544822 78054
rect 544586 77498 544822 77734
rect 544586 41818 544822 42054
rect 544586 41498 544822 41734
rect 544586 5818 544822 6054
rect 544586 5498 544822 5734
rect 544586 -2422 544822 -2186
rect 544586 -2742 544822 -2506
rect 548186 693418 548422 693654
rect 548186 693098 548422 693334
rect 548186 657418 548422 657654
rect 548186 657098 548422 657334
rect 548186 621418 548422 621654
rect 548186 621098 548422 621334
rect 548186 585418 548422 585654
rect 548186 585098 548422 585334
rect 548186 549418 548422 549654
rect 548186 549098 548422 549334
rect 548186 513418 548422 513654
rect 548186 513098 548422 513334
rect 548186 477418 548422 477654
rect 548186 477098 548422 477334
rect 548186 441418 548422 441654
rect 548186 441098 548422 441334
rect 548186 405418 548422 405654
rect 548186 405098 548422 405334
rect 548186 369418 548422 369654
rect 548186 369098 548422 369334
rect 548186 333418 548422 333654
rect 548186 333098 548422 333334
rect 569786 711042 570022 711278
rect 569786 710722 570022 710958
rect 566186 709202 566422 709438
rect 566186 708882 566422 709118
rect 562586 707362 562822 707598
rect 562586 707042 562822 707278
rect 551786 697018 552022 697254
rect 551786 696698 552022 696934
rect 551786 661018 552022 661254
rect 551786 660698 552022 660934
rect 551786 625018 552022 625254
rect 551786 624698 552022 624934
rect 551786 589018 552022 589254
rect 551786 588698 552022 588934
rect 551786 553018 552022 553254
rect 551786 552698 552022 552934
rect 551786 517018 552022 517254
rect 551786 516698 552022 516934
rect 551786 481018 552022 481254
rect 551786 480698 552022 480934
rect 551786 445018 552022 445254
rect 551786 444698 552022 444934
rect 551786 409018 552022 409254
rect 551786 408698 552022 408934
rect 551786 373018 552022 373254
rect 551786 372698 552022 372934
rect 551786 337018 552022 337254
rect 551786 336698 552022 336934
rect 548186 297418 548422 297654
rect 548186 297098 548422 297334
rect 548186 261418 548422 261654
rect 548186 261098 548422 261334
rect 548186 225418 548422 225654
rect 548186 225098 548422 225334
rect 548186 189418 548422 189654
rect 548186 189098 548422 189334
rect 548186 153418 548422 153654
rect 548186 153098 548422 153334
rect 548186 117418 548422 117654
rect 548186 117098 548422 117334
rect 548186 81418 548422 81654
rect 548186 81098 548422 81334
rect 548186 45418 548422 45654
rect 548186 45098 548422 45334
rect 548186 9418 548422 9654
rect 548186 9098 548422 9334
rect 548186 -4262 548422 -4026
rect 548186 -4582 548422 -4346
rect 551786 301018 552022 301254
rect 551786 300698 552022 300934
rect 551786 265018 552022 265254
rect 551786 264698 552022 264934
rect 551786 229018 552022 229254
rect 551786 228698 552022 228934
rect 551786 193018 552022 193254
rect 551786 192698 552022 192934
rect 551786 157018 552022 157254
rect 551786 156698 552022 156934
rect 551786 121018 552022 121254
rect 551786 120698 552022 120934
rect 551786 85018 552022 85254
rect 551786 84698 552022 84934
rect 551786 49018 552022 49254
rect 551786 48698 552022 48934
rect 551786 13018 552022 13254
rect 551786 12698 552022 12934
rect 533786 -7022 534022 -6786
rect 533786 -7342 534022 -7106
rect 558986 705522 559222 705758
rect 558986 705202 559222 705438
rect 558986 668218 559222 668454
rect 558986 667898 559222 668134
rect 558986 632218 559222 632454
rect 558986 631898 559222 632134
rect 558986 596218 559222 596454
rect 558986 595898 559222 596134
rect 558986 560218 559222 560454
rect 558986 559898 559222 560134
rect 558986 524218 559222 524454
rect 558986 523898 559222 524134
rect 558986 488218 559222 488454
rect 558986 487898 559222 488134
rect 558986 452218 559222 452454
rect 558986 451898 559222 452134
rect 558986 416218 559222 416454
rect 558986 415898 559222 416134
rect 558986 380218 559222 380454
rect 558986 379898 559222 380134
rect 558986 344218 559222 344454
rect 558986 343898 559222 344134
rect 562586 671818 562822 672054
rect 562586 671498 562822 671734
rect 562586 635818 562822 636054
rect 562586 635498 562822 635734
rect 562586 599818 562822 600054
rect 562586 599498 562822 599734
rect 562586 563818 562822 564054
rect 562586 563498 562822 563734
rect 562586 527818 562822 528054
rect 562586 527498 562822 527734
rect 562586 491818 562822 492054
rect 562586 491498 562822 491734
rect 562586 455818 562822 456054
rect 562586 455498 562822 455734
rect 562586 419818 562822 420054
rect 562586 419498 562822 419734
rect 562586 383818 562822 384054
rect 562586 383498 562822 383734
rect 562586 347818 562822 348054
rect 562586 347498 562822 347734
rect 562586 311818 562822 312054
rect 562586 311498 562822 311734
rect 558986 308218 559222 308454
rect 558986 307898 559222 308134
rect 558986 272218 559222 272454
rect 558986 271898 559222 272134
rect 558986 236218 559222 236454
rect 558986 235898 559222 236134
rect 558986 200218 559222 200454
rect 558986 199898 559222 200134
rect 558986 164218 559222 164454
rect 558986 163898 559222 164134
rect 558986 128218 559222 128454
rect 558986 127898 559222 128134
rect 558986 92218 559222 92454
rect 558986 91898 559222 92134
rect 558986 56218 559222 56454
rect 558986 55898 559222 56134
rect 558986 20218 559222 20454
rect 558986 19898 559222 20134
rect 558986 -1502 559222 -1266
rect 558986 -1822 559222 -1586
rect 562586 275818 562822 276054
rect 562586 275498 562822 275734
rect 562586 239818 562822 240054
rect 562586 239498 562822 239734
rect 562586 203818 562822 204054
rect 562586 203498 562822 203734
rect 562586 167818 562822 168054
rect 562586 167498 562822 167734
rect 562586 131818 562822 132054
rect 562586 131498 562822 131734
rect 562586 95818 562822 96054
rect 562586 95498 562822 95734
rect 562586 59818 562822 60054
rect 562586 59498 562822 59734
rect 562586 23818 562822 24054
rect 562586 23498 562822 23734
rect 562586 -3342 562822 -3106
rect 562586 -3662 562822 -3426
rect 566186 675418 566422 675654
rect 566186 675098 566422 675334
rect 566186 639418 566422 639654
rect 566186 639098 566422 639334
rect 566186 603418 566422 603654
rect 566186 603098 566422 603334
rect 566186 567418 566422 567654
rect 566186 567098 566422 567334
rect 566186 531418 566422 531654
rect 566186 531098 566422 531334
rect 566186 495418 566422 495654
rect 566186 495098 566422 495334
rect 566186 459418 566422 459654
rect 566186 459098 566422 459334
rect 566186 423418 566422 423654
rect 566186 423098 566422 423334
rect 566186 387418 566422 387654
rect 566186 387098 566422 387334
rect 566186 351418 566422 351654
rect 566186 351098 566422 351334
rect 566186 315418 566422 315654
rect 566186 315098 566422 315334
rect 566186 279418 566422 279654
rect 566186 279098 566422 279334
rect 566186 243418 566422 243654
rect 566186 243098 566422 243334
rect 566186 207418 566422 207654
rect 566186 207098 566422 207334
rect 566186 171418 566422 171654
rect 566186 171098 566422 171334
rect 566186 135418 566422 135654
rect 566186 135098 566422 135334
rect 566186 99418 566422 99654
rect 566186 99098 566422 99334
rect 566186 63418 566422 63654
rect 566186 63098 566422 63334
rect 566186 27418 566422 27654
rect 566186 27098 566422 27334
rect 566186 -5182 566422 -4946
rect 566186 -5502 566422 -5266
rect 591942 711042 592178 711278
rect 591942 710722 592178 710958
rect 591022 710122 591258 710358
rect 591022 709802 591258 710038
rect 590102 709202 590338 709438
rect 590102 708882 590338 709118
rect 589182 708282 589418 708518
rect 589182 707962 589418 708198
rect 588262 707362 588498 707598
rect 588262 707042 588498 707278
rect 580586 706442 580822 706678
rect 580586 706122 580822 706358
rect 569786 679018 570022 679254
rect 569786 678698 570022 678934
rect 569786 643018 570022 643254
rect 569786 642698 570022 642934
rect 569786 607018 570022 607254
rect 569786 606698 570022 606934
rect 569786 571018 570022 571254
rect 569786 570698 570022 570934
rect 569786 535018 570022 535254
rect 569786 534698 570022 534934
rect 569786 499018 570022 499254
rect 569786 498698 570022 498934
rect 569786 463018 570022 463254
rect 569786 462698 570022 462934
rect 569786 427018 570022 427254
rect 569786 426698 570022 426934
rect 569786 391018 570022 391254
rect 569786 390698 570022 390934
rect 569786 355018 570022 355254
rect 569786 354698 570022 354934
rect 569786 319018 570022 319254
rect 569786 318698 570022 318934
rect 569786 283018 570022 283254
rect 569786 282698 570022 282934
rect 569786 247018 570022 247254
rect 569786 246698 570022 246934
rect 569786 211018 570022 211254
rect 569786 210698 570022 210934
rect 569786 175018 570022 175254
rect 569786 174698 570022 174934
rect 569786 139018 570022 139254
rect 569786 138698 570022 138934
rect 569786 103018 570022 103254
rect 569786 102698 570022 102934
rect 569786 67018 570022 67254
rect 569786 66698 570022 66934
rect 569786 31018 570022 31254
rect 569786 30698 570022 30934
rect 551786 -6102 552022 -5866
rect 551786 -6422 552022 -6186
rect 576986 704602 577222 704838
rect 576986 704282 577222 704518
rect 576986 686218 577222 686454
rect 576986 685898 577222 686134
rect 576986 650218 577222 650454
rect 576986 649898 577222 650134
rect 576986 614218 577222 614454
rect 576986 613898 577222 614134
rect 576986 578218 577222 578454
rect 576986 577898 577222 578134
rect 576986 542218 577222 542454
rect 576986 541898 577222 542134
rect 576986 506218 577222 506454
rect 576986 505898 577222 506134
rect 576986 470218 577222 470454
rect 576986 469898 577222 470134
rect 576986 434218 577222 434454
rect 576986 433898 577222 434134
rect 576986 398218 577222 398454
rect 576986 397898 577222 398134
rect 576986 362218 577222 362454
rect 576986 361898 577222 362134
rect 576986 326218 577222 326454
rect 576986 325898 577222 326134
rect 576986 290218 577222 290454
rect 576986 289898 577222 290134
rect 576986 254218 577222 254454
rect 576986 253898 577222 254134
rect 576986 218218 577222 218454
rect 576986 217898 577222 218134
rect 576986 182218 577222 182454
rect 576986 181898 577222 182134
rect 576986 146218 577222 146454
rect 576986 145898 577222 146134
rect 576986 110218 577222 110454
rect 576986 109898 577222 110134
rect 576986 74218 577222 74454
rect 576986 73898 577222 74134
rect 576986 38218 577222 38454
rect 576986 37898 577222 38134
rect 576986 2218 577222 2454
rect 576986 1898 577222 2134
rect 576986 -582 577222 -346
rect 576986 -902 577222 -666
rect 587342 706442 587578 706678
rect 587342 706122 587578 706358
rect 586422 705522 586658 705758
rect 586422 705202 586658 705438
rect 580586 689818 580822 690054
rect 580586 689498 580822 689734
rect 580586 653818 580822 654054
rect 580586 653498 580822 653734
rect 580586 617818 580822 618054
rect 580586 617498 580822 617734
rect 580586 581818 580822 582054
rect 580586 581498 580822 581734
rect 580586 545818 580822 546054
rect 580586 545498 580822 545734
rect 580586 509818 580822 510054
rect 580586 509498 580822 509734
rect 580586 473818 580822 474054
rect 580586 473498 580822 473734
rect 580586 437818 580822 438054
rect 580586 437498 580822 437734
rect 580586 401818 580822 402054
rect 580586 401498 580822 401734
rect 580586 365818 580822 366054
rect 580586 365498 580822 365734
rect 580586 329818 580822 330054
rect 580586 329498 580822 329734
rect 580586 293818 580822 294054
rect 580586 293498 580822 293734
rect 580586 257818 580822 258054
rect 580586 257498 580822 257734
rect 580586 221818 580822 222054
rect 580586 221498 580822 221734
rect 580586 185818 580822 186054
rect 580586 185498 580822 185734
rect 580586 149818 580822 150054
rect 580586 149498 580822 149734
rect 580586 113818 580822 114054
rect 580586 113498 580822 113734
rect 580586 77818 580822 78054
rect 580586 77498 580822 77734
rect 580586 41818 580822 42054
rect 580586 41498 580822 41734
rect 580586 5818 580822 6054
rect 580586 5498 580822 5734
rect 585502 704602 585738 704838
rect 585502 704282 585738 704518
rect 585502 686218 585738 686454
rect 585502 685898 585738 686134
rect 585502 650218 585738 650454
rect 585502 649898 585738 650134
rect 585502 614218 585738 614454
rect 585502 613898 585738 614134
rect 585502 578218 585738 578454
rect 585502 577898 585738 578134
rect 585502 542218 585738 542454
rect 585502 541898 585738 542134
rect 585502 506218 585738 506454
rect 585502 505898 585738 506134
rect 585502 470218 585738 470454
rect 585502 469898 585738 470134
rect 585502 434218 585738 434454
rect 585502 433898 585738 434134
rect 585502 398218 585738 398454
rect 585502 397898 585738 398134
rect 585502 362218 585738 362454
rect 585502 361898 585738 362134
rect 585502 326218 585738 326454
rect 585502 325898 585738 326134
rect 585502 290218 585738 290454
rect 585502 289898 585738 290134
rect 585502 254218 585738 254454
rect 585502 253898 585738 254134
rect 585502 218218 585738 218454
rect 585502 217898 585738 218134
rect 585502 182218 585738 182454
rect 585502 181898 585738 182134
rect 585502 146218 585738 146454
rect 585502 145898 585738 146134
rect 585502 110218 585738 110454
rect 585502 109898 585738 110134
rect 585502 74218 585738 74454
rect 585502 73898 585738 74134
rect 585502 38218 585738 38454
rect 585502 37898 585738 38134
rect 585502 2218 585738 2454
rect 585502 1898 585738 2134
rect 585502 -582 585738 -346
rect 585502 -902 585738 -666
rect 586422 668218 586658 668454
rect 586422 667898 586658 668134
rect 586422 632218 586658 632454
rect 586422 631898 586658 632134
rect 586422 596218 586658 596454
rect 586422 595898 586658 596134
rect 586422 560218 586658 560454
rect 586422 559898 586658 560134
rect 586422 524218 586658 524454
rect 586422 523898 586658 524134
rect 586422 488218 586658 488454
rect 586422 487898 586658 488134
rect 586422 452218 586658 452454
rect 586422 451898 586658 452134
rect 586422 416218 586658 416454
rect 586422 415898 586658 416134
rect 586422 380218 586658 380454
rect 586422 379898 586658 380134
rect 586422 344218 586658 344454
rect 586422 343898 586658 344134
rect 586422 308218 586658 308454
rect 586422 307898 586658 308134
rect 586422 272218 586658 272454
rect 586422 271898 586658 272134
rect 586422 236218 586658 236454
rect 586422 235898 586658 236134
rect 586422 200218 586658 200454
rect 586422 199898 586658 200134
rect 586422 164218 586658 164454
rect 586422 163898 586658 164134
rect 586422 128218 586658 128454
rect 586422 127898 586658 128134
rect 586422 92218 586658 92454
rect 586422 91898 586658 92134
rect 586422 56218 586658 56454
rect 586422 55898 586658 56134
rect 586422 20218 586658 20454
rect 586422 19898 586658 20134
rect 586422 -1502 586658 -1266
rect 586422 -1822 586658 -1586
rect 587342 689818 587578 690054
rect 587342 689498 587578 689734
rect 587342 653818 587578 654054
rect 587342 653498 587578 653734
rect 587342 617818 587578 618054
rect 587342 617498 587578 617734
rect 587342 581818 587578 582054
rect 587342 581498 587578 581734
rect 587342 545818 587578 546054
rect 587342 545498 587578 545734
rect 587342 509818 587578 510054
rect 587342 509498 587578 509734
rect 587342 473818 587578 474054
rect 587342 473498 587578 473734
rect 587342 437818 587578 438054
rect 587342 437498 587578 437734
rect 587342 401818 587578 402054
rect 587342 401498 587578 401734
rect 587342 365818 587578 366054
rect 587342 365498 587578 365734
rect 587342 329818 587578 330054
rect 587342 329498 587578 329734
rect 587342 293818 587578 294054
rect 587342 293498 587578 293734
rect 587342 257818 587578 258054
rect 587342 257498 587578 257734
rect 587342 221818 587578 222054
rect 587342 221498 587578 221734
rect 587342 185818 587578 186054
rect 587342 185498 587578 185734
rect 587342 149818 587578 150054
rect 587342 149498 587578 149734
rect 587342 113818 587578 114054
rect 587342 113498 587578 113734
rect 587342 77818 587578 78054
rect 587342 77498 587578 77734
rect 587342 41818 587578 42054
rect 587342 41498 587578 41734
rect 587342 5818 587578 6054
rect 587342 5498 587578 5734
rect 580586 -2422 580822 -2186
rect 580586 -2742 580822 -2506
rect 587342 -2422 587578 -2186
rect 587342 -2742 587578 -2506
rect 588262 671818 588498 672054
rect 588262 671498 588498 671734
rect 588262 635818 588498 636054
rect 588262 635498 588498 635734
rect 588262 599818 588498 600054
rect 588262 599498 588498 599734
rect 588262 563818 588498 564054
rect 588262 563498 588498 563734
rect 588262 527818 588498 528054
rect 588262 527498 588498 527734
rect 588262 491818 588498 492054
rect 588262 491498 588498 491734
rect 588262 455818 588498 456054
rect 588262 455498 588498 455734
rect 588262 419818 588498 420054
rect 588262 419498 588498 419734
rect 588262 383818 588498 384054
rect 588262 383498 588498 383734
rect 588262 347818 588498 348054
rect 588262 347498 588498 347734
rect 588262 311818 588498 312054
rect 588262 311498 588498 311734
rect 588262 275818 588498 276054
rect 588262 275498 588498 275734
rect 588262 239818 588498 240054
rect 588262 239498 588498 239734
rect 588262 203818 588498 204054
rect 588262 203498 588498 203734
rect 588262 167818 588498 168054
rect 588262 167498 588498 167734
rect 588262 131818 588498 132054
rect 588262 131498 588498 131734
rect 588262 95818 588498 96054
rect 588262 95498 588498 95734
rect 588262 59818 588498 60054
rect 588262 59498 588498 59734
rect 588262 23818 588498 24054
rect 588262 23498 588498 23734
rect 588262 -3342 588498 -3106
rect 588262 -3662 588498 -3426
rect 589182 693418 589418 693654
rect 589182 693098 589418 693334
rect 589182 657418 589418 657654
rect 589182 657098 589418 657334
rect 589182 621418 589418 621654
rect 589182 621098 589418 621334
rect 589182 585418 589418 585654
rect 589182 585098 589418 585334
rect 589182 549418 589418 549654
rect 589182 549098 589418 549334
rect 589182 513418 589418 513654
rect 589182 513098 589418 513334
rect 589182 477418 589418 477654
rect 589182 477098 589418 477334
rect 589182 441418 589418 441654
rect 589182 441098 589418 441334
rect 589182 405418 589418 405654
rect 589182 405098 589418 405334
rect 589182 369418 589418 369654
rect 589182 369098 589418 369334
rect 589182 333418 589418 333654
rect 589182 333098 589418 333334
rect 589182 297418 589418 297654
rect 589182 297098 589418 297334
rect 589182 261418 589418 261654
rect 589182 261098 589418 261334
rect 589182 225418 589418 225654
rect 589182 225098 589418 225334
rect 589182 189418 589418 189654
rect 589182 189098 589418 189334
rect 589182 153418 589418 153654
rect 589182 153098 589418 153334
rect 589182 117418 589418 117654
rect 589182 117098 589418 117334
rect 589182 81418 589418 81654
rect 589182 81098 589418 81334
rect 589182 45418 589418 45654
rect 589182 45098 589418 45334
rect 589182 9418 589418 9654
rect 589182 9098 589418 9334
rect 589182 -4262 589418 -4026
rect 589182 -4582 589418 -4346
rect 590102 675418 590338 675654
rect 590102 675098 590338 675334
rect 590102 639418 590338 639654
rect 590102 639098 590338 639334
rect 590102 603418 590338 603654
rect 590102 603098 590338 603334
rect 590102 567418 590338 567654
rect 590102 567098 590338 567334
rect 590102 531418 590338 531654
rect 590102 531098 590338 531334
rect 590102 495418 590338 495654
rect 590102 495098 590338 495334
rect 590102 459418 590338 459654
rect 590102 459098 590338 459334
rect 590102 423418 590338 423654
rect 590102 423098 590338 423334
rect 590102 387418 590338 387654
rect 590102 387098 590338 387334
rect 590102 351418 590338 351654
rect 590102 351098 590338 351334
rect 590102 315418 590338 315654
rect 590102 315098 590338 315334
rect 590102 279418 590338 279654
rect 590102 279098 590338 279334
rect 590102 243418 590338 243654
rect 590102 243098 590338 243334
rect 590102 207418 590338 207654
rect 590102 207098 590338 207334
rect 590102 171418 590338 171654
rect 590102 171098 590338 171334
rect 590102 135418 590338 135654
rect 590102 135098 590338 135334
rect 590102 99418 590338 99654
rect 590102 99098 590338 99334
rect 590102 63418 590338 63654
rect 590102 63098 590338 63334
rect 590102 27418 590338 27654
rect 590102 27098 590338 27334
rect 590102 -5182 590338 -4946
rect 590102 -5502 590338 -5266
rect 591022 697018 591258 697254
rect 591022 696698 591258 696934
rect 591022 661018 591258 661254
rect 591022 660698 591258 660934
rect 591022 625018 591258 625254
rect 591022 624698 591258 624934
rect 591022 589018 591258 589254
rect 591022 588698 591258 588934
rect 591022 553018 591258 553254
rect 591022 552698 591258 552934
rect 591022 517018 591258 517254
rect 591022 516698 591258 516934
rect 591022 481018 591258 481254
rect 591022 480698 591258 480934
rect 591022 445018 591258 445254
rect 591022 444698 591258 444934
rect 591022 409018 591258 409254
rect 591022 408698 591258 408934
rect 591022 373018 591258 373254
rect 591022 372698 591258 372934
rect 591022 337018 591258 337254
rect 591022 336698 591258 336934
rect 591022 301018 591258 301254
rect 591022 300698 591258 300934
rect 591022 265018 591258 265254
rect 591022 264698 591258 264934
rect 591022 229018 591258 229254
rect 591022 228698 591258 228934
rect 591022 193018 591258 193254
rect 591022 192698 591258 192934
rect 591022 157018 591258 157254
rect 591022 156698 591258 156934
rect 591022 121018 591258 121254
rect 591022 120698 591258 120934
rect 591022 85018 591258 85254
rect 591022 84698 591258 84934
rect 591022 49018 591258 49254
rect 591022 48698 591258 48934
rect 591022 13018 591258 13254
rect 591022 12698 591258 12934
rect 591022 -6102 591258 -5866
rect 591022 -6422 591258 -6186
rect 591942 679018 592178 679254
rect 591942 678698 592178 678934
rect 591942 643018 592178 643254
rect 591942 642698 592178 642934
rect 591942 607018 592178 607254
rect 591942 606698 592178 606934
rect 591942 571018 592178 571254
rect 591942 570698 592178 570934
rect 591942 535018 592178 535254
rect 591942 534698 592178 534934
rect 591942 499018 592178 499254
rect 591942 498698 592178 498934
rect 591942 463018 592178 463254
rect 591942 462698 592178 462934
rect 591942 427018 592178 427254
rect 591942 426698 592178 426934
rect 591942 391018 592178 391254
rect 591942 390698 592178 390934
rect 591942 355018 592178 355254
rect 591942 354698 592178 354934
rect 591942 319018 592178 319254
rect 591942 318698 592178 318934
rect 591942 283018 592178 283254
rect 591942 282698 592178 282934
rect 591942 247018 592178 247254
rect 591942 246698 592178 246934
rect 591942 211018 592178 211254
rect 591942 210698 592178 210934
rect 591942 175018 592178 175254
rect 591942 174698 592178 174934
rect 591942 139018 592178 139254
rect 591942 138698 592178 138934
rect 591942 103018 592178 103254
rect 591942 102698 592178 102934
rect 591942 67018 592178 67254
rect 591942 66698 592178 66934
rect 591942 31018 592178 31254
rect 591942 30698 592178 30934
rect 569786 -7022 570022 -6786
rect 569786 -7342 570022 -7106
rect 591942 -7022 592178 -6786
rect 591942 -7342 592178 -7106
<< metal5 >>
rect -8436 711300 -7836 711302
rect 29604 711300 30204 711302
rect 65604 711300 66204 711302
rect 101604 711300 102204 711302
rect 137604 711300 138204 711302
rect 173604 711300 174204 711302
rect 209604 711300 210204 711302
rect 245604 711300 246204 711302
rect 281604 711300 282204 711302
rect 317604 711300 318204 711302
rect 353604 711300 354204 711302
rect 389604 711300 390204 711302
rect 425604 711300 426204 711302
rect 461604 711300 462204 711302
rect 497604 711300 498204 711302
rect 533604 711300 534204 711302
rect 569604 711300 570204 711302
rect 591760 711300 592360 711302
rect -8436 711278 592360 711300
rect -8436 711042 -8254 711278
rect -8018 711042 29786 711278
rect 30022 711042 65786 711278
rect 66022 711042 101786 711278
rect 102022 711042 137786 711278
rect 138022 711042 173786 711278
rect 174022 711042 209786 711278
rect 210022 711042 245786 711278
rect 246022 711042 281786 711278
rect 282022 711042 317786 711278
rect 318022 711042 353786 711278
rect 354022 711042 389786 711278
rect 390022 711042 425786 711278
rect 426022 711042 461786 711278
rect 462022 711042 497786 711278
rect 498022 711042 533786 711278
rect 534022 711042 569786 711278
rect 570022 711042 591942 711278
rect 592178 711042 592360 711278
rect -8436 710958 592360 711042
rect -8436 710722 -8254 710958
rect -8018 710722 29786 710958
rect 30022 710722 65786 710958
rect 66022 710722 101786 710958
rect 102022 710722 137786 710958
rect 138022 710722 173786 710958
rect 174022 710722 209786 710958
rect 210022 710722 245786 710958
rect 246022 710722 281786 710958
rect 282022 710722 317786 710958
rect 318022 710722 353786 710958
rect 354022 710722 389786 710958
rect 390022 710722 425786 710958
rect 426022 710722 461786 710958
rect 462022 710722 497786 710958
rect 498022 710722 533786 710958
rect 534022 710722 569786 710958
rect 570022 710722 591942 710958
rect 592178 710722 592360 710958
rect -8436 710700 592360 710722
rect -8436 710698 -7836 710700
rect 29604 710698 30204 710700
rect 65604 710698 66204 710700
rect 101604 710698 102204 710700
rect 137604 710698 138204 710700
rect 173604 710698 174204 710700
rect 209604 710698 210204 710700
rect 245604 710698 246204 710700
rect 281604 710698 282204 710700
rect 317604 710698 318204 710700
rect 353604 710698 354204 710700
rect 389604 710698 390204 710700
rect 425604 710698 426204 710700
rect 461604 710698 462204 710700
rect 497604 710698 498204 710700
rect 533604 710698 534204 710700
rect 569604 710698 570204 710700
rect 591760 710698 592360 710700
rect -7516 710380 -6916 710382
rect 11604 710380 12204 710382
rect 47604 710380 48204 710382
rect 83604 710380 84204 710382
rect 119604 710380 120204 710382
rect 155604 710380 156204 710382
rect 191604 710380 192204 710382
rect 227604 710380 228204 710382
rect 263604 710380 264204 710382
rect 299604 710380 300204 710382
rect 335604 710380 336204 710382
rect 371604 710380 372204 710382
rect 407604 710380 408204 710382
rect 443604 710380 444204 710382
rect 479604 710380 480204 710382
rect 515604 710380 516204 710382
rect 551604 710380 552204 710382
rect 590840 710380 591440 710382
rect -7516 710358 591440 710380
rect -7516 710122 -7334 710358
rect -7098 710122 11786 710358
rect 12022 710122 47786 710358
rect 48022 710122 83786 710358
rect 84022 710122 119786 710358
rect 120022 710122 155786 710358
rect 156022 710122 191786 710358
rect 192022 710122 227786 710358
rect 228022 710122 263786 710358
rect 264022 710122 299786 710358
rect 300022 710122 335786 710358
rect 336022 710122 371786 710358
rect 372022 710122 407786 710358
rect 408022 710122 443786 710358
rect 444022 710122 479786 710358
rect 480022 710122 515786 710358
rect 516022 710122 551786 710358
rect 552022 710122 591022 710358
rect 591258 710122 591440 710358
rect -7516 710038 591440 710122
rect -7516 709802 -7334 710038
rect -7098 709802 11786 710038
rect 12022 709802 47786 710038
rect 48022 709802 83786 710038
rect 84022 709802 119786 710038
rect 120022 709802 155786 710038
rect 156022 709802 191786 710038
rect 192022 709802 227786 710038
rect 228022 709802 263786 710038
rect 264022 709802 299786 710038
rect 300022 709802 335786 710038
rect 336022 709802 371786 710038
rect 372022 709802 407786 710038
rect 408022 709802 443786 710038
rect 444022 709802 479786 710038
rect 480022 709802 515786 710038
rect 516022 709802 551786 710038
rect 552022 709802 591022 710038
rect 591258 709802 591440 710038
rect -7516 709780 591440 709802
rect -7516 709778 -6916 709780
rect 11604 709778 12204 709780
rect 47604 709778 48204 709780
rect 83604 709778 84204 709780
rect 119604 709778 120204 709780
rect 155604 709778 156204 709780
rect 191604 709778 192204 709780
rect 227604 709778 228204 709780
rect 263604 709778 264204 709780
rect 299604 709778 300204 709780
rect 335604 709778 336204 709780
rect 371604 709778 372204 709780
rect 407604 709778 408204 709780
rect 443604 709778 444204 709780
rect 479604 709778 480204 709780
rect 515604 709778 516204 709780
rect 551604 709778 552204 709780
rect 590840 709778 591440 709780
rect -6596 709460 -5996 709462
rect 26004 709460 26604 709462
rect 62004 709460 62604 709462
rect 98004 709460 98604 709462
rect 134004 709460 134604 709462
rect 170004 709460 170604 709462
rect 206004 709460 206604 709462
rect 242004 709460 242604 709462
rect 278004 709460 278604 709462
rect 314004 709460 314604 709462
rect 350004 709460 350604 709462
rect 386004 709460 386604 709462
rect 422004 709460 422604 709462
rect 458004 709460 458604 709462
rect 494004 709460 494604 709462
rect 530004 709460 530604 709462
rect 566004 709460 566604 709462
rect 589920 709460 590520 709462
rect -6596 709438 590520 709460
rect -6596 709202 -6414 709438
rect -6178 709202 26186 709438
rect 26422 709202 62186 709438
rect 62422 709202 98186 709438
rect 98422 709202 134186 709438
rect 134422 709202 170186 709438
rect 170422 709202 206186 709438
rect 206422 709202 242186 709438
rect 242422 709202 278186 709438
rect 278422 709202 314186 709438
rect 314422 709202 350186 709438
rect 350422 709202 386186 709438
rect 386422 709202 422186 709438
rect 422422 709202 458186 709438
rect 458422 709202 494186 709438
rect 494422 709202 530186 709438
rect 530422 709202 566186 709438
rect 566422 709202 590102 709438
rect 590338 709202 590520 709438
rect -6596 709118 590520 709202
rect -6596 708882 -6414 709118
rect -6178 708882 26186 709118
rect 26422 708882 62186 709118
rect 62422 708882 98186 709118
rect 98422 708882 134186 709118
rect 134422 708882 170186 709118
rect 170422 708882 206186 709118
rect 206422 708882 242186 709118
rect 242422 708882 278186 709118
rect 278422 708882 314186 709118
rect 314422 708882 350186 709118
rect 350422 708882 386186 709118
rect 386422 708882 422186 709118
rect 422422 708882 458186 709118
rect 458422 708882 494186 709118
rect 494422 708882 530186 709118
rect 530422 708882 566186 709118
rect 566422 708882 590102 709118
rect 590338 708882 590520 709118
rect -6596 708860 590520 708882
rect -6596 708858 -5996 708860
rect 26004 708858 26604 708860
rect 62004 708858 62604 708860
rect 98004 708858 98604 708860
rect 134004 708858 134604 708860
rect 170004 708858 170604 708860
rect 206004 708858 206604 708860
rect 242004 708858 242604 708860
rect 278004 708858 278604 708860
rect 314004 708858 314604 708860
rect 350004 708858 350604 708860
rect 386004 708858 386604 708860
rect 422004 708858 422604 708860
rect 458004 708858 458604 708860
rect 494004 708858 494604 708860
rect 530004 708858 530604 708860
rect 566004 708858 566604 708860
rect 589920 708858 590520 708860
rect -5676 708540 -5076 708542
rect 8004 708540 8604 708542
rect 44004 708540 44604 708542
rect 80004 708540 80604 708542
rect 116004 708540 116604 708542
rect 152004 708540 152604 708542
rect 188004 708540 188604 708542
rect 224004 708540 224604 708542
rect 260004 708540 260604 708542
rect 296004 708540 296604 708542
rect 332004 708540 332604 708542
rect 368004 708540 368604 708542
rect 404004 708540 404604 708542
rect 440004 708540 440604 708542
rect 476004 708540 476604 708542
rect 512004 708540 512604 708542
rect 548004 708540 548604 708542
rect 589000 708540 589600 708542
rect -5676 708518 589600 708540
rect -5676 708282 -5494 708518
rect -5258 708282 8186 708518
rect 8422 708282 44186 708518
rect 44422 708282 80186 708518
rect 80422 708282 116186 708518
rect 116422 708282 152186 708518
rect 152422 708282 188186 708518
rect 188422 708282 224186 708518
rect 224422 708282 260186 708518
rect 260422 708282 296186 708518
rect 296422 708282 332186 708518
rect 332422 708282 368186 708518
rect 368422 708282 404186 708518
rect 404422 708282 440186 708518
rect 440422 708282 476186 708518
rect 476422 708282 512186 708518
rect 512422 708282 548186 708518
rect 548422 708282 589182 708518
rect 589418 708282 589600 708518
rect -5676 708198 589600 708282
rect -5676 707962 -5494 708198
rect -5258 707962 8186 708198
rect 8422 707962 44186 708198
rect 44422 707962 80186 708198
rect 80422 707962 116186 708198
rect 116422 707962 152186 708198
rect 152422 707962 188186 708198
rect 188422 707962 224186 708198
rect 224422 707962 260186 708198
rect 260422 707962 296186 708198
rect 296422 707962 332186 708198
rect 332422 707962 368186 708198
rect 368422 707962 404186 708198
rect 404422 707962 440186 708198
rect 440422 707962 476186 708198
rect 476422 707962 512186 708198
rect 512422 707962 548186 708198
rect 548422 707962 589182 708198
rect 589418 707962 589600 708198
rect -5676 707940 589600 707962
rect -5676 707938 -5076 707940
rect 8004 707938 8604 707940
rect 44004 707938 44604 707940
rect 80004 707938 80604 707940
rect 116004 707938 116604 707940
rect 152004 707938 152604 707940
rect 188004 707938 188604 707940
rect 224004 707938 224604 707940
rect 260004 707938 260604 707940
rect 296004 707938 296604 707940
rect 332004 707938 332604 707940
rect 368004 707938 368604 707940
rect 404004 707938 404604 707940
rect 440004 707938 440604 707940
rect 476004 707938 476604 707940
rect 512004 707938 512604 707940
rect 548004 707938 548604 707940
rect 589000 707938 589600 707940
rect -4756 707620 -4156 707622
rect 22404 707620 23004 707622
rect 58404 707620 59004 707622
rect 94404 707620 95004 707622
rect 130404 707620 131004 707622
rect 166404 707620 167004 707622
rect 202404 707620 203004 707622
rect 238404 707620 239004 707622
rect 274404 707620 275004 707622
rect 310404 707620 311004 707622
rect 346404 707620 347004 707622
rect 382404 707620 383004 707622
rect 418404 707620 419004 707622
rect 454404 707620 455004 707622
rect 490404 707620 491004 707622
rect 526404 707620 527004 707622
rect 562404 707620 563004 707622
rect 588080 707620 588680 707622
rect -4756 707598 588680 707620
rect -4756 707362 -4574 707598
rect -4338 707362 22586 707598
rect 22822 707362 58586 707598
rect 58822 707362 94586 707598
rect 94822 707362 130586 707598
rect 130822 707362 166586 707598
rect 166822 707362 202586 707598
rect 202822 707362 238586 707598
rect 238822 707362 274586 707598
rect 274822 707362 310586 707598
rect 310822 707362 346586 707598
rect 346822 707362 382586 707598
rect 382822 707362 418586 707598
rect 418822 707362 454586 707598
rect 454822 707362 490586 707598
rect 490822 707362 526586 707598
rect 526822 707362 562586 707598
rect 562822 707362 588262 707598
rect 588498 707362 588680 707598
rect -4756 707278 588680 707362
rect -4756 707042 -4574 707278
rect -4338 707042 22586 707278
rect 22822 707042 58586 707278
rect 58822 707042 94586 707278
rect 94822 707042 130586 707278
rect 130822 707042 166586 707278
rect 166822 707042 202586 707278
rect 202822 707042 238586 707278
rect 238822 707042 274586 707278
rect 274822 707042 310586 707278
rect 310822 707042 346586 707278
rect 346822 707042 382586 707278
rect 382822 707042 418586 707278
rect 418822 707042 454586 707278
rect 454822 707042 490586 707278
rect 490822 707042 526586 707278
rect 526822 707042 562586 707278
rect 562822 707042 588262 707278
rect 588498 707042 588680 707278
rect -4756 707020 588680 707042
rect -4756 707018 -4156 707020
rect 22404 707018 23004 707020
rect 58404 707018 59004 707020
rect 94404 707018 95004 707020
rect 130404 707018 131004 707020
rect 166404 707018 167004 707020
rect 202404 707018 203004 707020
rect 238404 707018 239004 707020
rect 274404 707018 275004 707020
rect 310404 707018 311004 707020
rect 346404 707018 347004 707020
rect 382404 707018 383004 707020
rect 418404 707018 419004 707020
rect 454404 707018 455004 707020
rect 490404 707018 491004 707020
rect 526404 707018 527004 707020
rect 562404 707018 563004 707020
rect 588080 707018 588680 707020
rect -3836 706700 -3236 706702
rect 4404 706700 5004 706702
rect 40404 706700 41004 706702
rect 76404 706700 77004 706702
rect 112404 706700 113004 706702
rect 148404 706700 149004 706702
rect 184404 706700 185004 706702
rect 220404 706700 221004 706702
rect 256404 706700 257004 706702
rect 292404 706700 293004 706702
rect 328404 706700 329004 706702
rect 364404 706700 365004 706702
rect 400404 706700 401004 706702
rect 436404 706700 437004 706702
rect 472404 706700 473004 706702
rect 508404 706700 509004 706702
rect 544404 706700 545004 706702
rect 580404 706700 581004 706702
rect 587160 706700 587760 706702
rect -3836 706678 587760 706700
rect -3836 706442 -3654 706678
rect -3418 706442 4586 706678
rect 4822 706442 40586 706678
rect 40822 706442 76586 706678
rect 76822 706442 112586 706678
rect 112822 706442 148586 706678
rect 148822 706442 184586 706678
rect 184822 706442 220586 706678
rect 220822 706442 256586 706678
rect 256822 706442 292586 706678
rect 292822 706442 328586 706678
rect 328822 706442 364586 706678
rect 364822 706442 400586 706678
rect 400822 706442 436586 706678
rect 436822 706442 472586 706678
rect 472822 706442 508586 706678
rect 508822 706442 544586 706678
rect 544822 706442 580586 706678
rect 580822 706442 587342 706678
rect 587578 706442 587760 706678
rect -3836 706358 587760 706442
rect -3836 706122 -3654 706358
rect -3418 706122 4586 706358
rect 4822 706122 40586 706358
rect 40822 706122 76586 706358
rect 76822 706122 112586 706358
rect 112822 706122 148586 706358
rect 148822 706122 184586 706358
rect 184822 706122 220586 706358
rect 220822 706122 256586 706358
rect 256822 706122 292586 706358
rect 292822 706122 328586 706358
rect 328822 706122 364586 706358
rect 364822 706122 400586 706358
rect 400822 706122 436586 706358
rect 436822 706122 472586 706358
rect 472822 706122 508586 706358
rect 508822 706122 544586 706358
rect 544822 706122 580586 706358
rect 580822 706122 587342 706358
rect 587578 706122 587760 706358
rect -3836 706100 587760 706122
rect -3836 706098 -3236 706100
rect 4404 706098 5004 706100
rect 40404 706098 41004 706100
rect 76404 706098 77004 706100
rect 112404 706098 113004 706100
rect 148404 706098 149004 706100
rect 184404 706098 185004 706100
rect 220404 706098 221004 706100
rect 256404 706098 257004 706100
rect 292404 706098 293004 706100
rect 328404 706098 329004 706100
rect 364404 706098 365004 706100
rect 400404 706098 401004 706100
rect 436404 706098 437004 706100
rect 472404 706098 473004 706100
rect 508404 706098 509004 706100
rect 544404 706098 545004 706100
rect 580404 706098 581004 706100
rect 587160 706098 587760 706100
rect -2916 705780 -2316 705782
rect 18804 705780 19404 705782
rect 54804 705780 55404 705782
rect 90804 705780 91404 705782
rect 126804 705780 127404 705782
rect 162804 705780 163404 705782
rect 198804 705780 199404 705782
rect 234804 705780 235404 705782
rect 270804 705780 271404 705782
rect 306804 705780 307404 705782
rect 342804 705780 343404 705782
rect 378804 705780 379404 705782
rect 414804 705780 415404 705782
rect 450804 705780 451404 705782
rect 486804 705780 487404 705782
rect 522804 705780 523404 705782
rect 558804 705780 559404 705782
rect 586240 705780 586840 705782
rect -2916 705758 586840 705780
rect -2916 705522 -2734 705758
rect -2498 705522 18986 705758
rect 19222 705522 54986 705758
rect 55222 705522 90986 705758
rect 91222 705522 126986 705758
rect 127222 705522 162986 705758
rect 163222 705522 198986 705758
rect 199222 705522 234986 705758
rect 235222 705522 270986 705758
rect 271222 705522 306986 705758
rect 307222 705522 342986 705758
rect 343222 705522 378986 705758
rect 379222 705522 414986 705758
rect 415222 705522 450986 705758
rect 451222 705522 486986 705758
rect 487222 705522 522986 705758
rect 523222 705522 558986 705758
rect 559222 705522 586422 705758
rect 586658 705522 586840 705758
rect -2916 705438 586840 705522
rect -2916 705202 -2734 705438
rect -2498 705202 18986 705438
rect 19222 705202 54986 705438
rect 55222 705202 90986 705438
rect 91222 705202 126986 705438
rect 127222 705202 162986 705438
rect 163222 705202 198986 705438
rect 199222 705202 234986 705438
rect 235222 705202 270986 705438
rect 271222 705202 306986 705438
rect 307222 705202 342986 705438
rect 343222 705202 378986 705438
rect 379222 705202 414986 705438
rect 415222 705202 450986 705438
rect 451222 705202 486986 705438
rect 487222 705202 522986 705438
rect 523222 705202 558986 705438
rect 559222 705202 586422 705438
rect 586658 705202 586840 705438
rect -2916 705180 586840 705202
rect -2916 705178 -2316 705180
rect 18804 705178 19404 705180
rect 54804 705178 55404 705180
rect 90804 705178 91404 705180
rect 126804 705178 127404 705180
rect 162804 705178 163404 705180
rect 198804 705178 199404 705180
rect 234804 705178 235404 705180
rect 270804 705178 271404 705180
rect 306804 705178 307404 705180
rect 342804 705178 343404 705180
rect 378804 705178 379404 705180
rect 414804 705178 415404 705180
rect 450804 705178 451404 705180
rect 486804 705178 487404 705180
rect 522804 705178 523404 705180
rect 558804 705178 559404 705180
rect 586240 705178 586840 705180
rect -1996 704860 -1396 704862
rect 804 704860 1404 704862
rect 36804 704860 37404 704862
rect 72804 704860 73404 704862
rect 108804 704860 109404 704862
rect 144804 704860 145404 704862
rect 180804 704860 181404 704862
rect 216804 704860 217404 704862
rect 252804 704860 253404 704862
rect 288804 704860 289404 704862
rect 324804 704860 325404 704862
rect 360804 704860 361404 704862
rect 396804 704860 397404 704862
rect 432804 704860 433404 704862
rect 468804 704860 469404 704862
rect 504804 704860 505404 704862
rect 540804 704860 541404 704862
rect 576804 704860 577404 704862
rect 585320 704860 585920 704862
rect -1996 704838 585920 704860
rect -1996 704602 -1814 704838
rect -1578 704602 986 704838
rect 1222 704602 36986 704838
rect 37222 704602 72986 704838
rect 73222 704602 108986 704838
rect 109222 704602 144986 704838
rect 145222 704602 180986 704838
rect 181222 704602 216986 704838
rect 217222 704602 252986 704838
rect 253222 704602 288986 704838
rect 289222 704602 324986 704838
rect 325222 704602 360986 704838
rect 361222 704602 396986 704838
rect 397222 704602 432986 704838
rect 433222 704602 468986 704838
rect 469222 704602 504986 704838
rect 505222 704602 540986 704838
rect 541222 704602 576986 704838
rect 577222 704602 585502 704838
rect 585738 704602 585920 704838
rect -1996 704518 585920 704602
rect -1996 704282 -1814 704518
rect -1578 704282 986 704518
rect 1222 704282 36986 704518
rect 37222 704282 72986 704518
rect 73222 704282 108986 704518
rect 109222 704282 144986 704518
rect 145222 704282 180986 704518
rect 181222 704282 216986 704518
rect 217222 704282 252986 704518
rect 253222 704282 288986 704518
rect 289222 704282 324986 704518
rect 325222 704282 360986 704518
rect 361222 704282 396986 704518
rect 397222 704282 432986 704518
rect 433222 704282 468986 704518
rect 469222 704282 504986 704518
rect 505222 704282 540986 704518
rect 541222 704282 576986 704518
rect 577222 704282 585502 704518
rect 585738 704282 585920 704518
rect -1996 704260 585920 704282
rect -1996 704258 -1396 704260
rect 804 704258 1404 704260
rect 36804 704258 37404 704260
rect 72804 704258 73404 704260
rect 108804 704258 109404 704260
rect 144804 704258 145404 704260
rect 180804 704258 181404 704260
rect 216804 704258 217404 704260
rect 252804 704258 253404 704260
rect 288804 704258 289404 704260
rect 324804 704258 325404 704260
rect 360804 704258 361404 704260
rect 396804 704258 397404 704260
rect 432804 704258 433404 704260
rect 468804 704258 469404 704260
rect 504804 704258 505404 704260
rect 540804 704258 541404 704260
rect 576804 704258 577404 704260
rect 585320 704258 585920 704260
rect -7516 697276 -6916 697278
rect 11604 697276 12204 697278
rect 47604 697276 48204 697278
rect 83604 697276 84204 697278
rect 119604 697276 120204 697278
rect 155604 697276 156204 697278
rect 191604 697276 192204 697278
rect 227604 697276 228204 697278
rect 263604 697276 264204 697278
rect 299604 697276 300204 697278
rect 335604 697276 336204 697278
rect 371604 697276 372204 697278
rect 407604 697276 408204 697278
rect 443604 697276 444204 697278
rect 479604 697276 480204 697278
rect 515604 697276 516204 697278
rect 551604 697276 552204 697278
rect 590840 697276 591440 697278
rect -8436 697254 592360 697276
rect -8436 697018 -7334 697254
rect -7098 697018 11786 697254
rect 12022 697018 47786 697254
rect 48022 697018 83786 697254
rect 84022 697018 119786 697254
rect 120022 697018 155786 697254
rect 156022 697018 191786 697254
rect 192022 697018 227786 697254
rect 228022 697018 263786 697254
rect 264022 697018 299786 697254
rect 300022 697018 335786 697254
rect 336022 697018 371786 697254
rect 372022 697018 407786 697254
rect 408022 697018 443786 697254
rect 444022 697018 479786 697254
rect 480022 697018 515786 697254
rect 516022 697018 551786 697254
rect 552022 697018 591022 697254
rect 591258 697018 592360 697254
rect -8436 696934 592360 697018
rect -8436 696698 -7334 696934
rect -7098 696698 11786 696934
rect 12022 696698 47786 696934
rect 48022 696698 83786 696934
rect 84022 696698 119786 696934
rect 120022 696698 155786 696934
rect 156022 696698 191786 696934
rect 192022 696698 227786 696934
rect 228022 696698 263786 696934
rect 264022 696698 299786 696934
rect 300022 696698 335786 696934
rect 336022 696698 371786 696934
rect 372022 696698 407786 696934
rect 408022 696698 443786 696934
rect 444022 696698 479786 696934
rect 480022 696698 515786 696934
rect 516022 696698 551786 696934
rect 552022 696698 591022 696934
rect 591258 696698 592360 696934
rect -8436 696676 592360 696698
rect -7516 696674 -6916 696676
rect 11604 696674 12204 696676
rect 47604 696674 48204 696676
rect 83604 696674 84204 696676
rect 119604 696674 120204 696676
rect 155604 696674 156204 696676
rect 191604 696674 192204 696676
rect 227604 696674 228204 696676
rect 263604 696674 264204 696676
rect 299604 696674 300204 696676
rect 335604 696674 336204 696676
rect 371604 696674 372204 696676
rect 407604 696674 408204 696676
rect 443604 696674 444204 696676
rect 479604 696674 480204 696676
rect 515604 696674 516204 696676
rect 551604 696674 552204 696676
rect 590840 696674 591440 696676
rect -5676 693676 -5076 693678
rect 8004 693676 8604 693678
rect 44004 693676 44604 693678
rect 80004 693676 80604 693678
rect 116004 693676 116604 693678
rect 152004 693676 152604 693678
rect 188004 693676 188604 693678
rect 224004 693676 224604 693678
rect 260004 693676 260604 693678
rect 296004 693676 296604 693678
rect 332004 693676 332604 693678
rect 368004 693676 368604 693678
rect 404004 693676 404604 693678
rect 440004 693676 440604 693678
rect 476004 693676 476604 693678
rect 512004 693676 512604 693678
rect 548004 693676 548604 693678
rect 589000 693676 589600 693678
rect -6596 693654 590520 693676
rect -6596 693418 -5494 693654
rect -5258 693418 8186 693654
rect 8422 693418 44186 693654
rect 44422 693418 80186 693654
rect 80422 693418 116186 693654
rect 116422 693418 152186 693654
rect 152422 693418 188186 693654
rect 188422 693418 224186 693654
rect 224422 693418 260186 693654
rect 260422 693418 296186 693654
rect 296422 693418 332186 693654
rect 332422 693418 368186 693654
rect 368422 693418 404186 693654
rect 404422 693418 440186 693654
rect 440422 693418 476186 693654
rect 476422 693418 512186 693654
rect 512422 693418 548186 693654
rect 548422 693418 589182 693654
rect 589418 693418 590520 693654
rect -6596 693334 590520 693418
rect -6596 693098 -5494 693334
rect -5258 693098 8186 693334
rect 8422 693098 44186 693334
rect 44422 693098 80186 693334
rect 80422 693098 116186 693334
rect 116422 693098 152186 693334
rect 152422 693098 188186 693334
rect 188422 693098 224186 693334
rect 224422 693098 260186 693334
rect 260422 693098 296186 693334
rect 296422 693098 332186 693334
rect 332422 693098 368186 693334
rect 368422 693098 404186 693334
rect 404422 693098 440186 693334
rect 440422 693098 476186 693334
rect 476422 693098 512186 693334
rect 512422 693098 548186 693334
rect 548422 693098 589182 693334
rect 589418 693098 590520 693334
rect -6596 693076 590520 693098
rect -5676 693074 -5076 693076
rect 8004 693074 8604 693076
rect 44004 693074 44604 693076
rect 80004 693074 80604 693076
rect 116004 693074 116604 693076
rect 152004 693074 152604 693076
rect 188004 693074 188604 693076
rect 224004 693074 224604 693076
rect 260004 693074 260604 693076
rect 296004 693074 296604 693076
rect 332004 693074 332604 693076
rect 368004 693074 368604 693076
rect 404004 693074 404604 693076
rect 440004 693074 440604 693076
rect 476004 693074 476604 693076
rect 512004 693074 512604 693076
rect 548004 693074 548604 693076
rect 589000 693074 589600 693076
rect -3836 690076 -3236 690078
rect 4404 690076 5004 690078
rect 40404 690076 41004 690078
rect 76404 690076 77004 690078
rect 112404 690076 113004 690078
rect 148404 690076 149004 690078
rect 184404 690076 185004 690078
rect 220404 690076 221004 690078
rect 256404 690076 257004 690078
rect 292404 690076 293004 690078
rect 328404 690076 329004 690078
rect 364404 690076 365004 690078
rect 400404 690076 401004 690078
rect 436404 690076 437004 690078
rect 472404 690076 473004 690078
rect 508404 690076 509004 690078
rect 544404 690076 545004 690078
rect 580404 690076 581004 690078
rect 587160 690076 587760 690078
rect -4756 690054 588680 690076
rect -4756 689818 -3654 690054
rect -3418 689818 4586 690054
rect 4822 689818 40586 690054
rect 40822 689818 76586 690054
rect 76822 689818 112586 690054
rect 112822 689818 148586 690054
rect 148822 689818 184586 690054
rect 184822 689818 220586 690054
rect 220822 689818 256586 690054
rect 256822 689818 292586 690054
rect 292822 689818 328586 690054
rect 328822 689818 364586 690054
rect 364822 689818 400586 690054
rect 400822 689818 436586 690054
rect 436822 689818 472586 690054
rect 472822 689818 508586 690054
rect 508822 689818 544586 690054
rect 544822 689818 580586 690054
rect 580822 689818 587342 690054
rect 587578 689818 588680 690054
rect -4756 689734 588680 689818
rect -4756 689498 -3654 689734
rect -3418 689498 4586 689734
rect 4822 689498 40586 689734
rect 40822 689498 76586 689734
rect 76822 689498 112586 689734
rect 112822 689498 148586 689734
rect 148822 689498 184586 689734
rect 184822 689498 220586 689734
rect 220822 689498 256586 689734
rect 256822 689498 292586 689734
rect 292822 689498 328586 689734
rect 328822 689498 364586 689734
rect 364822 689498 400586 689734
rect 400822 689498 436586 689734
rect 436822 689498 472586 689734
rect 472822 689498 508586 689734
rect 508822 689498 544586 689734
rect 544822 689498 580586 689734
rect 580822 689498 587342 689734
rect 587578 689498 588680 689734
rect -4756 689476 588680 689498
rect -3836 689474 -3236 689476
rect 4404 689474 5004 689476
rect 40404 689474 41004 689476
rect 76404 689474 77004 689476
rect 112404 689474 113004 689476
rect 148404 689474 149004 689476
rect 184404 689474 185004 689476
rect 220404 689474 221004 689476
rect 256404 689474 257004 689476
rect 292404 689474 293004 689476
rect 328404 689474 329004 689476
rect 364404 689474 365004 689476
rect 400404 689474 401004 689476
rect 436404 689474 437004 689476
rect 472404 689474 473004 689476
rect 508404 689474 509004 689476
rect 544404 689474 545004 689476
rect 580404 689474 581004 689476
rect 587160 689474 587760 689476
rect -1996 686476 -1396 686478
rect 804 686476 1404 686478
rect 36804 686476 37404 686478
rect 72804 686476 73404 686478
rect 108804 686476 109404 686478
rect 144804 686476 145404 686478
rect 180804 686476 181404 686478
rect 216804 686476 217404 686478
rect 252804 686476 253404 686478
rect 288804 686476 289404 686478
rect 324804 686476 325404 686478
rect 360804 686476 361404 686478
rect 396804 686476 397404 686478
rect 432804 686476 433404 686478
rect 468804 686476 469404 686478
rect 504804 686476 505404 686478
rect 540804 686476 541404 686478
rect 576804 686476 577404 686478
rect 585320 686476 585920 686478
rect -2916 686454 586840 686476
rect -2916 686218 -1814 686454
rect -1578 686218 986 686454
rect 1222 686218 36986 686454
rect 37222 686218 72986 686454
rect 73222 686218 108986 686454
rect 109222 686218 144986 686454
rect 145222 686218 180986 686454
rect 181222 686218 216986 686454
rect 217222 686218 252986 686454
rect 253222 686218 288986 686454
rect 289222 686218 324986 686454
rect 325222 686218 360986 686454
rect 361222 686218 396986 686454
rect 397222 686218 432986 686454
rect 433222 686218 468986 686454
rect 469222 686218 504986 686454
rect 505222 686218 540986 686454
rect 541222 686218 576986 686454
rect 577222 686218 585502 686454
rect 585738 686218 586840 686454
rect -2916 686134 586840 686218
rect -2916 685898 -1814 686134
rect -1578 685898 986 686134
rect 1222 685898 36986 686134
rect 37222 685898 72986 686134
rect 73222 685898 108986 686134
rect 109222 685898 144986 686134
rect 145222 685898 180986 686134
rect 181222 685898 216986 686134
rect 217222 685898 252986 686134
rect 253222 685898 288986 686134
rect 289222 685898 324986 686134
rect 325222 685898 360986 686134
rect 361222 685898 396986 686134
rect 397222 685898 432986 686134
rect 433222 685898 468986 686134
rect 469222 685898 504986 686134
rect 505222 685898 540986 686134
rect 541222 685898 576986 686134
rect 577222 685898 585502 686134
rect 585738 685898 586840 686134
rect -2916 685876 586840 685898
rect -1996 685874 -1396 685876
rect 804 685874 1404 685876
rect 36804 685874 37404 685876
rect 72804 685874 73404 685876
rect 108804 685874 109404 685876
rect 144804 685874 145404 685876
rect 180804 685874 181404 685876
rect 216804 685874 217404 685876
rect 252804 685874 253404 685876
rect 288804 685874 289404 685876
rect 324804 685874 325404 685876
rect 360804 685874 361404 685876
rect 396804 685874 397404 685876
rect 432804 685874 433404 685876
rect 468804 685874 469404 685876
rect 504804 685874 505404 685876
rect 540804 685874 541404 685876
rect 576804 685874 577404 685876
rect 585320 685874 585920 685876
rect -8436 679276 -7836 679278
rect 29604 679276 30204 679278
rect 65604 679276 66204 679278
rect 101604 679276 102204 679278
rect 137604 679276 138204 679278
rect 173604 679276 174204 679278
rect 209604 679276 210204 679278
rect 245604 679276 246204 679278
rect 281604 679276 282204 679278
rect 317604 679276 318204 679278
rect 353604 679276 354204 679278
rect 389604 679276 390204 679278
rect 425604 679276 426204 679278
rect 461604 679276 462204 679278
rect 497604 679276 498204 679278
rect 533604 679276 534204 679278
rect 569604 679276 570204 679278
rect 591760 679276 592360 679278
rect -8436 679254 592360 679276
rect -8436 679018 -8254 679254
rect -8018 679018 29786 679254
rect 30022 679018 65786 679254
rect 66022 679018 101786 679254
rect 102022 679018 137786 679254
rect 138022 679018 173786 679254
rect 174022 679018 209786 679254
rect 210022 679018 245786 679254
rect 246022 679018 281786 679254
rect 282022 679018 317786 679254
rect 318022 679018 353786 679254
rect 354022 679018 389786 679254
rect 390022 679018 425786 679254
rect 426022 679018 461786 679254
rect 462022 679018 497786 679254
rect 498022 679018 533786 679254
rect 534022 679018 569786 679254
rect 570022 679018 591942 679254
rect 592178 679018 592360 679254
rect -8436 678934 592360 679018
rect -8436 678698 -8254 678934
rect -8018 678698 29786 678934
rect 30022 678698 65786 678934
rect 66022 678698 101786 678934
rect 102022 678698 137786 678934
rect 138022 678698 173786 678934
rect 174022 678698 209786 678934
rect 210022 678698 245786 678934
rect 246022 678698 281786 678934
rect 282022 678698 317786 678934
rect 318022 678698 353786 678934
rect 354022 678698 389786 678934
rect 390022 678698 425786 678934
rect 426022 678698 461786 678934
rect 462022 678698 497786 678934
rect 498022 678698 533786 678934
rect 534022 678698 569786 678934
rect 570022 678698 591942 678934
rect 592178 678698 592360 678934
rect -8436 678676 592360 678698
rect -8436 678674 -7836 678676
rect 29604 678674 30204 678676
rect 65604 678674 66204 678676
rect 101604 678674 102204 678676
rect 137604 678674 138204 678676
rect 173604 678674 174204 678676
rect 209604 678674 210204 678676
rect 245604 678674 246204 678676
rect 281604 678674 282204 678676
rect 317604 678674 318204 678676
rect 353604 678674 354204 678676
rect 389604 678674 390204 678676
rect 425604 678674 426204 678676
rect 461604 678674 462204 678676
rect 497604 678674 498204 678676
rect 533604 678674 534204 678676
rect 569604 678674 570204 678676
rect 591760 678674 592360 678676
rect -6596 675676 -5996 675678
rect 26004 675676 26604 675678
rect 62004 675676 62604 675678
rect 98004 675676 98604 675678
rect 134004 675676 134604 675678
rect 170004 675676 170604 675678
rect 206004 675676 206604 675678
rect 242004 675676 242604 675678
rect 278004 675676 278604 675678
rect 314004 675676 314604 675678
rect 350004 675676 350604 675678
rect 386004 675676 386604 675678
rect 422004 675676 422604 675678
rect 458004 675676 458604 675678
rect 494004 675676 494604 675678
rect 530004 675676 530604 675678
rect 566004 675676 566604 675678
rect 589920 675676 590520 675678
rect -6596 675654 590520 675676
rect -6596 675418 -6414 675654
rect -6178 675418 26186 675654
rect 26422 675418 62186 675654
rect 62422 675418 98186 675654
rect 98422 675418 134186 675654
rect 134422 675418 170186 675654
rect 170422 675418 206186 675654
rect 206422 675418 242186 675654
rect 242422 675418 278186 675654
rect 278422 675418 314186 675654
rect 314422 675418 350186 675654
rect 350422 675418 386186 675654
rect 386422 675418 422186 675654
rect 422422 675418 458186 675654
rect 458422 675418 494186 675654
rect 494422 675418 530186 675654
rect 530422 675418 566186 675654
rect 566422 675418 590102 675654
rect 590338 675418 590520 675654
rect -6596 675334 590520 675418
rect -6596 675098 -6414 675334
rect -6178 675098 26186 675334
rect 26422 675098 62186 675334
rect 62422 675098 98186 675334
rect 98422 675098 134186 675334
rect 134422 675098 170186 675334
rect 170422 675098 206186 675334
rect 206422 675098 242186 675334
rect 242422 675098 278186 675334
rect 278422 675098 314186 675334
rect 314422 675098 350186 675334
rect 350422 675098 386186 675334
rect 386422 675098 422186 675334
rect 422422 675098 458186 675334
rect 458422 675098 494186 675334
rect 494422 675098 530186 675334
rect 530422 675098 566186 675334
rect 566422 675098 590102 675334
rect 590338 675098 590520 675334
rect -6596 675076 590520 675098
rect -6596 675074 -5996 675076
rect 26004 675074 26604 675076
rect 62004 675074 62604 675076
rect 98004 675074 98604 675076
rect 134004 675074 134604 675076
rect 170004 675074 170604 675076
rect 206004 675074 206604 675076
rect 242004 675074 242604 675076
rect 278004 675074 278604 675076
rect 314004 675074 314604 675076
rect 350004 675074 350604 675076
rect 386004 675074 386604 675076
rect 422004 675074 422604 675076
rect 458004 675074 458604 675076
rect 494004 675074 494604 675076
rect 530004 675074 530604 675076
rect 566004 675074 566604 675076
rect 589920 675074 590520 675076
rect -4756 672076 -4156 672078
rect 22404 672076 23004 672078
rect 58404 672076 59004 672078
rect 94404 672076 95004 672078
rect 130404 672076 131004 672078
rect 166404 672076 167004 672078
rect 202404 672076 203004 672078
rect 238404 672076 239004 672078
rect 274404 672076 275004 672078
rect 310404 672076 311004 672078
rect 346404 672076 347004 672078
rect 382404 672076 383004 672078
rect 418404 672076 419004 672078
rect 454404 672076 455004 672078
rect 490404 672076 491004 672078
rect 526404 672076 527004 672078
rect 562404 672076 563004 672078
rect 588080 672076 588680 672078
rect -4756 672054 588680 672076
rect -4756 671818 -4574 672054
rect -4338 671818 22586 672054
rect 22822 671818 58586 672054
rect 58822 671818 94586 672054
rect 94822 671818 130586 672054
rect 130822 671818 166586 672054
rect 166822 671818 202586 672054
rect 202822 671818 238586 672054
rect 238822 671818 274586 672054
rect 274822 671818 310586 672054
rect 310822 671818 346586 672054
rect 346822 671818 382586 672054
rect 382822 671818 418586 672054
rect 418822 671818 454586 672054
rect 454822 671818 490586 672054
rect 490822 671818 526586 672054
rect 526822 671818 562586 672054
rect 562822 671818 588262 672054
rect 588498 671818 588680 672054
rect -4756 671734 588680 671818
rect -4756 671498 -4574 671734
rect -4338 671498 22586 671734
rect 22822 671498 58586 671734
rect 58822 671498 94586 671734
rect 94822 671498 130586 671734
rect 130822 671498 166586 671734
rect 166822 671498 202586 671734
rect 202822 671498 238586 671734
rect 238822 671498 274586 671734
rect 274822 671498 310586 671734
rect 310822 671498 346586 671734
rect 346822 671498 382586 671734
rect 382822 671498 418586 671734
rect 418822 671498 454586 671734
rect 454822 671498 490586 671734
rect 490822 671498 526586 671734
rect 526822 671498 562586 671734
rect 562822 671498 588262 671734
rect 588498 671498 588680 671734
rect -4756 671476 588680 671498
rect -4756 671474 -4156 671476
rect 22404 671474 23004 671476
rect 58404 671474 59004 671476
rect 94404 671474 95004 671476
rect 130404 671474 131004 671476
rect 166404 671474 167004 671476
rect 202404 671474 203004 671476
rect 238404 671474 239004 671476
rect 274404 671474 275004 671476
rect 310404 671474 311004 671476
rect 346404 671474 347004 671476
rect 382404 671474 383004 671476
rect 418404 671474 419004 671476
rect 454404 671474 455004 671476
rect 490404 671474 491004 671476
rect 526404 671474 527004 671476
rect 562404 671474 563004 671476
rect 588080 671474 588680 671476
rect -2916 668476 -2316 668478
rect 18804 668476 19404 668478
rect 54804 668476 55404 668478
rect 90804 668476 91404 668478
rect 126804 668476 127404 668478
rect 162804 668476 163404 668478
rect 198804 668476 199404 668478
rect 234804 668476 235404 668478
rect 270804 668476 271404 668478
rect 306804 668476 307404 668478
rect 342804 668476 343404 668478
rect 378804 668476 379404 668478
rect 414804 668476 415404 668478
rect 450804 668476 451404 668478
rect 486804 668476 487404 668478
rect 522804 668476 523404 668478
rect 558804 668476 559404 668478
rect 586240 668476 586840 668478
rect -2916 668454 586840 668476
rect -2916 668218 -2734 668454
rect -2498 668218 18986 668454
rect 19222 668218 54986 668454
rect 55222 668218 90986 668454
rect 91222 668218 126986 668454
rect 127222 668218 162986 668454
rect 163222 668218 198986 668454
rect 199222 668218 234986 668454
rect 235222 668218 270986 668454
rect 271222 668218 306986 668454
rect 307222 668218 342986 668454
rect 343222 668218 378986 668454
rect 379222 668218 414986 668454
rect 415222 668218 450986 668454
rect 451222 668218 486986 668454
rect 487222 668218 522986 668454
rect 523222 668218 558986 668454
rect 559222 668218 586422 668454
rect 586658 668218 586840 668454
rect -2916 668134 586840 668218
rect -2916 667898 -2734 668134
rect -2498 667898 18986 668134
rect 19222 667898 54986 668134
rect 55222 667898 90986 668134
rect 91222 667898 126986 668134
rect 127222 667898 162986 668134
rect 163222 667898 198986 668134
rect 199222 667898 234986 668134
rect 235222 667898 270986 668134
rect 271222 667898 306986 668134
rect 307222 667898 342986 668134
rect 343222 667898 378986 668134
rect 379222 667898 414986 668134
rect 415222 667898 450986 668134
rect 451222 667898 486986 668134
rect 487222 667898 522986 668134
rect 523222 667898 558986 668134
rect 559222 667898 586422 668134
rect 586658 667898 586840 668134
rect -2916 667876 586840 667898
rect -2916 667874 -2316 667876
rect 18804 667874 19404 667876
rect 54804 667874 55404 667876
rect 90804 667874 91404 667876
rect 126804 667874 127404 667876
rect 162804 667874 163404 667876
rect 198804 667874 199404 667876
rect 234804 667874 235404 667876
rect 270804 667874 271404 667876
rect 306804 667874 307404 667876
rect 342804 667874 343404 667876
rect 378804 667874 379404 667876
rect 414804 667874 415404 667876
rect 450804 667874 451404 667876
rect 486804 667874 487404 667876
rect 522804 667874 523404 667876
rect 558804 667874 559404 667876
rect 586240 667874 586840 667876
rect -7516 661276 -6916 661278
rect 11604 661276 12204 661278
rect 47604 661276 48204 661278
rect 83604 661276 84204 661278
rect 119604 661276 120204 661278
rect 155604 661276 156204 661278
rect 191604 661276 192204 661278
rect 227604 661276 228204 661278
rect 263604 661276 264204 661278
rect 299604 661276 300204 661278
rect 335604 661276 336204 661278
rect 371604 661276 372204 661278
rect 407604 661276 408204 661278
rect 443604 661276 444204 661278
rect 479604 661276 480204 661278
rect 515604 661276 516204 661278
rect 551604 661276 552204 661278
rect 590840 661276 591440 661278
rect -8436 661254 592360 661276
rect -8436 661018 -7334 661254
rect -7098 661018 11786 661254
rect 12022 661018 47786 661254
rect 48022 661018 83786 661254
rect 84022 661018 119786 661254
rect 120022 661018 155786 661254
rect 156022 661018 191786 661254
rect 192022 661018 227786 661254
rect 228022 661018 263786 661254
rect 264022 661018 299786 661254
rect 300022 661018 335786 661254
rect 336022 661018 371786 661254
rect 372022 661018 407786 661254
rect 408022 661018 443786 661254
rect 444022 661018 479786 661254
rect 480022 661018 515786 661254
rect 516022 661018 551786 661254
rect 552022 661018 591022 661254
rect 591258 661018 592360 661254
rect -8436 660934 592360 661018
rect -8436 660698 -7334 660934
rect -7098 660698 11786 660934
rect 12022 660698 47786 660934
rect 48022 660698 83786 660934
rect 84022 660698 119786 660934
rect 120022 660698 155786 660934
rect 156022 660698 191786 660934
rect 192022 660698 227786 660934
rect 228022 660698 263786 660934
rect 264022 660698 299786 660934
rect 300022 660698 335786 660934
rect 336022 660698 371786 660934
rect 372022 660698 407786 660934
rect 408022 660698 443786 660934
rect 444022 660698 479786 660934
rect 480022 660698 515786 660934
rect 516022 660698 551786 660934
rect 552022 660698 591022 660934
rect 591258 660698 592360 660934
rect -8436 660676 592360 660698
rect -7516 660674 -6916 660676
rect 11604 660674 12204 660676
rect 47604 660674 48204 660676
rect 83604 660674 84204 660676
rect 119604 660674 120204 660676
rect 155604 660674 156204 660676
rect 191604 660674 192204 660676
rect 227604 660674 228204 660676
rect 263604 660674 264204 660676
rect 299604 660674 300204 660676
rect 335604 660674 336204 660676
rect 371604 660674 372204 660676
rect 407604 660674 408204 660676
rect 443604 660674 444204 660676
rect 479604 660674 480204 660676
rect 515604 660674 516204 660676
rect 551604 660674 552204 660676
rect 590840 660674 591440 660676
rect -5676 657676 -5076 657678
rect 8004 657676 8604 657678
rect 44004 657676 44604 657678
rect 80004 657676 80604 657678
rect 116004 657676 116604 657678
rect 152004 657676 152604 657678
rect 188004 657676 188604 657678
rect 224004 657676 224604 657678
rect 260004 657676 260604 657678
rect 296004 657676 296604 657678
rect 332004 657676 332604 657678
rect 368004 657676 368604 657678
rect 404004 657676 404604 657678
rect 440004 657676 440604 657678
rect 476004 657676 476604 657678
rect 512004 657676 512604 657678
rect 548004 657676 548604 657678
rect 589000 657676 589600 657678
rect -6596 657654 590520 657676
rect -6596 657418 -5494 657654
rect -5258 657418 8186 657654
rect 8422 657418 44186 657654
rect 44422 657418 80186 657654
rect 80422 657418 116186 657654
rect 116422 657418 152186 657654
rect 152422 657418 188186 657654
rect 188422 657418 224186 657654
rect 224422 657418 260186 657654
rect 260422 657418 296186 657654
rect 296422 657418 332186 657654
rect 332422 657418 368186 657654
rect 368422 657418 404186 657654
rect 404422 657418 440186 657654
rect 440422 657418 476186 657654
rect 476422 657418 512186 657654
rect 512422 657418 548186 657654
rect 548422 657418 589182 657654
rect 589418 657418 590520 657654
rect -6596 657334 590520 657418
rect -6596 657098 -5494 657334
rect -5258 657098 8186 657334
rect 8422 657098 44186 657334
rect 44422 657098 80186 657334
rect 80422 657098 116186 657334
rect 116422 657098 152186 657334
rect 152422 657098 188186 657334
rect 188422 657098 224186 657334
rect 224422 657098 260186 657334
rect 260422 657098 296186 657334
rect 296422 657098 332186 657334
rect 332422 657098 368186 657334
rect 368422 657098 404186 657334
rect 404422 657098 440186 657334
rect 440422 657098 476186 657334
rect 476422 657098 512186 657334
rect 512422 657098 548186 657334
rect 548422 657098 589182 657334
rect 589418 657098 590520 657334
rect -6596 657076 590520 657098
rect -5676 657074 -5076 657076
rect 8004 657074 8604 657076
rect 44004 657074 44604 657076
rect 80004 657074 80604 657076
rect 116004 657074 116604 657076
rect 152004 657074 152604 657076
rect 188004 657074 188604 657076
rect 224004 657074 224604 657076
rect 260004 657074 260604 657076
rect 296004 657074 296604 657076
rect 332004 657074 332604 657076
rect 368004 657074 368604 657076
rect 404004 657074 404604 657076
rect 440004 657074 440604 657076
rect 476004 657074 476604 657076
rect 512004 657074 512604 657076
rect 548004 657074 548604 657076
rect 589000 657074 589600 657076
rect -3836 654076 -3236 654078
rect 4404 654076 5004 654078
rect 40404 654076 41004 654078
rect 76404 654076 77004 654078
rect 112404 654076 113004 654078
rect 148404 654076 149004 654078
rect 184404 654076 185004 654078
rect 220404 654076 221004 654078
rect 256404 654076 257004 654078
rect 292404 654076 293004 654078
rect 328404 654076 329004 654078
rect 364404 654076 365004 654078
rect 400404 654076 401004 654078
rect 436404 654076 437004 654078
rect 472404 654076 473004 654078
rect 508404 654076 509004 654078
rect 544404 654076 545004 654078
rect 580404 654076 581004 654078
rect 587160 654076 587760 654078
rect -4756 654054 588680 654076
rect -4756 653818 -3654 654054
rect -3418 653818 4586 654054
rect 4822 653818 40586 654054
rect 40822 653818 76586 654054
rect 76822 653818 112586 654054
rect 112822 653818 148586 654054
rect 148822 653818 184586 654054
rect 184822 653818 220586 654054
rect 220822 653818 256586 654054
rect 256822 653818 292586 654054
rect 292822 653818 328586 654054
rect 328822 653818 364586 654054
rect 364822 653818 400586 654054
rect 400822 653818 436586 654054
rect 436822 653818 472586 654054
rect 472822 653818 508586 654054
rect 508822 653818 544586 654054
rect 544822 653818 580586 654054
rect 580822 653818 587342 654054
rect 587578 653818 588680 654054
rect -4756 653734 588680 653818
rect -4756 653498 -3654 653734
rect -3418 653498 4586 653734
rect 4822 653498 40586 653734
rect 40822 653498 76586 653734
rect 76822 653498 112586 653734
rect 112822 653498 148586 653734
rect 148822 653498 184586 653734
rect 184822 653498 220586 653734
rect 220822 653498 256586 653734
rect 256822 653498 292586 653734
rect 292822 653498 328586 653734
rect 328822 653498 364586 653734
rect 364822 653498 400586 653734
rect 400822 653498 436586 653734
rect 436822 653498 472586 653734
rect 472822 653498 508586 653734
rect 508822 653498 544586 653734
rect 544822 653498 580586 653734
rect 580822 653498 587342 653734
rect 587578 653498 588680 653734
rect -4756 653476 588680 653498
rect -3836 653474 -3236 653476
rect 4404 653474 5004 653476
rect 40404 653474 41004 653476
rect 76404 653474 77004 653476
rect 112404 653474 113004 653476
rect 148404 653474 149004 653476
rect 184404 653474 185004 653476
rect 220404 653474 221004 653476
rect 256404 653474 257004 653476
rect 292404 653474 293004 653476
rect 328404 653474 329004 653476
rect 364404 653474 365004 653476
rect 400404 653474 401004 653476
rect 436404 653474 437004 653476
rect 472404 653474 473004 653476
rect 508404 653474 509004 653476
rect 544404 653474 545004 653476
rect 580404 653474 581004 653476
rect 587160 653474 587760 653476
rect -1996 650476 -1396 650478
rect 804 650476 1404 650478
rect 36804 650476 37404 650478
rect 72804 650476 73404 650478
rect 108804 650476 109404 650478
rect 144804 650476 145404 650478
rect 180804 650476 181404 650478
rect 216804 650476 217404 650478
rect 252804 650476 253404 650478
rect 288804 650476 289404 650478
rect 324804 650476 325404 650478
rect 360804 650476 361404 650478
rect 396804 650476 397404 650478
rect 432804 650476 433404 650478
rect 468804 650476 469404 650478
rect 504804 650476 505404 650478
rect 540804 650476 541404 650478
rect 576804 650476 577404 650478
rect 585320 650476 585920 650478
rect -2916 650454 586840 650476
rect -2916 650218 -1814 650454
rect -1578 650218 986 650454
rect 1222 650218 36986 650454
rect 37222 650218 72986 650454
rect 73222 650218 108986 650454
rect 109222 650218 144986 650454
rect 145222 650218 180986 650454
rect 181222 650218 216986 650454
rect 217222 650218 252986 650454
rect 253222 650218 288986 650454
rect 289222 650218 324986 650454
rect 325222 650218 360986 650454
rect 361222 650218 396986 650454
rect 397222 650218 432986 650454
rect 433222 650218 468986 650454
rect 469222 650218 504986 650454
rect 505222 650218 540986 650454
rect 541222 650218 576986 650454
rect 577222 650218 585502 650454
rect 585738 650218 586840 650454
rect -2916 650134 586840 650218
rect -2916 649898 -1814 650134
rect -1578 649898 986 650134
rect 1222 649898 36986 650134
rect 37222 649898 72986 650134
rect 73222 649898 108986 650134
rect 109222 649898 144986 650134
rect 145222 649898 180986 650134
rect 181222 649898 216986 650134
rect 217222 649898 252986 650134
rect 253222 649898 288986 650134
rect 289222 649898 324986 650134
rect 325222 649898 360986 650134
rect 361222 649898 396986 650134
rect 397222 649898 432986 650134
rect 433222 649898 468986 650134
rect 469222 649898 504986 650134
rect 505222 649898 540986 650134
rect 541222 649898 576986 650134
rect 577222 649898 585502 650134
rect 585738 649898 586840 650134
rect -2916 649876 586840 649898
rect -1996 649874 -1396 649876
rect 804 649874 1404 649876
rect 36804 649874 37404 649876
rect 72804 649874 73404 649876
rect 108804 649874 109404 649876
rect 144804 649874 145404 649876
rect 180804 649874 181404 649876
rect 216804 649874 217404 649876
rect 252804 649874 253404 649876
rect 288804 649874 289404 649876
rect 324804 649874 325404 649876
rect 360804 649874 361404 649876
rect 396804 649874 397404 649876
rect 432804 649874 433404 649876
rect 468804 649874 469404 649876
rect 504804 649874 505404 649876
rect 540804 649874 541404 649876
rect 576804 649874 577404 649876
rect 585320 649874 585920 649876
rect -8436 643276 -7836 643278
rect 29604 643276 30204 643278
rect 65604 643276 66204 643278
rect 101604 643276 102204 643278
rect 137604 643276 138204 643278
rect 173604 643276 174204 643278
rect 209604 643276 210204 643278
rect 245604 643276 246204 643278
rect 281604 643276 282204 643278
rect 317604 643276 318204 643278
rect 353604 643276 354204 643278
rect 389604 643276 390204 643278
rect 425604 643276 426204 643278
rect 461604 643276 462204 643278
rect 497604 643276 498204 643278
rect 533604 643276 534204 643278
rect 569604 643276 570204 643278
rect 591760 643276 592360 643278
rect -8436 643254 592360 643276
rect -8436 643018 -8254 643254
rect -8018 643018 29786 643254
rect 30022 643018 65786 643254
rect 66022 643018 101786 643254
rect 102022 643018 137786 643254
rect 138022 643018 173786 643254
rect 174022 643018 209786 643254
rect 210022 643018 245786 643254
rect 246022 643018 281786 643254
rect 282022 643018 317786 643254
rect 318022 643018 353786 643254
rect 354022 643018 389786 643254
rect 390022 643018 425786 643254
rect 426022 643018 461786 643254
rect 462022 643018 497786 643254
rect 498022 643018 533786 643254
rect 534022 643018 569786 643254
rect 570022 643018 591942 643254
rect 592178 643018 592360 643254
rect -8436 642934 592360 643018
rect -8436 642698 -8254 642934
rect -8018 642698 29786 642934
rect 30022 642698 65786 642934
rect 66022 642698 101786 642934
rect 102022 642698 137786 642934
rect 138022 642698 173786 642934
rect 174022 642698 209786 642934
rect 210022 642698 245786 642934
rect 246022 642698 281786 642934
rect 282022 642698 317786 642934
rect 318022 642698 353786 642934
rect 354022 642698 389786 642934
rect 390022 642698 425786 642934
rect 426022 642698 461786 642934
rect 462022 642698 497786 642934
rect 498022 642698 533786 642934
rect 534022 642698 569786 642934
rect 570022 642698 591942 642934
rect 592178 642698 592360 642934
rect -8436 642676 592360 642698
rect -8436 642674 -7836 642676
rect 29604 642674 30204 642676
rect 65604 642674 66204 642676
rect 101604 642674 102204 642676
rect 137604 642674 138204 642676
rect 173604 642674 174204 642676
rect 209604 642674 210204 642676
rect 245604 642674 246204 642676
rect 281604 642674 282204 642676
rect 317604 642674 318204 642676
rect 353604 642674 354204 642676
rect 389604 642674 390204 642676
rect 425604 642674 426204 642676
rect 461604 642674 462204 642676
rect 497604 642674 498204 642676
rect 533604 642674 534204 642676
rect 569604 642674 570204 642676
rect 591760 642674 592360 642676
rect -6596 639676 -5996 639678
rect 26004 639676 26604 639678
rect 62004 639676 62604 639678
rect 98004 639676 98604 639678
rect 134004 639676 134604 639678
rect 170004 639676 170604 639678
rect 206004 639676 206604 639678
rect 242004 639676 242604 639678
rect 278004 639676 278604 639678
rect 314004 639676 314604 639678
rect 350004 639676 350604 639678
rect 386004 639676 386604 639678
rect 422004 639676 422604 639678
rect 458004 639676 458604 639678
rect 494004 639676 494604 639678
rect 530004 639676 530604 639678
rect 566004 639676 566604 639678
rect 589920 639676 590520 639678
rect -6596 639654 590520 639676
rect -6596 639418 -6414 639654
rect -6178 639418 26186 639654
rect 26422 639418 62186 639654
rect 62422 639418 98186 639654
rect 98422 639418 134186 639654
rect 134422 639418 170186 639654
rect 170422 639418 206186 639654
rect 206422 639418 242186 639654
rect 242422 639418 278186 639654
rect 278422 639418 314186 639654
rect 314422 639418 350186 639654
rect 350422 639418 386186 639654
rect 386422 639418 422186 639654
rect 422422 639418 458186 639654
rect 458422 639418 494186 639654
rect 494422 639418 530186 639654
rect 530422 639418 566186 639654
rect 566422 639418 590102 639654
rect 590338 639418 590520 639654
rect -6596 639334 590520 639418
rect -6596 639098 -6414 639334
rect -6178 639098 26186 639334
rect 26422 639098 62186 639334
rect 62422 639098 98186 639334
rect 98422 639098 134186 639334
rect 134422 639098 170186 639334
rect 170422 639098 206186 639334
rect 206422 639098 242186 639334
rect 242422 639098 278186 639334
rect 278422 639098 314186 639334
rect 314422 639098 350186 639334
rect 350422 639098 386186 639334
rect 386422 639098 422186 639334
rect 422422 639098 458186 639334
rect 458422 639098 494186 639334
rect 494422 639098 530186 639334
rect 530422 639098 566186 639334
rect 566422 639098 590102 639334
rect 590338 639098 590520 639334
rect -6596 639076 590520 639098
rect -6596 639074 -5996 639076
rect 26004 639074 26604 639076
rect 62004 639074 62604 639076
rect 98004 639074 98604 639076
rect 134004 639074 134604 639076
rect 170004 639074 170604 639076
rect 206004 639074 206604 639076
rect 242004 639074 242604 639076
rect 278004 639074 278604 639076
rect 314004 639074 314604 639076
rect 350004 639074 350604 639076
rect 386004 639074 386604 639076
rect 422004 639074 422604 639076
rect 458004 639074 458604 639076
rect 494004 639074 494604 639076
rect 530004 639074 530604 639076
rect 566004 639074 566604 639076
rect 589920 639074 590520 639076
rect -4756 636076 -4156 636078
rect 22404 636076 23004 636078
rect 58404 636076 59004 636078
rect 94404 636076 95004 636078
rect 130404 636076 131004 636078
rect 166404 636076 167004 636078
rect 202404 636076 203004 636078
rect 238404 636076 239004 636078
rect 274404 636076 275004 636078
rect 310404 636076 311004 636078
rect 346404 636076 347004 636078
rect 382404 636076 383004 636078
rect 418404 636076 419004 636078
rect 454404 636076 455004 636078
rect 490404 636076 491004 636078
rect 526404 636076 527004 636078
rect 562404 636076 563004 636078
rect 588080 636076 588680 636078
rect -4756 636054 588680 636076
rect -4756 635818 -4574 636054
rect -4338 635818 22586 636054
rect 22822 635818 58586 636054
rect 58822 635818 94586 636054
rect 94822 635818 130586 636054
rect 130822 635818 166586 636054
rect 166822 635818 202586 636054
rect 202822 635818 238586 636054
rect 238822 635818 274586 636054
rect 274822 635818 310586 636054
rect 310822 635818 346586 636054
rect 346822 635818 382586 636054
rect 382822 635818 418586 636054
rect 418822 635818 454586 636054
rect 454822 635818 490586 636054
rect 490822 635818 526586 636054
rect 526822 635818 562586 636054
rect 562822 635818 588262 636054
rect 588498 635818 588680 636054
rect -4756 635734 588680 635818
rect -4756 635498 -4574 635734
rect -4338 635498 22586 635734
rect 22822 635498 58586 635734
rect 58822 635498 94586 635734
rect 94822 635498 130586 635734
rect 130822 635498 166586 635734
rect 166822 635498 202586 635734
rect 202822 635498 238586 635734
rect 238822 635498 274586 635734
rect 274822 635498 310586 635734
rect 310822 635498 346586 635734
rect 346822 635498 382586 635734
rect 382822 635498 418586 635734
rect 418822 635498 454586 635734
rect 454822 635498 490586 635734
rect 490822 635498 526586 635734
rect 526822 635498 562586 635734
rect 562822 635498 588262 635734
rect 588498 635498 588680 635734
rect -4756 635476 588680 635498
rect -4756 635474 -4156 635476
rect 22404 635474 23004 635476
rect 58404 635474 59004 635476
rect 94404 635474 95004 635476
rect 130404 635474 131004 635476
rect 166404 635474 167004 635476
rect 202404 635474 203004 635476
rect 238404 635474 239004 635476
rect 274404 635474 275004 635476
rect 310404 635474 311004 635476
rect 346404 635474 347004 635476
rect 382404 635474 383004 635476
rect 418404 635474 419004 635476
rect 454404 635474 455004 635476
rect 490404 635474 491004 635476
rect 526404 635474 527004 635476
rect 562404 635474 563004 635476
rect 588080 635474 588680 635476
rect -2916 632476 -2316 632478
rect 18804 632476 19404 632478
rect 54804 632476 55404 632478
rect 90804 632476 91404 632478
rect 126804 632476 127404 632478
rect 162804 632476 163404 632478
rect 198804 632476 199404 632478
rect 234804 632476 235404 632478
rect 270804 632476 271404 632478
rect 306804 632476 307404 632478
rect 342804 632476 343404 632478
rect 378804 632476 379404 632478
rect 414804 632476 415404 632478
rect 450804 632476 451404 632478
rect 486804 632476 487404 632478
rect 522804 632476 523404 632478
rect 558804 632476 559404 632478
rect 586240 632476 586840 632478
rect -2916 632454 586840 632476
rect -2916 632218 -2734 632454
rect -2498 632218 18986 632454
rect 19222 632218 54986 632454
rect 55222 632218 90986 632454
rect 91222 632218 126986 632454
rect 127222 632218 162986 632454
rect 163222 632218 198986 632454
rect 199222 632218 234986 632454
rect 235222 632218 270986 632454
rect 271222 632218 306986 632454
rect 307222 632218 342986 632454
rect 343222 632218 378986 632454
rect 379222 632218 414986 632454
rect 415222 632218 450986 632454
rect 451222 632218 486986 632454
rect 487222 632218 522986 632454
rect 523222 632218 558986 632454
rect 559222 632218 586422 632454
rect 586658 632218 586840 632454
rect -2916 632134 586840 632218
rect -2916 631898 -2734 632134
rect -2498 631898 18986 632134
rect 19222 631898 54986 632134
rect 55222 631898 90986 632134
rect 91222 631898 126986 632134
rect 127222 631898 162986 632134
rect 163222 631898 198986 632134
rect 199222 631898 234986 632134
rect 235222 631898 270986 632134
rect 271222 631898 306986 632134
rect 307222 631898 342986 632134
rect 343222 631898 378986 632134
rect 379222 631898 414986 632134
rect 415222 631898 450986 632134
rect 451222 631898 486986 632134
rect 487222 631898 522986 632134
rect 523222 631898 558986 632134
rect 559222 631898 586422 632134
rect 586658 631898 586840 632134
rect -2916 631876 586840 631898
rect -2916 631874 -2316 631876
rect 18804 631874 19404 631876
rect 54804 631874 55404 631876
rect 90804 631874 91404 631876
rect 126804 631874 127404 631876
rect 162804 631874 163404 631876
rect 198804 631874 199404 631876
rect 234804 631874 235404 631876
rect 270804 631874 271404 631876
rect 306804 631874 307404 631876
rect 342804 631874 343404 631876
rect 378804 631874 379404 631876
rect 414804 631874 415404 631876
rect 450804 631874 451404 631876
rect 486804 631874 487404 631876
rect 522804 631874 523404 631876
rect 558804 631874 559404 631876
rect 586240 631874 586840 631876
rect -7516 625276 -6916 625278
rect 11604 625276 12204 625278
rect 47604 625276 48204 625278
rect 83604 625276 84204 625278
rect 119604 625276 120204 625278
rect 155604 625276 156204 625278
rect 191604 625276 192204 625278
rect 227604 625276 228204 625278
rect 263604 625276 264204 625278
rect 299604 625276 300204 625278
rect 335604 625276 336204 625278
rect 371604 625276 372204 625278
rect 407604 625276 408204 625278
rect 443604 625276 444204 625278
rect 479604 625276 480204 625278
rect 515604 625276 516204 625278
rect 551604 625276 552204 625278
rect 590840 625276 591440 625278
rect -8436 625254 592360 625276
rect -8436 625018 -7334 625254
rect -7098 625018 11786 625254
rect 12022 625018 47786 625254
rect 48022 625018 83786 625254
rect 84022 625018 119786 625254
rect 120022 625018 155786 625254
rect 156022 625018 191786 625254
rect 192022 625018 227786 625254
rect 228022 625018 263786 625254
rect 264022 625018 299786 625254
rect 300022 625018 335786 625254
rect 336022 625018 371786 625254
rect 372022 625018 407786 625254
rect 408022 625018 443786 625254
rect 444022 625018 479786 625254
rect 480022 625018 515786 625254
rect 516022 625018 551786 625254
rect 552022 625018 591022 625254
rect 591258 625018 592360 625254
rect -8436 624934 592360 625018
rect -8436 624698 -7334 624934
rect -7098 624698 11786 624934
rect 12022 624698 47786 624934
rect 48022 624698 83786 624934
rect 84022 624698 119786 624934
rect 120022 624698 155786 624934
rect 156022 624698 191786 624934
rect 192022 624698 227786 624934
rect 228022 624698 263786 624934
rect 264022 624698 299786 624934
rect 300022 624698 335786 624934
rect 336022 624698 371786 624934
rect 372022 624698 407786 624934
rect 408022 624698 443786 624934
rect 444022 624698 479786 624934
rect 480022 624698 515786 624934
rect 516022 624698 551786 624934
rect 552022 624698 591022 624934
rect 591258 624698 592360 624934
rect -8436 624676 592360 624698
rect -7516 624674 -6916 624676
rect 11604 624674 12204 624676
rect 47604 624674 48204 624676
rect 83604 624674 84204 624676
rect 119604 624674 120204 624676
rect 155604 624674 156204 624676
rect 191604 624674 192204 624676
rect 227604 624674 228204 624676
rect 263604 624674 264204 624676
rect 299604 624674 300204 624676
rect 335604 624674 336204 624676
rect 371604 624674 372204 624676
rect 407604 624674 408204 624676
rect 443604 624674 444204 624676
rect 479604 624674 480204 624676
rect 515604 624674 516204 624676
rect 551604 624674 552204 624676
rect 590840 624674 591440 624676
rect -5676 621676 -5076 621678
rect 8004 621676 8604 621678
rect 44004 621676 44604 621678
rect 80004 621676 80604 621678
rect 116004 621676 116604 621678
rect 152004 621676 152604 621678
rect 188004 621676 188604 621678
rect 224004 621676 224604 621678
rect 260004 621676 260604 621678
rect 296004 621676 296604 621678
rect 332004 621676 332604 621678
rect 368004 621676 368604 621678
rect 404004 621676 404604 621678
rect 440004 621676 440604 621678
rect 476004 621676 476604 621678
rect 512004 621676 512604 621678
rect 548004 621676 548604 621678
rect 589000 621676 589600 621678
rect -6596 621654 590520 621676
rect -6596 621418 -5494 621654
rect -5258 621418 8186 621654
rect 8422 621418 44186 621654
rect 44422 621418 80186 621654
rect 80422 621418 116186 621654
rect 116422 621418 152186 621654
rect 152422 621418 188186 621654
rect 188422 621418 224186 621654
rect 224422 621418 260186 621654
rect 260422 621418 296186 621654
rect 296422 621418 332186 621654
rect 332422 621418 368186 621654
rect 368422 621418 404186 621654
rect 404422 621418 440186 621654
rect 440422 621418 476186 621654
rect 476422 621418 512186 621654
rect 512422 621418 548186 621654
rect 548422 621418 589182 621654
rect 589418 621418 590520 621654
rect -6596 621334 590520 621418
rect -6596 621098 -5494 621334
rect -5258 621098 8186 621334
rect 8422 621098 44186 621334
rect 44422 621098 80186 621334
rect 80422 621098 116186 621334
rect 116422 621098 152186 621334
rect 152422 621098 188186 621334
rect 188422 621098 224186 621334
rect 224422 621098 260186 621334
rect 260422 621098 296186 621334
rect 296422 621098 332186 621334
rect 332422 621098 368186 621334
rect 368422 621098 404186 621334
rect 404422 621098 440186 621334
rect 440422 621098 476186 621334
rect 476422 621098 512186 621334
rect 512422 621098 548186 621334
rect 548422 621098 589182 621334
rect 589418 621098 590520 621334
rect -6596 621076 590520 621098
rect -5676 621074 -5076 621076
rect 8004 621074 8604 621076
rect 44004 621074 44604 621076
rect 80004 621074 80604 621076
rect 116004 621074 116604 621076
rect 152004 621074 152604 621076
rect 188004 621074 188604 621076
rect 224004 621074 224604 621076
rect 260004 621074 260604 621076
rect 296004 621074 296604 621076
rect 332004 621074 332604 621076
rect 368004 621074 368604 621076
rect 404004 621074 404604 621076
rect 440004 621074 440604 621076
rect 476004 621074 476604 621076
rect 512004 621074 512604 621076
rect 548004 621074 548604 621076
rect 589000 621074 589600 621076
rect -3836 618076 -3236 618078
rect 4404 618076 5004 618078
rect 40404 618076 41004 618078
rect 76404 618076 77004 618078
rect 112404 618076 113004 618078
rect 148404 618076 149004 618078
rect 184404 618076 185004 618078
rect 220404 618076 221004 618078
rect 256404 618076 257004 618078
rect 292404 618076 293004 618078
rect 328404 618076 329004 618078
rect 364404 618076 365004 618078
rect 400404 618076 401004 618078
rect 436404 618076 437004 618078
rect 472404 618076 473004 618078
rect 508404 618076 509004 618078
rect 544404 618076 545004 618078
rect 580404 618076 581004 618078
rect 587160 618076 587760 618078
rect -4756 618054 588680 618076
rect -4756 617818 -3654 618054
rect -3418 617818 4586 618054
rect 4822 617818 40586 618054
rect 40822 617818 76586 618054
rect 76822 617818 112586 618054
rect 112822 617818 148586 618054
rect 148822 617818 184586 618054
rect 184822 617818 220586 618054
rect 220822 617818 256586 618054
rect 256822 617818 292586 618054
rect 292822 617818 328586 618054
rect 328822 617818 364586 618054
rect 364822 617818 400586 618054
rect 400822 617818 436586 618054
rect 436822 617818 472586 618054
rect 472822 617818 508586 618054
rect 508822 617818 544586 618054
rect 544822 617818 580586 618054
rect 580822 617818 587342 618054
rect 587578 617818 588680 618054
rect -4756 617734 588680 617818
rect -4756 617498 -3654 617734
rect -3418 617498 4586 617734
rect 4822 617498 40586 617734
rect 40822 617498 76586 617734
rect 76822 617498 112586 617734
rect 112822 617498 148586 617734
rect 148822 617498 184586 617734
rect 184822 617498 220586 617734
rect 220822 617498 256586 617734
rect 256822 617498 292586 617734
rect 292822 617498 328586 617734
rect 328822 617498 364586 617734
rect 364822 617498 400586 617734
rect 400822 617498 436586 617734
rect 436822 617498 472586 617734
rect 472822 617498 508586 617734
rect 508822 617498 544586 617734
rect 544822 617498 580586 617734
rect 580822 617498 587342 617734
rect 587578 617498 588680 617734
rect -4756 617476 588680 617498
rect -3836 617474 -3236 617476
rect 4404 617474 5004 617476
rect 40404 617474 41004 617476
rect 76404 617474 77004 617476
rect 112404 617474 113004 617476
rect 148404 617474 149004 617476
rect 184404 617474 185004 617476
rect 220404 617474 221004 617476
rect 256404 617474 257004 617476
rect 292404 617474 293004 617476
rect 328404 617474 329004 617476
rect 364404 617474 365004 617476
rect 400404 617474 401004 617476
rect 436404 617474 437004 617476
rect 472404 617474 473004 617476
rect 508404 617474 509004 617476
rect 544404 617474 545004 617476
rect 580404 617474 581004 617476
rect 587160 617474 587760 617476
rect -1996 614476 -1396 614478
rect 804 614476 1404 614478
rect 36804 614476 37404 614478
rect 72804 614476 73404 614478
rect 108804 614476 109404 614478
rect 144804 614476 145404 614478
rect 180804 614476 181404 614478
rect 216804 614476 217404 614478
rect 252804 614476 253404 614478
rect 288804 614476 289404 614478
rect 324804 614476 325404 614478
rect 360804 614476 361404 614478
rect 396804 614476 397404 614478
rect 432804 614476 433404 614478
rect 468804 614476 469404 614478
rect 504804 614476 505404 614478
rect 540804 614476 541404 614478
rect 576804 614476 577404 614478
rect 585320 614476 585920 614478
rect -2916 614454 586840 614476
rect -2916 614218 -1814 614454
rect -1578 614218 986 614454
rect 1222 614218 36986 614454
rect 37222 614218 72986 614454
rect 73222 614218 108986 614454
rect 109222 614218 144986 614454
rect 145222 614218 180986 614454
rect 181222 614218 216986 614454
rect 217222 614218 252986 614454
rect 253222 614218 288986 614454
rect 289222 614218 324986 614454
rect 325222 614218 360986 614454
rect 361222 614218 396986 614454
rect 397222 614218 432986 614454
rect 433222 614218 468986 614454
rect 469222 614218 504986 614454
rect 505222 614218 540986 614454
rect 541222 614218 576986 614454
rect 577222 614218 585502 614454
rect 585738 614218 586840 614454
rect -2916 614134 586840 614218
rect -2916 613898 -1814 614134
rect -1578 613898 986 614134
rect 1222 613898 36986 614134
rect 37222 613898 72986 614134
rect 73222 613898 108986 614134
rect 109222 613898 144986 614134
rect 145222 613898 180986 614134
rect 181222 613898 216986 614134
rect 217222 613898 252986 614134
rect 253222 613898 288986 614134
rect 289222 613898 324986 614134
rect 325222 613898 360986 614134
rect 361222 613898 396986 614134
rect 397222 613898 432986 614134
rect 433222 613898 468986 614134
rect 469222 613898 504986 614134
rect 505222 613898 540986 614134
rect 541222 613898 576986 614134
rect 577222 613898 585502 614134
rect 585738 613898 586840 614134
rect -2916 613876 586840 613898
rect -1996 613874 -1396 613876
rect 804 613874 1404 613876
rect 36804 613874 37404 613876
rect 72804 613874 73404 613876
rect 108804 613874 109404 613876
rect 144804 613874 145404 613876
rect 180804 613874 181404 613876
rect 216804 613874 217404 613876
rect 252804 613874 253404 613876
rect 288804 613874 289404 613876
rect 324804 613874 325404 613876
rect 360804 613874 361404 613876
rect 396804 613874 397404 613876
rect 432804 613874 433404 613876
rect 468804 613874 469404 613876
rect 504804 613874 505404 613876
rect 540804 613874 541404 613876
rect 576804 613874 577404 613876
rect 585320 613874 585920 613876
rect -8436 607276 -7836 607278
rect 29604 607276 30204 607278
rect 65604 607276 66204 607278
rect 101604 607276 102204 607278
rect 137604 607276 138204 607278
rect 173604 607276 174204 607278
rect 209604 607276 210204 607278
rect 245604 607276 246204 607278
rect 281604 607276 282204 607278
rect 317604 607276 318204 607278
rect 353604 607276 354204 607278
rect 389604 607276 390204 607278
rect 425604 607276 426204 607278
rect 461604 607276 462204 607278
rect 497604 607276 498204 607278
rect 533604 607276 534204 607278
rect 569604 607276 570204 607278
rect 591760 607276 592360 607278
rect -8436 607254 592360 607276
rect -8436 607018 -8254 607254
rect -8018 607018 29786 607254
rect 30022 607018 65786 607254
rect 66022 607018 101786 607254
rect 102022 607018 137786 607254
rect 138022 607018 173786 607254
rect 174022 607018 209786 607254
rect 210022 607018 245786 607254
rect 246022 607018 281786 607254
rect 282022 607018 317786 607254
rect 318022 607018 353786 607254
rect 354022 607018 389786 607254
rect 390022 607018 425786 607254
rect 426022 607018 461786 607254
rect 462022 607018 497786 607254
rect 498022 607018 533786 607254
rect 534022 607018 569786 607254
rect 570022 607018 591942 607254
rect 592178 607018 592360 607254
rect -8436 606934 592360 607018
rect -8436 606698 -8254 606934
rect -8018 606698 29786 606934
rect 30022 606698 65786 606934
rect 66022 606698 101786 606934
rect 102022 606698 137786 606934
rect 138022 606698 173786 606934
rect 174022 606698 209786 606934
rect 210022 606698 245786 606934
rect 246022 606698 281786 606934
rect 282022 606698 317786 606934
rect 318022 606698 353786 606934
rect 354022 606698 389786 606934
rect 390022 606698 425786 606934
rect 426022 606698 461786 606934
rect 462022 606698 497786 606934
rect 498022 606698 533786 606934
rect 534022 606698 569786 606934
rect 570022 606698 591942 606934
rect 592178 606698 592360 606934
rect -8436 606676 592360 606698
rect -8436 606674 -7836 606676
rect 29604 606674 30204 606676
rect 65604 606674 66204 606676
rect 101604 606674 102204 606676
rect 137604 606674 138204 606676
rect 173604 606674 174204 606676
rect 209604 606674 210204 606676
rect 245604 606674 246204 606676
rect 281604 606674 282204 606676
rect 317604 606674 318204 606676
rect 353604 606674 354204 606676
rect 389604 606674 390204 606676
rect 425604 606674 426204 606676
rect 461604 606674 462204 606676
rect 497604 606674 498204 606676
rect 533604 606674 534204 606676
rect 569604 606674 570204 606676
rect 591760 606674 592360 606676
rect -6596 603676 -5996 603678
rect 26004 603676 26604 603678
rect 62004 603676 62604 603678
rect 98004 603676 98604 603678
rect 134004 603676 134604 603678
rect 170004 603676 170604 603678
rect 206004 603676 206604 603678
rect 242004 603676 242604 603678
rect 278004 603676 278604 603678
rect 314004 603676 314604 603678
rect 350004 603676 350604 603678
rect 386004 603676 386604 603678
rect 422004 603676 422604 603678
rect 458004 603676 458604 603678
rect 494004 603676 494604 603678
rect 530004 603676 530604 603678
rect 566004 603676 566604 603678
rect 589920 603676 590520 603678
rect -6596 603654 590520 603676
rect -6596 603418 -6414 603654
rect -6178 603418 26186 603654
rect 26422 603418 62186 603654
rect 62422 603418 98186 603654
rect 98422 603418 134186 603654
rect 134422 603418 170186 603654
rect 170422 603418 206186 603654
rect 206422 603418 242186 603654
rect 242422 603418 278186 603654
rect 278422 603418 314186 603654
rect 314422 603418 350186 603654
rect 350422 603418 386186 603654
rect 386422 603418 422186 603654
rect 422422 603418 458186 603654
rect 458422 603418 494186 603654
rect 494422 603418 530186 603654
rect 530422 603418 566186 603654
rect 566422 603418 590102 603654
rect 590338 603418 590520 603654
rect -6596 603334 590520 603418
rect -6596 603098 -6414 603334
rect -6178 603098 26186 603334
rect 26422 603098 62186 603334
rect 62422 603098 98186 603334
rect 98422 603098 134186 603334
rect 134422 603098 170186 603334
rect 170422 603098 206186 603334
rect 206422 603098 242186 603334
rect 242422 603098 278186 603334
rect 278422 603098 314186 603334
rect 314422 603098 350186 603334
rect 350422 603098 386186 603334
rect 386422 603098 422186 603334
rect 422422 603098 458186 603334
rect 458422 603098 494186 603334
rect 494422 603098 530186 603334
rect 530422 603098 566186 603334
rect 566422 603098 590102 603334
rect 590338 603098 590520 603334
rect -6596 603076 590520 603098
rect -6596 603074 -5996 603076
rect 26004 603074 26604 603076
rect 62004 603074 62604 603076
rect 98004 603074 98604 603076
rect 134004 603074 134604 603076
rect 170004 603074 170604 603076
rect 206004 603074 206604 603076
rect 242004 603074 242604 603076
rect 278004 603074 278604 603076
rect 314004 603074 314604 603076
rect 350004 603074 350604 603076
rect 386004 603074 386604 603076
rect 422004 603074 422604 603076
rect 458004 603074 458604 603076
rect 494004 603074 494604 603076
rect 530004 603074 530604 603076
rect 566004 603074 566604 603076
rect 589920 603074 590520 603076
rect -4756 600076 -4156 600078
rect 22404 600076 23004 600078
rect 58404 600076 59004 600078
rect 94404 600076 95004 600078
rect 130404 600076 131004 600078
rect 166404 600076 167004 600078
rect 202404 600076 203004 600078
rect 238404 600076 239004 600078
rect 274404 600076 275004 600078
rect 310404 600076 311004 600078
rect 346404 600076 347004 600078
rect 382404 600076 383004 600078
rect 418404 600076 419004 600078
rect 454404 600076 455004 600078
rect 490404 600076 491004 600078
rect 526404 600076 527004 600078
rect 562404 600076 563004 600078
rect 588080 600076 588680 600078
rect -4756 600054 588680 600076
rect -4756 599818 -4574 600054
rect -4338 599818 22586 600054
rect 22822 599818 58586 600054
rect 58822 599818 94586 600054
rect 94822 599818 130586 600054
rect 130822 599818 166586 600054
rect 166822 599818 202586 600054
rect 202822 599818 238586 600054
rect 238822 599818 274586 600054
rect 274822 599818 310586 600054
rect 310822 599818 346586 600054
rect 346822 599818 382586 600054
rect 382822 599818 418586 600054
rect 418822 599818 454586 600054
rect 454822 599818 490586 600054
rect 490822 599818 526586 600054
rect 526822 599818 562586 600054
rect 562822 599818 588262 600054
rect 588498 599818 588680 600054
rect -4756 599734 588680 599818
rect -4756 599498 -4574 599734
rect -4338 599498 22586 599734
rect 22822 599498 58586 599734
rect 58822 599498 94586 599734
rect 94822 599498 130586 599734
rect 130822 599498 166586 599734
rect 166822 599498 202586 599734
rect 202822 599498 238586 599734
rect 238822 599498 274586 599734
rect 274822 599498 310586 599734
rect 310822 599498 346586 599734
rect 346822 599498 382586 599734
rect 382822 599498 418586 599734
rect 418822 599498 454586 599734
rect 454822 599498 490586 599734
rect 490822 599498 526586 599734
rect 526822 599498 562586 599734
rect 562822 599498 588262 599734
rect 588498 599498 588680 599734
rect -4756 599476 588680 599498
rect -4756 599474 -4156 599476
rect 22404 599474 23004 599476
rect 58404 599474 59004 599476
rect 94404 599474 95004 599476
rect 130404 599474 131004 599476
rect 166404 599474 167004 599476
rect 202404 599474 203004 599476
rect 238404 599474 239004 599476
rect 274404 599474 275004 599476
rect 310404 599474 311004 599476
rect 346404 599474 347004 599476
rect 382404 599474 383004 599476
rect 418404 599474 419004 599476
rect 454404 599474 455004 599476
rect 490404 599474 491004 599476
rect 526404 599474 527004 599476
rect 562404 599474 563004 599476
rect 588080 599474 588680 599476
rect -2916 596476 -2316 596478
rect 18804 596476 19404 596478
rect 54804 596476 55404 596478
rect 90804 596476 91404 596478
rect 126804 596476 127404 596478
rect 162804 596476 163404 596478
rect 198804 596476 199404 596478
rect 234804 596476 235404 596478
rect 270804 596476 271404 596478
rect 306804 596476 307404 596478
rect 342804 596476 343404 596478
rect 378804 596476 379404 596478
rect 414804 596476 415404 596478
rect 450804 596476 451404 596478
rect 486804 596476 487404 596478
rect 522804 596476 523404 596478
rect 558804 596476 559404 596478
rect 586240 596476 586840 596478
rect -2916 596454 586840 596476
rect -2916 596218 -2734 596454
rect -2498 596218 18986 596454
rect 19222 596218 54986 596454
rect 55222 596218 90986 596454
rect 91222 596218 126986 596454
rect 127222 596218 162986 596454
rect 163222 596218 198986 596454
rect 199222 596218 234986 596454
rect 235222 596218 270986 596454
rect 271222 596218 306986 596454
rect 307222 596218 342986 596454
rect 343222 596218 378986 596454
rect 379222 596218 414986 596454
rect 415222 596218 450986 596454
rect 451222 596218 486986 596454
rect 487222 596218 522986 596454
rect 523222 596218 558986 596454
rect 559222 596218 586422 596454
rect 586658 596218 586840 596454
rect -2916 596134 586840 596218
rect -2916 595898 -2734 596134
rect -2498 595898 18986 596134
rect 19222 595898 54986 596134
rect 55222 595898 90986 596134
rect 91222 595898 126986 596134
rect 127222 595898 162986 596134
rect 163222 595898 198986 596134
rect 199222 595898 234986 596134
rect 235222 595898 270986 596134
rect 271222 595898 306986 596134
rect 307222 595898 342986 596134
rect 343222 595898 378986 596134
rect 379222 595898 414986 596134
rect 415222 595898 450986 596134
rect 451222 595898 486986 596134
rect 487222 595898 522986 596134
rect 523222 595898 558986 596134
rect 559222 595898 586422 596134
rect 586658 595898 586840 596134
rect -2916 595876 586840 595898
rect -2916 595874 -2316 595876
rect 18804 595874 19404 595876
rect 54804 595874 55404 595876
rect 90804 595874 91404 595876
rect 126804 595874 127404 595876
rect 162804 595874 163404 595876
rect 198804 595874 199404 595876
rect 234804 595874 235404 595876
rect 270804 595874 271404 595876
rect 306804 595874 307404 595876
rect 342804 595874 343404 595876
rect 378804 595874 379404 595876
rect 414804 595874 415404 595876
rect 450804 595874 451404 595876
rect 486804 595874 487404 595876
rect 522804 595874 523404 595876
rect 558804 595874 559404 595876
rect 586240 595874 586840 595876
rect -7516 589276 -6916 589278
rect 11604 589276 12204 589278
rect 47604 589276 48204 589278
rect 83604 589276 84204 589278
rect 119604 589276 120204 589278
rect 155604 589276 156204 589278
rect 191604 589276 192204 589278
rect 227604 589276 228204 589278
rect 263604 589276 264204 589278
rect 299604 589276 300204 589278
rect 335604 589276 336204 589278
rect 371604 589276 372204 589278
rect 407604 589276 408204 589278
rect 443604 589276 444204 589278
rect 479604 589276 480204 589278
rect 515604 589276 516204 589278
rect 551604 589276 552204 589278
rect 590840 589276 591440 589278
rect -8436 589254 592360 589276
rect -8436 589018 -7334 589254
rect -7098 589018 11786 589254
rect 12022 589018 47786 589254
rect 48022 589018 83786 589254
rect 84022 589018 119786 589254
rect 120022 589018 155786 589254
rect 156022 589018 191786 589254
rect 192022 589018 227786 589254
rect 228022 589018 263786 589254
rect 264022 589018 299786 589254
rect 300022 589018 335786 589254
rect 336022 589018 371786 589254
rect 372022 589018 407786 589254
rect 408022 589018 443786 589254
rect 444022 589018 479786 589254
rect 480022 589018 515786 589254
rect 516022 589018 551786 589254
rect 552022 589018 591022 589254
rect 591258 589018 592360 589254
rect -8436 588934 592360 589018
rect -8436 588698 -7334 588934
rect -7098 588698 11786 588934
rect 12022 588698 47786 588934
rect 48022 588698 83786 588934
rect 84022 588698 119786 588934
rect 120022 588698 155786 588934
rect 156022 588698 191786 588934
rect 192022 588698 227786 588934
rect 228022 588698 263786 588934
rect 264022 588698 299786 588934
rect 300022 588698 335786 588934
rect 336022 588698 371786 588934
rect 372022 588698 407786 588934
rect 408022 588698 443786 588934
rect 444022 588698 479786 588934
rect 480022 588698 515786 588934
rect 516022 588698 551786 588934
rect 552022 588698 591022 588934
rect 591258 588698 592360 588934
rect -8436 588676 592360 588698
rect -7516 588674 -6916 588676
rect 11604 588674 12204 588676
rect 47604 588674 48204 588676
rect 83604 588674 84204 588676
rect 119604 588674 120204 588676
rect 155604 588674 156204 588676
rect 191604 588674 192204 588676
rect 227604 588674 228204 588676
rect 263604 588674 264204 588676
rect 299604 588674 300204 588676
rect 335604 588674 336204 588676
rect 371604 588674 372204 588676
rect 407604 588674 408204 588676
rect 443604 588674 444204 588676
rect 479604 588674 480204 588676
rect 515604 588674 516204 588676
rect 551604 588674 552204 588676
rect 590840 588674 591440 588676
rect -5676 585676 -5076 585678
rect 8004 585676 8604 585678
rect 44004 585676 44604 585678
rect 80004 585676 80604 585678
rect 116004 585676 116604 585678
rect 152004 585676 152604 585678
rect 188004 585676 188604 585678
rect 224004 585676 224604 585678
rect 260004 585676 260604 585678
rect 296004 585676 296604 585678
rect 332004 585676 332604 585678
rect 368004 585676 368604 585678
rect 404004 585676 404604 585678
rect 440004 585676 440604 585678
rect 476004 585676 476604 585678
rect 512004 585676 512604 585678
rect 548004 585676 548604 585678
rect 589000 585676 589600 585678
rect -6596 585654 590520 585676
rect -6596 585418 -5494 585654
rect -5258 585418 8186 585654
rect 8422 585418 44186 585654
rect 44422 585418 80186 585654
rect 80422 585418 116186 585654
rect 116422 585418 152186 585654
rect 152422 585418 188186 585654
rect 188422 585418 224186 585654
rect 224422 585418 260186 585654
rect 260422 585418 296186 585654
rect 296422 585418 332186 585654
rect 332422 585418 368186 585654
rect 368422 585418 404186 585654
rect 404422 585418 440186 585654
rect 440422 585418 476186 585654
rect 476422 585418 512186 585654
rect 512422 585418 548186 585654
rect 548422 585418 589182 585654
rect 589418 585418 590520 585654
rect -6596 585334 590520 585418
rect -6596 585098 -5494 585334
rect -5258 585098 8186 585334
rect 8422 585098 44186 585334
rect 44422 585098 80186 585334
rect 80422 585098 116186 585334
rect 116422 585098 152186 585334
rect 152422 585098 188186 585334
rect 188422 585098 224186 585334
rect 224422 585098 260186 585334
rect 260422 585098 296186 585334
rect 296422 585098 332186 585334
rect 332422 585098 368186 585334
rect 368422 585098 404186 585334
rect 404422 585098 440186 585334
rect 440422 585098 476186 585334
rect 476422 585098 512186 585334
rect 512422 585098 548186 585334
rect 548422 585098 589182 585334
rect 589418 585098 590520 585334
rect -6596 585076 590520 585098
rect -5676 585074 -5076 585076
rect 8004 585074 8604 585076
rect 44004 585074 44604 585076
rect 80004 585074 80604 585076
rect 116004 585074 116604 585076
rect 152004 585074 152604 585076
rect 188004 585074 188604 585076
rect 224004 585074 224604 585076
rect 260004 585074 260604 585076
rect 296004 585074 296604 585076
rect 332004 585074 332604 585076
rect 368004 585074 368604 585076
rect 404004 585074 404604 585076
rect 440004 585074 440604 585076
rect 476004 585074 476604 585076
rect 512004 585074 512604 585076
rect 548004 585074 548604 585076
rect 589000 585074 589600 585076
rect -3836 582076 -3236 582078
rect 4404 582076 5004 582078
rect 40404 582076 41004 582078
rect 76404 582076 77004 582078
rect 112404 582076 113004 582078
rect 148404 582076 149004 582078
rect 184404 582076 185004 582078
rect 220404 582076 221004 582078
rect 256404 582076 257004 582078
rect 292404 582076 293004 582078
rect 328404 582076 329004 582078
rect 364404 582076 365004 582078
rect 400404 582076 401004 582078
rect 436404 582076 437004 582078
rect 472404 582076 473004 582078
rect 508404 582076 509004 582078
rect 544404 582076 545004 582078
rect 580404 582076 581004 582078
rect 587160 582076 587760 582078
rect -4756 582054 588680 582076
rect -4756 581818 -3654 582054
rect -3418 581818 4586 582054
rect 4822 581818 40586 582054
rect 40822 581818 76586 582054
rect 76822 581818 112586 582054
rect 112822 581818 148586 582054
rect 148822 581818 184586 582054
rect 184822 581818 220586 582054
rect 220822 581818 256586 582054
rect 256822 581818 292586 582054
rect 292822 581818 328586 582054
rect 328822 581818 364586 582054
rect 364822 581818 400586 582054
rect 400822 581818 436586 582054
rect 436822 581818 472586 582054
rect 472822 581818 508586 582054
rect 508822 581818 544586 582054
rect 544822 581818 580586 582054
rect 580822 581818 587342 582054
rect 587578 581818 588680 582054
rect -4756 581734 588680 581818
rect -4756 581498 -3654 581734
rect -3418 581498 4586 581734
rect 4822 581498 40586 581734
rect 40822 581498 76586 581734
rect 76822 581498 112586 581734
rect 112822 581498 148586 581734
rect 148822 581498 184586 581734
rect 184822 581498 220586 581734
rect 220822 581498 256586 581734
rect 256822 581498 292586 581734
rect 292822 581498 328586 581734
rect 328822 581498 364586 581734
rect 364822 581498 400586 581734
rect 400822 581498 436586 581734
rect 436822 581498 472586 581734
rect 472822 581498 508586 581734
rect 508822 581498 544586 581734
rect 544822 581498 580586 581734
rect 580822 581498 587342 581734
rect 587578 581498 588680 581734
rect -4756 581476 588680 581498
rect -3836 581474 -3236 581476
rect 4404 581474 5004 581476
rect 40404 581474 41004 581476
rect 76404 581474 77004 581476
rect 112404 581474 113004 581476
rect 148404 581474 149004 581476
rect 184404 581474 185004 581476
rect 220404 581474 221004 581476
rect 256404 581474 257004 581476
rect 292404 581474 293004 581476
rect 328404 581474 329004 581476
rect 364404 581474 365004 581476
rect 400404 581474 401004 581476
rect 436404 581474 437004 581476
rect 472404 581474 473004 581476
rect 508404 581474 509004 581476
rect 544404 581474 545004 581476
rect 580404 581474 581004 581476
rect 587160 581474 587760 581476
rect -1996 578476 -1396 578478
rect 804 578476 1404 578478
rect 36804 578476 37404 578478
rect 72804 578476 73404 578478
rect 108804 578476 109404 578478
rect 144804 578476 145404 578478
rect 180804 578476 181404 578478
rect 216804 578476 217404 578478
rect 252804 578476 253404 578478
rect 288804 578476 289404 578478
rect 324804 578476 325404 578478
rect 360804 578476 361404 578478
rect 396804 578476 397404 578478
rect 432804 578476 433404 578478
rect 468804 578476 469404 578478
rect 504804 578476 505404 578478
rect 540804 578476 541404 578478
rect 576804 578476 577404 578478
rect 585320 578476 585920 578478
rect -2916 578454 586840 578476
rect -2916 578218 -1814 578454
rect -1578 578218 986 578454
rect 1222 578218 36986 578454
rect 37222 578218 72986 578454
rect 73222 578218 108986 578454
rect 109222 578218 144986 578454
rect 145222 578218 180986 578454
rect 181222 578218 216986 578454
rect 217222 578218 252986 578454
rect 253222 578218 288986 578454
rect 289222 578218 324986 578454
rect 325222 578218 360986 578454
rect 361222 578218 396986 578454
rect 397222 578218 432986 578454
rect 433222 578218 468986 578454
rect 469222 578218 504986 578454
rect 505222 578218 540986 578454
rect 541222 578218 576986 578454
rect 577222 578218 585502 578454
rect 585738 578218 586840 578454
rect -2916 578134 586840 578218
rect -2916 577898 -1814 578134
rect -1578 577898 986 578134
rect 1222 577898 36986 578134
rect 37222 577898 72986 578134
rect 73222 577898 108986 578134
rect 109222 577898 144986 578134
rect 145222 577898 180986 578134
rect 181222 577898 216986 578134
rect 217222 577898 252986 578134
rect 253222 577898 288986 578134
rect 289222 577898 324986 578134
rect 325222 577898 360986 578134
rect 361222 577898 396986 578134
rect 397222 577898 432986 578134
rect 433222 577898 468986 578134
rect 469222 577898 504986 578134
rect 505222 577898 540986 578134
rect 541222 577898 576986 578134
rect 577222 577898 585502 578134
rect 585738 577898 586840 578134
rect -2916 577876 586840 577898
rect -1996 577874 -1396 577876
rect 804 577874 1404 577876
rect 36804 577874 37404 577876
rect 72804 577874 73404 577876
rect 108804 577874 109404 577876
rect 144804 577874 145404 577876
rect 180804 577874 181404 577876
rect 216804 577874 217404 577876
rect 252804 577874 253404 577876
rect 288804 577874 289404 577876
rect 324804 577874 325404 577876
rect 360804 577874 361404 577876
rect 396804 577874 397404 577876
rect 432804 577874 433404 577876
rect 468804 577874 469404 577876
rect 504804 577874 505404 577876
rect 540804 577874 541404 577876
rect 576804 577874 577404 577876
rect 585320 577874 585920 577876
rect -8436 571276 -7836 571278
rect 29604 571276 30204 571278
rect 65604 571276 66204 571278
rect 101604 571276 102204 571278
rect 137604 571276 138204 571278
rect 173604 571276 174204 571278
rect 209604 571276 210204 571278
rect 245604 571276 246204 571278
rect 281604 571276 282204 571278
rect 317604 571276 318204 571278
rect 353604 571276 354204 571278
rect 389604 571276 390204 571278
rect 425604 571276 426204 571278
rect 461604 571276 462204 571278
rect 497604 571276 498204 571278
rect 533604 571276 534204 571278
rect 569604 571276 570204 571278
rect 591760 571276 592360 571278
rect -8436 571254 592360 571276
rect -8436 571018 -8254 571254
rect -8018 571018 29786 571254
rect 30022 571018 65786 571254
rect 66022 571018 101786 571254
rect 102022 571018 137786 571254
rect 138022 571018 173786 571254
rect 174022 571018 209786 571254
rect 210022 571018 245786 571254
rect 246022 571018 281786 571254
rect 282022 571018 317786 571254
rect 318022 571018 353786 571254
rect 354022 571018 389786 571254
rect 390022 571018 425786 571254
rect 426022 571018 461786 571254
rect 462022 571018 497786 571254
rect 498022 571018 533786 571254
rect 534022 571018 569786 571254
rect 570022 571018 591942 571254
rect 592178 571018 592360 571254
rect -8436 570934 592360 571018
rect -8436 570698 -8254 570934
rect -8018 570698 29786 570934
rect 30022 570698 65786 570934
rect 66022 570698 101786 570934
rect 102022 570698 137786 570934
rect 138022 570698 173786 570934
rect 174022 570698 209786 570934
rect 210022 570698 245786 570934
rect 246022 570698 281786 570934
rect 282022 570698 317786 570934
rect 318022 570698 353786 570934
rect 354022 570698 389786 570934
rect 390022 570698 425786 570934
rect 426022 570698 461786 570934
rect 462022 570698 497786 570934
rect 498022 570698 533786 570934
rect 534022 570698 569786 570934
rect 570022 570698 591942 570934
rect 592178 570698 592360 570934
rect -8436 570676 592360 570698
rect -8436 570674 -7836 570676
rect 29604 570674 30204 570676
rect 65604 570674 66204 570676
rect 101604 570674 102204 570676
rect 137604 570674 138204 570676
rect 173604 570674 174204 570676
rect 209604 570674 210204 570676
rect 245604 570674 246204 570676
rect 281604 570674 282204 570676
rect 317604 570674 318204 570676
rect 353604 570674 354204 570676
rect 389604 570674 390204 570676
rect 425604 570674 426204 570676
rect 461604 570674 462204 570676
rect 497604 570674 498204 570676
rect 533604 570674 534204 570676
rect 569604 570674 570204 570676
rect 591760 570674 592360 570676
rect -6596 567676 -5996 567678
rect 26004 567676 26604 567678
rect 62004 567676 62604 567678
rect 98004 567676 98604 567678
rect 134004 567676 134604 567678
rect 170004 567676 170604 567678
rect 206004 567676 206604 567678
rect 242004 567676 242604 567678
rect 278004 567676 278604 567678
rect 314004 567676 314604 567678
rect 350004 567676 350604 567678
rect 386004 567676 386604 567678
rect 422004 567676 422604 567678
rect 458004 567676 458604 567678
rect 494004 567676 494604 567678
rect 530004 567676 530604 567678
rect 566004 567676 566604 567678
rect 589920 567676 590520 567678
rect -6596 567654 590520 567676
rect -6596 567418 -6414 567654
rect -6178 567418 26186 567654
rect 26422 567418 62186 567654
rect 62422 567418 98186 567654
rect 98422 567418 134186 567654
rect 134422 567418 170186 567654
rect 170422 567418 206186 567654
rect 206422 567418 242186 567654
rect 242422 567418 278186 567654
rect 278422 567418 314186 567654
rect 314422 567418 350186 567654
rect 350422 567418 386186 567654
rect 386422 567418 422186 567654
rect 422422 567418 458186 567654
rect 458422 567418 494186 567654
rect 494422 567418 530186 567654
rect 530422 567418 566186 567654
rect 566422 567418 590102 567654
rect 590338 567418 590520 567654
rect -6596 567334 590520 567418
rect -6596 567098 -6414 567334
rect -6178 567098 26186 567334
rect 26422 567098 62186 567334
rect 62422 567098 98186 567334
rect 98422 567098 134186 567334
rect 134422 567098 170186 567334
rect 170422 567098 206186 567334
rect 206422 567098 242186 567334
rect 242422 567098 278186 567334
rect 278422 567098 314186 567334
rect 314422 567098 350186 567334
rect 350422 567098 386186 567334
rect 386422 567098 422186 567334
rect 422422 567098 458186 567334
rect 458422 567098 494186 567334
rect 494422 567098 530186 567334
rect 530422 567098 566186 567334
rect 566422 567098 590102 567334
rect 590338 567098 590520 567334
rect -6596 567076 590520 567098
rect -6596 567074 -5996 567076
rect 26004 567074 26604 567076
rect 62004 567074 62604 567076
rect 98004 567074 98604 567076
rect 134004 567074 134604 567076
rect 170004 567074 170604 567076
rect 206004 567074 206604 567076
rect 242004 567074 242604 567076
rect 278004 567074 278604 567076
rect 314004 567074 314604 567076
rect 350004 567074 350604 567076
rect 386004 567074 386604 567076
rect 422004 567074 422604 567076
rect 458004 567074 458604 567076
rect 494004 567074 494604 567076
rect 530004 567074 530604 567076
rect 566004 567074 566604 567076
rect 589920 567074 590520 567076
rect -4756 564076 -4156 564078
rect 22404 564076 23004 564078
rect 58404 564076 59004 564078
rect 94404 564076 95004 564078
rect 130404 564076 131004 564078
rect 166404 564076 167004 564078
rect 202404 564076 203004 564078
rect 238404 564076 239004 564078
rect 274404 564076 275004 564078
rect 310404 564076 311004 564078
rect 346404 564076 347004 564078
rect 382404 564076 383004 564078
rect 418404 564076 419004 564078
rect 454404 564076 455004 564078
rect 490404 564076 491004 564078
rect 526404 564076 527004 564078
rect 562404 564076 563004 564078
rect 588080 564076 588680 564078
rect -4756 564054 588680 564076
rect -4756 563818 -4574 564054
rect -4338 563818 22586 564054
rect 22822 563818 58586 564054
rect 58822 563818 94586 564054
rect 94822 563818 130586 564054
rect 130822 563818 166586 564054
rect 166822 563818 202586 564054
rect 202822 563818 238586 564054
rect 238822 563818 274586 564054
rect 274822 563818 310586 564054
rect 310822 563818 346586 564054
rect 346822 563818 382586 564054
rect 382822 563818 418586 564054
rect 418822 563818 454586 564054
rect 454822 563818 490586 564054
rect 490822 563818 526586 564054
rect 526822 563818 562586 564054
rect 562822 563818 588262 564054
rect 588498 563818 588680 564054
rect -4756 563734 588680 563818
rect -4756 563498 -4574 563734
rect -4338 563498 22586 563734
rect 22822 563498 58586 563734
rect 58822 563498 94586 563734
rect 94822 563498 130586 563734
rect 130822 563498 166586 563734
rect 166822 563498 202586 563734
rect 202822 563498 238586 563734
rect 238822 563498 274586 563734
rect 274822 563498 310586 563734
rect 310822 563498 346586 563734
rect 346822 563498 382586 563734
rect 382822 563498 418586 563734
rect 418822 563498 454586 563734
rect 454822 563498 490586 563734
rect 490822 563498 526586 563734
rect 526822 563498 562586 563734
rect 562822 563498 588262 563734
rect 588498 563498 588680 563734
rect -4756 563476 588680 563498
rect -4756 563474 -4156 563476
rect 22404 563474 23004 563476
rect 58404 563474 59004 563476
rect 94404 563474 95004 563476
rect 130404 563474 131004 563476
rect 166404 563474 167004 563476
rect 202404 563474 203004 563476
rect 238404 563474 239004 563476
rect 274404 563474 275004 563476
rect 310404 563474 311004 563476
rect 346404 563474 347004 563476
rect 382404 563474 383004 563476
rect 418404 563474 419004 563476
rect 454404 563474 455004 563476
rect 490404 563474 491004 563476
rect 526404 563474 527004 563476
rect 562404 563474 563004 563476
rect 588080 563474 588680 563476
rect -2916 560476 -2316 560478
rect 18804 560476 19404 560478
rect 54804 560476 55404 560478
rect 90804 560476 91404 560478
rect 126804 560476 127404 560478
rect 162804 560476 163404 560478
rect 198804 560476 199404 560478
rect 234804 560476 235404 560478
rect 270804 560476 271404 560478
rect 306804 560476 307404 560478
rect 342804 560476 343404 560478
rect 378804 560476 379404 560478
rect 414804 560476 415404 560478
rect 450804 560476 451404 560478
rect 486804 560476 487404 560478
rect 522804 560476 523404 560478
rect 558804 560476 559404 560478
rect 586240 560476 586840 560478
rect -2916 560454 586840 560476
rect -2916 560218 -2734 560454
rect -2498 560218 18986 560454
rect 19222 560218 54986 560454
rect 55222 560218 90986 560454
rect 91222 560218 126986 560454
rect 127222 560218 162986 560454
rect 163222 560218 198986 560454
rect 199222 560218 234986 560454
rect 235222 560218 270986 560454
rect 271222 560218 306986 560454
rect 307222 560218 342986 560454
rect 343222 560218 378986 560454
rect 379222 560218 414986 560454
rect 415222 560218 450986 560454
rect 451222 560218 486986 560454
rect 487222 560218 522986 560454
rect 523222 560218 558986 560454
rect 559222 560218 586422 560454
rect 586658 560218 586840 560454
rect -2916 560134 586840 560218
rect -2916 559898 -2734 560134
rect -2498 559898 18986 560134
rect 19222 559898 54986 560134
rect 55222 559898 90986 560134
rect 91222 559898 126986 560134
rect 127222 559898 162986 560134
rect 163222 559898 198986 560134
rect 199222 559898 234986 560134
rect 235222 559898 270986 560134
rect 271222 559898 306986 560134
rect 307222 559898 342986 560134
rect 343222 559898 378986 560134
rect 379222 559898 414986 560134
rect 415222 559898 450986 560134
rect 451222 559898 486986 560134
rect 487222 559898 522986 560134
rect 523222 559898 558986 560134
rect 559222 559898 586422 560134
rect 586658 559898 586840 560134
rect -2916 559876 586840 559898
rect -2916 559874 -2316 559876
rect 18804 559874 19404 559876
rect 54804 559874 55404 559876
rect 90804 559874 91404 559876
rect 126804 559874 127404 559876
rect 162804 559874 163404 559876
rect 198804 559874 199404 559876
rect 234804 559874 235404 559876
rect 270804 559874 271404 559876
rect 306804 559874 307404 559876
rect 342804 559874 343404 559876
rect 378804 559874 379404 559876
rect 414804 559874 415404 559876
rect 450804 559874 451404 559876
rect 486804 559874 487404 559876
rect 522804 559874 523404 559876
rect 558804 559874 559404 559876
rect 586240 559874 586840 559876
rect -7516 553276 -6916 553278
rect 11604 553276 12204 553278
rect 47604 553276 48204 553278
rect 83604 553276 84204 553278
rect 119604 553276 120204 553278
rect 155604 553276 156204 553278
rect 191604 553276 192204 553278
rect 227604 553276 228204 553278
rect 263604 553276 264204 553278
rect 299604 553276 300204 553278
rect 335604 553276 336204 553278
rect 371604 553276 372204 553278
rect 407604 553276 408204 553278
rect 443604 553276 444204 553278
rect 479604 553276 480204 553278
rect 515604 553276 516204 553278
rect 551604 553276 552204 553278
rect 590840 553276 591440 553278
rect -8436 553254 592360 553276
rect -8436 553018 -7334 553254
rect -7098 553018 11786 553254
rect 12022 553018 47786 553254
rect 48022 553018 83786 553254
rect 84022 553018 119786 553254
rect 120022 553018 155786 553254
rect 156022 553018 191786 553254
rect 192022 553018 227786 553254
rect 228022 553018 263786 553254
rect 264022 553018 299786 553254
rect 300022 553018 335786 553254
rect 336022 553018 371786 553254
rect 372022 553018 407786 553254
rect 408022 553018 443786 553254
rect 444022 553018 479786 553254
rect 480022 553018 515786 553254
rect 516022 553018 551786 553254
rect 552022 553018 591022 553254
rect 591258 553018 592360 553254
rect -8436 552934 592360 553018
rect -8436 552698 -7334 552934
rect -7098 552698 11786 552934
rect 12022 552698 47786 552934
rect 48022 552698 83786 552934
rect 84022 552698 119786 552934
rect 120022 552698 155786 552934
rect 156022 552698 191786 552934
rect 192022 552698 227786 552934
rect 228022 552698 263786 552934
rect 264022 552698 299786 552934
rect 300022 552698 335786 552934
rect 336022 552698 371786 552934
rect 372022 552698 407786 552934
rect 408022 552698 443786 552934
rect 444022 552698 479786 552934
rect 480022 552698 515786 552934
rect 516022 552698 551786 552934
rect 552022 552698 591022 552934
rect 591258 552698 592360 552934
rect -8436 552676 592360 552698
rect -7516 552674 -6916 552676
rect 11604 552674 12204 552676
rect 47604 552674 48204 552676
rect 83604 552674 84204 552676
rect 119604 552674 120204 552676
rect 155604 552674 156204 552676
rect 191604 552674 192204 552676
rect 227604 552674 228204 552676
rect 263604 552674 264204 552676
rect 299604 552674 300204 552676
rect 335604 552674 336204 552676
rect 371604 552674 372204 552676
rect 407604 552674 408204 552676
rect 443604 552674 444204 552676
rect 479604 552674 480204 552676
rect 515604 552674 516204 552676
rect 551604 552674 552204 552676
rect 590840 552674 591440 552676
rect -5676 549676 -5076 549678
rect 8004 549676 8604 549678
rect 44004 549676 44604 549678
rect 80004 549676 80604 549678
rect 116004 549676 116604 549678
rect 152004 549676 152604 549678
rect 188004 549676 188604 549678
rect 224004 549676 224604 549678
rect 260004 549676 260604 549678
rect 296004 549676 296604 549678
rect 332004 549676 332604 549678
rect 368004 549676 368604 549678
rect 404004 549676 404604 549678
rect 440004 549676 440604 549678
rect 476004 549676 476604 549678
rect 512004 549676 512604 549678
rect 548004 549676 548604 549678
rect 589000 549676 589600 549678
rect -6596 549654 590520 549676
rect -6596 549418 -5494 549654
rect -5258 549418 8186 549654
rect 8422 549418 44186 549654
rect 44422 549418 80186 549654
rect 80422 549418 116186 549654
rect 116422 549418 152186 549654
rect 152422 549418 188186 549654
rect 188422 549418 224186 549654
rect 224422 549418 260186 549654
rect 260422 549418 296186 549654
rect 296422 549418 332186 549654
rect 332422 549418 368186 549654
rect 368422 549418 404186 549654
rect 404422 549418 440186 549654
rect 440422 549418 476186 549654
rect 476422 549418 512186 549654
rect 512422 549418 548186 549654
rect 548422 549418 589182 549654
rect 589418 549418 590520 549654
rect -6596 549334 590520 549418
rect -6596 549098 -5494 549334
rect -5258 549098 8186 549334
rect 8422 549098 44186 549334
rect 44422 549098 80186 549334
rect 80422 549098 116186 549334
rect 116422 549098 152186 549334
rect 152422 549098 188186 549334
rect 188422 549098 224186 549334
rect 224422 549098 260186 549334
rect 260422 549098 296186 549334
rect 296422 549098 332186 549334
rect 332422 549098 368186 549334
rect 368422 549098 404186 549334
rect 404422 549098 440186 549334
rect 440422 549098 476186 549334
rect 476422 549098 512186 549334
rect 512422 549098 548186 549334
rect 548422 549098 589182 549334
rect 589418 549098 590520 549334
rect -6596 549076 590520 549098
rect -5676 549074 -5076 549076
rect 8004 549074 8604 549076
rect 44004 549074 44604 549076
rect 80004 549074 80604 549076
rect 116004 549074 116604 549076
rect 152004 549074 152604 549076
rect 188004 549074 188604 549076
rect 224004 549074 224604 549076
rect 260004 549074 260604 549076
rect 296004 549074 296604 549076
rect 332004 549074 332604 549076
rect 368004 549074 368604 549076
rect 404004 549074 404604 549076
rect 440004 549074 440604 549076
rect 476004 549074 476604 549076
rect 512004 549074 512604 549076
rect 548004 549074 548604 549076
rect 589000 549074 589600 549076
rect -3836 546076 -3236 546078
rect 4404 546076 5004 546078
rect 40404 546076 41004 546078
rect 76404 546076 77004 546078
rect 112404 546076 113004 546078
rect 148404 546076 149004 546078
rect 184404 546076 185004 546078
rect 220404 546076 221004 546078
rect 256404 546076 257004 546078
rect 292404 546076 293004 546078
rect 328404 546076 329004 546078
rect 364404 546076 365004 546078
rect 400404 546076 401004 546078
rect 436404 546076 437004 546078
rect 472404 546076 473004 546078
rect 508404 546076 509004 546078
rect 544404 546076 545004 546078
rect 580404 546076 581004 546078
rect 587160 546076 587760 546078
rect -4756 546054 588680 546076
rect -4756 545818 -3654 546054
rect -3418 545818 4586 546054
rect 4822 545818 40586 546054
rect 40822 545818 76586 546054
rect 76822 545818 112586 546054
rect 112822 545818 148586 546054
rect 148822 545818 184586 546054
rect 184822 545818 220586 546054
rect 220822 545818 256586 546054
rect 256822 545818 292586 546054
rect 292822 545818 328586 546054
rect 328822 545818 364586 546054
rect 364822 545818 400586 546054
rect 400822 545818 436586 546054
rect 436822 545818 472586 546054
rect 472822 545818 508586 546054
rect 508822 545818 544586 546054
rect 544822 545818 580586 546054
rect 580822 545818 587342 546054
rect 587578 545818 588680 546054
rect -4756 545734 588680 545818
rect -4756 545498 -3654 545734
rect -3418 545498 4586 545734
rect 4822 545498 40586 545734
rect 40822 545498 76586 545734
rect 76822 545498 112586 545734
rect 112822 545498 148586 545734
rect 148822 545498 184586 545734
rect 184822 545498 220586 545734
rect 220822 545498 256586 545734
rect 256822 545498 292586 545734
rect 292822 545498 328586 545734
rect 328822 545498 364586 545734
rect 364822 545498 400586 545734
rect 400822 545498 436586 545734
rect 436822 545498 472586 545734
rect 472822 545498 508586 545734
rect 508822 545498 544586 545734
rect 544822 545498 580586 545734
rect 580822 545498 587342 545734
rect 587578 545498 588680 545734
rect -4756 545476 588680 545498
rect -3836 545474 -3236 545476
rect 4404 545474 5004 545476
rect 40404 545474 41004 545476
rect 76404 545474 77004 545476
rect 112404 545474 113004 545476
rect 148404 545474 149004 545476
rect 184404 545474 185004 545476
rect 220404 545474 221004 545476
rect 256404 545474 257004 545476
rect 292404 545474 293004 545476
rect 328404 545474 329004 545476
rect 364404 545474 365004 545476
rect 400404 545474 401004 545476
rect 436404 545474 437004 545476
rect 472404 545474 473004 545476
rect 508404 545474 509004 545476
rect 544404 545474 545004 545476
rect 580404 545474 581004 545476
rect 587160 545474 587760 545476
rect -1996 542476 -1396 542478
rect 804 542476 1404 542478
rect 36804 542476 37404 542478
rect 72804 542476 73404 542478
rect 108804 542476 109404 542478
rect 144804 542476 145404 542478
rect 180804 542476 181404 542478
rect 216804 542476 217404 542478
rect 252804 542476 253404 542478
rect 288804 542476 289404 542478
rect 324804 542476 325404 542478
rect 360804 542476 361404 542478
rect 396804 542476 397404 542478
rect 432804 542476 433404 542478
rect 468804 542476 469404 542478
rect 504804 542476 505404 542478
rect 540804 542476 541404 542478
rect 576804 542476 577404 542478
rect 585320 542476 585920 542478
rect -2916 542454 586840 542476
rect -2916 542218 -1814 542454
rect -1578 542218 986 542454
rect 1222 542218 36986 542454
rect 37222 542218 72986 542454
rect 73222 542218 108986 542454
rect 109222 542218 144986 542454
rect 145222 542218 180986 542454
rect 181222 542218 216986 542454
rect 217222 542218 252986 542454
rect 253222 542218 288986 542454
rect 289222 542218 324986 542454
rect 325222 542218 360986 542454
rect 361222 542218 396986 542454
rect 397222 542218 432986 542454
rect 433222 542218 468986 542454
rect 469222 542218 504986 542454
rect 505222 542218 540986 542454
rect 541222 542218 576986 542454
rect 577222 542218 585502 542454
rect 585738 542218 586840 542454
rect -2916 542134 586840 542218
rect -2916 541898 -1814 542134
rect -1578 541898 986 542134
rect 1222 541898 36986 542134
rect 37222 541898 72986 542134
rect 73222 541898 108986 542134
rect 109222 541898 144986 542134
rect 145222 541898 180986 542134
rect 181222 541898 216986 542134
rect 217222 541898 252986 542134
rect 253222 541898 288986 542134
rect 289222 541898 324986 542134
rect 325222 541898 360986 542134
rect 361222 541898 396986 542134
rect 397222 541898 432986 542134
rect 433222 541898 468986 542134
rect 469222 541898 504986 542134
rect 505222 541898 540986 542134
rect 541222 541898 576986 542134
rect 577222 541898 585502 542134
rect 585738 541898 586840 542134
rect -2916 541876 586840 541898
rect -1996 541874 -1396 541876
rect 804 541874 1404 541876
rect 36804 541874 37404 541876
rect 72804 541874 73404 541876
rect 108804 541874 109404 541876
rect 144804 541874 145404 541876
rect 180804 541874 181404 541876
rect 216804 541874 217404 541876
rect 252804 541874 253404 541876
rect 288804 541874 289404 541876
rect 324804 541874 325404 541876
rect 360804 541874 361404 541876
rect 396804 541874 397404 541876
rect 432804 541874 433404 541876
rect 468804 541874 469404 541876
rect 504804 541874 505404 541876
rect 540804 541874 541404 541876
rect 576804 541874 577404 541876
rect 585320 541874 585920 541876
rect -8436 535276 -7836 535278
rect 29604 535276 30204 535278
rect 65604 535276 66204 535278
rect 101604 535276 102204 535278
rect 137604 535276 138204 535278
rect 173604 535276 174204 535278
rect 209604 535276 210204 535278
rect 245604 535276 246204 535278
rect 281604 535276 282204 535278
rect 317604 535276 318204 535278
rect 353604 535276 354204 535278
rect 389604 535276 390204 535278
rect 425604 535276 426204 535278
rect 461604 535276 462204 535278
rect 497604 535276 498204 535278
rect 533604 535276 534204 535278
rect 569604 535276 570204 535278
rect 591760 535276 592360 535278
rect -8436 535254 592360 535276
rect -8436 535018 -8254 535254
rect -8018 535018 29786 535254
rect 30022 535018 65786 535254
rect 66022 535018 101786 535254
rect 102022 535018 137786 535254
rect 138022 535018 173786 535254
rect 174022 535018 209786 535254
rect 210022 535018 245786 535254
rect 246022 535018 281786 535254
rect 282022 535018 317786 535254
rect 318022 535018 353786 535254
rect 354022 535018 389786 535254
rect 390022 535018 425786 535254
rect 426022 535018 461786 535254
rect 462022 535018 497786 535254
rect 498022 535018 533786 535254
rect 534022 535018 569786 535254
rect 570022 535018 591942 535254
rect 592178 535018 592360 535254
rect -8436 534934 592360 535018
rect -8436 534698 -8254 534934
rect -8018 534698 29786 534934
rect 30022 534698 65786 534934
rect 66022 534698 101786 534934
rect 102022 534698 137786 534934
rect 138022 534698 173786 534934
rect 174022 534698 209786 534934
rect 210022 534698 245786 534934
rect 246022 534698 281786 534934
rect 282022 534698 317786 534934
rect 318022 534698 353786 534934
rect 354022 534698 389786 534934
rect 390022 534698 425786 534934
rect 426022 534698 461786 534934
rect 462022 534698 497786 534934
rect 498022 534698 533786 534934
rect 534022 534698 569786 534934
rect 570022 534698 591942 534934
rect 592178 534698 592360 534934
rect -8436 534676 592360 534698
rect -8436 534674 -7836 534676
rect 29604 534674 30204 534676
rect 65604 534674 66204 534676
rect 101604 534674 102204 534676
rect 137604 534674 138204 534676
rect 173604 534674 174204 534676
rect 209604 534674 210204 534676
rect 245604 534674 246204 534676
rect 281604 534674 282204 534676
rect 317604 534674 318204 534676
rect 353604 534674 354204 534676
rect 389604 534674 390204 534676
rect 425604 534674 426204 534676
rect 461604 534674 462204 534676
rect 497604 534674 498204 534676
rect 533604 534674 534204 534676
rect 569604 534674 570204 534676
rect 591760 534674 592360 534676
rect -6596 531676 -5996 531678
rect 26004 531676 26604 531678
rect 62004 531676 62604 531678
rect 98004 531676 98604 531678
rect 134004 531676 134604 531678
rect 170004 531676 170604 531678
rect 206004 531676 206604 531678
rect 242004 531676 242604 531678
rect 278004 531676 278604 531678
rect 314004 531676 314604 531678
rect 350004 531676 350604 531678
rect 386004 531676 386604 531678
rect 422004 531676 422604 531678
rect 458004 531676 458604 531678
rect 494004 531676 494604 531678
rect 530004 531676 530604 531678
rect 566004 531676 566604 531678
rect 589920 531676 590520 531678
rect -6596 531654 590520 531676
rect -6596 531418 -6414 531654
rect -6178 531418 26186 531654
rect 26422 531418 62186 531654
rect 62422 531418 98186 531654
rect 98422 531418 134186 531654
rect 134422 531418 170186 531654
rect 170422 531418 206186 531654
rect 206422 531418 242186 531654
rect 242422 531418 278186 531654
rect 278422 531418 314186 531654
rect 314422 531418 350186 531654
rect 350422 531418 386186 531654
rect 386422 531418 422186 531654
rect 422422 531418 458186 531654
rect 458422 531418 494186 531654
rect 494422 531418 530186 531654
rect 530422 531418 566186 531654
rect 566422 531418 590102 531654
rect 590338 531418 590520 531654
rect -6596 531334 590520 531418
rect -6596 531098 -6414 531334
rect -6178 531098 26186 531334
rect 26422 531098 62186 531334
rect 62422 531098 98186 531334
rect 98422 531098 134186 531334
rect 134422 531098 170186 531334
rect 170422 531098 206186 531334
rect 206422 531098 242186 531334
rect 242422 531098 278186 531334
rect 278422 531098 314186 531334
rect 314422 531098 350186 531334
rect 350422 531098 386186 531334
rect 386422 531098 422186 531334
rect 422422 531098 458186 531334
rect 458422 531098 494186 531334
rect 494422 531098 530186 531334
rect 530422 531098 566186 531334
rect 566422 531098 590102 531334
rect 590338 531098 590520 531334
rect -6596 531076 590520 531098
rect -6596 531074 -5996 531076
rect 26004 531074 26604 531076
rect 62004 531074 62604 531076
rect 98004 531074 98604 531076
rect 134004 531074 134604 531076
rect 170004 531074 170604 531076
rect 206004 531074 206604 531076
rect 242004 531074 242604 531076
rect 278004 531074 278604 531076
rect 314004 531074 314604 531076
rect 350004 531074 350604 531076
rect 386004 531074 386604 531076
rect 422004 531074 422604 531076
rect 458004 531074 458604 531076
rect 494004 531074 494604 531076
rect 530004 531074 530604 531076
rect 566004 531074 566604 531076
rect 589920 531074 590520 531076
rect -4756 528076 -4156 528078
rect 22404 528076 23004 528078
rect 58404 528076 59004 528078
rect 94404 528076 95004 528078
rect 130404 528076 131004 528078
rect 166404 528076 167004 528078
rect 202404 528076 203004 528078
rect 238404 528076 239004 528078
rect 274404 528076 275004 528078
rect 310404 528076 311004 528078
rect 346404 528076 347004 528078
rect 382404 528076 383004 528078
rect 418404 528076 419004 528078
rect 454404 528076 455004 528078
rect 490404 528076 491004 528078
rect 526404 528076 527004 528078
rect 562404 528076 563004 528078
rect 588080 528076 588680 528078
rect -4756 528054 588680 528076
rect -4756 527818 -4574 528054
rect -4338 527818 22586 528054
rect 22822 527818 58586 528054
rect 58822 527818 94586 528054
rect 94822 527818 130586 528054
rect 130822 527818 166586 528054
rect 166822 527818 202586 528054
rect 202822 527818 238586 528054
rect 238822 527818 274586 528054
rect 274822 527818 310586 528054
rect 310822 527818 346586 528054
rect 346822 527818 382586 528054
rect 382822 527818 418586 528054
rect 418822 527818 454586 528054
rect 454822 527818 490586 528054
rect 490822 527818 526586 528054
rect 526822 527818 562586 528054
rect 562822 527818 588262 528054
rect 588498 527818 588680 528054
rect -4756 527734 588680 527818
rect -4756 527498 -4574 527734
rect -4338 527498 22586 527734
rect 22822 527498 58586 527734
rect 58822 527498 94586 527734
rect 94822 527498 130586 527734
rect 130822 527498 166586 527734
rect 166822 527498 202586 527734
rect 202822 527498 238586 527734
rect 238822 527498 274586 527734
rect 274822 527498 310586 527734
rect 310822 527498 346586 527734
rect 346822 527498 382586 527734
rect 382822 527498 418586 527734
rect 418822 527498 454586 527734
rect 454822 527498 490586 527734
rect 490822 527498 526586 527734
rect 526822 527498 562586 527734
rect 562822 527498 588262 527734
rect 588498 527498 588680 527734
rect -4756 527476 588680 527498
rect -4756 527474 -4156 527476
rect 22404 527474 23004 527476
rect 58404 527474 59004 527476
rect 94404 527474 95004 527476
rect 130404 527474 131004 527476
rect 166404 527474 167004 527476
rect 202404 527474 203004 527476
rect 238404 527474 239004 527476
rect 274404 527474 275004 527476
rect 310404 527474 311004 527476
rect 346404 527474 347004 527476
rect 382404 527474 383004 527476
rect 418404 527474 419004 527476
rect 454404 527474 455004 527476
rect 490404 527474 491004 527476
rect 526404 527474 527004 527476
rect 562404 527474 563004 527476
rect 588080 527474 588680 527476
rect -2916 524476 -2316 524478
rect 18804 524476 19404 524478
rect 54804 524476 55404 524478
rect 90804 524476 91404 524478
rect 126804 524476 127404 524478
rect 162804 524476 163404 524478
rect 198804 524476 199404 524478
rect 234804 524476 235404 524478
rect 270804 524476 271404 524478
rect 306804 524476 307404 524478
rect 342804 524476 343404 524478
rect 378804 524476 379404 524478
rect 414804 524476 415404 524478
rect 450804 524476 451404 524478
rect 486804 524476 487404 524478
rect 522804 524476 523404 524478
rect 558804 524476 559404 524478
rect 586240 524476 586840 524478
rect -2916 524454 586840 524476
rect -2916 524218 -2734 524454
rect -2498 524218 18986 524454
rect 19222 524218 54986 524454
rect 55222 524218 90986 524454
rect 91222 524218 126986 524454
rect 127222 524218 162986 524454
rect 163222 524218 198986 524454
rect 199222 524218 234986 524454
rect 235222 524218 270986 524454
rect 271222 524218 306986 524454
rect 307222 524218 342986 524454
rect 343222 524218 378986 524454
rect 379222 524218 414986 524454
rect 415222 524218 450986 524454
rect 451222 524218 486986 524454
rect 487222 524218 522986 524454
rect 523222 524218 558986 524454
rect 559222 524218 586422 524454
rect 586658 524218 586840 524454
rect -2916 524134 586840 524218
rect -2916 523898 -2734 524134
rect -2498 523898 18986 524134
rect 19222 523898 54986 524134
rect 55222 523898 90986 524134
rect 91222 523898 126986 524134
rect 127222 523898 162986 524134
rect 163222 523898 198986 524134
rect 199222 523898 234986 524134
rect 235222 523898 270986 524134
rect 271222 523898 306986 524134
rect 307222 523898 342986 524134
rect 343222 523898 378986 524134
rect 379222 523898 414986 524134
rect 415222 523898 450986 524134
rect 451222 523898 486986 524134
rect 487222 523898 522986 524134
rect 523222 523898 558986 524134
rect 559222 523898 586422 524134
rect 586658 523898 586840 524134
rect -2916 523876 586840 523898
rect -2916 523874 -2316 523876
rect 18804 523874 19404 523876
rect 54804 523874 55404 523876
rect 90804 523874 91404 523876
rect 126804 523874 127404 523876
rect 162804 523874 163404 523876
rect 198804 523874 199404 523876
rect 234804 523874 235404 523876
rect 270804 523874 271404 523876
rect 306804 523874 307404 523876
rect 342804 523874 343404 523876
rect 378804 523874 379404 523876
rect 414804 523874 415404 523876
rect 450804 523874 451404 523876
rect 486804 523874 487404 523876
rect 522804 523874 523404 523876
rect 558804 523874 559404 523876
rect 586240 523874 586840 523876
rect -7516 517276 -6916 517278
rect 11604 517276 12204 517278
rect 47604 517276 48204 517278
rect 83604 517276 84204 517278
rect 119604 517276 120204 517278
rect 155604 517276 156204 517278
rect 191604 517276 192204 517278
rect 227604 517276 228204 517278
rect 263604 517276 264204 517278
rect 299604 517276 300204 517278
rect 335604 517276 336204 517278
rect 371604 517276 372204 517278
rect 407604 517276 408204 517278
rect 443604 517276 444204 517278
rect 479604 517276 480204 517278
rect 515604 517276 516204 517278
rect 551604 517276 552204 517278
rect 590840 517276 591440 517278
rect -8436 517254 592360 517276
rect -8436 517018 -7334 517254
rect -7098 517018 11786 517254
rect 12022 517018 47786 517254
rect 48022 517018 83786 517254
rect 84022 517018 119786 517254
rect 120022 517018 155786 517254
rect 156022 517018 191786 517254
rect 192022 517018 227786 517254
rect 228022 517018 263786 517254
rect 264022 517018 299786 517254
rect 300022 517018 335786 517254
rect 336022 517018 371786 517254
rect 372022 517018 407786 517254
rect 408022 517018 443786 517254
rect 444022 517018 479786 517254
rect 480022 517018 515786 517254
rect 516022 517018 551786 517254
rect 552022 517018 591022 517254
rect 591258 517018 592360 517254
rect -8436 516934 592360 517018
rect -8436 516698 -7334 516934
rect -7098 516698 11786 516934
rect 12022 516698 47786 516934
rect 48022 516698 83786 516934
rect 84022 516698 119786 516934
rect 120022 516698 155786 516934
rect 156022 516698 191786 516934
rect 192022 516698 227786 516934
rect 228022 516698 263786 516934
rect 264022 516698 299786 516934
rect 300022 516698 335786 516934
rect 336022 516698 371786 516934
rect 372022 516698 407786 516934
rect 408022 516698 443786 516934
rect 444022 516698 479786 516934
rect 480022 516698 515786 516934
rect 516022 516698 551786 516934
rect 552022 516698 591022 516934
rect 591258 516698 592360 516934
rect -8436 516676 592360 516698
rect -7516 516674 -6916 516676
rect 11604 516674 12204 516676
rect 47604 516674 48204 516676
rect 83604 516674 84204 516676
rect 119604 516674 120204 516676
rect 155604 516674 156204 516676
rect 191604 516674 192204 516676
rect 227604 516674 228204 516676
rect 263604 516674 264204 516676
rect 299604 516674 300204 516676
rect 335604 516674 336204 516676
rect 371604 516674 372204 516676
rect 407604 516674 408204 516676
rect 443604 516674 444204 516676
rect 479604 516674 480204 516676
rect 515604 516674 516204 516676
rect 551604 516674 552204 516676
rect 590840 516674 591440 516676
rect -5676 513676 -5076 513678
rect 8004 513676 8604 513678
rect 44004 513676 44604 513678
rect 80004 513676 80604 513678
rect 116004 513676 116604 513678
rect 152004 513676 152604 513678
rect 188004 513676 188604 513678
rect 224004 513676 224604 513678
rect 260004 513676 260604 513678
rect 296004 513676 296604 513678
rect 332004 513676 332604 513678
rect 368004 513676 368604 513678
rect 404004 513676 404604 513678
rect 440004 513676 440604 513678
rect 476004 513676 476604 513678
rect 512004 513676 512604 513678
rect 548004 513676 548604 513678
rect 589000 513676 589600 513678
rect -6596 513654 590520 513676
rect -6596 513418 -5494 513654
rect -5258 513418 8186 513654
rect 8422 513418 44186 513654
rect 44422 513418 80186 513654
rect 80422 513418 116186 513654
rect 116422 513418 152186 513654
rect 152422 513418 188186 513654
rect 188422 513418 224186 513654
rect 224422 513418 260186 513654
rect 260422 513418 296186 513654
rect 296422 513418 332186 513654
rect 332422 513418 368186 513654
rect 368422 513418 404186 513654
rect 404422 513418 440186 513654
rect 440422 513418 476186 513654
rect 476422 513418 512186 513654
rect 512422 513418 548186 513654
rect 548422 513418 589182 513654
rect 589418 513418 590520 513654
rect -6596 513334 590520 513418
rect -6596 513098 -5494 513334
rect -5258 513098 8186 513334
rect 8422 513098 44186 513334
rect 44422 513098 80186 513334
rect 80422 513098 116186 513334
rect 116422 513098 152186 513334
rect 152422 513098 188186 513334
rect 188422 513098 224186 513334
rect 224422 513098 260186 513334
rect 260422 513098 296186 513334
rect 296422 513098 332186 513334
rect 332422 513098 368186 513334
rect 368422 513098 404186 513334
rect 404422 513098 440186 513334
rect 440422 513098 476186 513334
rect 476422 513098 512186 513334
rect 512422 513098 548186 513334
rect 548422 513098 589182 513334
rect 589418 513098 590520 513334
rect -6596 513076 590520 513098
rect -5676 513074 -5076 513076
rect 8004 513074 8604 513076
rect 44004 513074 44604 513076
rect 80004 513074 80604 513076
rect 116004 513074 116604 513076
rect 152004 513074 152604 513076
rect 188004 513074 188604 513076
rect 224004 513074 224604 513076
rect 260004 513074 260604 513076
rect 296004 513074 296604 513076
rect 332004 513074 332604 513076
rect 368004 513074 368604 513076
rect 404004 513074 404604 513076
rect 440004 513074 440604 513076
rect 476004 513074 476604 513076
rect 512004 513074 512604 513076
rect 548004 513074 548604 513076
rect 589000 513074 589600 513076
rect -3836 510076 -3236 510078
rect 4404 510076 5004 510078
rect 40404 510076 41004 510078
rect 76404 510076 77004 510078
rect 112404 510076 113004 510078
rect 148404 510076 149004 510078
rect 184404 510076 185004 510078
rect 220404 510076 221004 510078
rect 256404 510076 257004 510078
rect 292404 510076 293004 510078
rect 328404 510076 329004 510078
rect 364404 510076 365004 510078
rect 400404 510076 401004 510078
rect 436404 510076 437004 510078
rect 472404 510076 473004 510078
rect 508404 510076 509004 510078
rect 544404 510076 545004 510078
rect 580404 510076 581004 510078
rect 587160 510076 587760 510078
rect -4756 510054 588680 510076
rect -4756 509818 -3654 510054
rect -3418 509818 4586 510054
rect 4822 509818 40586 510054
rect 40822 509818 76586 510054
rect 76822 509818 112586 510054
rect 112822 509818 148586 510054
rect 148822 509818 184586 510054
rect 184822 509818 220586 510054
rect 220822 509818 256586 510054
rect 256822 509818 292586 510054
rect 292822 509818 328586 510054
rect 328822 509818 364586 510054
rect 364822 509818 400586 510054
rect 400822 509818 436586 510054
rect 436822 509818 472586 510054
rect 472822 509818 508586 510054
rect 508822 509818 544586 510054
rect 544822 509818 580586 510054
rect 580822 509818 587342 510054
rect 587578 509818 588680 510054
rect -4756 509734 588680 509818
rect -4756 509498 -3654 509734
rect -3418 509498 4586 509734
rect 4822 509498 40586 509734
rect 40822 509498 76586 509734
rect 76822 509498 112586 509734
rect 112822 509498 148586 509734
rect 148822 509498 184586 509734
rect 184822 509498 220586 509734
rect 220822 509498 256586 509734
rect 256822 509498 292586 509734
rect 292822 509498 328586 509734
rect 328822 509498 364586 509734
rect 364822 509498 400586 509734
rect 400822 509498 436586 509734
rect 436822 509498 472586 509734
rect 472822 509498 508586 509734
rect 508822 509498 544586 509734
rect 544822 509498 580586 509734
rect 580822 509498 587342 509734
rect 587578 509498 588680 509734
rect -4756 509476 588680 509498
rect -3836 509474 -3236 509476
rect 4404 509474 5004 509476
rect 40404 509474 41004 509476
rect 76404 509474 77004 509476
rect 112404 509474 113004 509476
rect 148404 509474 149004 509476
rect 184404 509474 185004 509476
rect 220404 509474 221004 509476
rect 256404 509474 257004 509476
rect 292404 509474 293004 509476
rect 328404 509474 329004 509476
rect 364404 509474 365004 509476
rect 400404 509474 401004 509476
rect 436404 509474 437004 509476
rect 472404 509474 473004 509476
rect 508404 509474 509004 509476
rect 544404 509474 545004 509476
rect 580404 509474 581004 509476
rect 587160 509474 587760 509476
rect -1996 506476 -1396 506478
rect 804 506476 1404 506478
rect 36804 506476 37404 506478
rect 72804 506476 73404 506478
rect 108804 506476 109404 506478
rect 144804 506476 145404 506478
rect 180804 506476 181404 506478
rect 216804 506476 217404 506478
rect 252804 506476 253404 506478
rect 288804 506476 289404 506478
rect 324804 506476 325404 506478
rect 360804 506476 361404 506478
rect 396804 506476 397404 506478
rect 432804 506476 433404 506478
rect 468804 506476 469404 506478
rect 504804 506476 505404 506478
rect 540804 506476 541404 506478
rect 576804 506476 577404 506478
rect 585320 506476 585920 506478
rect -2916 506454 586840 506476
rect -2916 506218 -1814 506454
rect -1578 506218 986 506454
rect 1222 506218 36986 506454
rect 37222 506218 72986 506454
rect 73222 506218 108986 506454
rect 109222 506218 144986 506454
rect 145222 506218 180986 506454
rect 181222 506218 216986 506454
rect 217222 506218 252986 506454
rect 253222 506218 288986 506454
rect 289222 506218 324986 506454
rect 325222 506218 360986 506454
rect 361222 506218 396986 506454
rect 397222 506218 432986 506454
rect 433222 506218 468986 506454
rect 469222 506218 504986 506454
rect 505222 506218 540986 506454
rect 541222 506218 576986 506454
rect 577222 506218 585502 506454
rect 585738 506218 586840 506454
rect -2916 506134 586840 506218
rect -2916 505898 -1814 506134
rect -1578 505898 986 506134
rect 1222 505898 36986 506134
rect 37222 505898 72986 506134
rect 73222 505898 108986 506134
rect 109222 505898 144986 506134
rect 145222 505898 180986 506134
rect 181222 505898 216986 506134
rect 217222 505898 252986 506134
rect 253222 505898 288986 506134
rect 289222 505898 324986 506134
rect 325222 505898 360986 506134
rect 361222 505898 396986 506134
rect 397222 505898 432986 506134
rect 433222 505898 468986 506134
rect 469222 505898 504986 506134
rect 505222 505898 540986 506134
rect 541222 505898 576986 506134
rect 577222 505898 585502 506134
rect 585738 505898 586840 506134
rect -2916 505876 586840 505898
rect -1996 505874 -1396 505876
rect 804 505874 1404 505876
rect 36804 505874 37404 505876
rect 72804 505874 73404 505876
rect 108804 505874 109404 505876
rect 144804 505874 145404 505876
rect 180804 505874 181404 505876
rect 216804 505874 217404 505876
rect 252804 505874 253404 505876
rect 288804 505874 289404 505876
rect 324804 505874 325404 505876
rect 360804 505874 361404 505876
rect 396804 505874 397404 505876
rect 432804 505874 433404 505876
rect 468804 505874 469404 505876
rect 504804 505874 505404 505876
rect 540804 505874 541404 505876
rect 576804 505874 577404 505876
rect 585320 505874 585920 505876
rect -8436 499276 -7836 499278
rect 29604 499276 30204 499278
rect 65604 499276 66204 499278
rect 101604 499276 102204 499278
rect 137604 499276 138204 499278
rect 173604 499276 174204 499278
rect 209604 499276 210204 499278
rect 245604 499276 246204 499278
rect 281604 499276 282204 499278
rect 317604 499276 318204 499278
rect 353604 499276 354204 499278
rect 389604 499276 390204 499278
rect 425604 499276 426204 499278
rect 461604 499276 462204 499278
rect 497604 499276 498204 499278
rect 533604 499276 534204 499278
rect 569604 499276 570204 499278
rect 591760 499276 592360 499278
rect -8436 499254 592360 499276
rect -8436 499018 -8254 499254
rect -8018 499018 29786 499254
rect 30022 499018 65786 499254
rect 66022 499018 101786 499254
rect 102022 499018 137786 499254
rect 138022 499018 173786 499254
rect 174022 499018 209786 499254
rect 210022 499018 245786 499254
rect 246022 499018 281786 499254
rect 282022 499018 317786 499254
rect 318022 499018 353786 499254
rect 354022 499018 389786 499254
rect 390022 499018 425786 499254
rect 426022 499018 461786 499254
rect 462022 499018 497786 499254
rect 498022 499018 533786 499254
rect 534022 499018 569786 499254
rect 570022 499018 591942 499254
rect 592178 499018 592360 499254
rect -8436 498934 592360 499018
rect -8436 498698 -8254 498934
rect -8018 498698 29786 498934
rect 30022 498698 65786 498934
rect 66022 498698 101786 498934
rect 102022 498698 137786 498934
rect 138022 498698 173786 498934
rect 174022 498698 209786 498934
rect 210022 498698 245786 498934
rect 246022 498698 281786 498934
rect 282022 498698 317786 498934
rect 318022 498698 353786 498934
rect 354022 498698 389786 498934
rect 390022 498698 425786 498934
rect 426022 498698 461786 498934
rect 462022 498698 497786 498934
rect 498022 498698 533786 498934
rect 534022 498698 569786 498934
rect 570022 498698 591942 498934
rect 592178 498698 592360 498934
rect -8436 498676 592360 498698
rect -8436 498674 -7836 498676
rect 29604 498674 30204 498676
rect 65604 498674 66204 498676
rect 101604 498674 102204 498676
rect 137604 498674 138204 498676
rect 173604 498674 174204 498676
rect 209604 498674 210204 498676
rect 245604 498674 246204 498676
rect 281604 498674 282204 498676
rect 317604 498674 318204 498676
rect 353604 498674 354204 498676
rect 389604 498674 390204 498676
rect 425604 498674 426204 498676
rect 461604 498674 462204 498676
rect 497604 498674 498204 498676
rect 533604 498674 534204 498676
rect 569604 498674 570204 498676
rect 591760 498674 592360 498676
rect -6596 495676 -5996 495678
rect 26004 495676 26604 495678
rect 62004 495676 62604 495678
rect 98004 495676 98604 495678
rect 134004 495676 134604 495678
rect 170004 495676 170604 495678
rect 206004 495676 206604 495678
rect 242004 495676 242604 495678
rect 278004 495676 278604 495678
rect 314004 495676 314604 495678
rect 350004 495676 350604 495678
rect 386004 495676 386604 495678
rect 422004 495676 422604 495678
rect 458004 495676 458604 495678
rect 494004 495676 494604 495678
rect 530004 495676 530604 495678
rect 566004 495676 566604 495678
rect 589920 495676 590520 495678
rect -6596 495654 590520 495676
rect -6596 495418 -6414 495654
rect -6178 495418 26186 495654
rect 26422 495418 62186 495654
rect 62422 495418 98186 495654
rect 98422 495418 134186 495654
rect 134422 495418 170186 495654
rect 170422 495418 206186 495654
rect 206422 495418 242186 495654
rect 242422 495418 278186 495654
rect 278422 495418 314186 495654
rect 314422 495418 350186 495654
rect 350422 495418 386186 495654
rect 386422 495418 422186 495654
rect 422422 495418 458186 495654
rect 458422 495418 494186 495654
rect 494422 495418 530186 495654
rect 530422 495418 566186 495654
rect 566422 495418 590102 495654
rect 590338 495418 590520 495654
rect -6596 495334 590520 495418
rect -6596 495098 -6414 495334
rect -6178 495098 26186 495334
rect 26422 495098 62186 495334
rect 62422 495098 98186 495334
rect 98422 495098 134186 495334
rect 134422 495098 170186 495334
rect 170422 495098 206186 495334
rect 206422 495098 242186 495334
rect 242422 495098 278186 495334
rect 278422 495098 314186 495334
rect 314422 495098 350186 495334
rect 350422 495098 386186 495334
rect 386422 495098 422186 495334
rect 422422 495098 458186 495334
rect 458422 495098 494186 495334
rect 494422 495098 530186 495334
rect 530422 495098 566186 495334
rect 566422 495098 590102 495334
rect 590338 495098 590520 495334
rect -6596 495076 590520 495098
rect -6596 495074 -5996 495076
rect 26004 495074 26604 495076
rect 62004 495074 62604 495076
rect 98004 495074 98604 495076
rect 134004 495074 134604 495076
rect 170004 495074 170604 495076
rect 206004 495074 206604 495076
rect 242004 495074 242604 495076
rect 278004 495074 278604 495076
rect 314004 495074 314604 495076
rect 350004 495074 350604 495076
rect 386004 495074 386604 495076
rect 422004 495074 422604 495076
rect 458004 495074 458604 495076
rect 494004 495074 494604 495076
rect 530004 495074 530604 495076
rect 566004 495074 566604 495076
rect 589920 495074 590520 495076
rect -4756 492076 -4156 492078
rect 22404 492076 23004 492078
rect 58404 492076 59004 492078
rect 94404 492076 95004 492078
rect 130404 492076 131004 492078
rect 166404 492076 167004 492078
rect 202404 492076 203004 492078
rect 238404 492076 239004 492078
rect 274404 492076 275004 492078
rect 310404 492076 311004 492078
rect 346404 492076 347004 492078
rect 382404 492076 383004 492078
rect 418404 492076 419004 492078
rect 454404 492076 455004 492078
rect 490404 492076 491004 492078
rect 526404 492076 527004 492078
rect 562404 492076 563004 492078
rect 588080 492076 588680 492078
rect -4756 492054 588680 492076
rect -4756 491818 -4574 492054
rect -4338 491818 22586 492054
rect 22822 491818 58586 492054
rect 58822 491818 94586 492054
rect 94822 491818 130586 492054
rect 130822 491818 166586 492054
rect 166822 491818 202586 492054
rect 202822 491818 238586 492054
rect 238822 491818 274586 492054
rect 274822 491818 310586 492054
rect 310822 491818 346586 492054
rect 346822 491818 382586 492054
rect 382822 491818 418586 492054
rect 418822 491818 454586 492054
rect 454822 491818 490586 492054
rect 490822 491818 526586 492054
rect 526822 491818 562586 492054
rect 562822 491818 588262 492054
rect 588498 491818 588680 492054
rect -4756 491734 588680 491818
rect -4756 491498 -4574 491734
rect -4338 491498 22586 491734
rect 22822 491498 58586 491734
rect 58822 491498 94586 491734
rect 94822 491498 130586 491734
rect 130822 491498 166586 491734
rect 166822 491498 202586 491734
rect 202822 491498 238586 491734
rect 238822 491498 274586 491734
rect 274822 491498 310586 491734
rect 310822 491498 346586 491734
rect 346822 491498 382586 491734
rect 382822 491498 418586 491734
rect 418822 491498 454586 491734
rect 454822 491498 490586 491734
rect 490822 491498 526586 491734
rect 526822 491498 562586 491734
rect 562822 491498 588262 491734
rect 588498 491498 588680 491734
rect -4756 491476 588680 491498
rect -4756 491474 -4156 491476
rect 22404 491474 23004 491476
rect 58404 491474 59004 491476
rect 94404 491474 95004 491476
rect 130404 491474 131004 491476
rect 166404 491474 167004 491476
rect 202404 491474 203004 491476
rect 238404 491474 239004 491476
rect 274404 491474 275004 491476
rect 310404 491474 311004 491476
rect 346404 491474 347004 491476
rect 382404 491474 383004 491476
rect 418404 491474 419004 491476
rect 454404 491474 455004 491476
rect 490404 491474 491004 491476
rect 526404 491474 527004 491476
rect 562404 491474 563004 491476
rect 588080 491474 588680 491476
rect -2916 488476 -2316 488478
rect 18804 488476 19404 488478
rect 54804 488476 55404 488478
rect 90804 488476 91404 488478
rect 126804 488476 127404 488478
rect 162804 488476 163404 488478
rect 198804 488476 199404 488478
rect 234804 488476 235404 488478
rect 270804 488476 271404 488478
rect 306804 488476 307404 488478
rect 342804 488476 343404 488478
rect 378804 488476 379404 488478
rect 414804 488476 415404 488478
rect 450804 488476 451404 488478
rect 486804 488476 487404 488478
rect 522804 488476 523404 488478
rect 558804 488476 559404 488478
rect 586240 488476 586840 488478
rect -2916 488454 586840 488476
rect -2916 488218 -2734 488454
rect -2498 488218 18986 488454
rect 19222 488218 54986 488454
rect 55222 488218 90986 488454
rect 91222 488218 126986 488454
rect 127222 488218 162986 488454
rect 163222 488218 198986 488454
rect 199222 488218 234986 488454
rect 235222 488218 270986 488454
rect 271222 488218 306986 488454
rect 307222 488218 342986 488454
rect 343222 488218 378986 488454
rect 379222 488218 414986 488454
rect 415222 488218 450986 488454
rect 451222 488218 486986 488454
rect 487222 488218 522986 488454
rect 523222 488218 558986 488454
rect 559222 488218 586422 488454
rect 586658 488218 586840 488454
rect -2916 488134 586840 488218
rect -2916 487898 -2734 488134
rect -2498 487898 18986 488134
rect 19222 487898 54986 488134
rect 55222 487898 90986 488134
rect 91222 487898 126986 488134
rect 127222 487898 162986 488134
rect 163222 487898 198986 488134
rect 199222 487898 234986 488134
rect 235222 487898 270986 488134
rect 271222 487898 306986 488134
rect 307222 487898 342986 488134
rect 343222 487898 378986 488134
rect 379222 487898 414986 488134
rect 415222 487898 450986 488134
rect 451222 487898 486986 488134
rect 487222 487898 522986 488134
rect 523222 487898 558986 488134
rect 559222 487898 586422 488134
rect 586658 487898 586840 488134
rect -2916 487876 586840 487898
rect -2916 487874 -2316 487876
rect 18804 487874 19404 487876
rect 54804 487874 55404 487876
rect 90804 487874 91404 487876
rect 126804 487874 127404 487876
rect 162804 487874 163404 487876
rect 198804 487874 199404 487876
rect 234804 487874 235404 487876
rect 270804 487874 271404 487876
rect 306804 487874 307404 487876
rect 342804 487874 343404 487876
rect 378804 487874 379404 487876
rect 414804 487874 415404 487876
rect 450804 487874 451404 487876
rect 486804 487874 487404 487876
rect 522804 487874 523404 487876
rect 558804 487874 559404 487876
rect 586240 487874 586840 487876
rect -7516 481276 -6916 481278
rect 11604 481276 12204 481278
rect 47604 481276 48204 481278
rect 83604 481276 84204 481278
rect 119604 481276 120204 481278
rect 155604 481276 156204 481278
rect 191604 481276 192204 481278
rect 227604 481276 228204 481278
rect 263604 481276 264204 481278
rect 299604 481276 300204 481278
rect 335604 481276 336204 481278
rect 371604 481276 372204 481278
rect 407604 481276 408204 481278
rect 443604 481276 444204 481278
rect 479604 481276 480204 481278
rect 515604 481276 516204 481278
rect 551604 481276 552204 481278
rect 590840 481276 591440 481278
rect -8436 481254 592360 481276
rect -8436 481018 -7334 481254
rect -7098 481018 11786 481254
rect 12022 481018 47786 481254
rect 48022 481018 83786 481254
rect 84022 481018 119786 481254
rect 120022 481018 155786 481254
rect 156022 481018 191786 481254
rect 192022 481018 227786 481254
rect 228022 481018 263786 481254
rect 264022 481018 299786 481254
rect 300022 481018 335786 481254
rect 336022 481018 371786 481254
rect 372022 481018 407786 481254
rect 408022 481018 443786 481254
rect 444022 481018 479786 481254
rect 480022 481018 515786 481254
rect 516022 481018 551786 481254
rect 552022 481018 591022 481254
rect 591258 481018 592360 481254
rect -8436 480934 592360 481018
rect -8436 480698 -7334 480934
rect -7098 480698 11786 480934
rect 12022 480698 47786 480934
rect 48022 480698 83786 480934
rect 84022 480698 119786 480934
rect 120022 480698 155786 480934
rect 156022 480698 191786 480934
rect 192022 480698 227786 480934
rect 228022 480698 263786 480934
rect 264022 480698 299786 480934
rect 300022 480698 335786 480934
rect 336022 480698 371786 480934
rect 372022 480698 407786 480934
rect 408022 480698 443786 480934
rect 444022 480698 479786 480934
rect 480022 480698 515786 480934
rect 516022 480698 551786 480934
rect 552022 480698 591022 480934
rect 591258 480698 592360 480934
rect -8436 480676 592360 480698
rect -7516 480674 -6916 480676
rect 11604 480674 12204 480676
rect 47604 480674 48204 480676
rect 83604 480674 84204 480676
rect 119604 480674 120204 480676
rect 155604 480674 156204 480676
rect 191604 480674 192204 480676
rect 227604 480674 228204 480676
rect 263604 480674 264204 480676
rect 299604 480674 300204 480676
rect 335604 480674 336204 480676
rect 371604 480674 372204 480676
rect 407604 480674 408204 480676
rect 443604 480674 444204 480676
rect 479604 480674 480204 480676
rect 515604 480674 516204 480676
rect 551604 480674 552204 480676
rect 590840 480674 591440 480676
rect -5676 477676 -5076 477678
rect 8004 477676 8604 477678
rect 44004 477676 44604 477678
rect 80004 477676 80604 477678
rect 116004 477676 116604 477678
rect 152004 477676 152604 477678
rect 188004 477676 188604 477678
rect 224004 477676 224604 477678
rect 260004 477676 260604 477678
rect 296004 477676 296604 477678
rect 332004 477676 332604 477678
rect 368004 477676 368604 477678
rect 404004 477676 404604 477678
rect 440004 477676 440604 477678
rect 476004 477676 476604 477678
rect 512004 477676 512604 477678
rect 548004 477676 548604 477678
rect 589000 477676 589600 477678
rect -6596 477654 590520 477676
rect -6596 477418 -5494 477654
rect -5258 477418 8186 477654
rect 8422 477418 44186 477654
rect 44422 477418 80186 477654
rect 80422 477418 116186 477654
rect 116422 477418 152186 477654
rect 152422 477418 188186 477654
rect 188422 477418 224186 477654
rect 224422 477418 260186 477654
rect 260422 477418 296186 477654
rect 296422 477418 332186 477654
rect 332422 477418 368186 477654
rect 368422 477418 404186 477654
rect 404422 477418 440186 477654
rect 440422 477418 476186 477654
rect 476422 477418 512186 477654
rect 512422 477418 548186 477654
rect 548422 477418 589182 477654
rect 589418 477418 590520 477654
rect -6596 477334 590520 477418
rect -6596 477098 -5494 477334
rect -5258 477098 8186 477334
rect 8422 477098 44186 477334
rect 44422 477098 80186 477334
rect 80422 477098 116186 477334
rect 116422 477098 152186 477334
rect 152422 477098 188186 477334
rect 188422 477098 224186 477334
rect 224422 477098 260186 477334
rect 260422 477098 296186 477334
rect 296422 477098 332186 477334
rect 332422 477098 368186 477334
rect 368422 477098 404186 477334
rect 404422 477098 440186 477334
rect 440422 477098 476186 477334
rect 476422 477098 512186 477334
rect 512422 477098 548186 477334
rect 548422 477098 589182 477334
rect 589418 477098 590520 477334
rect -6596 477076 590520 477098
rect -5676 477074 -5076 477076
rect 8004 477074 8604 477076
rect 44004 477074 44604 477076
rect 80004 477074 80604 477076
rect 116004 477074 116604 477076
rect 152004 477074 152604 477076
rect 188004 477074 188604 477076
rect 224004 477074 224604 477076
rect 260004 477074 260604 477076
rect 296004 477074 296604 477076
rect 332004 477074 332604 477076
rect 368004 477074 368604 477076
rect 404004 477074 404604 477076
rect 440004 477074 440604 477076
rect 476004 477074 476604 477076
rect 512004 477074 512604 477076
rect 548004 477074 548604 477076
rect 589000 477074 589600 477076
rect -3836 474076 -3236 474078
rect 4404 474076 5004 474078
rect 40404 474076 41004 474078
rect 76404 474076 77004 474078
rect 112404 474076 113004 474078
rect 148404 474076 149004 474078
rect 184404 474076 185004 474078
rect 220404 474076 221004 474078
rect 256404 474076 257004 474078
rect 292404 474076 293004 474078
rect 328404 474076 329004 474078
rect 364404 474076 365004 474078
rect 400404 474076 401004 474078
rect 436404 474076 437004 474078
rect 472404 474076 473004 474078
rect 508404 474076 509004 474078
rect 544404 474076 545004 474078
rect 580404 474076 581004 474078
rect 587160 474076 587760 474078
rect -4756 474054 588680 474076
rect -4756 473818 -3654 474054
rect -3418 473818 4586 474054
rect 4822 473818 40586 474054
rect 40822 473818 76586 474054
rect 76822 473818 112586 474054
rect 112822 473818 148586 474054
rect 148822 473818 184586 474054
rect 184822 473818 220586 474054
rect 220822 473818 256586 474054
rect 256822 473818 292586 474054
rect 292822 473818 328586 474054
rect 328822 473818 364586 474054
rect 364822 473818 400586 474054
rect 400822 473818 436586 474054
rect 436822 473818 472586 474054
rect 472822 473818 508586 474054
rect 508822 473818 544586 474054
rect 544822 473818 580586 474054
rect 580822 473818 587342 474054
rect 587578 473818 588680 474054
rect -4756 473734 588680 473818
rect -4756 473498 -3654 473734
rect -3418 473498 4586 473734
rect 4822 473498 40586 473734
rect 40822 473498 76586 473734
rect 76822 473498 112586 473734
rect 112822 473498 148586 473734
rect 148822 473498 184586 473734
rect 184822 473498 220586 473734
rect 220822 473498 256586 473734
rect 256822 473498 292586 473734
rect 292822 473498 328586 473734
rect 328822 473498 364586 473734
rect 364822 473498 400586 473734
rect 400822 473498 436586 473734
rect 436822 473498 472586 473734
rect 472822 473498 508586 473734
rect 508822 473498 544586 473734
rect 544822 473498 580586 473734
rect 580822 473498 587342 473734
rect 587578 473498 588680 473734
rect -4756 473476 588680 473498
rect -3836 473474 -3236 473476
rect 4404 473474 5004 473476
rect 40404 473474 41004 473476
rect 76404 473474 77004 473476
rect 112404 473474 113004 473476
rect 148404 473474 149004 473476
rect 184404 473474 185004 473476
rect 220404 473474 221004 473476
rect 256404 473474 257004 473476
rect 292404 473474 293004 473476
rect 328404 473474 329004 473476
rect 364404 473474 365004 473476
rect 400404 473474 401004 473476
rect 436404 473474 437004 473476
rect 472404 473474 473004 473476
rect 508404 473474 509004 473476
rect 544404 473474 545004 473476
rect 580404 473474 581004 473476
rect 587160 473474 587760 473476
rect -1996 470476 -1396 470478
rect 804 470476 1404 470478
rect 36804 470476 37404 470478
rect 72804 470476 73404 470478
rect 108804 470476 109404 470478
rect 144804 470476 145404 470478
rect 180804 470476 181404 470478
rect 216804 470476 217404 470478
rect 252804 470476 253404 470478
rect 288804 470476 289404 470478
rect 324804 470476 325404 470478
rect 360804 470476 361404 470478
rect 396804 470476 397404 470478
rect 432804 470476 433404 470478
rect 468804 470476 469404 470478
rect 504804 470476 505404 470478
rect 540804 470476 541404 470478
rect 576804 470476 577404 470478
rect 585320 470476 585920 470478
rect -2916 470454 586840 470476
rect -2916 470218 -1814 470454
rect -1578 470218 986 470454
rect 1222 470218 36986 470454
rect 37222 470218 72986 470454
rect 73222 470218 108986 470454
rect 109222 470218 144986 470454
rect 145222 470218 180986 470454
rect 181222 470218 216986 470454
rect 217222 470218 252986 470454
rect 253222 470218 288986 470454
rect 289222 470218 324986 470454
rect 325222 470218 360986 470454
rect 361222 470218 396986 470454
rect 397222 470218 432986 470454
rect 433222 470218 468986 470454
rect 469222 470218 504986 470454
rect 505222 470218 540986 470454
rect 541222 470218 576986 470454
rect 577222 470218 585502 470454
rect 585738 470218 586840 470454
rect -2916 470134 586840 470218
rect -2916 469898 -1814 470134
rect -1578 469898 986 470134
rect 1222 469898 36986 470134
rect 37222 469898 72986 470134
rect 73222 469898 108986 470134
rect 109222 469898 144986 470134
rect 145222 469898 180986 470134
rect 181222 469898 216986 470134
rect 217222 469898 252986 470134
rect 253222 469898 288986 470134
rect 289222 469898 324986 470134
rect 325222 469898 360986 470134
rect 361222 469898 396986 470134
rect 397222 469898 432986 470134
rect 433222 469898 468986 470134
rect 469222 469898 504986 470134
rect 505222 469898 540986 470134
rect 541222 469898 576986 470134
rect 577222 469898 585502 470134
rect 585738 469898 586840 470134
rect -2916 469876 586840 469898
rect -1996 469874 -1396 469876
rect 804 469874 1404 469876
rect 36804 469874 37404 469876
rect 72804 469874 73404 469876
rect 108804 469874 109404 469876
rect 144804 469874 145404 469876
rect 180804 469874 181404 469876
rect 216804 469874 217404 469876
rect 252804 469874 253404 469876
rect 288804 469874 289404 469876
rect 324804 469874 325404 469876
rect 360804 469874 361404 469876
rect 396804 469874 397404 469876
rect 432804 469874 433404 469876
rect 468804 469874 469404 469876
rect 504804 469874 505404 469876
rect 540804 469874 541404 469876
rect 576804 469874 577404 469876
rect 585320 469874 585920 469876
rect -8436 463276 -7836 463278
rect 29604 463276 30204 463278
rect 65604 463276 66204 463278
rect 101604 463276 102204 463278
rect 137604 463276 138204 463278
rect 173604 463276 174204 463278
rect 209604 463276 210204 463278
rect 245604 463276 246204 463278
rect 281604 463276 282204 463278
rect 317604 463276 318204 463278
rect 353604 463276 354204 463278
rect 389604 463276 390204 463278
rect 425604 463276 426204 463278
rect 461604 463276 462204 463278
rect 497604 463276 498204 463278
rect 533604 463276 534204 463278
rect 569604 463276 570204 463278
rect 591760 463276 592360 463278
rect -8436 463254 592360 463276
rect -8436 463018 -8254 463254
rect -8018 463018 29786 463254
rect 30022 463018 65786 463254
rect 66022 463018 101786 463254
rect 102022 463018 137786 463254
rect 138022 463018 173786 463254
rect 174022 463018 209786 463254
rect 210022 463018 245786 463254
rect 246022 463018 281786 463254
rect 282022 463018 317786 463254
rect 318022 463018 353786 463254
rect 354022 463018 389786 463254
rect 390022 463018 425786 463254
rect 426022 463018 461786 463254
rect 462022 463018 497786 463254
rect 498022 463018 533786 463254
rect 534022 463018 569786 463254
rect 570022 463018 591942 463254
rect 592178 463018 592360 463254
rect -8436 462934 592360 463018
rect -8436 462698 -8254 462934
rect -8018 462698 29786 462934
rect 30022 462698 65786 462934
rect 66022 462698 101786 462934
rect 102022 462698 137786 462934
rect 138022 462698 173786 462934
rect 174022 462698 209786 462934
rect 210022 462698 245786 462934
rect 246022 462698 281786 462934
rect 282022 462698 317786 462934
rect 318022 462698 353786 462934
rect 354022 462698 389786 462934
rect 390022 462698 425786 462934
rect 426022 462698 461786 462934
rect 462022 462698 497786 462934
rect 498022 462698 533786 462934
rect 534022 462698 569786 462934
rect 570022 462698 591942 462934
rect 592178 462698 592360 462934
rect -8436 462676 592360 462698
rect -8436 462674 -7836 462676
rect 29604 462674 30204 462676
rect 65604 462674 66204 462676
rect 101604 462674 102204 462676
rect 137604 462674 138204 462676
rect 173604 462674 174204 462676
rect 209604 462674 210204 462676
rect 245604 462674 246204 462676
rect 281604 462674 282204 462676
rect 317604 462674 318204 462676
rect 353604 462674 354204 462676
rect 389604 462674 390204 462676
rect 425604 462674 426204 462676
rect 461604 462674 462204 462676
rect 497604 462674 498204 462676
rect 533604 462674 534204 462676
rect 569604 462674 570204 462676
rect 591760 462674 592360 462676
rect -6596 459676 -5996 459678
rect 26004 459676 26604 459678
rect 62004 459676 62604 459678
rect 98004 459676 98604 459678
rect 134004 459676 134604 459678
rect 170004 459676 170604 459678
rect 206004 459676 206604 459678
rect 242004 459676 242604 459678
rect 278004 459676 278604 459678
rect 314004 459676 314604 459678
rect 350004 459676 350604 459678
rect 386004 459676 386604 459678
rect 422004 459676 422604 459678
rect 458004 459676 458604 459678
rect 494004 459676 494604 459678
rect 530004 459676 530604 459678
rect 566004 459676 566604 459678
rect 589920 459676 590520 459678
rect -6596 459654 590520 459676
rect -6596 459418 -6414 459654
rect -6178 459418 26186 459654
rect 26422 459418 62186 459654
rect 62422 459418 98186 459654
rect 98422 459418 134186 459654
rect 134422 459418 170186 459654
rect 170422 459418 206186 459654
rect 206422 459418 242186 459654
rect 242422 459418 278186 459654
rect 278422 459418 314186 459654
rect 314422 459418 350186 459654
rect 350422 459418 386186 459654
rect 386422 459418 422186 459654
rect 422422 459418 458186 459654
rect 458422 459418 494186 459654
rect 494422 459418 530186 459654
rect 530422 459418 566186 459654
rect 566422 459418 590102 459654
rect 590338 459418 590520 459654
rect -6596 459334 590520 459418
rect -6596 459098 -6414 459334
rect -6178 459098 26186 459334
rect 26422 459098 62186 459334
rect 62422 459098 98186 459334
rect 98422 459098 134186 459334
rect 134422 459098 170186 459334
rect 170422 459098 206186 459334
rect 206422 459098 242186 459334
rect 242422 459098 278186 459334
rect 278422 459098 314186 459334
rect 314422 459098 350186 459334
rect 350422 459098 386186 459334
rect 386422 459098 422186 459334
rect 422422 459098 458186 459334
rect 458422 459098 494186 459334
rect 494422 459098 530186 459334
rect 530422 459098 566186 459334
rect 566422 459098 590102 459334
rect 590338 459098 590520 459334
rect -6596 459076 590520 459098
rect -6596 459074 -5996 459076
rect 26004 459074 26604 459076
rect 62004 459074 62604 459076
rect 98004 459074 98604 459076
rect 134004 459074 134604 459076
rect 170004 459074 170604 459076
rect 206004 459074 206604 459076
rect 242004 459074 242604 459076
rect 278004 459074 278604 459076
rect 314004 459074 314604 459076
rect 350004 459074 350604 459076
rect 386004 459074 386604 459076
rect 422004 459074 422604 459076
rect 458004 459074 458604 459076
rect 494004 459074 494604 459076
rect 530004 459074 530604 459076
rect 566004 459074 566604 459076
rect 589920 459074 590520 459076
rect -4756 456076 -4156 456078
rect 22404 456076 23004 456078
rect 58404 456076 59004 456078
rect 94404 456076 95004 456078
rect 130404 456076 131004 456078
rect 166404 456076 167004 456078
rect 202404 456076 203004 456078
rect 238404 456076 239004 456078
rect 274404 456076 275004 456078
rect 310404 456076 311004 456078
rect 346404 456076 347004 456078
rect 382404 456076 383004 456078
rect 418404 456076 419004 456078
rect 454404 456076 455004 456078
rect 490404 456076 491004 456078
rect 526404 456076 527004 456078
rect 562404 456076 563004 456078
rect 588080 456076 588680 456078
rect -4756 456054 588680 456076
rect -4756 455818 -4574 456054
rect -4338 455818 22586 456054
rect 22822 455818 58586 456054
rect 58822 455818 94586 456054
rect 94822 455818 130586 456054
rect 130822 455818 166586 456054
rect 166822 455818 202586 456054
rect 202822 455818 238586 456054
rect 238822 455818 274586 456054
rect 274822 455818 310586 456054
rect 310822 455818 346586 456054
rect 346822 455818 382586 456054
rect 382822 455818 418586 456054
rect 418822 455818 454586 456054
rect 454822 455818 490586 456054
rect 490822 455818 526586 456054
rect 526822 455818 562586 456054
rect 562822 455818 588262 456054
rect 588498 455818 588680 456054
rect -4756 455734 588680 455818
rect -4756 455498 -4574 455734
rect -4338 455498 22586 455734
rect 22822 455498 58586 455734
rect 58822 455498 94586 455734
rect 94822 455498 130586 455734
rect 130822 455498 166586 455734
rect 166822 455498 202586 455734
rect 202822 455498 238586 455734
rect 238822 455498 274586 455734
rect 274822 455498 310586 455734
rect 310822 455498 346586 455734
rect 346822 455498 382586 455734
rect 382822 455498 418586 455734
rect 418822 455498 454586 455734
rect 454822 455498 490586 455734
rect 490822 455498 526586 455734
rect 526822 455498 562586 455734
rect 562822 455498 588262 455734
rect 588498 455498 588680 455734
rect -4756 455476 588680 455498
rect -4756 455474 -4156 455476
rect 22404 455474 23004 455476
rect 58404 455474 59004 455476
rect 94404 455474 95004 455476
rect 130404 455474 131004 455476
rect 166404 455474 167004 455476
rect 202404 455474 203004 455476
rect 238404 455474 239004 455476
rect 274404 455474 275004 455476
rect 310404 455474 311004 455476
rect 346404 455474 347004 455476
rect 382404 455474 383004 455476
rect 418404 455474 419004 455476
rect 454404 455474 455004 455476
rect 490404 455474 491004 455476
rect 526404 455474 527004 455476
rect 562404 455474 563004 455476
rect 588080 455474 588680 455476
rect -2916 452476 -2316 452478
rect 18804 452476 19404 452478
rect 54804 452476 55404 452478
rect 90804 452476 91404 452478
rect 126804 452476 127404 452478
rect 162804 452476 163404 452478
rect 198804 452476 199404 452478
rect 234804 452476 235404 452478
rect 270804 452476 271404 452478
rect 306804 452476 307404 452478
rect 342804 452476 343404 452478
rect 378804 452476 379404 452478
rect 414804 452476 415404 452478
rect 450804 452476 451404 452478
rect 486804 452476 487404 452478
rect 522804 452476 523404 452478
rect 558804 452476 559404 452478
rect 586240 452476 586840 452478
rect -2916 452454 586840 452476
rect -2916 452218 -2734 452454
rect -2498 452218 18986 452454
rect 19222 452218 54986 452454
rect 55222 452218 90986 452454
rect 91222 452218 126986 452454
rect 127222 452218 162986 452454
rect 163222 452218 198986 452454
rect 199222 452218 234986 452454
rect 235222 452218 270986 452454
rect 271222 452218 306986 452454
rect 307222 452218 342986 452454
rect 343222 452218 378986 452454
rect 379222 452218 414986 452454
rect 415222 452218 450986 452454
rect 451222 452218 486986 452454
rect 487222 452218 522986 452454
rect 523222 452218 558986 452454
rect 559222 452218 586422 452454
rect 586658 452218 586840 452454
rect -2916 452134 586840 452218
rect -2916 451898 -2734 452134
rect -2498 451898 18986 452134
rect 19222 451898 54986 452134
rect 55222 451898 90986 452134
rect 91222 451898 126986 452134
rect 127222 451898 162986 452134
rect 163222 451898 198986 452134
rect 199222 451898 234986 452134
rect 235222 451898 270986 452134
rect 271222 451898 306986 452134
rect 307222 451898 342986 452134
rect 343222 451898 378986 452134
rect 379222 451898 414986 452134
rect 415222 451898 450986 452134
rect 451222 451898 486986 452134
rect 487222 451898 522986 452134
rect 523222 451898 558986 452134
rect 559222 451898 586422 452134
rect 586658 451898 586840 452134
rect -2916 451876 586840 451898
rect -2916 451874 -2316 451876
rect 18804 451874 19404 451876
rect 54804 451874 55404 451876
rect 90804 451874 91404 451876
rect 126804 451874 127404 451876
rect 162804 451874 163404 451876
rect 198804 451874 199404 451876
rect 234804 451874 235404 451876
rect 270804 451874 271404 451876
rect 306804 451874 307404 451876
rect 342804 451874 343404 451876
rect 378804 451874 379404 451876
rect 414804 451874 415404 451876
rect 450804 451874 451404 451876
rect 486804 451874 487404 451876
rect 522804 451874 523404 451876
rect 558804 451874 559404 451876
rect 586240 451874 586840 451876
rect -7516 445276 -6916 445278
rect 11604 445276 12204 445278
rect 47604 445276 48204 445278
rect 83604 445276 84204 445278
rect 119604 445276 120204 445278
rect 155604 445276 156204 445278
rect 191604 445276 192204 445278
rect 227604 445276 228204 445278
rect 263604 445276 264204 445278
rect 299604 445276 300204 445278
rect 335604 445276 336204 445278
rect 371604 445276 372204 445278
rect 407604 445276 408204 445278
rect 443604 445276 444204 445278
rect 479604 445276 480204 445278
rect 515604 445276 516204 445278
rect 551604 445276 552204 445278
rect 590840 445276 591440 445278
rect -8436 445254 592360 445276
rect -8436 445018 -7334 445254
rect -7098 445018 11786 445254
rect 12022 445018 47786 445254
rect 48022 445018 83786 445254
rect 84022 445018 119786 445254
rect 120022 445018 155786 445254
rect 156022 445018 191786 445254
rect 192022 445018 227786 445254
rect 228022 445018 263786 445254
rect 264022 445018 299786 445254
rect 300022 445018 335786 445254
rect 336022 445018 371786 445254
rect 372022 445018 407786 445254
rect 408022 445018 443786 445254
rect 444022 445018 479786 445254
rect 480022 445018 515786 445254
rect 516022 445018 551786 445254
rect 552022 445018 591022 445254
rect 591258 445018 592360 445254
rect -8436 444934 592360 445018
rect -8436 444698 -7334 444934
rect -7098 444698 11786 444934
rect 12022 444698 47786 444934
rect 48022 444698 83786 444934
rect 84022 444698 119786 444934
rect 120022 444698 155786 444934
rect 156022 444698 191786 444934
rect 192022 444698 227786 444934
rect 228022 444698 263786 444934
rect 264022 444698 299786 444934
rect 300022 444698 335786 444934
rect 336022 444698 371786 444934
rect 372022 444698 407786 444934
rect 408022 444698 443786 444934
rect 444022 444698 479786 444934
rect 480022 444698 515786 444934
rect 516022 444698 551786 444934
rect 552022 444698 591022 444934
rect 591258 444698 592360 444934
rect -8436 444676 592360 444698
rect -7516 444674 -6916 444676
rect 11604 444674 12204 444676
rect 47604 444674 48204 444676
rect 83604 444674 84204 444676
rect 119604 444674 120204 444676
rect 155604 444674 156204 444676
rect 191604 444674 192204 444676
rect 227604 444674 228204 444676
rect 263604 444674 264204 444676
rect 299604 444674 300204 444676
rect 335604 444674 336204 444676
rect 371604 444674 372204 444676
rect 407604 444674 408204 444676
rect 443604 444674 444204 444676
rect 479604 444674 480204 444676
rect 515604 444674 516204 444676
rect 551604 444674 552204 444676
rect 590840 444674 591440 444676
rect -5676 441676 -5076 441678
rect 8004 441676 8604 441678
rect 44004 441676 44604 441678
rect 80004 441676 80604 441678
rect 116004 441676 116604 441678
rect 152004 441676 152604 441678
rect 188004 441676 188604 441678
rect 224004 441676 224604 441678
rect 260004 441676 260604 441678
rect 296004 441676 296604 441678
rect 332004 441676 332604 441678
rect 368004 441676 368604 441678
rect 404004 441676 404604 441678
rect 440004 441676 440604 441678
rect 476004 441676 476604 441678
rect 512004 441676 512604 441678
rect 548004 441676 548604 441678
rect 589000 441676 589600 441678
rect -6596 441654 590520 441676
rect -6596 441418 -5494 441654
rect -5258 441418 8186 441654
rect 8422 441418 44186 441654
rect 44422 441418 80186 441654
rect 80422 441418 116186 441654
rect 116422 441418 152186 441654
rect 152422 441418 188186 441654
rect 188422 441418 224186 441654
rect 224422 441418 260186 441654
rect 260422 441418 296186 441654
rect 296422 441418 332186 441654
rect 332422 441418 368186 441654
rect 368422 441418 404186 441654
rect 404422 441418 440186 441654
rect 440422 441418 476186 441654
rect 476422 441418 512186 441654
rect 512422 441418 548186 441654
rect 548422 441418 589182 441654
rect 589418 441418 590520 441654
rect -6596 441334 590520 441418
rect -6596 441098 -5494 441334
rect -5258 441098 8186 441334
rect 8422 441098 44186 441334
rect 44422 441098 80186 441334
rect 80422 441098 116186 441334
rect 116422 441098 152186 441334
rect 152422 441098 188186 441334
rect 188422 441098 224186 441334
rect 224422 441098 260186 441334
rect 260422 441098 296186 441334
rect 296422 441098 332186 441334
rect 332422 441098 368186 441334
rect 368422 441098 404186 441334
rect 404422 441098 440186 441334
rect 440422 441098 476186 441334
rect 476422 441098 512186 441334
rect 512422 441098 548186 441334
rect 548422 441098 589182 441334
rect 589418 441098 590520 441334
rect -6596 441076 590520 441098
rect -5676 441074 -5076 441076
rect 8004 441074 8604 441076
rect 44004 441074 44604 441076
rect 80004 441074 80604 441076
rect 116004 441074 116604 441076
rect 152004 441074 152604 441076
rect 188004 441074 188604 441076
rect 224004 441074 224604 441076
rect 260004 441074 260604 441076
rect 296004 441074 296604 441076
rect 332004 441074 332604 441076
rect 368004 441074 368604 441076
rect 404004 441074 404604 441076
rect 440004 441074 440604 441076
rect 476004 441074 476604 441076
rect 512004 441074 512604 441076
rect 548004 441074 548604 441076
rect 589000 441074 589600 441076
rect -3836 438076 -3236 438078
rect 4404 438076 5004 438078
rect 40404 438076 41004 438078
rect 76404 438076 77004 438078
rect 112404 438076 113004 438078
rect 148404 438076 149004 438078
rect 184404 438076 185004 438078
rect 220404 438076 221004 438078
rect 256404 438076 257004 438078
rect 292404 438076 293004 438078
rect 328404 438076 329004 438078
rect 364404 438076 365004 438078
rect 400404 438076 401004 438078
rect 436404 438076 437004 438078
rect 472404 438076 473004 438078
rect 508404 438076 509004 438078
rect 544404 438076 545004 438078
rect 580404 438076 581004 438078
rect 587160 438076 587760 438078
rect -4756 438054 588680 438076
rect -4756 437818 -3654 438054
rect -3418 437818 4586 438054
rect 4822 437818 40586 438054
rect 40822 437818 76586 438054
rect 76822 437818 112586 438054
rect 112822 437818 148586 438054
rect 148822 437818 184586 438054
rect 184822 437818 220586 438054
rect 220822 437818 256586 438054
rect 256822 437818 292586 438054
rect 292822 437818 328586 438054
rect 328822 437818 364586 438054
rect 364822 437818 400586 438054
rect 400822 437818 436586 438054
rect 436822 437818 472586 438054
rect 472822 437818 508586 438054
rect 508822 437818 544586 438054
rect 544822 437818 580586 438054
rect 580822 437818 587342 438054
rect 587578 437818 588680 438054
rect -4756 437734 588680 437818
rect -4756 437498 -3654 437734
rect -3418 437498 4586 437734
rect 4822 437498 40586 437734
rect 40822 437498 76586 437734
rect 76822 437498 112586 437734
rect 112822 437498 148586 437734
rect 148822 437498 184586 437734
rect 184822 437498 220586 437734
rect 220822 437498 256586 437734
rect 256822 437498 292586 437734
rect 292822 437498 328586 437734
rect 328822 437498 364586 437734
rect 364822 437498 400586 437734
rect 400822 437498 436586 437734
rect 436822 437498 472586 437734
rect 472822 437498 508586 437734
rect 508822 437498 544586 437734
rect 544822 437498 580586 437734
rect 580822 437498 587342 437734
rect 587578 437498 588680 437734
rect -4756 437476 588680 437498
rect -3836 437474 -3236 437476
rect 4404 437474 5004 437476
rect 40404 437474 41004 437476
rect 76404 437474 77004 437476
rect 112404 437474 113004 437476
rect 148404 437474 149004 437476
rect 184404 437474 185004 437476
rect 220404 437474 221004 437476
rect 256404 437474 257004 437476
rect 292404 437474 293004 437476
rect 328404 437474 329004 437476
rect 364404 437474 365004 437476
rect 400404 437474 401004 437476
rect 436404 437474 437004 437476
rect 472404 437474 473004 437476
rect 508404 437474 509004 437476
rect 544404 437474 545004 437476
rect 580404 437474 581004 437476
rect 587160 437474 587760 437476
rect -1996 434476 -1396 434478
rect 804 434476 1404 434478
rect 36804 434476 37404 434478
rect 72804 434476 73404 434478
rect 108804 434476 109404 434478
rect 144804 434476 145404 434478
rect 180804 434476 181404 434478
rect 216804 434476 217404 434478
rect 252804 434476 253404 434478
rect 288804 434476 289404 434478
rect 324804 434476 325404 434478
rect 360804 434476 361404 434478
rect 396804 434476 397404 434478
rect 432804 434476 433404 434478
rect 468804 434476 469404 434478
rect 504804 434476 505404 434478
rect 540804 434476 541404 434478
rect 576804 434476 577404 434478
rect 585320 434476 585920 434478
rect -2916 434454 586840 434476
rect -2916 434218 -1814 434454
rect -1578 434218 986 434454
rect 1222 434218 36986 434454
rect 37222 434218 72986 434454
rect 73222 434218 108986 434454
rect 109222 434218 144986 434454
rect 145222 434218 180986 434454
rect 181222 434218 216986 434454
rect 217222 434218 252986 434454
rect 253222 434218 288986 434454
rect 289222 434218 324986 434454
rect 325222 434218 360986 434454
rect 361222 434218 396986 434454
rect 397222 434218 432986 434454
rect 433222 434218 468986 434454
rect 469222 434218 504986 434454
rect 505222 434218 540986 434454
rect 541222 434218 576986 434454
rect 577222 434218 585502 434454
rect 585738 434218 586840 434454
rect -2916 434134 586840 434218
rect -2916 433898 -1814 434134
rect -1578 433898 986 434134
rect 1222 433898 36986 434134
rect 37222 433898 72986 434134
rect 73222 433898 108986 434134
rect 109222 433898 144986 434134
rect 145222 433898 180986 434134
rect 181222 433898 216986 434134
rect 217222 433898 252986 434134
rect 253222 433898 288986 434134
rect 289222 433898 324986 434134
rect 325222 433898 360986 434134
rect 361222 433898 396986 434134
rect 397222 433898 432986 434134
rect 433222 433898 468986 434134
rect 469222 433898 504986 434134
rect 505222 433898 540986 434134
rect 541222 433898 576986 434134
rect 577222 433898 585502 434134
rect 585738 433898 586840 434134
rect -2916 433876 586840 433898
rect -1996 433874 -1396 433876
rect 804 433874 1404 433876
rect 36804 433874 37404 433876
rect 72804 433874 73404 433876
rect 108804 433874 109404 433876
rect 144804 433874 145404 433876
rect 180804 433874 181404 433876
rect 216804 433874 217404 433876
rect 252804 433874 253404 433876
rect 288804 433874 289404 433876
rect 324804 433874 325404 433876
rect 360804 433874 361404 433876
rect 396804 433874 397404 433876
rect 432804 433874 433404 433876
rect 468804 433874 469404 433876
rect 504804 433874 505404 433876
rect 540804 433874 541404 433876
rect 576804 433874 577404 433876
rect 585320 433874 585920 433876
rect -8436 427276 -7836 427278
rect 29604 427276 30204 427278
rect 65604 427276 66204 427278
rect 101604 427276 102204 427278
rect 137604 427276 138204 427278
rect 173604 427276 174204 427278
rect 209604 427276 210204 427278
rect 245604 427276 246204 427278
rect 281604 427276 282204 427278
rect 317604 427276 318204 427278
rect 353604 427276 354204 427278
rect 389604 427276 390204 427278
rect 425604 427276 426204 427278
rect 461604 427276 462204 427278
rect 497604 427276 498204 427278
rect 533604 427276 534204 427278
rect 569604 427276 570204 427278
rect 591760 427276 592360 427278
rect -8436 427254 592360 427276
rect -8436 427018 -8254 427254
rect -8018 427018 29786 427254
rect 30022 427018 65786 427254
rect 66022 427018 101786 427254
rect 102022 427018 137786 427254
rect 138022 427018 173786 427254
rect 174022 427018 209786 427254
rect 210022 427018 245786 427254
rect 246022 427018 281786 427254
rect 282022 427018 317786 427254
rect 318022 427018 353786 427254
rect 354022 427018 389786 427254
rect 390022 427018 425786 427254
rect 426022 427018 461786 427254
rect 462022 427018 497786 427254
rect 498022 427018 533786 427254
rect 534022 427018 569786 427254
rect 570022 427018 591942 427254
rect 592178 427018 592360 427254
rect -8436 426934 592360 427018
rect -8436 426698 -8254 426934
rect -8018 426698 29786 426934
rect 30022 426698 65786 426934
rect 66022 426698 101786 426934
rect 102022 426698 137786 426934
rect 138022 426698 173786 426934
rect 174022 426698 209786 426934
rect 210022 426698 245786 426934
rect 246022 426698 281786 426934
rect 282022 426698 317786 426934
rect 318022 426698 353786 426934
rect 354022 426698 389786 426934
rect 390022 426698 425786 426934
rect 426022 426698 461786 426934
rect 462022 426698 497786 426934
rect 498022 426698 533786 426934
rect 534022 426698 569786 426934
rect 570022 426698 591942 426934
rect 592178 426698 592360 426934
rect -8436 426676 592360 426698
rect -8436 426674 -7836 426676
rect 29604 426674 30204 426676
rect 65604 426674 66204 426676
rect 101604 426674 102204 426676
rect 137604 426674 138204 426676
rect 173604 426674 174204 426676
rect 209604 426674 210204 426676
rect 245604 426674 246204 426676
rect 281604 426674 282204 426676
rect 317604 426674 318204 426676
rect 353604 426674 354204 426676
rect 389604 426674 390204 426676
rect 425604 426674 426204 426676
rect 461604 426674 462204 426676
rect 497604 426674 498204 426676
rect 533604 426674 534204 426676
rect 569604 426674 570204 426676
rect 591760 426674 592360 426676
rect -6596 423676 -5996 423678
rect 26004 423676 26604 423678
rect 62004 423676 62604 423678
rect 98004 423676 98604 423678
rect 134004 423676 134604 423678
rect 170004 423676 170604 423678
rect 206004 423676 206604 423678
rect 242004 423676 242604 423678
rect 278004 423676 278604 423678
rect 314004 423676 314604 423678
rect 350004 423676 350604 423678
rect 386004 423676 386604 423678
rect 422004 423676 422604 423678
rect 458004 423676 458604 423678
rect 494004 423676 494604 423678
rect 530004 423676 530604 423678
rect 566004 423676 566604 423678
rect 589920 423676 590520 423678
rect -6596 423654 590520 423676
rect -6596 423418 -6414 423654
rect -6178 423418 26186 423654
rect 26422 423418 62186 423654
rect 62422 423418 98186 423654
rect 98422 423418 134186 423654
rect 134422 423418 170186 423654
rect 170422 423418 206186 423654
rect 206422 423418 242186 423654
rect 242422 423418 278186 423654
rect 278422 423418 314186 423654
rect 314422 423418 350186 423654
rect 350422 423418 386186 423654
rect 386422 423418 422186 423654
rect 422422 423418 458186 423654
rect 458422 423418 494186 423654
rect 494422 423418 530186 423654
rect 530422 423418 566186 423654
rect 566422 423418 590102 423654
rect 590338 423418 590520 423654
rect -6596 423334 590520 423418
rect -6596 423098 -6414 423334
rect -6178 423098 26186 423334
rect 26422 423098 62186 423334
rect 62422 423098 98186 423334
rect 98422 423098 134186 423334
rect 134422 423098 170186 423334
rect 170422 423098 206186 423334
rect 206422 423098 242186 423334
rect 242422 423098 278186 423334
rect 278422 423098 314186 423334
rect 314422 423098 350186 423334
rect 350422 423098 386186 423334
rect 386422 423098 422186 423334
rect 422422 423098 458186 423334
rect 458422 423098 494186 423334
rect 494422 423098 530186 423334
rect 530422 423098 566186 423334
rect 566422 423098 590102 423334
rect 590338 423098 590520 423334
rect -6596 423076 590520 423098
rect -6596 423074 -5996 423076
rect 26004 423074 26604 423076
rect 62004 423074 62604 423076
rect 98004 423074 98604 423076
rect 134004 423074 134604 423076
rect 170004 423074 170604 423076
rect 206004 423074 206604 423076
rect 242004 423074 242604 423076
rect 278004 423074 278604 423076
rect 314004 423074 314604 423076
rect 350004 423074 350604 423076
rect 386004 423074 386604 423076
rect 422004 423074 422604 423076
rect 458004 423074 458604 423076
rect 494004 423074 494604 423076
rect 530004 423074 530604 423076
rect 566004 423074 566604 423076
rect 589920 423074 590520 423076
rect -4756 420076 -4156 420078
rect 22404 420076 23004 420078
rect 58404 420076 59004 420078
rect 94404 420076 95004 420078
rect 130404 420076 131004 420078
rect 166404 420076 167004 420078
rect 202404 420076 203004 420078
rect 238404 420076 239004 420078
rect 274404 420076 275004 420078
rect 310404 420076 311004 420078
rect 346404 420076 347004 420078
rect 382404 420076 383004 420078
rect 418404 420076 419004 420078
rect 454404 420076 455004 420078
rect 490404 420076 491004 420078
rect 526404 420076 527004 420078
rect 562404 420076 563004 420078
rect 588080 420076 588680 420078
rect -4756 420054 588680 420076
rect -4756 419818 -4574 420054
rect -4338 419818 22586 420054
rect 22822 419818 58586 420054
rect 58822 419818 94586 420054
rect 94822 419818 130586 420054
rect 130822 419818 166586 420054
rect 166822 419818 202586 420054
rect 202822 419818 238586 420054
rect 238822 419818 274586 420054
rect 274822 419818 310586 420054
rect 310822 419818 346586 420054
rect 346822 419818 382586 420054
rect 382822 419818 418586 420054
rect 418822 419818 454586 420054
rect 454822 419818 490586 420054
rect 490822 419818 526586 420054
rect 526822 419818 562586 420054
rect 562822 419818 588262 420054
rect 588498 419818 588680 420054
rect -4756 419734 588680 419818
rect -4756 419498 -4574 419734
rect -4338 419498 22586 419734
rect 22822 419498 58586 419734
rect 58822 419498 94586 419734
rect 94822 419498 130586 419734
rect 130822 419498 166586 419734
rect 166822 419498 202586 419734
rect 202822 419498 238586 419734
rect 238822 419498 274586 419734
rect 274822 419498 310586 419734
rect 310822 419498 346586 419734
rect 346822 419498 382586 419734
rect 382822 419498 418586 419734
rect 418822 419498 454586 419734
rect 454822 419498 490586 419734
rect 490822 419498 526586 419734
rect 526822 419498 562586 419734
rect 562822 419498 588262 419734
rect 588498 419498 588680 419734
rect -4756 419476 588680 419498
rect -4756 419474 -4156 419476
rect 22404 419474 23004 419476
rect 58404 419474 59004 419476
rect 94404 419474 95004 419476
rect 130404 419474 131004 419476
rect 166404 419474 167004 419476
rect 202404 419474 203004 419476
rect 238404 419474 239004 419476
rect 274404 419474 275004 419476
rect 310404 419474 311004 419476
rect 346404 419474 347004 419476
rect 382404 419474 383004 419476
rect 418404 419474 419004 419476
rect 454404 419474 455004 419476
rect 490404 419474 491004 419476
rect 526404 419474 527004 419476
rect 562404 419474 563004 419476
rect 588080 419474 588680 419476
rect -2916 416476 -2316 416478
rect 18804 416476 19404 416478
rect 54804 416476 55404 416478
rect 90804 416476 91404 416478
rect 126804 416476 127404 416478
rect 162804 416476 163404 416478
rect 198804 416476 199404 416478
rect 234804 416476 235404 416478
rect 270804 416476 271404 416478
rect 306804 416476 307404 416478
rect 342804 416476 343404 416478
rect 378804 416476 379404 416478
rect 414804 416476 415404 416478
rect 450804 416476 451404 416478
rect 486804 416476 487404 416478
rect 522804 416476 523404 416478
rect 558804 416476 559404 416478
rect 586240 416476 586840 416478
rect -2916 416454 586840 416476
rect -2916 416218 -2734 416454
rect -2498 416218 18986 416454
rect 19222 416218 54986 416454
rect 55222 416218 90986 416454
rect 91222 416218 126986 416454
rect 127222 416218 162986 416454
rect 163222 416218 198986 416454
rect 199222 416218 234986 416454
rect 235222 416218 270986 416454
rect 271222 416218 306986 416454
rect 307222 416218 342986 416454
rect 343222 416218 378986 416454
rect 379222 416218 414986 416454
rect 415222 416218 450986 416454
rect 451222 416218 486986 416454
rect 487222 416218 522986 416454
rect 523222 416218 558986 416454
rect 559222 416218 586422 416454
rect 586658 416218 586840 416454
rect -2916 416134 586840 416218
rect -2916 415898 -2734 416134
rect -2498 415898 18986 416134
rect 19222 415898 54986 416134
rect 55222 415898 90986 416134
rect 91222 415898 126986 416134
rect 127222 415898 162986 416134
rect 163222 415898 198986 416134
rect 199222 415898 234986 416134
rect 235222 415898 270986 416134
rect 271222 415898 306986 416134
rect 307222 415898 342986 416134
rect 343222 415898 378986 416134
rect 379222 415898 414986 416134
rect 415222 415898 450986 416134
rect 451222 415898 486986 416134
rect 487222 415898 522986 416134
rect 523222 415898 558986 416134
rect 559222 415898 586422 416134
rect 586658 415898 586840 416134
rect -2916 415876 586840 415898
rect -2916 415874 -2316 415876
rect 18804 415874 19404 415876
rect 54804 415874 55404 415876
rect 90804 415874 91404 415876
rect 126804 415874 127404 415876
rect 162804 415874 163404 415876
rect 198804 415874 199404 415876
rect 234804 415874 235404 415876
rect 270804 415874 271404 415876
rect 306804 415874 307404 415876
rect 342804 415874 343404 415876
rect 378804 415874 379404 415876
rect 414804 415874 415404 415876
rect 450804 415874 451404 415876
rect 486804 415874 487404 415876
rect 522804 415874 523404 415876
rect 558804 415874 559404 415876
rect 586240 415874 586840 415876
rect -7516 409276 -6916 409278
rect 11604 409276 12204 409278
rect 47604 409276 48204 409278
rect 83604 409276 84204 409278
rect 119604 409276 120204 409278
rect 155604 409276 156204 409278
rect 191604 409276 192204 409278
rect 227604 409276 228204 409278
rect 263604 409276 264204 409278
rect 299604 409276 300204 409278
rect 335604 409276 336204 409278
rect 371604 409276 372204 409278
rect 407604 409276 408204 409278
rect 443604 409276 444204 409278
rect 479604 409276 480204 409278
rect 515604 409276 516204 409278
rect 551604 409276 552204 409278
rect 590840 409276 591440 409278
rect -8436 409254 592360 409276
rect -8436 409018 -7334 409254
rect -7098 409018 11786 409254
rect 12022 409018 47786 409254
rect 48022 409018 83786 409254
rect 84022 409018 119786 409254
rect 120022 409018 155786 409254
rect 156022 409018 191786 409254
rect 192022 409018 227786 409254
rect 228022 409018 263786 409254
rect 264022 409018 299786 409254
rect 300022 409018 335786 409254
rect 336022 409018 371786 409254
rect 372022 409018 407786 409254
rect 408022 409018 443786 409254
rect 444022 409018 479786 409254
rect 480022 409018 515786 409254
rect 516022 409018 551786 409254
rect 552022 409018 591022 409254
rect 591258 409018 592360 409254
rect -8436 408934 592360 409018
rect -8436 408698 -7334 408934
rect -7098 408698 11786 408934
rect 12022 408698 47786 408934
rect 48022 408698 83786 408934
rect 84022 408698 119786 408934
rect 120022 408698 155786 408934
rect 156022 408698 191786 408934
rect 192022 408698 227786 408934
rect 228022 408698 263786 408934
rect 264022 408698 299786 408934
rect 300022 408698 335786 408934
rect 336022 408698 371786 408934
rect 372022 408698 407786 408934
rect 408022 408698 443786 408934
rect 444022 408698 479786 408934
rect 480022 408698 515786 408934
rect 516022 408698 551786 408934
rect 552022 408698 591022 408934
rect 591258 408698 592360 408934
rect -8436 408676 592360 408698
rect -7516 408674 -6916 408676
rect 11604 408674 12204 408676
rect 47604 408674 48204 408676
rect 83604 408674 84204 408676
rect 119604 408674 120204 408676
rect 155604 408674 156204 408676
rect 191604 408674 192204 408676
rect 227604 408674 228204 408676
rect 263604 408674 264204 408676
rect 299604 408674 300204 408676
rect 335604 408674 336204 408676
rect 371604 408674 372204 408676
rect 407604 408674 408204 408676
rect 443604 408674 444204 408676
rect 479604 408674 480204 408676
rect 515604 408674 516204 408676
rect 551604 408674 552204 408676
rect 590840 408674 591440 408676
rect -5676 405676 -5076 405678
rect 8004 405676 8604 405678
rect 44004 405676 44604 405678
rect 80004 405676 80604 405678
rect 116004 405676 116604 405678
rect 152004 405676 152604 405678
rect 188004 405676 188604 405678
rect 224004 405676 224604 405678
rect 260004 405676 260604 405678
rect 296004 405676 296604 405678
rect 332004 405676 332604 405678
rect 368004 405676 368604 405678
rect 404004 405676 404604 405678
rect 440004 405676 440604 405678
rect 476004 405676 476604 405678
rect 512004 405676 512604 405678
rect 548004 405676 548604 405678
rect 589000 405676 589600 405678
rect -6596 405654 590520 405676
rect -6596 405418 -5494 405654
rect -5258 405418 8186 405654
rect 8422 405418 44186 405654
rect 44422 405418 80186 405654
rect 80422 405418 116186 405654
rect 116422 405418 152186 405654
rect 152422 405418 188186 405654
rect 188422 405418 224186 405654
rect 224422 405418 260186 405654
rect 260422 405418 296186 405654
rect 296422 405418 332186 405654
rect 332422 405418 368186 405654
rect 368422 405418 404186 405654
rect 404422 405418 440186 405654
rect 440422 405418 476186 405654
rect 476422 405418 512186 405654
rect 512422 405418 548186 405654
rect 548422 405418 589182 405654
rect 589418 405418 590520 405654
rect -6596 405334 590520 405418
rect -6596 405098 -5494 405334
rect -5258 405098 8186 405334
rect 8422 405098 44186 405334
rect 44422 405098 80186 405334
rect 80422 405098 116186 405334
rect 116422 405098 152186 405334
rect 152422 405098 188186 405334
rect 188422 405098 224186 405334
rect 224422 405098 260186 405334
rect 260422 405098 296186 405334
rect 296422 405098 332186 405334
rect 332422 405098 368186 405334
rect 368422 405098 404186 405334
rect 404422 405098 440186 405334
rect 440422 405098 476186 405334
rect 476422 405098 512186 405334
rect 512422 405098 548186 405334
rect 548422 405098 589182 405334
rect 589418 405098 590520 405334
rect -6596 405076 590520 405098
rect -5676 405074 -5076 405076
rect 8004 405074 8604 405076
rect 44004 405074 44604 405076
rect 80004 405074 80604 405076
rect 116004 405074 116604 405076
rect 152004 405074 152604 405076
rect 188004 405074 188604 405076
rect 224004 405074 224604 405076
rect 260004 405074 260604 405076
rect 296004 405074 296604 405076
rect 332004 405074 332604 405076
rect 368004 405074 368604 405076
rect 404004 405074 404604 405076
rect 440004 405074 440604 405076
rect 476004 405074 476604 405076
rect 512004 405074 512604 405076
rect 548004 405074 548604 405076
rect 589000 405074 589600 405076
rect -3836 402076 -3236 402078
rect 4404 402076 5004 402078
rect 40404 402076 41004 402078
rect 76404 402076 77004 402078
rect 112404 402076 113004 402078
rect 148404 402076 149004 402078
rect 184404 402076 185004 402078
rect 220404 402076 221004 402078
rect 256404 402076 257004 402078
rect 292404 402076 293004 402078
rect 328404 402076 329004 402078
rect 364404 402076 365004 402078
rect 400404 402076 401004 402078
rect 436404 402076 437004 402078
rect 472404 402076 473004 402078
rect 508404 402076 509004 402078
rect 544404 402076 545004 402078
rect 580404 402076 581004 402078
rect 587160 402076 587760 402078
rect -4756 402054 588680 402076
rect -4756 401818 -3654 402054
rect -3418 401818 4586 402054
rect 4822 401818 40586 402054
rect 40822 401818 76586 402054
rect 76822 401818 112586 402054
rect 112822 401818 148586 402054
rect 148822 401818 184586 402054
rect 184822 401818 220586 402054
rect 220822 401818 256586 402054
rect 256822 401818 292586 402054
rect 292822 401818 328586 402054
rect 328822 401818 364586 402054
rect 364822 401818 400586 402054
rect 400822 401818 436586 402054
rect 436822 401818 472586 402054
rect 472822 401818 508586 402054
rect 508822 401818 544586 402054
rect 544822 401818 580586 402054
rect 580822 401818 587342 402054
rect 587578 401818 588680 402054
rect -4756 401734 588680 401818
rect -4756 401498 -3654 401734
rect -3418 401498 4586 401734
rect 4822 401498 40586 401734
rect 40822 401498 76586 401734
rect 76822 401498 112586 401734
rect 112822 401498 148586 401734
rect 148822 401498 184586 401734
rect 184822 401498 220586 401734
rect 220822 401498 256586 401734
rect 256822 401498 292586 401734
rect 292822 401498 328586 401734
rect 328822 401498 364586 401734
rect 364822 401498 400586 401734
rect 400822 401498 436586 401734
rect 436822 401498 472586 401734
rect 472822 401498 508586 401734
rect 508822 401498 544586 401734
rect 544822 401498 580586 401734
rect 580822 401498 587342 401734
rect 587578 401498 588680 401734
rect -4756 401476 588680 401498
rect -3836 401474 -3236 401476
rect 4404 401474 5004 401476
rect 40404 401474 41004 401476
rect 76404 401474 77004 401476
rect 112404 401474 113004 401476
rect 148404 401474 149004 401476
rect 184404 401474 185004 401476
rect 220404 401474 221004 401476
rect 256404 401474 257004 401476
rect 292404 401474 293004 401476
rect 328404 401474 329004 401476
rect 364404 401474 365004 401476
rect 400404 401474 401004 401476
rect 436404 401474 437004 401476
rect 472404 401474 473004 401476
rect 508404 401474 509004 401476
rect 544404 401474 545004 401476
rect 580404 401474 581004 401476
rect 587160 401474 587760 401476
rect -1996 398476 -1396 398478
rect 804 398476 1404 398478
rect 36804 398476 37404 398478
rect 72804 398476 73404 398478
rect 108804 398476 109404 398478
rect 144804 398476 145404 398478
rect 180804 398476 181404 398478
rect 216804 398476 217404 398478
rect 252804 398476 253404 398478
rect 288804 398476 289404 398478
rect 324804 398476 325404 398478
rect 360804 398476 361404 398478
rect 396804 398476 397404 398478
rect 432804 398476 433404 398478
rect 468804 398476 469404 398478
rect 504804 398476 505404 398478
rect 540804 398476 541404 398478
rect 576804 398476 577404 398478
rect 585320 398476 585920 398478
rect -2916 398454 586840 398476
rect -2916 398218 -1814 398454
rect -1578 398218 986 398454
rect 1222 398218 36986 398454
rect 37222 398218 72986 398454
rect 73222 398218 108986 398454
rect 109222 398218 144986 398454
rect 145222 398218 180986 398454
rect 181222 398218 216986 398454
rect 217222 398218 252986 398454
rect 253222 398218 288986 398454
rect 289222 398218 324986 398454
rect 325222 398218 360986 398454
rect 361222 398218 396986 398454
rect 397222 398218 432986 398454
rect 433222 398218 468986 398454
rect 469222 398218 504986 398454
rect 505222 398218 540986 398454
rect 541222 398218 576986 398454
rect 577222 398218 585502 398454
rect 585738 398218 586840 398454
rect -2916 398134 586840 398218
rect -2916 397898 -1814 398134
rect -1578 397898 986 398134
rect 1222 397898 36986 398134
rect 37222 397898 72986 398134
rect 73222 397898 108986 398134
rect 109222 397898 144986 398134
rect 145222 397898 180986 398134
rect 181222 397898 216986 398134
rect 217222 397898 252986 398134
rect 253222 397898 288986 398134
rect 289222 397898 324986 398134
rect 325222 397898 360986 398134
rect 361222 397898 396986 398134
rect 397222 397898 432986 398134
rect 433222 397898 468986 398134
rect 469222 397898 504986 398134
rect 505222 397898 540986 398134
rect 541222 397898 576986 398134
rect 577222 397898 585502 398134
rect 585738 397898 586840 398134
rect -2916 397876 586840 397898
rect -1996 397874 -1396 397876
rect 804 397874 1404 397876
rect 36804 397874 37404 397876
rect 72804 397874 73404 397876
rect 108804 397874 109404 397876
rect 144804 397874 145404 397876
rect 180804 397874 181404 397876
rect 216804 397874 217404 397876
rect 252804 397874 253404 397876
rect 288804 397874 289404 397876
rect 324804 397874 325404 397876
rect 360804 397874 361404 397876
rect 396804 397874 397404 397876
rect 432804 397874 433404 397876
rect 468804 397874 469404 397876
rect 504804 397874 505404 397876
rect 540804 397874 541404 397876
rect 576804 397874 577404 397876
rect 585320 397874 585920 397876
rect -8436 391276 -7836 391278
rect 29604 391276 30204 391278
rect 65604 391276 66204 391278
rect 101604 391276 102204 391278
rect 137604 391276 138204 391278
rect 173604 391276 174204 391278
rect 209604 391276 210204 391278
rect 245604 391276 246204 391278
rect 281604 391276 282204 391278
rect 317604 391276 318204 391278
rect 353604 391276 354204 391278
rect 389604 391276 390204 391278
rect 425604 391276 426204 391278
rect 461604 391276 462204 391278
rect 497604 391276 498204 391278
rect 533604 391276 534204 391278
rect 569604 391276 570204 391278
rect 591760 391276 592360 391278
rect -8436 391254 592360 391276
rect -8436 391018 -8254 391254
rect -8018 391018 29786 391254
rect 30022 391018 65786 391254
rect 66022 391018 101786 391254
rect 102022 391018 137786 391254
rect 138022 391018 173786 391254
rect 174022 391018 209786 391254
rect 210022 391018 245786 391254
rect 246022 391018 281786 391254
rect 282022 391018 317786 391254
rect 318022 391018 353786 391254
rect 354022 391018 389786 391254
rect 390022 391018 425786 391254
rect 426022 391018 461786 391254
rect 462022 391018 497786 391254
rect 498022 391018 533786 391254
rect 534022 391018 569786 391254
rect 570022 391018 591942 391254
rect 592178 391018 592360 391254
rect -8436 390934 592360 391018
rect -8436 390698 -8254 390934
rect -8018 390698 29786 390934
rect 30022 390698 65786 390934
rect 66022 390698 101786 390934
rect 102022 390698 137786 390934
rect 138022 390698 173786 390934
rect 174022 390698 209786 390934
rect 210022 390698 245786 390934
rect 246022 390698 281786 390934
rect 282022 390698 317786 390934
rect 318022 390698 353786 390934
rect 354022 390698 389786 390934
rect 390022 390698 425786 390934
rect 426022 390698 461786 390934
rect 462022 390698 497786 390934
rect 498022 390698 533786 390934
rect 534022 390698 569786 390934
rect 570022 390698 591942 390934
rect 592178 390698 592360 390934
rect -8436 390676 592360 390698
rect -8436 390674 -7836 390676
rect 29604 390674 30204 390676
rect 65604 390674 66204 390676
rect 101604 390674 102204 390676
rect 137604 390674 138204 390676
rect 173604 390674 174204 390676
rect 209604 390674 210204 390676
rect 245604 390674 246204 390676
rect 281604 390674 282204 390676
rect 317604 390674 318204 390676
rect 353604 390674 354204 390676
rect 389604 390674 390204 390676
rect 425604 390674 426204 390676
rect 461604 390674 462204 390676
rect 497604 390674 498204 390676
rect 533604 390674 534204 390676
rect 569604 390674 570204 390676
rect 591760 390674 592360 390676
rect -6596 387676 -5996 387678
rect 26004 387676 26604 387678
rect 62004 387676 62604 387678
rect 98004 387676 98604 387678
rect 134004 387676 134604 387678
rect 170004 387676 170604 387678
rect 206004 387676 206604 387678
rect 242004 387676 242604 387678
rect 278004 387676 278604 387678
rect 314004 387676 314604 387678
rect 350004 387676 350604 387678
rect 386004 387676 386604 387678
rect 422004 387676 422604 387678
rect 458004 387676 458604 387678
rect 494004 387676 494604 387678
rect 530004 387676 530604 387678
rect 566004 387676 566604 387678
rect 589920 387676 590520 387678
rect -6596 387654 590520 387676
rect -6596 387418 -6414 387654
rect -6178 387418 26186 387654
rect 26422 387418 62186 387654
rect 62422 387418 98186 387654
rect 98422 387418 134186 387654
rect 134422 387418 170186 387654
rect 170422 387418 206186 387654
rect 206422 387418 242186 387654
rect 242422 387418 278186 387654
rect 278422 387418 314186 387654
rect 314422 387418 350186 387654
rect 350422 387418 386186 387654
rect 386422 387418 422186 387654
rect 422422 387418 458186 387654
rect 458422 387418 494186 387654
rect 494422 387418 530186 387654
rect 530422 387418 566186 387654
rect 566422 387418 590102 387654
rect 590338 387418 590520 387654
rect -6596 387334 590520 387418
rect -6596 387098 -6414 387334
rect -6178 387098 26186 387334
rect 26422 387098 62186 387334
rect 62422 387098 98186 387334
rect 98422 387098 134186 387334
rect 134422 387098 170186 387334
rect 170422 387098 206186 387334
rect 206422 387098 242186 387334
rect 242422 387098 278186 387334
rect 278422 387098 314186 387334
rect 314422 387098 350186 387334
rect 350422 387098 386186 387334
rect 386422 387098 422186 387334
rect 422422 387098 458186 387334
rect 458422 387098 494186 387334
rect 494422 387098 530186 387334
rect 530422 387098 566186 387334
rect 566422 387098 590102 387334
rect 590338 387098 590520 387334
rect -6596 387076 590520 387098
rect -6596 387074 -5996 387076
rect 26004 387074 26604 387076
rect 62004 387074 62604 387076
rect 98004 387074 98604 387076
rect 134004 387074 134604 387076
rect 170004 387074 170604 387076
rect 206004 387074 206604 387076
rect 242004 387074 242604 387076
rect 278004 387074 278604 387076
rect 314004 387074 314604 387076
rect 350004 387074 350604 387076
rect 386004 387074 386604 387076
rect 422004 387074 422604 387076
rect 458004 387074 458604 387076
rect 494004 387074 494604 387076
rect 530004 387074 530604 387076
rect 566004 387074 566604 387076
rect 589920 387074 590520 387076
rect -4756 384076 -4156 384078
rect 22404 384076 23004 384078
rect 58404 384076 59004 384078
rect 94404 384076 95004 384078
rect 130404 384076 131004 384078
rect 166404 384076 167004 384078
rect 202404 384076 203004 384078
rect 238404 384076 239004 384078
rect 274404 384076 275004 384078
rect 310404 384076 311004 384078
rect 346404 384076 347004 384078
rect 382404 384076 383004 384078
rect 418404 384076 419004 384078
rect 454404 384076 455004 384078
rect 490404 384076 491004 384078
rect 526404 384076 527004 384078
rect 562404 384076 563004 384078
rect 588080 384076 588680 384078
rect -4756 384054 588680 384076
rect -4756 383818 -4574 384054
rect -4338 383818 22586 384054
rect 22822 383818 58586 384054
rect 58822 383818 94586 384054
rect 94822 383818 130586 384054
rect 130822 383818 166586 384054
rect 166822 383818 202586 384054
rect 202822 383818 238586 384054
rect 238822 383818 274586 384054
rect 274822 383818 310586 384054
rect 310822 383818 346586 384054
rect 346822 383818 382586 384054
rect 382822 383818 418586 384054
rect 418822 383818 454586 384054
rect 454822 383818 490586 384054
rect 490822 383818 526586 384054
rect 526822 383818 562586 384054
rect 562822 383818 588262 384054
rect 588498 383818 588680 384054
rect -4756 383734 588680 383818
rect -4756 383498 -4574 383734
rect -4338 383498 22586 383734
rect 22822 383498 58586 383734
rect 58822 383498 94586 383734
rect 94822 383498 130586 383734
rect 130822 383498 166586 383734
rect 166822 383498 202586 383734
rect 202822 383498 238586 383734
rect 238822 383498 274586 383734
rect 274822 383498 310586 383734
rect 310822 383498 346586 383734
rect 346822 383498 382586 383734
rect 382822 383498 418586 383734
rect 418822 383498 454586 383734
rect 454822 383498 490586 383734
rect 490822 383498 526586 383734
rect 526822 383498 562586 383734
rect 562822 383498 588262 383734
rect 588498 383498 588680 383734
rect -4756 383476 588680 383498
rect -4756 383474 -4156 383476
rect 22404 383474 23004 383476
rect 58404 383474 59004 383476
rect 94404 383474 95004 383476
rect 130404 383474 131004 383476
rect 166404 383474 167004 383476
rect 202404 383474 203004 383476
rect 238404 383474 239004 383476
rect 274404 383474 275004 383476
rect 310404 383474 311004 383476
rect 346404 383474 347004 383476
rect 382404 383474 383004 383476
rect 418404 383474 419004 383476
rect 454404 383474 455004 383476
rect 490404 383474 491004 383476
rect 526404 383474 527004 383476
rect 562404 383474 563004 383476
rect 588080 383474 588680 383476
rect -2916 380476 -2316 380478
rect 18804 380476 19404 380478
rect 54804 380476 55404 380478
rect 90804 380476 91404 380478
rect 126804 380476 127404 380478
rect 162804 380476 163404 380478
rect 198804 380476 199404 380478
rect 234804 380476 235404 380478
rect 270804 380476 271404 380478
rect 306804 380476 307404 380478
rect 342804 380476 343404 380478
rect 378804 380476 379404 380478
rect 414804 380476 415404 380478
rect 450804 380476 451404 380478
rect 486804 380476 487404 380478
rect 522804 380476 523404 380478
rect 558804 380476 559404 380478
rect 586240 380476 586840 380478
rect -2916 380454 586840 380476
rect -2916 380218 -2734 380454
rect -2498 380218 18986 380454
rect 19222 380218 54986 380454
rect 55222 380218 90986 380454
rect 91222 380218 126986 380454
rect 127222 380218 162986 380454
rect 163222 380218 198986 380454
rect 199222 380218 234986 380454
rect 235222 380218 270986 380454
rect 271222 380218 306986 380454
rect 307222 380218 342986 380454
rect 343222 380218 378986 380454
rect 379222 380218 414986 380454
rect 415222 380218 450986 380454
rect 451222 380218 486986 380454
rect 487222 380218 522986 380454
rect 523222 380218 558986 380454
rect 559222 380218 586422 380454
rect 586658 380218 586840 380454
rect -2916 380134 586840 380218
rect -2916 379898 -2734 380134
rect -2498 379898 18986 380134
rect 19222 379898 54986 380134
rect 55222 379898 90986 380134
rect 91222 379898 126986 380134
rect 127222 379898 162986 380134
rect 163222 379898 198986 380134
rect 199222 379898 234986 380134
rect 235222 379898 270986 380134
rect 271222 379898 306986 380134
rect 307222 379898 342986 380134
rect 343222 379898 378986 380134
rect 379222 379898 414986 380134
rect 415222 379898 450986 380134
rect 451222 379898 486986 380134
rect 487222 379898 522986 380134
rect 523222 379898 558986 380134
rect 559222 379898 586422 380134
rect 586658 379898 586840 380134
rect -2916 379876 586840 379898
rect -2916 379874 -2316 379876
rect 18804 379874 19404 379876
rect 54804 379874 55404 379876
rect 90804 379874 91404 379876
rect 126804 379874 127404 379876
rect 162804 379874 163404 379876
rect 198804 379874 199404 379876
rect 234804 379874 235404 379876
rect 270804 379874 271404 379876
rect 306804 379874 307404 379876
rect 342804 379874 343404 379876
rect 378804 379874 379404 379876
rect 414804 379874 415404 379876
rect 450804 379874 451404 379876
rect 486804 379874 487404 379876
rect 522804 379874 523404 379876
rect 558804 379874 559404 379876
rect 586240 379874 586840 379876
rect -7516 373276 -6916 373278
rect 11604 373276 12204 373278
rect 47604 373276 48204 373278
rect 83604 373276 84204 373278
rect 119604 373276 120204 373278
rect 155604 373276 156204 373278
rect 191604 373276 192204 373278
rect 227604 373276 228204 373278
rect 263604 373276 264204 373278
rect 299604 373276 300204 373278
rect 335604 373276 336204 373278
rect 371604 373276 372204 373278
rect 407604 373276 408204 373278
rect 443604 373276 444204 373278
rect 479604 373276 480204 373278
rect 515604 373276 516204 373278
rect 551604 373276 552204 373278
rect 590840 373276 591440 373278
rect -8436 373254 592360 373276
rect -8436 373018 -7334 373254
rect -7098 373018 11786 373254
rect 12022 373018 47786 373254
rect 48022 373018 83786 373254
rect 84022 373018 119786 373254
rect 120022 373018 155786 373254
rect 156022 373018 191786 373254
rect 192022 373018 227786 373254
rect 228022 373018 263786 373254
rect 264022 373018 299786 373254
rect 300022 373018 335786 373254
rect 336022 373018 371786 373254
rect 372022 373018 407786 373254
rect 408022 373018 443786 373254
rect 444022 373018 479786 373254
rect 480022 373018 515786 373254
rect 516022 373018 551786 373254
rect 552022 373018 591022 373254
rect 591258 373018 592360 373254
rect -8436 372934 592360 373018
rect -8436 372698 -7334 372934
rect -7098 372698 11786 372934
rect 12022 372698 47786 372934
rect 48022 372698 83786 372934
rect 84022 372698 119786 372934
rect 120022 372698 155786 372934
rect 156022 372698 191786 372934
rect 192022 372698 227786 372934
rect 228022 372698 263786 372934
rect 264022 372698 299786 372934
rect 300022 372698 335786 372934
rect 336022 372698 371786 372934
rect 372022 372698 407786 372934
rect 408022 372698 443786 372934
rect 444022 372698 479786 372934
rect 480022 372698 515786 372934
rect 516022 372698 551786 372934
rect 552022 372698 591022 372934
rect 591258 372698 592360 372934
rect -8436 372676 592360 372698
rect -7516 372674 -6916 372676
rect 11604 372674 12204 372676
rect 47604 372674 48204 372676
rect 83604 372674 84204 372676
rect 119604 372674 120204 372676
rect 155604 372674 156204 372676
rect 191604 372674 192204 372676
rect 227604 372674 228204 372676
rect 263604 372674 264204 372676
rect 299604 372674 300204 372676
rect 335604 372674 336204 372676
rect 371604 372674 372204 372676
rect 407604 372674 408204 372676
rect 443604 372674 444204 372676
rect 479604 372674 480204 372676
rect 515604 372674 516204 372676
rect 551604 372674 552204 372676
rect 590840 372674 591440 372676
rect -5676 369676 -5076 369678
rect 8004 369676 8604 369678
rect 44004 369676 44604 369678
rect 80004 369676 80604 369678
rect 116004 369676 116604 369678
rect 152004 369676 152604 369678
rect 188004 369676 188604 369678
rect 224004 369676 224604 369678
rect 260004 369676 260604 369678
rect 296004 369676 296604 369678
rect 332004 369676 332604 369678
rect 368004 369676 368604 369678
rect 404004 369676 404604 369678
rect 440004 369676 440604 369678
rect 476004 369676 476604 369678
rect 512004 369676 512604 369678
rect 548004 369676 548604 369678
rect 589000 369676 589600 369678
rect -6596 369654 590520 369676
rect -6596 369418 -5494 369654
rect -5258 369418 8186 369654
rect 8422 369418 44186 369654
rect 44422 369418 80186 369654
rect 80422 369418 116186 369654
rect 116422 369418 152186 369654
rect 152422 369418 188186 369654
rect 188422 369418 224186 369654
rect 224422 369418 260186 369654
rect 260422 369418 296186 369654
rect 296422 369418 332186 369654
rect 332422 369418 368186 369654
rect 368422 369418 404186 369654
rect 404422 369418 440186 369654
rect 440422 369418 476186 369654
rect 476422 369418 512186 369654
rect 512422 369418 548186 369654
rect 548422 369418 589182 369654
rect 589418 369418 590520 369654
rect -6596 369334 590520 369418
rect -6596 369098 -5494 369334
rect -5258 369098 8186 369334
rect 8422 369098 44186 369334
rect 44422 369098 80186 369334
rect 80422 369098 116186 369334
rect 116422 369098 152186 369334
rect 152422 369098 188186 369334
rect 188422 369098 224186 369334
rect 224422 369098 260186 369334
rect 260422 369098 296186 369334
rect 296422 369098 332186 369334
rect 332422 369098 368186 369334
rect 368422 369098 404186 369334
rect 404422 369098 440186 369334
rect 440422 369098 476186 369334
rect 476422 369098 512186 369334
rect 512422 369098 548186 369334
rect 548422 369098 589182 369334
rect 589418 369098 590520 369334
rect -6596 369076 590520 369098
rect -5676 369074 -5076 369076
rect 8004 369074 8604 369076
rect 44004 369074 44604 369076
rect 80004 369074 80604 369076
rect 116004 369074 116604 369076
rect 152004 369074 152604 369076
rect 188004 369074 188604 369076
rect 224004 369074 224604 369076
rect 260004 369074 260604 369076
rect 296004 369074 296604 369076
rect 332004 369074 332604 369076
rect 368004 369074 368604 369076
rect 404004 369074 404604 369076
rect 440004 369074 440604 369076
rect 476004 369074 476604 369076
rect 512004 369074 512604 369076
rect 548004 369074 548604 369076
rect 589000 369074 589600 369076
rect -3836 366076 -3236 366078
rect 4404 366076 5004 366078
rect 40404 366076 41004 366078
rect 76404 366076 77004 366078
rect 112404 366076 113004 366078
rect 148404 366076 149004 366078
rect 184404 366076 185004 366078
rect 220404 366076 221004 366078
rect 256404 366076 257004 366078
rect 292404 366076 293004 366078
rect 328404 366076 329004 366078
rect 364404 366076 365004 366078
rect 400404 366076 401004 366078
rect 436404 366076 437004 366078
rect 472404 366076 473004 366078
rect 508404 366076 509004 366078
rect 544404 366076 545004 366078
rect 580404 366076 581004 366078
rect 587160 366076 587760 366078
rect -4756 366054 588680 366076
rect -4756 365818 -3654 366054
rect -3418 365818 4586 366054
rect 4822 365818 40586 366054
rect 40822 365818 76586 366054
rect 76822 365818 112586 366054
rect 112822 365818 148586 366054
rect 148822 365818 184586 366054
rect 184822 365818 220586 366054
rect 220822 365818 256586 366054
rect 256822 365818 292586 366054
rect 292822 365818 328586 366054
rect 328822 365818 364586 366054
rect 364822 365818 400586 366054
rect 400822 365818 436586 366054
rect 436822 365818 472586 366054
rect 472822 365818 508586 366054
rect 508822 365818 544586 366054
rect 544822 365818 580586 366054
rect 580822 365818 587342 366054
rect 587578 365818 588680 366054
rect -4756 365734 588680 365818
rect -4756 365498 -3654 365734
rect -3418 365498 4586 365734
rect 4822 365498 40586 365734
rect 40822 365498 76586 365734
rect 76822 365498 112586 365734
rect 112822 365498 148586 365734
rect 148822 365498 184586 365734
rect 184822 365498 220586 365734
rect 220822 365498 256586 365734
rect 256822 365498 292586 365734
rect 292822 365498 328586 365734
rect 328822 365498 364586 365734
rect 364822 365498 400586 365734
rect 400822 365498 436586 365734
rect 436822 365498 472586 365734
rect 472822 365498 508586 365734
rect 508822 365498 544586 365734
rect 544822 365498 580586 365734
rect 580822 365498 587342 365734
rect 587578 365498 588680 365734
rect -4756 365476 588680 365498
rect -3836 365474 -3236 365476
rect 4404 365474 5004 365476
rect 40404 365474 41004 365476
rect 76404 365474 77004 365476
rect 112404 365474 113004 365476
rect 148404 365474 149004 365476
rect 184404 365474 185004 365476
rect 220404 365474 221004 365476
rect 256404 365474 257004 365476
rect 292404 365474 293004 365476
rect 328404 365474 329004 365476
rect 364404 365474 365004 365476
rect 400404 365474 401004 365476
rect 436404 365474 437004 365476
rect 472404 365474 473004 365476
rect 508404 365474 509004 365476
rect 544404 365474 545004 365476
rect 580404 365474 581004 365476
rect 587160 365474 587760 365476
rect -1996 362476 -1396 362478
rect 804 362476 1404 362478
rect 36804 362476 37404 362478
rect 72804 362476 73404 362478
rect 108804 362476 109404 362478
rect 144804 362476 145404 362478
rect 180804 362476 181404 362478
rect 216804 362476 217404 362478
rect 252804 362476 253404 362478
rect 288804 362476 289404 362478
rect 324804 362476 325404 362478
rect 360804 362476 361404 362478
rect 396804 362476 397404 362478
rect 432804 362476 433404 362478
rect 468804 362476 469404 362478
rect 504804 362476 505404 362478
rect 540804 362476 541404 362478
rect 576804 362476 577404 362478
rect 585320 362476 585920 362478
rect -2916 362454 586840 362476
rect -2916 362218 -1814 362454
rect -1578 362218 986 362454
rect 1222 362218 36986 362454
rect 37222 362218 72986 362454
rect 73222 362218 108986 362454
rect 109222 362218 144986 362454
rect 145222 362218 180986 362454
rect 181222 362218 216986 362454
rect 217222 362218 252986 362454
rect 253222 362218 288986 362454
rect 289222 362218 324986 362454
rect 325222 362218 360986 362454
rect 361222 362218 396986 362454
rect 397222 362218 432986 362454
rect 433222 362218 468986 362454
rect 469222 362218 504986 362454
rect 505222 362218 540986 362454
rect 541222 362218 576986 362454
rect 577222 362218 585502 362454
rect 585738 362218 586840 362454
rect -2916 362134 586840 362218
rect -2916 361898 -1814 362134
rect -1578 361898 986 362134
rect 1222 361898 36986 362134
rect 37222 361898 72986 362134
rect 73222 361898 108986 362134
rect 109222 361898 144986 362134
rect 145222 361898 180986 362134
rect 181222 361898 216986 362134
rect 217222 361898 252986 362134
rect 253222 361898 288986 362134
rect 289222 361898 324986 362134
rect 325222 361898 360986 362134
rect 361222 361898 396986 362134
rect 397222 361898 432986 362134
rect 433222 361898 468986 362134
rect 469222 361898 504986 362134
rect 505222 361898 540986 362134
rect 541222 361898 576986 362134
rect 577222 361898 585502 362134
rect 585738 361898 586840 362134
rect -2916 361876 586840 361898
rect -1996 361874 -1396 361876
rect 804 361874 1404 361876
rect 36804 361874 37404 361876
rect 72804 361874 73404 361876
rect 108804 361874 109404 361876
rect 144804 361874 145404 361876
rect 180804 361874 181404 361876
rect 216804 361874 217404 361876
rect 252804 361874 253404 361876
rect 288804 361874 289404 361876
rect 324804 361874 325404 361876
rect 360804 361874 361404 361876
rect 396804 361874 397404 361876
rect 432804 361874 433404 361876
rect 468804 361874 469404 361876
rect 504804 361874 505404 361876
rect 540804 361874 541404 361876
rect 576804 361874 577404 361876
rect 585320 361874 585920 361876
rect -8436 355276 -7836 355278
rect 29604 355276 30204 355278
rect 65604 355276 66204 355278
rect 101604 355276 102204 355278
rect 137604 355276 138204 355278
rect 173604 355276 174204 355278
rect 209604 355276 210204 355278
rect 245604 355276 246204 355278
rect 281604 355276 282204 355278
rect 317604 355276 318204 355278
rect 353604 355276 354204 355278
rect 389604 355276 390204 355278
rect 425604 355276 426204 355278
rect 461604 355276 462204 355278
rect 497604 355276 498204 355278
rect 533604 355276 534204 355278
rect 569604 355276 570204 355278
rect 591760 355276 592360 355278
rect -8436 355254 592360 355276
rect -8436 355018 -8254 355254
rect -8018 355018 29786 355254
rect 30022 355018 65786 355254
rect 66022 355018 101786 355254
rect 102022 355018 137786 355254
rect 138022 355018 173786 355254
rect 174022 355018 209786 355254
rect 210022 355018 245786 355254
rect 246022 355018 281786 355254
rect 282022 355018 317786 355254
rect 318022 355018 353786 355254
rect 354022 355018 389786 355254
rect 390022 355018 425786 355254
rect 426022 355018 461786 355254
rect 462022 355018 497786 355254
rect 498022 355018 533786 355254
rect 534022 355018 569786 355254
rect 570022 355018 591942 355254
rect 592178 355018 592360 355254
rect -8436 354934 592360 355018
rect -8436 354698 -8254 354934
rect -8018 354698 29786 354934
rect 30022 354698 65786 354934
rect 66022 354698 101786 354934
rect 102022 354698 137786 354934
rect 138022 354698 173786 354934
rect 174022 354698 209786 354934
rect 210022 354698 245786 354934
rect 246022 354698 281786 354934
rect 282022 354698 317786 354934
rect 318022 354698 353786 354934
rect 354022 354698 389786 354934
rect 390022 354698 425786 354934
rect 426022 354698 461786 354934
rect 462022 354698 497786 354934
rect 498022 354698 533786 354934
rect 534022 354698 569786 354934
rect 570022 354698 591942 354934
rect 592178 354698 592360 354934
rect -8436 354676 592360 354698
rect -8436 354674 -7836 354676
rect 29604 354674 30204 354676
rect 65604 354674 66204 354676
rect 101604 354674 102204 354676
rect 137604 354674 138204 354676
rect 173604 354674 174204 354676
rect 209604 354674 210204 354676
rect 245604 354674 246204 354676
rect 281604 354674 282204 354676
rect 317604 354674 318204 354676
rect 353604 354674 354204 354676
rect 389604 354674 390204 354676
rect 425604 354674 426204 354676
rect 461604 354674 462204 354676
rect 497604 354674 498204 354676
rect 533604 354674 534204 354676
rect 569604 354674 570204 354676
rect 591760 354674 592360 354676
rect -6596 351676 -5996 351678
rect 26004 351676 26604 351678
rect 62004 351676 62604 351678
rect 98004 351676 98604 351678
rect 134004 351676 134604 351678
rect 170004 351676 170604 351678
rect 206004 351676 206604 351678
rect 242004 351676 242604 351678
rect 278004 351676 278604 351678
rect 314004 351676 314604 351678
rect 350004 351676 350604 351678
rect 386004 351676 386604 351678
rect 422004 351676 422604 351678
rect 458004 351676 458604 351678
rect 494004 351676 494604 351678
rect 530004 351676 530604 351678
rect 566004 351676 566604 351678
rect 589920 351676 590520 351678
rect -6596 351654 590520 351676
rect -6596 351418 -6414 351654
rect -6178 351418 26186 351654
rect 26422 351418 62186 351654
rect 62422 351418 98186 351654
rect 98422 351418 134186 351654
rect 134422 351418 170186 351654
rect 170422 351418 206186 351654
rect 206422 351418 242186 351654
rect 242422 351418 278186 351654
rect 278422 351418 314186 351654
rect 314422 351418 350186 351654
rect 350422 351418 386186 351654
rect 386422 351418 422186 351654
rect 422422 351418 458186 351654
rect 458422 351418 494186 351654
rect 494422 351418 530186 351654
rect 530422 351418 566186 351654
rect 566422 351418 590102 351654
rect 590338 351418 590520 351654
rect -6596 351334 590520 351418
rect -6596 351098 -6414 351334
rect -6178 351098 26186 351334
rect 26422 351098 62186 351334
rect 62422 351098 98186 351334
rect 98422 351098 134186 351334
rect 134422 351098 170186 351334
rect 170422 351098 206186 351334
rect 206422 351098 242186 351334
rect 242422 351098 278186 351334
rect 278422 351098 314186 351334
rect 314422 351098 350186 351334
rect 350422 351098 386186 351334
rect 386422 351098 422186 351334
rect 422422 351098 458186 351334
rect 458422 351098 494186 351334
rect 494422 351098 530186 351334
rect 530422 351098 566186 351334
rect 566422 351098 590102 351334
rect 590338 351098 590520 351334
rect -6596 351076 590520 351098
rect -6596 351074 -5996 351076
rect 26004 351074 26604 351076
rect 62004 351074 62604 351076
rect 98004 351074 98604 351076
rect 134004 351074 134604 351076
rect 170004 351074 170604 351076
rect 206004 351074 206604 351076
rect 242004 351074 242604 351076
rect 278004 351074 278604 351076
rect 314004 351074 314604 351076
rect 350004 351074 350604 351076
rect 386004 351074 386604 351076
rect 422004 351074 422604 351076
rect 458004 351074 458604 351076
rect 494004 351074 494604 351076
rect 530004 351074 530604 351076
rect 566004 351074 566604 351076
rect 589920 351074 590520 351076
rect -4756 348076 -4156 348078
rect 22404 348076 23004 348078
rect 58404 348076 59004 348078
rect 94404 348076 95004 348078
rect 130404 348076 131004 348078
rect 166404 348076 167004 348078
rect 202404 348076 203004 348078
rect 238404 348076 239004 348078
rect 274404 348076 275004 348078
rect 310404 348076 311004 348078
rect 346404 348076 347004 348078
rect 382404 348076 383004 348078
rect 418404 348076 419004 348078
rect 454404 348076 455004 348078
rect 490404 348076 491004 348078
rect 526404 348076 527004 348078
rect 562404 348076 563004 348078
rect 588080 348076 588680 348078
rect -4756 348054 588680 348076
rect -4756 347818 -4574 348054
rect -4338 347818 22586 348054
rect 22822 347818 58586 348054
rect 58822 347818 94586 348054
rect 94822 347818 130586 348054
rect 130822 347818 166586 348054
rect 166822 347818 202586 348054
rect 202822 347818 238586 348054
rect 238822 347818 274586 348054
rect 274822 347818 310586 348054
rect 310822 347818 346586 348054
rect 346822 347818 382586 348054
rect 382822 347818 418586 348054
rect 418822 347818 454586 348054
rect 454822 347818 490586 348054
rect 490822 347818 526586 348054
rect 526822 347818 562586 348054
rect 562822 347818 588262 348054
rect 588498 347818 588680 348054
rect -4756 347734 588680 347818
rect -4756 347498 -4574 347734
rect -4338 347498 22586 347734
rect 22822 347498 58586 347734
rect 58822 347498 94586 347734
rect 94822 347498 130586 347734
rect 130822 347498 166586 347734
rect 166822 347498 202586 347734
rect 202822 347498 238586 347734
rect 238822 347498 274586 347734
rect 274822 347498 310586 347734
rect 310822 347498 346586 347734
rect 346822 347498 382586 347734
rect 382822 347498 418586 347734
rect 418822 347498 454586 347734
rect 454822 347498 490586 347734
rect 490822 347498 526586 347734
rect 526822 347498 562586 347734
rect 562822 347498 588262 347734
rect 588498 347498 588680 347734
rect -4756 347476 588680 347498
rect -4756 347474 -4156 347476
rect 22404 347474 23004 347476
rect 58404 347474 59004 347476
rect 94404 347474 95004 347476
rect 130404 347474 131004 347476
rect 166404 347474 167004 347476
rect 202404 347474 203004 347476
rect 238404 347474 239004 347476
rect 274404 347474 275004 347476
rect 310404 347474 311004 347476
rect 346404 347474 347004 347476
rect 382404 347474 383004 347476
rect 418404 347474 419004 347476
rect 454404 347474 455004 347476
rect 490404 347474 491004 347476
rect 526404 347474 527004 347476
rect 562404 347474 563004 347476
rect 588080 347474 588680 347476
rect -2916 344476 -2316 344478
rect 18804 344476 19404 344478
rect 54804 344476 55404 344478
rect 90804 344476 91404 344478
rect 126804 344476 127404 344478
rect 162804 344476 163404 344478
rect 198804 344476 199404 344478
rect 234804 344476 235404 344478
rect 270804 344476 271404 344478
rect 306804 344476 307404 344478
rect 342804 344476 343404 344478
rect 378804 344476 379404 344478
rect 414804 344476 415404 344478
rect 450804 344476 451404 344478
rect 486804 344476 487404 344478
rect 522804 344476 523404 344478
rect 558804 344476 559404 344478
rect 586240 344476 586840 344478
rect -2916 344454 586840 344476
rect -2916 344218 -2734 344454
rect -2498 344218 18986 344454
rect 19222 344218 54986 344454
rect 55222 344218 90986 344454
rect 91222 344218 126986 344454
rect 127222 344218 162986 344454
rect 163222 344218 198986 344454
rect 199222 344218 234986 344454
rect 235222 344218 270986 344454
rect 271222 344218 306986 344454
rect 307222 344218 342986 344454
rect 343222 344218 378986 344454
rect 379222 344218 414986 344454
rect 415222 344218 450986 344454
rect 451222 344218 486986 344454
rect 487222 344218 522986 344454
rect 523222 344218 558986 344454
rect 559222 344218 586422 344454
rect 586658 344218 586840 344454
rect -2916 344134 586840 344218
rect -2916 343898 -2734 344134
rect -2498 343898 18986 344134
rect 19222 343898 54986 344134
rect 55222 343898 90986 344134
rect 91222 343898 126986 344134
rect 127222 343898 162986 344134
rect 163222 343898 198986 344134
rect 199222 343898 234986 344134
rect 235222 343898 270986 344134
rect 271222 343898 306986 344134
rect 307222 343898 342986 344134
rect 343222 343898 378986 344134
rect 379222 343898 414986 344134
rect 415222 343898 450986 344134
rect 451222 343898 486986 344134
rect 487222 343898 522986 344134
rect 523222 343898 558986 344134
rect 559222 343898 586422 344134
rect 586658 343898 586840 344134
rect -2916 343876 586840 343898
rect -2916 343874 -2316 343876
rect 18804 343874 19404 343876
rect 54804 343874 55404 343876
rect 90804 343874 91404 343876
rect 126804 343874 127404 343876
rect 162804 343874 163404 343876
rect 198804 343874 199404 343876
rect 234804 343874 235404 343876
rect 270804 343874 271404 343876
rect 306804 343874 307404 343876
rect 342804 343874 343404 343876
rect 378804 343874 379404 343876
rect 414804 343874 415404 343876
rect 450804 343874 451404 343876
rect 486804 343874 487404 343876
rect 522804 343874 523404 343876
rect 558804 343874 559404 343876
rect 586240 343874 586840 343876
rect -7516 337276 -6916 337278
rect 11604 337276 12204 337278
rect 47604 337276 48204 337278
rect 83604 337276 84204 337278
rect 119604 337276 120204 337278
rect 155604 337276 156204 337278
rect 191604 337276 192204 337278
rect 227604 337276 228204 337278
rect 263604 337276 264204 337278
rect 299604 337276 300204 337278
rect 335604 337276 336204 337278
rect 371604 337276 372204 337278
rect 407604 337276 408204 337278
rect 443604 337276 444204 337278
rect 479604 337276 480204 337278
rect 515604 337276 516204 337278
rect 551604 337276 552204 337278
rect 590840 337276 591440 337278
rect -8436 337254 592360 337276
rect -8436 337018 -7334 337254
rect -7098 337018 11786 337254
rect 12022 337018 47786 337254
rect 48022 337018 83786 337254
rect 84022 337018 119786 337254
rect 120022 337018 155786 337254
rect 156022 337018 191786 337254
rect 192022 337018 227786 337254
rect 228022 337018 263786 337254
rect 264022 337018 299786 337254
rect 300022 337018 335786 337254
rect 336022 337018 371786 337254
rect 372022 337018 407786 337254
rect 408022 337018 443786 337254
rect 444022 337018 479786 337254
rect 480022 337018 515786 337254
rect 516022 337018 551786 337254
rect 552022 337018 591022 337254
rect 591258 337018 592360 337254
rect -8436 336934 592360 337018
rect -8436 336698 -7334 336934
rect -7098 336698 11786 336934
rect 12022 336698 47786 336934
rect 48022 336698 83786 336934
rect 84022 336698 119786 336934
rect 120022 336698 155786 336934
rect 156022 336698 191786 336934
rect 192022 336698 227786 336934
rect 228022 336698 263786 336934
rect 264022 336698 299786 336934
rect 300022 336698 335786 336934
rect 336022 336698 371786 336934
rect 372022 336698 407786 336934
rect 408022 336698 443786 336934
rect 444022 336698 479786 336934
rect 480022 336698 515786 336934
rect 516022 336698 551786 336934
rect 552022 336698 591022 336934
rect 591258 336698 592360 336934
rect -8436 336676 592360 336698
rect -7516 336674 -6916 336676
rect 11604 336674 12204 336676
rect 47604 336674 48204 336676
rect 83604 336674 84204 336676
rect 119604 336674 120204 336676
rect 155604 336674 156204 336676
rect 191604 336674 192204 336676
rect 227604 336674 228204 336676
rect 263604 336674 264204 336676
rect 299604 336674 300204 336676
rect 335604 336674 336204 336676
rect 371604 336674 372204 336676
rect 407604 336674 408204 336676
rect 443604 336674 444204 336676
rect 479604 336674 480204 336676
rect 515604 336674 516204 336676
rect 551604 336674 552204 336676
rect 590840 336674 591440 336676
rect -5676 333676 -5076 333678
rect 8004 333676 8604 333678
rect 44004 333676 44604 333678
rect 80004 333676 80604 333678
rect 116004 333676 116604 333678
rect 152004 333676 152604 333678
rect 188004 333676 188604 333678
rect 224004 333676 224604 333678
rect 260004 333676 260604 333678
rect 296004 333676 296604 333678
rect 332004 333676 332604 333678
rect 368004 333676 368604 333678
rect 404004 333676 404604 333678
rect 440004 333676 440604 333678
rect 476004 333676 476604 333678
rect 512004 333676 512604 333678
rect 548004 333676 548604 333678
rect 589000 333676 589600 333678
rect -6596 333654 590520 333676
rect -6596 333418 -5494 333654
rect -5258 333418 8186 333654
rect 8422 333418 44186 333654
rect 44422 333418 80186 333654
rect 80422 333418 116186 333654
rect 116422 333418 152186 333654
rect 152422 333418 188186 333654
rect 188422 333418 224186 333654
rect 224422 333418 260186 333654
rect 260422 333418 296186 333654
rect 296422 333418 332186 333654
rect 332422 333418 368186 333654
rect 368422 333418 404186 333654
rect 404422 333418 440186 333654
rect 440422 333418 476186 333654
rect 476422 333418 512186 333654
rect 512422 333418 548186 333654
rect 548422 333418 589182 333654
rect 589418 333418 590520 333654
rect -6596 333334 590520 333418
rect -6596 333098 -5494 333334
rect -5258 333098 8186 333334
rect 8422 333098 44186 333334
rect 44422 333098 80186 333334
rect 80422 333098 116186 333334
rect 116422 333098 152186 333334
rect 152422 333098 188186 333334
rect 188422 333098 224186 333334
rect 224422 333098 260186 333334
rect 260422 333098 296186 333334
rect 296422 333098 332186 333334
rect 332422 333098 368186 333334
rect 368422 333098 404186 333334
rect 404422 333098 440186 333334
rect 440422 333098 476186 333334
rect 476422 333098 512186 333334
rect 512422 333098 548186 333334
rect 548422 333098 589182 333334
rect 589418 333098 590520 333334
rect -6596 333076 590520 333098
rect -5676 333074 -5076 333076
rect 8004 333074 8604 333076
rect 44004 333074 44604 333076
rect 80004 333074 80604 333076
rect 116004 333074 116604 333076
rect 152004 333074 152604 333076
rect 188004 333074 188604 333076
rect 224004 333074 224604 333076
rect 260004 333074 260604 333076
rect 296004 333074 296604 333076
rect 332004 333074 332604 333076
rect 368004 333074 368604 333076
rect 404004 333074 404604 333076
rect 440004 333074 440604 333076
rect 476004 333074 476604 333076
rect 512004 333074 512604 333076
rect 548004 333074 548604 333076
rect 589000 333074 589600 333076
rect -3836 330076 -3236 330078
rect 4404 330076 5004 330078
rect 40404 330076 41004 330078
rect 76404 330076 77004 330078
rect 112404 330076 113004 330078
rect 148404 330076 149004 330078
rect 184404 330076 185004 330078
rect 220404 330076 221004 330078
rect 256404 330076 257004 330078
rect 292404 330076 293004 330078
rect 328404 330076 329004 330078
rect 364404 330076 365004 330078
rect 400404 330076 401004 330078
rect 436404 330076 437004 330078
rect 472404 330076 473004 330078
rect 508404 330076 509004 330078
rect 544404 330076 545004 330078
rect 580404 330076 581004 330078
rect 587160 330076 587760 330078
rect -4756 330054 588680 330076
rect -4756 329818 -3654 330054
rect -3418 329818 4586 330054
rect 4822 329818 40586 330054
rect 40822 329818 76586 330054
rect 76822 329818 112586 330054
rect 112822 329818 148586 330054
rect 148822 329818 184586 330054
rect 184822 329818 220586 330054
rect 220822 329818 256586 330054
rect 256822 329818 292586 330054
rect 292822 329818 328586 330054
rect 328822 329818 364586 330054
rect 364822 329818 400586 330054
rect 400822 329818 436586 330054
rect 436822 329818 472586 330054
rect 472822 329818 508586 330054
rect 508822 329818 544586 330054
rect 544822 329818 580586 330054
rect 580822 329818 587342 330054
rect 587578 329818 588680 330054
rect -4756 329734 588680 329818
rect -4756 329498 -3654 329734
rect -3418 329498 4586 329734
rect 4822 329498 40586 329734
rect 40822 329498 76586 329734
rect 76822 329498 112586 329734
rect 112822 329498 148586 329734
rect 148822 329498 184586 329734
rect 184822 329498 220586 329734
rect 220822 329498 256586 329734
rect 256822 329498 292586 329734
rect 292822 329498 328586 329734
rect 328822 329498 364586 329734
rect 364822 329498 400586 329734
rect 400822 329498 436586 329734
rect 436822 329498 472586 329734
rect 472822 329498 508586 329734
rect 508822 329498 544586 329734
rect 544822 329498 580586 329734
rect 580822 329498 587342 329734
rect 587578 329498 588680 329734
rect -4756 329476 588680 329498
rect -3836 329474 -3236 329476
rect 4404 329474 5004 329476
rect 40404 329474 41004 329476
rect 76404 329474 77004 329476
rect 112404 329474 113004 329476
rect 148404 329474 149004 329476
rect 184404 329474 185004 329476
rect 220404 329474 221004 329476
rect 256404 329474 257004 329476
rect 292404 329474 293004 329476
rect 328404 329474 329004 329476
rect 364404 329474 365004 329476
rect 400404 329474 401004 329476
rect 436404 329474 437004 329476
rect 472404 329474 473004 329476
rect 508404 329474 509004 329476
rect 544404 329474 545004 329476
rect 580404 329474 581004 329476
rect 587160 329474 587760 329476
rect -1996 326476 -1396 326478
rect 804 326476 1404 326478
rect 36804 326476 37404 326478
rect 72804 326476 73404 326478
rect 108804 326476 109404 326478
rect 144804 326476 145404 326478
rect 180804 326476 181404 326478
rect 216804 326476 217404 326478
rect 252804 326476 253404 326478
rect 288804 326476 289404 326478
rect 324804 326476 325404 326478
rect 360804 326476 361404 326478
rect 396804 326476 397404 326478
rect 432804 326476 433404 326478
rect 468804 326476 469404 326478
rect 504804 326476 505404 326478
rect 540804 326476 541404 326478
rect 576804 326476 577404 326478
rect 585320 326476 585920 326478
rect -2916 326454 586840 326476
rect -2916 326218 -1814 326454
rect -1578 326218 986 326454
rect 1222 326218 36986 326454
rect 37222 326218 72986 326454
rect 73222 326218 108986 326454
rect 109222 326218 144986 326454
rect 145222 326218 180986 326454
rect 181222 326218 216986 326454
rect 217222 326218 252986 326454
rect 253222 326218 288986 326454
rect 289222 326218 324986 326454
rect 325222 326218 360986 326454
rect 361222 326218 396986 326454
rect 397222 326218 432986 326454
rect 433222 326218 468986 326454
rect 469222 326218 504986 326454
rect 505222 326218 540986 326454
rect 541222 326218 576986 326454
rect 577222 326218 585502 326454
rect 585738 326218 586840 326454
rect -2916 326134 586840 326218
rect -2916 325898 -1814 326134
rect -1578 325898 986 326134
rect 1222 325898 36986 326134
rect 37222 325898 72986 326134
rect 73222 325898 108986 326134
rect 109222 325898 144986 326134
rect 145222 325898 180986 326134
rect 181222 325898 216986 326134
rect 217222 325898 252986 326134
rect 253222 325898 288986 326134
rect 289222 325898 324986 326134
rect 325222 325898 360986 326134
rect 361222 325898 396986 326134
rect 397222 325898 432986 326134
rect 433222 325898 468986 326134
rect 469222 325898 504986 326134
rect 505222 325898 540986 326134
rect 541222 325898 576986 326134
rect 577222 325898 585502 326134
rect 585738 325898 586840 326134
rect -2916 325876 586840 325898
rect -1996 325874 -1396 325876
rect 804 325874 1404 325876
rect 36804 325874 37404 325876
rect 72804 325874 73404 325876
rect 108804 325874 109404 325876
rect 144804 325874 145404 325876
rect 180804 325874 181404 325876
rect 216804 325874 217404 325876
rect 252804 325874 253404 325876
rect 288804 325874 289404 325876
rect 324804 325874 325404 325876
rect 360804 325874 361404 325876
rect 396804 325874 397404 325876
rect 432804 325874 433404 325876
rect 468804 325874 469404 325876
rect 504804 325874 505404 325876
rect 540804 325874 541404 325876
rect 576804 325874 577404 325876
rect 585320 325874 585920 325876
rect -8436 319276 -7836 319278
rect 29604 319276 30204 319278
rect 65604 319276 66204 319278
rect 101604 319276 102204 319278
rect 137604 319276 138204 319278
rect 173604 319276 174204 319278
rect 209604 319276 210204 319278
rect 245604 319276 246204 319278
rect 281604 319276 282204 319278
rect 317604 319276 318204 319278
rect 353604 319276 354204 319278
rect 389604 319276 390204 319278
rect 425604 319276 426204 319278
rect 461604 319276 462204 319278
rect 497604 319276 498204 319278
rect 533604 319276 534204 319278
rect 569604 319276 570204 319278
rect 591760 319276 592360 319278
rect -8436 319254 592360 319276
rect -8436 319018 -8254 319254
rect -8018 319018 29786 319254
rect 30022 319018 65786 319254
rect 66022 319018 101786 319254
rect 102022 319018 137786 319254
rect 138022 319018 173786 319254
rect 174022 319018 209786 319254
rect 210022 319018 245786 319254
rect 246022 319018 281786 319254
rect 282022 319018 317786 319254
rect 318022 319018 353786 319254
rect 354022 319018 389786 319254
rect 390022 319018 425786 319254
rect 426022 319018 461786 319254
rect 462022 319018 497786 319254
rect 498022 319018 533786 319254
rect 534022 319018 569786 319254
rect 570022 319018 591942 319254
rect 592178 319018 592360 319254
rect -8436 318934 592360 319018
rect -8436 318698 -8254 318934
rect -8018 318698 29786 318934
rect 30022 318698 65786 318934
rect 66022 318698 101786 318934
rect 102022 318698 137786 318934
rect 138022 318698 173786 318934
rect 174022 318698 209786 318934
rect 210022 318698 245786 318934
rect 246022 318698 281786 318934
rect 282022 318698 317786 318934
rect 318022 318698 353786 318934
rect 354022 318698 389786 318934
rect 390022 318698 425786 318934
rect 426022 318698 461786 318934
rect 462022 318698 497786 318934
rect 498022 318698 533786 318934
rect 534022 318698 569786 318934
rect 570022 318698 591942 318934
rect 592178 318698 592360 318934
rect -8436 318676 592360 318698
rect -8436 318674 -7836 318676
rect 29604 318674 30204 318676
rect 65604 318674 66204 318676
rect 101604 318674 102204 318676
rect 137604 318674 138204 318676
rect 173604 318674 174204 318676
rect 209604 318674 210204 318676
rect 245604 318674 246204 318676
rect 281604 318674 282204 318676
rect 317604 318674 318204 318676
rect 353604 318674 354204 318676
rect 389604 318674 390204 318676
rect 425604 318674 426204 318676
rect 461604 318674 462204 318676
rect 497604 318674 498204 318676
rect 533604 318674 534204 318676
rect 569604 318674 570204 318676
rect 591760 318674 592360 318676
rect -6596 315676 -5996 315678
rect 26004 315676 26604 315678
rect 62004 315676 62604 315678
rect 98004 315676 98604 315678
rect 134004 315676 134604 315678
rect 170004 315676 170604 315678
rect 206004 315676 206604 315678
rect 242004 315676 242604 315678
rect 278004 315676 278604 315678
rect 314004 315676 314604 315678
rect 350004 315676 350604 315678
rect 386004 315676 386604 315678
rect 422004 315676 422604 315678
rect 458004 315676 458604 315678
rect 494004 315676 494604 315678
rect 530004 315676 530604 315678
rect 566004 315676 566604 315678
rect 589920 315676 590520 315678
rect -6596 315654 590520 315676
rect -6596 315418 -6414 315654
rect -6178 315418 26186 315654
rect 26422 315418 62186 315654
rect 62422 315418 98186 315654
rect 98422 315418 134186 315654
rect 134422 315418 170186 315654
rect 170422 315418 206186 315654
rect 206422 315418 242186 315654
rect 242422 315418 278186 315654
rect 278422 315418 314186 315654
rect 314422 315418 350186 315654
rect 350422 315418 386186 315654
rect 386422 315418 422186 315654
rect 422422 315418 458186 315654
rect 458422 315418 494186 315654
rect 494422 315418 530186 315654
rect 530422 315418 566186 315654
rect 566422 315418 590102 315654
rect 590338 315418 590520 315654
rect -6596 315334 590520 315418
rect -6596 315098 -6414 315334
rect -6178 315098 26186 315334
rect 26422 315098 62186 315334
rect 62422 315098 98186 315334
rect 98422 315098 134186 315334
rect 134422 315098 170186 315334
rect 170422 315098 206186 315334
rect 206422 315098 242186 315334
rect 242422 315098 278186 315334
rect 278422 315098 314186 315334
rect 314422 315098 350186 315334
rect 350422 315098 386186 315334
rect 386422 315098 422186 315334
rect 422422 315098 458186 315334
rect 458422 315098 494186 315334
rect 494422 315098 530186 315334
rect 530422 315098 566186 315334
rect 566422 315098 590102 315334
rect 590338 315098 590520 315334
rect -6596 315076 590520 315098
rect -6596 315074 -5996 315076
rect 26004 315074 26604 315076
rect 62004 315074 62604 315076
rect 98004 315074 98604 315076
rect 134004 315074 134604 315076
rect 170004 315074 170604 315076
rect 206004 315074 206604 315076
rect 242004 315074 242604 315076
rect 278004 315074 278604 315076
rect 314004 315074 314604 315076
rect 350004 315074 350604 315076
rect 386004 315074 386604 315076
rect 422004 315074 422604 315076
rect 458004 315074 458604 315076
rect 494004 315074 494604 315076
rect 530004 315074 530604 315076
rect 566004 315074 566604 315076
rect 589920 315074 590520 315076
rect -4756 312076 -4156 312078
rect 22404 312076 23004 312078
rect 58404 312076 59004 312078
rect 94404 312076 95004 312078
rect 130404 312076 131004 312078
rect 166404 312076 167004 312078
rect 202404 312076 203004 312078
rect 238404 312076 239004 312078
rect 274404 312076 275004 312078
rect 310404 312076 311004 312078
rect 346404 312076 347004 312078
rect 382404 312076 383004 312078
rect 418404 312076 419004 312078
rect 454404 312076 455004 312078
rect 490404 312076 491004 312078
rect 526404 312076 527004 312078
rect 562404 312076 563004 312078
rect 588080 312076 588680 312078
rect -4756 312054 588680 312076
rect -4756 311818 -4574 312054
rect -4338 311818 22586 312054
rect 22822 311818 58586 312054
rect 58822 311818 94586 312054
rect 94822 311818 130586 312054
rect 130822 311818 166586 312054
rect 166822 311818 202586 312054
rect 202822 311818 238586 312054
rect 238822 311818 274586 312054
rect 274822 311818 310586 312054
rect 310822 311818 346586 312054
rect 346822 311818 382586 312054
rect 382822 311818 418586 312054
rect 418822 311818 454586 312054
rect 454822 311818 490586 312054
rect 490822 311818 526586 312054
rect 526822 311818 562586 312054
rect 562822 311818 588262 312054
rect 588498 311818 588680 312054
rect -4756 311734 588680 311818
rect -4756 311498 -4574 311734
rect -4338 311498 22586 311734
rect 22822 311498 58586 311734
rect 58822 311498 94586 311734
rect 94822 311498 130586 311734
rect 130822 311498 166586 311734
rect 166822 311498 202586 311734
rect 202822 311498 238586 311734
rect 238822 311498 274586 311734
rect 274822 311498 310586 311734
rect 310822 311498 346586 311734
rect 346822 311498 382586 311734
rect 382822 311498 418586 311734
rect 418822 311498 454586 311734
rect 454822 311498 490586 311734
rect 490822 311498 526586 311734
rect 526822 311498 562586 311734
rect 562822 311498 588262 311734
rect 588498 311498 588680 311734
rect -4756 311476 588680 311498
rect -4756 311474 -4156 311476
rect 22404 311474 23004 311476
rect 58404 311474 59004 311476
rect 94404 311474 95004 311476
rect 130404 311474 131004 311476
rect 166404 311474 167004 311476
rect 202404 311474 203004 311476
rect 238404 311474 239004 311476
rect 274404 311474 275004 311476
rect 310404 311474 311004 311476
rect 346404 311474 347004 311476
rect 382404 311474 383004 311476
rect 418404 311474 419004 311476
rect 454404 311474 455004 311476
rect 490404 311474 491004 311476
rect 526404 311474 527004 311476
rect 562404 311474 563004 311476
rect 588080 311474 588680 311476
rect -2916 308476 -2316 308478
rect 18804 308476 19404 308478
rect 54804 308476 55404 308478
rect 90804 308476 91404 308478
rect 126804 308476 127404 308478
rect 162804 308476 163404 308478
rect 198804 308476 199404 308478
rect 234804 308476 235404 308478
rect 270804 308476 271404 308478
rect 306804 308476 307404 308478
rect 342804 308476 343404 308478
rect 378804 308476 379404 308478
rect 414804 308476 415404 308478
rect 450804 308476 451404 308478
rect 486804 308476 487404 308478
rect 522804 308476 523404 308478
rect 558804 308476 559404 308478
rect 586240 308476 586840 308478
rect -2916 308454 586840 308476
rect -2916 308218 -2734 308454
rect -2498 308218 18986 308454
rect 19222 308218 54986 308454
rect 55222 308218 90986 308454
rect 91222 308218 126986 308454
rect 127222 308218 162986 308454
rect 163222 308218 198986 308454
rect 199222 308218 234986 308454
rect 235222 308218 270986 308454
rect 271222 308218 306986 308454
rect 307222 308218 342986 308454
rect 343222 308218 378986 308454
rect 379222 308218 414986 308454
rect 415222 308218 450986 308454
rect 451222 308218 486986 308454
rect 487222 308218 522986 308454
rect 523222 308218 558986 308454
rect 559222 308218 586422 308454
rect 586658 308218 586840 308454
rect -2916 308134 586840 308218
rect -2916 307898 -2734 308134
rect -2498 307898 18986 308134
rect 19222 307898 54986 308134
rect 55222 307898 90986 308134
rect 91222 307898 126986 308134
rect 127222 307898 162986 308134
rect 163222 307898 198986 308134
rect 199222 307898 234986 308134
rect 235222 307898 270986 308134
rect 271222 307898 306986 308134
rect 307222 307898 342986 308134
rect 343222 307898 378986 308134
rect 379222 307898 414986 308134
rect 415222 307898 450986 308134
rect 451222 307898 486986 308134
rect 487222 307898 522986 308134
rect 523222 307898 558986 308134
rect 559222 307898 586422 308134
rect 586658 307898 586840 308134
rect -2916 307876 586840 307898
rect -2916 307874 -2316 307876
rect 18804 307874 19404 307876
rect 54804 307874 55404 307876
rect 90804 307874 91404 307876
rect 126804 307874 127404 307876
rect 162804 307874 163404 307876
rect 198804 307874 199404 307876
rect 234804 307874 235404 307876
rect 270804 307874 271404 307876
rect 306804 307874 307404 307876
rect 342804 307874 343404 307876
rect 378804 307874 379404 307876
rect 414804 307874 415404 307876
rect 450804 307874 451404 307876
rect 486804 307874 487404 307876
rect 522804 307874 523404 307876
rect 558804 307874 559404 307876
rect 586240 307874 586840 307876
rect -7516 301276 -6916 301278
rect 11604 301276 12204 301278
rect 47604 301276 48204 301278
rect 83604 301276 84204 301278
rect 119604 301276 120204 301278
rect 155604 301276 156204 301278
rect 191604 301276 192204 301278
rect 227604 301276 228204 301278
rect 263604 301276 264204 301278
rect 299604 301276 300204 301278
rect 335604 301276 336204 301278
rect 371604 301276 372204 301278
rect 407604 301276 408204 301278
rect 443604 301276 444204 301278
rect 479604 301276 480204 301278
rect 515604 301276 516204 301278
rect 551604 301276 552204 301278
rect 590840 301276 591440 301278
rect -8436 301254 592360 301276
rect -8436 301018 -7334 301254
rect -7098 301018 11786 301254
rect 12022 301018 47786 301254
rect 48022 301018 83786 301254
rect 84022 301018 119786 301254
rect 120022 301018 155786 301254
rect 156022 301018 191786 301254
rect 192022 301018 227786 301254
rect 228022 301018 263786 301254
rect 264022 301018 299786 301254
rect 300022 301018 335786 301254
rect 336022 301018 371786 301254
rect 372022 301018 407786 301254
rect 408022 301018 443786 301254
rect 444022 301018 479786 301254
rect 480022 301018 515786 301254
rect 516022 301018 551786 301254
rect 552022 301018 591022 301254
rect 591258 301018 592360 301254
rect -8436 300934 592360 301018
rect -8436 300698 -7334 300934
rect -7098 300698 11786 300934
rect 12022 300698 47786 300934
rect 48022 300698 83786 300934
rect 84022 300698 119786 300934
rect 120022 300698 155786 300934
rect 156022 300698 191786 300934
rect 192022 300698 227786 300934
rect 228022 300698 263786 300934
rect 264022 300698 299786 300934
rect 300022 300698 335786 300934
rect 336022 300698 371786 300934
rect 372022 300698 407786 300934
rect 408022 300698 443786 300934
rect 444022 300698 479786 300934
rect 480022 300698 515786 300934
rect 516022 300698 551786 300934
rect 552022 300698 591022 300934
rect 591258 300698 592360 300934
rect -8436 300676 592360 300698
rect -7516 300674 -6916 300676
rect 11604 300674 12204 300676
rect 47604 300674 48204 300676
rect 83604 300674 84204 300676
rect 119604 300674 120204 300676
rect 155604 300674 156204 300676
rect 191604 300674 192204 300676
rect 227604 300674 228204 300676
rect 263604 300674 264204 300676
rect 299604 300674 300204 300676
rect 335604 300674 336204 300676
rect 371604 300674 372204 300676
rect 407604 300674 408204 300676
rect 443604 300674 444204 300676
rect 479604 300674 480204 300676
rect 515604 300674 516204 300676
rect 551604 300674 552204 300676
rect 590840 300674 591440 300676
rect -5676 297676 -5076 297678
rect 8004 297676 8604 297678
rect 44004 297676 44604 297678
rect 80004 297676 80604 297678
rect 116004 297676 116604 297678
rect 152004 297676 152604 297678
rect 188004 297676 188604 297678
rect 224004 297676 224604 297678
rect 260004 297676 260604 297678
rect 296004 297676 296604 297678
rect 332004 297676 332604 297678
rect 368004 297676 368604 297678
rect 404004 297676 404604 297678
rect 440004 297676 440604 297678
rect 476004 297676 476604 297678
rect 512004 297676 512604 297678
rect 548004 297676 548604 297678
rect 589000 297676 589600 297678
rect -6596 297654 590520 297676
rect -6596 297418 -5494 297654
rect -5258 297418 8186 297654
rect 8422 297418 44186 297654
rect 44422 297418 80186 297654
rect 80422 297418 116186 297654
rect 116422 297418 152186 297654
rect 152422 297418 188186 297654
rect 188422 297418 224186 297654
rect 224422 297418 260186 297654
rect 260422 297418 296186 297654
rect 296422 297418 332186 297654
rect 332422 297418 368186 297654
rect 368422 297418 404186 297654
rect 404422 297418 440186 297654
rect 440422 297418 476186 297654
rect 476422 297418 512186 297654
rect 512422 297418 548186 297654
rect 548422 297418 589182 297654
rect 589418 297418 590520 297654
rect -6596 297334 590520 297418
rect -6596 297098 -5494 297334
rect -5258 297098 8186 297334
rect 8422 297098 44186 297334
rect 44422 297098 80186 297334
rect 80422 297098 116186 297334
rect 116422 297098 152186 297334
rect 152422 297098 188186 297334
rect 188422 297098 224186 297334
rect 224422 297098 260186 297334
rect 260422 297098 296186 297334
rect 296422 297098 332186 297334
rect 332422 297098 368186 297334
rect 368422 297098 404186 297334
rect 404422 297098 440186 297334
rect 440422 297098 476186 297334
rect 476422 297098 512186 297334
rect 512422 297098 548186 297334
rect 548422 297098 589182 297334
rect 589418 297098 590520 297334
rect -6596 297076 590520 297098
rect -5676 297074 -5076 297076
rect 8004 297074 8604 297076
rect 44004 297074 44604 297076
rect 80004 297074 80604 297076
rect 116004 297074 116604 297076
rect 152004 297074 152604 297076
rect 188004 297074 188604 297076
rect 224004 297074 224604 297076
rect 260004 297074 260604 297076
rect 296004 297074 296604 297076
rect 332004 297074 332604 297076
rect 368004 297074 368604 297076
rect 404004 297074 404604 297076
rect 440004 297074 440604 297076
rect 476004 297074 476604 297076
rect 512004 297074 512604 297076
rect 548004 297074 548604 297076
rect 589000 297074 589600 297076
rect -3836 294076 -3236 294078
rect 4404 294076 5004 294078
rect 40404 294076 41004 294078
rect 76404 294076 77004 294078
rect 112404 294076 113004 294078
rect 148404 294076 149004 294078
rect 184404 294076 185004 294078
rect 220404 294076 221004 294078
rect 256404 294076 257004 294078
rect 292404 294076 293004 294078
rect 328404 294076 329004 294078
rect 364404 294076 365004 294078
rect 400404 294076 401004 294078
rect 436404 294076 437004 294078
rect 472404 294076 473004 294078
rect 508404 294076 509004 294078
rect 544404 294076 545004 294078
rect 580404 294076 581004 294078
rect 587160 294076 587760 294078
rect -4756 294054 588680 294076
rect -4756 293818 -3654 294054
rect -3418 293818 4586 294054
rect 4822 293818 40586 294054
rect 40822 293818 76586 294054
rect 76822 293818 112586 294054
rect 112822 293818 148586 294054
rect 148822 293818 184586 294054
rect 184822 293818 220586 294054
rect 220822 293818 256586 294054
rect 256822 293818 292586 294054
rect 292822 293818 328586 294054
rect 328822 293818 364586 294054
rect 364822 293818 400586 294054
rect 400822 293818 436586 294054
rect 436822 293818 472586 294054
rect 472822 293818 508586 294054
rect 508822 293818 544586 294054
rect 544822 293818 580586 294054
rect 580822 293818 587342 294054
rect 587578 293818 588680 294054
rect -4756 293734 588680 293818
rect -4756 293498 -3654 293734
rect -3418 293498 4586 293734
rect 4822 293498 40586 293734
rect 40822 293498 76586 293734
rect 76822 293498 112586 293734
rect 112822 293498 148586 293734
rect 148822 293498 184586 293734
rect 184822 293498 220586 293734
rect 220822 293498 256586 293734
rect 256822 293498 292586 293734
rect 292822 293498 328586 293734
rect 328822 293498 364586 293734
rect 364822 293498 400586 293734
rect 400822 293498 436586 293734
rect 436822 293498 472586 293734
rect 472822 293498 508586 293734
rect 508822 293498 544586 293734
rect 544822 293498 580586 293734
rect 580822 293498 587342 293734
rect 587578 293498 588680 293734
rect -4756 293476 588680 293498
rect -3836 293474 -3236 293476
rect 4404 293474 5004 293476
rect 40404 293474 41004 293476
rect 76404 293474 77004 293476
rect 112404 293474 113004 293476
rect 148404 293474 149004 293476
rect 184404 293474 185004 293476
rect 220404 293474 221004 293476
rect 256404 293474 257004 293476
rect 292404 293474 293004 293476
rect 328404 293474 329004 293476
rect 364404 293474 365004 293476
rect 400404 293474 401004 293476
rect 436404 293474 437004 293476
rect 472404 293474 473004 293476
rect 508404 293474 509004 293476
rect 544404 293474 545004 293476
rect 580404 293474 581004 293476
rect 587160 293474 587760 293476
rect -1996 290476 -1396 290478
rect 804 290476 1404 290478
rect 36804 290476 37404 290478
rect 72804 290476 73404 290478
rect 108804 290476 109404 290478
rect 144804 290476 145404 290478
rect 180804 290476 181404 290478
rect 216804 290476 217404 290478
rect 252804 290476 253404 290478
rect 288804 290476 289404 290478
rect 324804 290476 325404 290478
rect 360804 290476 361404 290478
rect 396804 290476 397404 290478
rect 432804 290476 433404 290478
rect 468804 290476 469404 290478
rect 504804 290476 505404 290478
rect 540804 290476 541404 290478
rect 576804 290476 577404 290478
rect 585320 290476 585920 290478
rect -2916 290454 586840 290476
rect -2916 290218 -1814 290454
rect -1578 290218 986 290454
rect 1222 290218 36986 290454
rect 37222 290218 72986 290454
rect 73222 290218 108986 290454
rect 109222 290218 144986 290454
rect 145222 290218 180986 290454
rect 181222 290218 216986 290454
rect 217222 290218 252986 290454
rect 253222 290218 288986 290454
rect 289222 290218 324986 290454
rect 325222 290218 360986 290454
rect 361222 290218 396986 290454
rect 397222 290218 432986 290454
rect 433222 290218 468986 290454
rect 469222 290218 504986 290454
rect 505222 290218 540986 290454
rect 541222 290218 576986 290454
rect 577222 290218 585502 290454
rect 585738 290218 586840 290454
rect -2916 290134 586840 290218
rect -2916 289898 -1814 290134
rect -1578 289898 986 290134
rect 1222 289898 36986 290134
rect 37222 289898 72986 290134
rect 73222 289898 108986 290134
rect 109222 289898 144986 290134
rect 145222 289898 180986 290134
rect 181222 289898 216986 290134
rect 217222 289898 252986 290134
rect 253222 289898 288986 290134
rect 289222 289898 324986 290134
rect 325222 289898 360986 290134
rect 361222 289898 396986 290134
rect 397222 289898 432986 290134
rect 433222 289898 468986 290134
rect 469222 289898 504986 290134
rect 505222 289898 540986 290134
rect 541222 289898 576986 290134
rect 577222 289898 585502 290134
rect 585738 289898 586840 290134
rect -2916 289876 586840 289898
rect -1996 289874 -1396 289876
rect 804 289874 1404 289876
rect 36804 289874 37404 289876
rect 72804 289874 73404 289876
rect 108804 289874 109404 289876
rect 144804 289874 145404 289876
rect 180804 289874 181404 289876
rect 216804 289874 217404 289876
rect 252804 289874 253404 289876
rect 288804 289874 289404 289876
rect 324804 289874 325404 289876
rect 360804 289874 361404 289876
rect 396804 289874 397404 289876
rect 432804 289874 433404 289876
rect 468804 289874 469404 289876
rect 504804 289874 505404 289876
rect 540804 289874 541404 289876
rect 576804 289874 577404 289876
rect 585320 289874 585920 289876
rect -8436 283276 -7836 283278
rect 29604 283276 30204 283278
rect 65604 283276 66204 283278
rect 101604 283276 102204 283278
rect 137604 283276 138204 283278
rect 173604 283276 174204 283278
rect 209604 283276 210204 283278
rect 245604 283276 246204 283278
rect 281604 283276 282204 283278
rect 317604 283276 318204 283278
rect 353604 283276 354204 283278
rect 389604 283276 390204 283278
rect 425604 283276 426204 283278
rect 461604 283276 462204 283278
rect 497604 283276 498204 283278
rect 533604 283276 534204 283278
rect 569604 283276 570204 283278
rect 591760 283276 592360 283278
rect -8436 283254 592360 283276
rect -8436 283018 -8254 283254
rect -8018 283018 29786 283254
rect 30022 283018 65786 283254
rect 66022 283018 101786 283254
rect 102022 283018 137786 283254
rect 138022 283018 173786 283254
rect 174022 283018 209786 283254
rect 210022 283018 245786 283254
rect 246022 283018 281786 283254
rect 282022 283018 317786 283254
rect 318022 283018 353786 283254
rect 354022 283018 389786 283254
rect 390022 283018 425786 283254
rect 426022 283018 461786 283254
rect 462022 283018 497786 283254
rect 498022 283018 533786 283254
rect 534022 283018 569786 283254
rect 570022 283018 591942 283254
rect 592178 283018 592360 283254
rect -8436 282934 592360 283018
rect -8436 282698 -8254 282934
rect -8018 282698 29786 282934
rect 30022 282698 65786 282934
rect 66022 282698 101786 282934
rect 102022 282698 137786 282934
rect 138022 282698 173786 282934
rect 174022 282698 209786 282934
rect 210022 282698 245786 282934
rect 246022 282698 281786 282934
rect 282022 282698 317786 282934
rect 318022 282698 353786 282934
rect 354022 282698 389786 282934
rect 390022 282698 425786 282934
rect 426022 282698 461786 282934
rect 462022 282698 497786 282934
rect 498022 282698 533786 282934
rect 534022 282698 569786 282934
rect 570022 282698 591942 282934
rect 592178 282698 592360 282934
rect -8436 282676 592360 282698
rect -8436 282674 -7836 282676
rect 29604 282674 30204 282676
rect 65604 282674 66204 282676
rect 101604 282674 102204 282676
rect 137604 282674 138204 282676
rect 173604 282674 174204 282676
rect 209604 282674 210204 282676
rect 245604 282674 246204 282676
rect 281604 282674 282204 282676
rect 317604 282674 318204 282676
rect 353604 282674 354204 282676
rect 389604 282674 390204 282676
rect 425604 282674 426204 282676
rect 461604 282674 462204 282676
rect 497604 282674 498204 282676
rect 533604 282674 534204 282676
rect 569604 282674 570204 282676
rect 591760 282674 592360 282676
rect -6596 279676 -5996 279678
rect 26004 279676 26604 279678
rect 62004 279676 62604 279678
rect 98004 279676 98604 279678
rect 134004 279676 134604 279678
rect 170004 279676 170604 279678
rect 206004 279676 206604 279678
rect 242004 279676 242604 279678
rect 278004 279676 278604 279678
rect 314004 279676 314604 279678
rect 350004 279676 350604 279678
rect 386004 279676 386604 279678
rect 422004 279676 422604 279678
rect 458004 279676 458604 279678
rect 494004 279676 494604 279678
rect 530004 279676 530604 279678
rect 566004 279676 566604 279678
rect 589920 279676 590520 279678
rect -6596 279654 590520 279676
rect -6596 279418 -6414 279654
rect -6178 279418 26186 279654
rect 26422 279418 62186 279654
rect 62422 279418 98186 279654
rect 98422 279418 134186 279654
rect 134422 279418 170186 279654
rect 170422 279418 206186 279654
rect 206422 279418 242186 279654
rect 242422 279418 278186 279654
rect 278422 279418 314186 279654
rect 314422 279418 350186 279654
rect 350422 279418 386186 279654
rect 386422 279418 422186 279654
rect 422422 279418 458186 279654
rect 458422 279418 494186 279654
rect 494422 279418 530186 279654
rect 530422 279418 566186 279654
rect 566422 279418 590102 279654
rect 590338 279418 590520 279654
rect -6596 279334 590520 279418
rect -6596 279098 -6414 279334
rect -6178 279098 26186 279334
rect 26422 279098 62186 279334
rect 62422 279098 98186 279334
rect 98422 279098 134186 279334
rect 134422 279098 170186 279334
rect 170422 279098 206186 279334
rect 206422 279098 242186 279334
rect 242422 279098 278186 279334
rect 278422 279098 314186 279334
rect 314422 279098 350186 279334
rect 350422 279098 386186 279334
rect 386422 279098 422186 279334
rect 422422 279098 458186 279334
rect 458422 279098 494186 279334
rect 494422 279098 530186 279334
rect 530422 279098 566186 279334
rect 566422 279098 590102 279334
rect 590338 279098 590520 279334
rect -6596 279076 590520 279098
rect -6596 279074 -5996 279076
rect 26004 279074 26604 279076
rect 62004 279074 62604 279076
rect 98004 279074 98604 279076
rect 134004 279074 134604 279076
rect 170004 279074 170604 279076
rect 206004 279074 206604 279076
rect 242004 279074 242604 279076
rect 278004 279074 278604 279076
rect 314004 279074 314604 279076
rect 350004 279074 350604 279076
rect 386004 279074 386604 279076
rect 422004 279074 422604 279076
rect 458004 279074 458604 279076
rect 494004 279074 494604 279076
rect 530004 279074 530604 279076
rect 566004 279074 566604 279076
rect 589920 279074 590520 279076
rect -4756 276076 -4156 276078
rect 22404 276076 23004 276078
rect 58404 276076 59004 276078
rect 94404 276076 95004 276078
rect 130404 276076 131004 276078
rect 166404 276076 167004 276078
rect 202404 276076 203004 276078
rect 238404 276076 239004 276078
rect 274404 276076 275004 276078
rect 310404 276076 311004 276078
rect 346404 276076 347004 276078
rect 382404 276076 383004 276078
rect 418404 276076 419004 276078
rect 454404 276076 455004 276078
rect 490404 276076 491004 276078
rect 526404 276076 527004 276078
rect 562404 276076 563004 276078
rect 588080 276076 588680 276078
rect -4756 276054 588680 276076
rect -4756 275818 -4574 276054
rect -4338 275818 22586 276054
rect 22822 275818 58586 276054
rect 58822 275818 94586 276054
rect 94822 275818 130586 276054
rect 130822 275818 166586 276054
rect 166822 275818 202586 276054
rect 202822 275818 238586 276054
rect 238822 275818 274586 276054
rect 274822 275818 310586 276054
rect 310822 275818 346586 276054
rect 346822 275818 382586 276054
rect 382822 275818 418586 276054
rect 418822 275818 454586 276054
rect 454822 275818 490586 276054
rect 490822 275818 526586 276054
rect 526822 275818 562586 276054
rect 562822 275818 588262 276054
rect 588498 275818 588680 276054
rect -4756 275734 588680 275818
rect -4756 275498 -4574 275734
rect -4338 275498 22586 275734
rect 22822 275498 58586 275734
rect 58822 275498 94586 275734
rect 94822 275498 130586 275734
rect 130822 275498 166586 275734
rect 166822 275498 202586 275734
rect 202822 275498 238586 275734
rect 238822 275498 274586 275734
rect 274822 275498 310586 275734
rect 310822 275498 346586 275734
rect 346822 275498 382586 275734
rect 382822 275498 418586 275734
rect 418822 275498 454586 275734
rect 454822 275498 490586 275734
rect 490822 275498 526586 275734
rect 526822 275498 562586 275734
rect 562822 275498 588262 275734
rect 588498 275498 588680 275734
rect -4756 275476 588680 275498
rect -4756 275474 -4156 275476
rect 22404 275474 23004 275476
rect 58404 275474 59004 275476
rect 94404 275474 95004 275476
rect 130404 275474 131004 275476
rect 166404 275474 167004 275476
rect 202404 275474 203004 275476
rect 238404 275474 239004 275476
rect 274404 275474 275004 275476
rect 310404 275474 311004 275476
rect 346404 275474 347004 275476
rect 382404 275474 383004 275476
rect 418404 275474 419004 275476
rect 454404 275474 455004 275476
rect 490404 275474 491004 275476
rect 526404 275474 527004 275476
rect 562404 275474 563004 275476
rect 588080 275474 588680 275476
rect -2916 272476 -2316 272478
rect 18804 272476 19404 272478
rect 54804 272476 55404 272478
rect 90804 272476 91404 272478
rect 126804 272476 127404 272478
rect 162804 272476 163404 272478
rect 198804 272476 199404 272478
rect 234804 272476 235404 272478
rect 270804 272476 271404 272478
rect 306804 272476 307404 272478
rect 342804 272476 343404 272478
rect 378804 272476 379404 272478
rect 414804 272476 415404 272478
rect 450804 272476 451404 272478
rect 486804 272476 487404 272478
rect 522804 272476 523404 272478
rect 558804 272476 559404 272478
rect 586240 272476 586840 272478
rect -2916 272454 586840 272476
rect -2916 272218 -2734 272454
rect -2498 272218 18986 272454
rect 19222 272218 54986 272454
rect 55222 272218 90986 272454
rect 91222 272218 126986 272454
rect 127222 272218 162986 272454
rect 163222 272218 198986 272454
rect 199222 272218 234986 272454
rect 235222 272218 270986 272454
rect 271222 272218 306986 272454
rect 307222 272218 342986 272454
rect 343222 272218 378986 272454
rect 379222 272218 414986 272454
rect 415222 272218 450986 272454
rect 451222 272218 486986 272454
rect 487222 272218 522986 272454
rect 523222 272218 558986 272454
rect 559222 272218 586422 272454
rect 586658 272218 586840 272454
rect -2916 272134 586840 272218
rect -2916 271898 -2734 272134
rect -2498 271898 18986 272134
rect 19222 271898 54986 272134
rect 55222 271898 90986 272134
rect 91222 271898 126986 272134
rect 127222 271898 162986 272134
rect 163222 271898 198986 272134
rect 199222 271898 234986 272134
rect 235222 271898 270986 272134
rect 271222 271898 306986 272134
rect 307222 271898 342986 272134
rect 343222 271898 378986 272134
rect 379222 271898 414986 272134
rect 415222 271898 450986 272134
rect 451222 271898 486986 272134
rect 487222 271898 522986 272134
rect 523222 271898 558986 272134
rect 559222 271898 586422 272134
rect 586658 271898 586840 272134
rect -2916 271876 586840 271898
rect -2916 271874 -2316 271876
rect 18804 271874 19404 271876
rect 54804 271874 55404 271876
rect 90804 271874 91404 271876
rect 126804 271874 127404 271876
rect 162804 271874 163404 271876
rect 198804 271874 199404 271876
rect 234804 271874 235404 271876
rect 270804 271874 271404 271876
rect 306804 271874 307404 271876
rect 342804 271874 343404 271876
rect 378804 271874 379404 271876
rect 414804 271874 415404 271876
rect 450804 271874 451404 271876
rect 486804 271874 487404 271876
rect 522804 271874 523404 271876
rect 558804 271874 559404 271876
rect 586240 271874 586840 271876
rect -7516 265276 -6916 265278
rect 11604 265276 12204 265278
rect 47604 265276 48204 265278
rect 83604 265276 84204 265278
rect 119604 265276 120204 265278
rect 155604 265276 156204 265278
rect 191604 265276 192204 265278
rect 227604 265276 228204 265278
rect 263604 265276 264204 265278
rect 299604 265276 300204 265278
rect 335604 265276 336204 265278
rect 371604 265276 372204 265278
rect 407604 265276 408204 265278
rect 443604 265276 444204 265278
rect 479604 265276 480204 265278
rect 515604 265276 516204 265278
rect 551604 265276 552204 265278
rect 590840 265276 591440 265278
rect -8436 265254 592360 265276
rect -8436 265018 -7334 265254
rect -7098 265018 11786 265254
rect 12022 265018 47786 265254
rect 48022 265018 83786 265254
rect 84022 265018 119786 265254
rect 120022 265018 155786 265254
rect 156022 265018 191786 265254
rect 192022 265018 227786 265254
rect 228022 265018 263786 265254
rect 264022 265018 299786 265254
rect 300022 265018 335786 265254
rect 336022 265018 371786 265254
rect 372022 265018 407786 265254
rect 408022 265018 443786 265254
rect 444022 265018 479786 265254
rect 480022 265018 515786 265254
rect 516022 265018 551786 265254
rect 552022 265018 591022 265254
rect 591258 265018 592360 265254
rect -8436 264934 592360 265018
rect -8436 264698 -7334 264934
rect -7098 264698 11786 264934
rect 12022 264698 47786 264934
rect 48022 264698 83786 264934
rect 84022 264698 119786 264934
rect 120022 264698 155786 264934
rect 156022 264698 191786 264934
rect 192022 264698 227786 264934
rect 228022 264698 263786 264934
rect 264022 264698 299786 264934
rect 300022 264698 335786 264934
rect 336022 264698 371786 264934
rect 372022 264698 407786 264934
rect 408022 264698 443786 264934
rect 444022 264698 479786 264934
rect 480022 264698 515786 264934
rect 516022 264698 551786 264934
rect 552022 264698 591022 264934
rect 591258 264698 592360 264934
rect -8436 264676 592360 264698
rect -7516 264674 -6916 264676
rect 11604 264674 12204 264676
rect 47604 264674 48204 264676
rect 83604 264674 84204 264676
rect 119604 264674 120204 264676
rect 155604 264674 156204 264676
rect 191604 264674 192204 264676
rect 227604 264674 228204 264676
rect 263604 264674 264204 264676
rect 299604 264674 300204 264676
rect 335604 264674 336204 264676
rect 371604 264674 372204 264676
rect 407604 264674 408204 264676
rect 443604 264674 444204 264676
rect 479604 264674 480204 264676
rect 515604 264674 516204 264676
rect 551604 264674 552204 264676
rect 590840 264674 591440 264676
rect -5676 261676 -5076 261678
rect 8004 261676 8604 261678
rect 44004 261676 44604 261678
rect 80004 261676 80604 261678
rect 116004 261676 116604 261678
rect 152004 261676 152604 261678
rect 188004 261676 188604 261678
rect 224004 261676 224604 261678
rect 260004 261676 260604 261678
rect 296004 261676 296604 261678
rect 332004 261676 332604 261678
rect 368004 261676 368604 261678
rect 404004 261676 404604 261678
rect 440004 261676 440604 261678
rect 476004 261676 476604 261678
rect 512004 261676 512604 261678
rect 548004 261676 548604 261678
rect 589000 261676 589600 261678
rect -6596 261654 590520 261676
rect -6596 261418 -5494 261654
rect -5258 261418 8186 261654
rect 8422 261418 44186 261654
rect 44422 261418 80186 261654
rect 80422 261418 116186 261654
rect 116422 261418 152186 261654
rect 152422 261418 188186 261654
rect 188422 261418 224186 261654
rect 224422 261418 260186 261654
rect 260422 261418 296186 261654
rect 296422 261418 332186 261654
rect 332422 261418 368186 261654
rect 368422 261418 404186 261654
rect 404422 261418 440186 261654
rect 440422 261418 476186 261654
rect 476422 261418 512186 261654
rect 512422 261418 548186 261654
rect 548422 261418 589182 261654
rect 589418 261418 590520 261654
rect -6596 261334 590520 261418
rect -6596 261098 -5494 261334
rect -5258 261098 8186 261334
rect 8422 261098 44186 261334
rect 44422 261098 80186 261334
rect 80422 261098 116186 261334
rect 116422 261098 152186 261334
rect 152422 261098 188186 261334
rect 188422 261098 224186 261334
rect 224422 261098 260186 261334
rect 260422 261098 296186 261334
rect 296422 261098 332186 261334
rect 332422 261098 368186 261334
rect 368422 261098 404186 261334
rect 404422 261098 440186 261334
rect 440422 261098 476186 261334
rect 476422 261098 512186 261334
rect 512422 261098 548186 261334
rect 548422 261098 589182 261334
rect 589418 261098 590520 261334
rect -6596 261076 590520 261098
rect -5676 261074 -5076 261076
rect 8004 261074 8604 261076
rect 44004 261074 44604 261076
rect 80004 261074 80604 261076
rect 116004 261074 116604 261076
rect 152004 261074 152604 261076
rect 188004 261074 188604 261076
rect 224004 261074 224604 261076
rect 260004 261074 260604 261076
rect 296004 261074 296604 261076
rect 332004 261074 332604 261076
rect 368004 261074 368604 261076
rect 404004 261074 404604 261076
rect 440004 261074 440604 261076
rect 476004 261074 476604 261076
rect 512004 261074 512604 261076
rect 548004 261074 548604 261076
rect 589000 261074 589600 261076
rect -3836 258076 -3236 258078
rect 4404 258076 5004 258078
rect 40404 258076 41004 258078
rect 76404 258076 77004 258078
rect 112404 258076 113004 258078
rect 148404 258076 149004 258078
rect 184404 258076 185004 258078
rect 220404 258076 221004 258078
rect 256404 258076 257004 258078
rect 292404 258076 293004 258078
rect 328404 258076 329004 258078
rect 364404 258076 365004 258078
rect 400404 258076 401004 258078
rect 436404 258076 437004 258078
rect 472404 258076 473004 258078
rect 508404 258076 509004 258078
rect 544404 258076 545004 258078
rect 580404 258076 581004 258078
rect 587160 258076 587760 258078
rect -4756 258054 588680 258076
rect -4756 257818 -3654 258054
rect -3418 257818 4586 258054
rect 4822 257818 40586 258054
rect 40822 257818 76586 258054
rect 76822 257818 112586 258054
rect 112822 257818 148586 258054
rect 148822 257818 184586 258054
rect 184822 257818 220586 258054
rect 220822 257818 256586 258054
rect 256822 257818 292586 258054
rect 292822 257818 328586 258054
rect 328822 257818 364586 258054
rect 364822 257818 400586 258054
rect 400822 257818 436586 258054
rect 436822 257818 472586 258054
rect 472822 257818 508586 258054
rect 508822 257818 544586 258054
rect 544822 257818 580586 258054
rect 580822 257818 587342 258054
rect 587578 257818 588680 258054
rect -4756 257734 588680 257818
rect -4756 257498 -3654 257734
rect -3418 257498 4586 257734
rect 4822 257498 40586 257734
rect 40822 257498 76586 257734
rect 76822 257498 112586 257734
rect 112822 257498 148586 257734
rect 148822 257498 184586 257734
rect 184822 257498 220586 257734
rect 220822 257498 256586 257734
rect 256822 257498 292586 257734
rect 292822 257498 328586 257734
rect 328822 257498 364586 257734
rect 364822 257498 400586 257734
rect 400822 257498 436586 257734
rect 436822 257498 472586 257734
rect 472822 257498 508586 257734
rect 508822 257498 544586 257734
rect 544822 257498 580586 257734
rect 580822 257498 587342 257734
rect 587578 257498 588680 257734
rect -4756 257476 588680 257498
rect -3836 257474 -3236 257476
rect 4404 257474 5004 257476
rect 40404 257474 41004 257476
rect 76404 257474 77004 257476
rect 112404 257474 113004 257476
rect 148404 257474 149004 257476
rect 184404 257474 185004 257476
rect 220404 257474 221004 257476
rect 256404 257474 257004 257476
rect 292404 257474 293004 257476
rect 328404 257474 329004 257476
rect 364404 257474 365004 257476
rect 400404 257474 401004 257476
rect 436404 257474 437004 257476
rect 472404 257474 473004 257476
rect 508404 257474 509004 257476
rect 544404 257474 545004 257476
rect 580404 257474 581004 257476
rect 587160 257474 587760 257476
rect -1996 254476 -1396 254478
rect 804 254476 1404 254478
rect 36804 254476 37404 254478
rect 72804 254476 73404 254478
rect 108804 254476 109404 254478
rect 144804 254476 145404 254478
rect 180804 254476 181404 254478
rect 216804 254476 217404 254478
rect 252804 254476 253404 254478
rect 288804 254476 289404 254478
rect 324804 254476 325404 254478
rect 360804 254476 361404 254478
rect 396804 254476 397404 254478
rect 432804 254476 433404 254478
rect 468804 254476 469404 254478
rect 504804 254476 505404 254478
rect 540804 254476 541404 254478
rect 576804 254476 577404 254478
rect 585320 254476 585920 254478
rect -2916 254454 586840 254476
rect -2916 254218 -1814 254454
rect -1578 254218 986 254454
rect 1222 254218 36986 254454
rect 37222 254218 72986 254454
rect 73222 254218 108986 254454
rect 109222 254218 144986 254454
rect 145222 254218 180986 254454
rect 181222 254218 216986 254454
rect 217222 254218 252986 254454
rect 253222 254218 288986 254454
rect 289222 254218 324986 254454
rect 325222 254218 360986 254454
rect 361222 254218 396986 254454
rect 397222 254218 432986 254454
rect 433222 254218 468986 254454
rect 469222 254218 504986 254454
rect 505222 254218 540986 254454
rect 541222 254218 576986 254454
rect 577222 254218 585502 254454
rect 585738 254218 586840 254454
rect -2916 254134 586840 254218
rect -2916 253898 -1814 254134
rect -1578 253898 986 254134
rect 1222 253898 36986 254134
rect 37222 253898 72986 254134
rect 73222 253898 108986 254134
rect 109222 253898 144986 254134
rect 145222 253898 180986 254134
rect 181222 253898 216986 254134
rect 217222 253898 252986 254134
rect 253222 253898 288986 254134
rect 289222 253898 324986 254134
rect 325222 253898 360986 254134
rect 361222 253898 396986 254134
rect 397222 253898 432986 254134
rect 433222 253898 468986 254134
rect 469222 253898 504986 254134
rect 505222 253898 540986 254134
rect 541222 253898 576986 254134
rect 577222 253898 585502 254134
rect 585738 253898 586840 254134
rect -2916 253876 586840 253898
rect -1996 253874 -1396 253876
rect 804 253874 1404 253876
rect 36804 253874 37404 253876
rect 72804 253874 73404 253876
rect 108804 253874 109404 253876
rect 144804 253874 145404 253876
rect 180804 253874 181404 253876
rect 216804 253874 217404 253876
rect 252804 253874 253404 253876
rect 288804 253874 289404 253876
rect 324804 253874 325404 253876
rect 360804 253874 361404 253876
rect 396804 253874 397404 253876
rect 432804 253874 433404 253876
rect 468804 253874 469404 253876
rect 504804 253874 505404 253876
rect 540804 253874 541404 253876
rect 576804 253874 577404 253876
rect 585320 253874 585920 253876
rect -8436 247276 -7836 247278
rect 29604 247276 30204 247278
rect 65604 247276 66204 247278
rect 101604 247276 102204 247278
rect 137604 247276 138204 247278
rect 173604 247276 174204 247278
rect 209604 247276 210204 247278
rect 245604 247276 246204 247278
rect 281604 247276 282204 247278
rect 317604 247276 318204 247278
rect 353604 247276 354204 247278
rect 389604 247276 390204 247278
rect 425604 247276 426204 247278
rect 461604 247276 462204 247278
rect 497604 247276 498204 247278
rect 533604 247276 534204 247278
rect 569604 247276 570204 247278
rect 591760 247276 592360 247278
rect -8436 247254 592360 247276
rect -8436 247018 -8254 247254
rect -8018 247018 29786 247254
rect 30022 247018 65786 247254
rect 66022 247018 101786 247254
rect 102022 247018 137786 247254
rect 138022 247018 173786 247254
rect 174022 247018 209786 247254
rect 210022 247018 245786 247254
rect 246022 247018 281786 247254
rect 282022 247018 317786 247254
rect 318022 247018 353786 247254
rect 354022 247018 389786 247254
rect 390022 247018 425786 247254
rect 426022 247018 461786 247254
rect 462022 247018 497786 247254
rect 498022 247018 533786 247254
rect 534022 247018 569786 247254
rect 570022 247018 591942 247254
rect 592178 247018 592360 247254
rect -8436 246934 592360 247018
rect -8436 246698 -8254 246934
rect -8018 246698 29786 246934
rect 30022 246698 65786 246934
rect 66022 246698 101786 246934
rect 102022 246698 137786 246934
rect 138022 246698 173786 246934
rect 174022 246698 209786 246934
rect 210022 246698 245786 246934
rect 246022 246698 281786 246934
rect 282022 246698 317786 246934
rect 318022 246698 353786 246934
rect 354022 246698 389786 246934
rect 390022 246698 425786 246934
rect 426022 246698 461786 246934
rect 462022 246698 497786 246934
rect 498022 246698 533786 246934
rect 534022 246698 569786 246934
rect 570022 246698 591942 246934
rect 592178 246698 592360 246934
rect -8436 246676 592360 246698
rect -8436 246674 -7836 246676
rect 29604 246674 30204 246676
rect 65604 246674 66204 246676
rect 101604 246674 102204 246676
rect 137604 246674 138204 246676
rect 173604 246674 174204 246676
rect 209604 246674 210204 246676
rect 245604 246674 246204 246676
rect 281604 246674 282204 246676
rect 317604 246674 318204 246676
rect 353604 246674 354204 246676
rect 389604 246674 390204 246676
rect 425604 246674 426204 246676
rect 461604 246674 462204 246676
rect 497604 246674 498204 246676
rect 533604 246674 534204 246676
rect 569604 246674 570204 246676
rect 591760 246674 592360 246676
rect -6596 243676 -5996 243678
rect 26004 243676 26604 243678
rect 62004 243676 62604 243678
rect 98004 243676 98604 243678
rect 134004 243676 134604 243678
rect 170004 243676 170604 243678
rect 206004 243676 206604 243678
rect 242004 243676 242604 243678
rect 278004 243676 278604 243678
rect 314004 243676 314604 243678
rect 350004 243676 350604 243678
rect 386004 243676 386604 243678
rect 422004 243676 422604 243678
rect 458004 243676 458604 243678
rect 494004 243676 494604 243678
rect 530004 243676 530604 243678
rect 566004 243676 566604 243678
rect 589920 243676 590520 243678
rect -6596 243654 590520 243676
rect -6596 243418 -6414 243654
rect -6178 243418 26186 243654
rect 26422 243418 62186 243654
rect 62422 243418 98186 243654
rect 98422 243418 134186 243654
rect 134422 243418 170186 243654
rect 170422 243418 206186 243654
rect 206422 243418 242186 243654
rect 242422 243418 278186 243654
rect 278422 243418 314186 243654
rect 314422 243418 350186 243654
rect 350422 243418 386186 243654
rect 386422 243418 422186 243654
rect 422422 243418 458186 243654
rect 458422 243418 494186 243654
rect 494422 243418 530186 243654
rect 530422 243418 566186 243654
rect 566422 243418 590102 243654
rect 590338 243418 590520 243654
rect -6596 243334 590520 243418
rect -6596 243098 -6414 243334
rect -6178 243098 26186 243334
rect 26422 243098 62186 243334
rect 62422 243098 98186 243334
rect 98422 243098 134186 243334
rect 134422 243098 170186 243334
rect 170422 243098 206186 243334
rect 206422 243098 242186 243334
rect 242422 243098 278186 243334
rect 278422 243098 314186 243334
rect 314422 243098 350186 243334
rect 350422 243098 386186 243334
rect 386422 243098 422186 243334
rect 422422 243098 458186 243334
rect 458422 243098 494186 243334
rect 494422 243098 530186 243334
rect 530422 243098 566186 243334
rect 566422 243098 590102 243334
rect 590338 243098 590520 243334
rect -6596 243076 590520 243098
rect -6596 243074 -5996 243076
rect 26004 243074 26604 243076
rect 62004 243074 62604 243076
rect 98004 243074 98604 243076
rect 134004 243074 134604 243076
rect 170004 243074 170604 243076
rect 206004 243074 206604 243076
rect 242004 243074 242604 243076
rect 278004 243074 278604 243076
rect 314004 243074 314604 243076
rect 350004 243074 350604 243076
rect 386004 243074 386604 243076
rect 422004 243074 422604 243076
rect 458004 243074 458604 243076
rect 494004 243074 494604 243076
rect 530004 243074 530604 243076
rect 566004 243074 566604 243076
rect 589920 243074 590520 243076
rect -4756 240076 -4156 240078
rect 22404 240076 23004 240078
rect 58404 240076 59004 240078
rect 94404 240076 95004 240078
rect 130404 240076 131004 240078
rect 166404 240076 167004 240078
rect 202404 240076 203004 240078
rect 238404 240076 239004 240078
rect 274404 240076 275004 240078
rect 310404 240076 311004 240078
rect 346404 240076 347004 240078
rect 382404 240076 383004 240078
rect 418404 240076 419004 240078
rect 454404 240076 455004 240078
rect 490404 240076 491004 240078
rect 526404 240076 527004 240078
rect 562404 240076 563004 240078
rect 588080 240076 588680 240078
rect -4756 240054 588680 240076
rect -4756 239818 -4574 240054
rect -4338 239818 22586 240054
rect 22822 239818 58586 240054
rect 58822 239818 94586 240054
rect 94822 239818 130586 240054
rect 130822 239818 166586 240054
rect 166822 239818 202586 240054
rect 202822 239818 238586 240054
rect 238822 239818 274586 240054
rect 274822 239818 310586 240054
rect 310822 239818 346586 240054
rect 346822 239818 382586 240054
rect 382822 239818 418586 240054
rect 418822 239818 454586 240054
rect 454822 239818 490586 240054
rect 490822 239818 526586 240054
rect 526822 239818 562586 240054
rect 562822 239818 588262 240054
rect 588498 239818 588680 240054
rect -4756 239734 588680 239818
rect -4756 239498 -4574 239734
rect -4338 239498 22586 239734
rect 22822 239498 58586 239734
rect 58822 239498 94586 239734
rect 94822 239498 130586 239734
rect 130822 239498 166586 239734
rect 166822 239498 202586 239734
rect 202822 239498 238586 239734
rect 238822 239498 274586 239734
rect 274822 239498 310586 239734
rect 310822 239498 346586 239734
rect 346822 239498 382586 239734
rect 382822 239498 418586 239734
rect 418822 239498 454586 239734
rect 454822 239498 490586 239734
rect 490822 239498 526586 239734
rect 526822 239498 562586 239734
rect 562822 239498 588262 239734
rect 588498 239498 588680 239734
rect -4756 239476 588680 239498
rect -4756 239474 -4156 239476
rect 22404 239474 23004 239476
rect 58404 239474 59004 239476
rect 94404 239474 95004 239476
rect 130404 239474 131004 239476
rect 166404 239474 167004 239476
rect 202404 239474 203004 239476
rect 238404 239474 239004 239476
rect 274404 239474 275004 239476
rect 310404 239474 311004 239476
rect 346404 239474 347004 239476
rect 382404 239474 383004 239476
rect 418404 239474 419004 239476
rect 454404 239474 455004 239476
rect 490404 239474 491004 239476
rect 526404 239474 527004 239476
rect 562404 239474 563004 239476
rect 588080 239474 588680 239476
rect -2916 236476 -2316 236478
rect 18804 236476 19404 236478
rect 54804 236476 55404 236478
rect 90804 236476 91404 236478
rect 126804 236476 127404 236478
rect 162804 236476 163404 236478
rect 198804 236476 199404 236478
rect 234804 236476 235404 236478
rect 270804 236476 271404 236478
rect 306804 236476 307404 236478
rect 342804 236476 343404 236478
rect 378804 236476 379404 236478
rect 414804 236476 415404 236478
rect 450804 236476 451404 236478
rect 486804 236476 487404 236478
rect 522804 236476 523404 236478
rect 558804 236476 559404 236478
rect 586240 236476 586840 236478
rect -2916 236454 586840 236476
rect -2916 236218 -2734 236454
rect -2498 236218 18986 236454
rect 19222 236218 54986 236454
rect 55222 236218 90986 236454
rect 91222 236218 126986 236454
rect 127222 236218 162986 236454
rect 163222 236218 198986 236454
rect 199222 236218 234986 236454
rect 235222 236218 270986 236454
rect 271222 236218 306986 236454
rect 307222 236218 342986 236454
rect 343222 236218 378986 236454
rect 379222 236218 414986 236454
rect 415222 236218 450986 236454
rect 451222 236218 486986 236454
rect 487222 236218 522986 236454
rect 523222 236218 558986 236454
rect 559222 236218 586422 236454
rect 586658 236218 586840 236454
rect -2916 236134 586840 236218
rect -2916 235898 -2734 236134
rect -2498 235898 18986 236134
rect 19222 235898 54986 236134
rect 55222 235898 90986 236134
rect 91222 235898 126986 236134
rect 127222 235898 162986 236134
rect 163222 235898 198986 236134
rect 199222 235898 234986 236134
rect 235222 235898 270986 236134
rect 271222 235898 306986 236134
rect 307222 235898 342986 236134
rect 343222 235898 378986 236134
rect 379222 235898 414986 236134
rect 415222 235898 450986 236134
rect 451222 235898 486986 236134
rect 487222 235898 522986 236134
rect 523222 235898 558986 236134
rect 559222 235898 586422 236134
rect 586658 235898 586840 236134
rect -2916 235876 586840 235898
rect -2916 235874 -2316 235876
rect 18804 235874 19404 235876
rect 54804 235874 55404 235876
rect 90804 235874 91404 235876
rect 126804 235874 127404 235876
rect 162804 235874 163404 235876
rect 198804 235874 199404 235876
rect 234804 235874 235404 235876
rect 270804 235874 271404 235876
rect 306804 235874 307404 235876
rect 342804 235874 343404 235876
rect 378804 235874 379404 235876
rect 414804 235874 415404 235876
rect 450804 235874 451404 235876
rect 486804 235874 487404 235876
rect 522804 235874 523404 235876
rect 558804 235874 559404 235876
rect 586240 235874 586840 235876
rect -7516 229276 -6916 229278
rect 11604 229276 12204 229278
rect 47604 229276 48204 229278
rect 83604 229276 84204 229278
rect 119604 229276 120204 229278
rect 155604 229276 156204 229278
rect 191604 229276 192204 229278
rect 227604 229276 228204 229278
rect 263604 229276 264204 229278
rect 299604 229276 300204 229278
rect 335604 229276 336204 229278
rect 371604 229276 372204 229278
rect 407604 229276 408204 229278
rect 443604 229276 444204 229278
rect 479604 229276 480204 229278
rect 515604 229276 516204 229278
rect 551604 229276 552204 229278
rect 590840 229276 591440 229278
rect -8436 229254 592360 229276
rect -8436 229018 -7334 229254
rect -7098 229018 11786 229254
rect 12022 229018 47786 229254
rect 48022 229018 83786 229254
rect 84022 229018 119786 229254
rect 120022 229018 155786 229254
rect 156022 229018 191786 229254
rect 192022 229018 227786 229254
rect 228022 229018 263786 229254
rect 264022 229018 299786 229254
rect 300022 229018 335786 229254
rect 336022 229018 371786 229254
rect 372022 229018 407786 229254
rect 408022 229018 443786 229254
rect 444022 229018 479786 229254
rect 480022 229018 515786 229254
rect 516022 229018 551786 229254
rect 552022 229018 591022 229254
rect 591258 229018 592360 229254
rect -8436 228934 592360 229018
rect -8436 228698 -7334 228934
rect -7098 228698 11786 228934
rect 12022 228698 47786 228934
rect 48022 228698 83786 228934
rect 84022 228698 119786 228934
rect 120022 228698 155786 228934
rect 156022 228698 191786 228934
rect 192022 228698 227786 228934
rect 228022 228698 263786 228934
rect 264022 228698 299786 228934
rect 300022 228698 335786 228934
rect 336022 228698 371786 228934
rect 372022 228698 407786 228934
rect 408022 228698 443786 228934
rect 444022 228698 479786 228934
rect 480022 228698 515786 228934
rect 516022 228698 551786 228934
rect 552022 228698 591022 228934
rect 591258 228698 592360 228934
rect -8436 228676 592360 228698
rect -7516 228674 -6916 228676
rect 11604 228674 12204 228676
rect 47604 228674 48204 228676
rect 83604 228674 84204 228676
rect 119604 228674 120204 228676
rect 155604 228674 156204 228676
rect 191604 228674 192204 228676
rect 227604 228674 228204 228676
rect 263604 228674 264204 228676
rect 299604 228674 300204 228676
rect 335604 228674 336204 228676
rect 371604 228674 372204 228676
rect 407604 228674 408204 228676
rect 443604 228674 444204 228676
rect 479604 228674 480204 228676
rect 515604 228674 516204 228676
rect 551604 228674 552204 228676
rect 590840 228674 591440 228676
rect -5676 225676 -5076 225678
rect 8004 225676 8604 225678
rect 44004 225676 44604 225678
rect 80004 225676 80604 225678
rect 116004 225676 116604 225678
rect 152004 225676 152604 225678
rect 188004 225676 188604 225678
rect 224004 225676 224604 225678
rect 260004 225676 260604 225678
rect 296004 225676 296604 225678
rect 332004 225676 332604 225678
rect 368004 225676 368604 225678
rect 404004 225676 404604 225678
rect 440004 225676 440604 225678
rect 476004 225676 476604 225678
rect 512004 225676 512604 225678
rect 548004 225676 548604 225678
rect 589000 225676 589600 225678
rect -6596 225654 590520 225676
rect -6596 225418 -5494 225654
rect -5258 225418 8186 225654
rect 8422 225418 44186 225654
rect 44422 225418 80186 225654
rect 80422 225418 116186 225654
rect 116422 225418 152186 225654
rect 152422 225418 188186 225654
rect 188422 225418 224186 225654
rect 224422 225418 260186 225654
rect 260422 225418 296186 225654
rect 296422 225418 332186 225654
rect 332422 225418 368186 225654
rect 368422 225418 404186 225654
rect 404422 225418 440186 225654
rect 440422 225418 476186 225654
rect 476422 225418 512186 225654
rect 512422 225418 548186 225654
rect 548422 225418 589182 225654
rect 589418 225418 590520 225654
rect -6596 225334 590520 225418
rect -6596 225098 -5494 225334
rect -5258 225098 8186 225334
rect 8422 225098 44186 225334
rect 44422 225098 80186 225334
rect 80422 225098 116186 225334
rect 116422 225098 152186 225334
rect 152422 225098 188186 225334
rect 188422 225098 224186 225334
rect 224422 225098 260186 225334
rect 260422 225098 296186 225334
rect 296422 225098 332186 225334
rect 332422 225098 368186 225334
rect 368422 225098 404186 225334
rect 404422 225098 440186 225334
rect 440422 225098 476186 225334
rect 476422 225098 512186 225334
rect 512422 225098 548186 225334
rect 548422 225098 589182 225334
rect 589418 225098 590520 225334
rect -6596 225076 590520 225098
rect -5676 225074 -5076 225076
rect 8004 225074 8604 225076
rect 44004 225074 44604 225076
rect 80004 225074 80604 225076
rect 116004 225074 116604 225076
rect 152004 225074 152604 225076
rect 188004 225074 188604 225076
rect 224004 225074 224604 225076
rect 260004 225074 260604 225076
rect 296004 225074 296604 225076
rect 332004 225074 332604 225076
rect 368004 225074 368604 225076
rect 404004 225074 404604 225076
rect 440004 225074 440604 225076
rect 476004 225074 476604 225076
rect 512004 225074 512604 225076
rect 548004 225074 548604 225076
rect 589000 225074 589600 225076
rect -3836 222076 -3236 222078
rect 4404 222076 5004 222078
rect 40404 222076 41004 222078
rect 76404 222076 77004 222078
rect 112404 222076 113004 222078
rect 148404 222076 149004 222078
rect 184404 222076 185004 222078
rect 220404 222076 221004 222078
rect 256404 222076 257004 222078
rect 292404 222076 293004 222078
rect 328404 222076 329004 222078
rect 364404 222076 365004 222078
rect 400404 222076 401004 222078
rect 436404 222076 437004 222078
rect 472404 222076 473004 222078
rect 508404 222076 509004 222078
rect 544404 222076 545004 222078
rect 580404 222076 581004 222078
rect 587160 222076 587760 222078
rect -4756 222054 588680 222076
rect -4756 221818 -3654 222054
rect -3418 221818 4586 222054
rect 4822 221818 40586 222054
rect 40822 221818 76586 222054
rect 76822 221818 112586 222054
rect 112822 221818 148586 222054
rect 148822 221818 184586 222054
rect 184822 221818 220586 222054
rect 220822 221818 256586 222054
rect 256822 221818 292586 222054
rect 292822 221818 328586 222054
rect 328822 221818 364586 222054
rect 364822 221818 400586 222054
rect 400822 221818 436586 222054
rect 436822 221818 472586 222054
rect 472822 221818 508586 222054
rect 508822 221818 544586 222054
rect 544822 221818 580586 222054
rect 580822 221818 587342 222054
rect 587578 221818 588680 222054
rect -4756 221734 588680 221818
rect -4756 221498 -3654 221734
rect -3418 221498 4586 221734
rect 4822 221498 40586 221734
rect 40822 221498 76586 221734
rect 76822 221498 112586 221734
rect 112822 221498 148586 221734
rect 148822 221498 184586 221734
rect 184822 221498 220586 221734
rect 220822 221498 256586 221734
rect 256822 221498 292586 221734
rect 292822 221498 328586 221734
rect 328822 221498 364586 221734
rect 364822 221498 400586 221734
rect 400822 221498 436586 221734
rect 436822 221498 472586 221734
rect 472822 221498 508586 221734
rect 508822 221498 544586 221734
rect 544822 221498 580586 221734
rect 580822 221498 587342 221734
rect 587578 221498 588680 221734
rect -4756 221476 588680 221498
rect -3836 221474 -3236 221476
rect 4404 221474 5004 221476
rect 40404 221474 41004 221476
rect 76404 221474 77004 221476
rect 112404 221474 113004 221476
rect 148404 221474 149004 221476
rect 184404 221474 185004 221476
rect 220404 221474 221004 221476
rect 256404 221474 257004 221476
rect 292404 221474 293004 221476
rect 328404 221474 329004 221476
rect 364404 221474 365004 221476
rect 400404 221474 401004 221476
rect 436404 221474 437004 221476
rect 472404 221474 473004 221476
rect 508404 221474 509004 221476
rect 544404 221474 545004 221476
rect 580404 221474 581004 221476
rect 587160 221474 587760 221476
rect -1996 218476 -1396 218478
rect 804 218476 1404 218478
rect 36804 218476 37404 218478
rect 72804 218476 73404 218478
rect 108804 218476 109404 218478
rect 144804 218476 145404 218478
rect 180804 218476 181404 218478
rect 216804 218476 217404 218478
rect 252804 218476 253404 218478
rect 288804 218476 289404 218478
rect 324804 218476 325404 218478
rect 360804 218476 361404 218478
rect 396804 218476 397404 218478
rect 432804 218476 433404 218478
rect 468804 218476 469404 218478
rect 504804 218476 505404 218478
rect 540804 218476 541404 218478
rect 576804 218476 577404 218478
rect 585320 218476 585920 218478
rect -2916 218454 586840 218476
rect -2916 218218 -1814 218454
rect -1578 218218 986 218454
rect 1222 218218 36986 218454
rect 37222 218218 72986 218454
rect 73222 218218 108986 218454
rect 109222 218218 144986 218454
rect 145222 218218 180986 218454
rect 181222 218218 216986 218454
rect 217222 218218 252986 218454
rect 253222 218218 288986 218454
rect 289222 218218 324986 218454
rect 325222 218218 360986 218454
rect 361222 218218 396986 218454
rect 397222 218218 432986 218454
rect 433222 218218 468986 218454
rect 469222 218218 504986 218454
rect 505222 218218 540986 218454
rect 541222 218218 576986 218454
rect 577222 218218 585502 218454
rect 585738 218218 586840 218454
rect -2916 218134 586840 218218
rect -2916 217898 -1814 218134
rect -1578 217898 986 218134
rect 1222 217898 36986 218134
rect 37222 217898 72986 218134
rect 73222 217898 108986 218134
rect 109222 217898 144986 218134
rect 145222 217898 180986 218134
rect 181222 217898 216986 218134
rect 217222 217898 252986 218134
rect 253222 217898 288986 218134
rect 289222 217898 324986 218134
rect 325222 217898 360986 218134
rect 361222 217898 396986 218134
rect 397222 217898 432986 218134
rect 433222 217898 468986 218134
rect 469222 217898 504986 218134
rect 505222 217898 540986 218134
rect 541222 217898 576986 218134
rect 577222 217898 585502 218134
rect 585738 217898 586840 218134
rect -2916 217876 586840 217898
rect -1996 217874 -1396 217876
rect 804 217874 1404 217876
rect 36804 217874 37404 217876
rect 72804 217874 73404 217876
rect 108804 217874 109404 217876
rect 144804 217874 145404 217876
rect 180804 217874 181404 217876
rect 216804 217874 217404 217876
rect 252804 217874 253404 217876
rect 288804 217874 289404 217876
rect 324804 217874 325404 217876
rect 360804 217874 361404 217876
rect 396804 217874 397404 217876
rect 432804 217874 433404 217876
rect 468804 217874 469404 217876
rect 504804 217874 505404 217876
rect 540804 217874 541404 217876
rect 576804 217874 577404 217876
rect 585320 217874 585920 217876
rect -8436 211276 -7836 211278
rect 29604 211276 30204 211278
rect 65604 211276 66204 211278
rect 101604 211276 102204 211278
rect 137604 211276 138204 211278
rect 173604 211276 174204 211278
rect 209604 211276 210204 211278
rect 245604 211276 246204 211278
rect 281604 211276 282204 211278
rect 317604 211276 318204 211278
rect 353604 211276 354204 211278
rect 389604 211276 390204 211278
rect 425604 211276 426204 211278
rect 461604 211276 462204 211278
rect 497604 211276 498204 211278
rect 533604 211276 534204 211278
rect 569604 211276 570204 211278
rect 591760 211276 592360 211278
rect -8436 211254 592360 211276
rect -8436 211018 -8254 211254
rect -8018 211018 29786 211254
rect 30022 211018 65786 211254
rect 66022 211018 101786 211254
rect 102022 211018 137786 211254
rect 138022 211018 173786 211254
rect 174022 211018 209786 211254
rect 210022 211018 245786 211254
rect 246022 211018 281786 211254
rect 282022 211018 317786 211254
rect 318022 211018 353786 211254
rect 354022 211018 389786 211254
rect 390022 211018 425786 211254
rect 426022 211018 461786 211254
rect 462022 211018 497786 211254
rect 498022 211018 533786 211254
rect 534022 211018 569786 211254
rect 570022 211018 591942 211254
rect 592178 211018 592360 211254
rect -8436 210934 592360 211018
rect -8436 210698 -8254 210934
rect -8018 210698 29786 210934
rect 30022 210698 65786 210934
rect 66022 210698 101786 210934
rect 102022 210698 137786 210934
rect 138022 210698 173786 210934
rect 174022 210698 209786 210934
rect 210022 210698 245786 210934
rect 246022 210698 281786 210934
rect 282022 210698 317786 210934
rect 318022 210698 353786 210934
rect 354022 210698 389786 210934
rect 390022 210698 425786 210934
rect 426022 210698 461786 210934
rect 462022 210698 497786 210934
rect 498022 210698 533786 210934
rect 534022 210698 569786 210934
rect 570022 210698 591942 210934
rect 592178 210698 592360 210934
rect -8436 210676 592360 210698
rect -8436 210674 -7836 210676
rect 29604 210674 30204 210676
rect 65604 210674 66204 210676
rect 101604 210674 102204 210676
rect 137604 210674 138204 210676
rect 173604 210674 174204 210676
rect 209604 210674 210204 210676
rect 245604 210674 246204 210676
rect 281604 210674 282204 210676
rect 317604 210674 318204 210676
rect 353604 210674 354204 210676
rect 389604 210674 390204 210676
rect 425604 210674 426204 210676
rect 461604 210674 462204 210676
rect 497604 210674 498204 210676
rect 533604 210674 534204 210676
rect 569604 210674 570204 210676
rect 591760 210674 592360 210676
rect -6596 207676 -5996 207678
rect 26004 207676 26604 207678
rect 62004 207676 62604 207678
rect 98004 207676 98604 207678
rect 134004 207676 134604 207678
rect 170004 207676 170604 207678
rect 206004 207676 206604 207678
rect 242004 207676 242604 207678
rect 278004 207676 278604 207678
rect 314004 207676 314604 207678
rect 350004 207676 350604 207678
rect 386004 207676 386604 207678
rect 422004 207676 422604 207678
rect 458004 207676 458604 207678
rect 494004 207676 494604 207678
rect 530004 207676 530604 207678
rect 566004 207676 566604 207678
rect 589920 207676 590520 207678
rect -6596 207654 590520 207676
rect -6596 207418 -6414 207654
rect -6178 207418 26186 207654
rect 26422 207418 62186 207654
rect 62422 207418 98186 207654
rect 98422 207418 134186 207654
rect 134422 207418 170186 207654
rect 170422 207418 206186 207654
rect 206422 207418 242186 207654
rect 242422 207418 278186 207654
rect 278422 207418 314186 207654
rect 314422 207418 350186 207654
rect 350422 207418 386186 207654
rect 386422 207418 422186 207654
rect 422422 207418 458186 207654
rect 458422 207418 494186 207654
rect 494422 207418 530186 207654
rect 530422 207418 566186 207654
rect 566422 207418 590102 207654
rect 590338 207418 590520 207654
rect -6596 207334 590520 207418
rect -6596 207098 -6414 207334
rect -6178 207098 26186 207334
rect 26422 207098 62186 207334
rect 62422 207098 98186 207334
rect 98422 207098 134186 207334
rect 134422 207098 170186 207334
rect 170422 207098 206186 207334
rect 206422 207098 242186 207334
rect 242422 207098 278186 207334
rect 278422 207098 314186 207334
rect 314422 207098 350186 207334
rect 350422 207098 386186 207334
rect 386422 207098 422186 207334
rect 422422 207098 458186 207334
rect 458422 207098 494186 207334
rect 494422 207098 530186 207334
rect 530422 207098 566186 207334
rect 566422 207098 590102 207334
rect 590338 207098 590520 207334
rect -6596 207076 590520 207098
rect -6596 207074 -5996 207076
rect 26004 207074 26604 207076
rect 62004 207074 62604 207076
rect 98004 207074 98604 207076
rect 134004 207074 134604 207076
rect 170004 207074 170604 207076
rect 206004 207074 206604 207076
rect 242004 207074 242604 207076
rect 278004 207074 278604 207076
rect 314004 207074 314604 207076
rect 350004 207074 350604 207076
rect 386004 207074 386604 207076
rect 422004 207074 422604 207076
rect 458004 207074 458604 207076
rect 494004 207074 494604 207076
rect 530004 207074 530604 207076
rect 566004 207074 566604 207076
rect 589920 207074 590520 207076
rect -4756 204076 -4156 204078
rect 22404 204076 23004 204078
rect 58404 204076 59004 204078
rect 94404 204076 95004 204078
rect 130404 204076 131004 204078
rect 166404 204076 167004 204078
rect 202404 204076 203004 204078
rect 238404 204076 239004 204078
rect 274404 204076 275004 204078
rect 310404 204076 311004 204078
rect 346404 204076 347004 204078
rect 382404 204076 383004 204078
rect 418404 204076 419004 204078
rect 454404 204076 455004 204078
rect 490404 204076 491004 204078
rect 526404 204076 527004 204078
rect 562404 204076 563004 204078
rect 588080 204076 588680 204078
rect -4756 204054 588680 204076
rect -4756 203818 -4574 204054
rect -4338 203818 22586 204054
rect 22822 203818 58586 204054
rect 58822 203818 94586 204054
rect 94822 203818 130586 204054
rect 130822 203818 166586 204054
rect 166822 203818 202586 204054
rect 202822 203818 238586 204054
rect 238822 203818 274586 204054
rect 274822 203818 310586 204054
rect 310822 203818 346586 204054
rect 346822 203818 382586 204054
rect 382822 203818 418586 204054
rect 418822 203818 454586 204054
rect 454822 203818 490586 204054
rect 490822 203818 526586 204054
rect 526822 203818 562586 204054
rect 562822 203818 588262 204054
rect 588498 203818 588680 204054
rect -4756 203734 588680 203818
rect -4756 203498 -4574 203734
rect -4338 203498 22586 203734
rect 22822 203498 58586 203734
rect 58822 203498 94586 203734
rect 94822 203498 130586 203734
rect 130822 203498 166586 203734
rect 166822 203498 202586 203734
rect 202822 203498 238586 203734
rect 238822 203498 274586 203734
rect 274822 203498 310586 203734
rect 310822 203498 346586 203734
rect 346822 203498 382586 203734
rect 382822 203498 418586 203734
rect 418822 203498 454586 203734
rect 454822 203498 490586 203734
rect 490822 203498 526586 203734
rect 526822 203498 562586 203734
rect 562822 203498 588262 203734
rect 588498 203498 588680 203734
rect -4756 203476 588680 203498
rect -4756 203474 -4156 203476
rect 22404 203474 23004 203476
rect 58404 203474 59004 203476
rect 94404 203474 95004 203476
rect 130404 203474 131004 203476
rect 166404 203474 167004 203476
rect 202404 203474 203004 203476
rect 238404 203474 239004 203476
rect 274404 203474 275004 203476
rect 310404 203474 311004 203476
rect 346404 203474 347004 203476
rect 382404 203474 383004 203476
rect 418404 203474 419004 203476
rect 454404 203474 455004 203476
rect 490404 203474 491004 203476
rect 526404 203474 527004 203476
rect 562404 203474 563004 203476
rect 588080 203474 588680 203476
rect -2916 200476 -2316 200478
rect 18804 200476 19404 200478
rect 54804 200476 55404 200478
rect 90804 200476 91404 200478
rect 126804 200476 127404 200478
rect 162804 200476 163404 200478
rect 198804 200476 199404 200478
rect 234804 200476 235404 200478
rect 270804 200476 271404 200478
rect 306804 200476 307404 200478
rect 342804 200476 343404 200478
rect 378804 200476 379404 200478
rect 414804 200476 415404 200478
rect 450804 200476 451404 200478
rect 486804 200476 487404 200478
rect 522804 200476 523404 200478
rect 558804 200476 559404 200478
rect 586240 200476 586840 200478
rect -2916 200454 586840 200476
rect -2916 200218 -2734 200454
rect -2498 200218 18986 200454
rect 19222 200218 54986 200454
rect 55222 200218 90986 200454
rect 91222 200218 126986 200454
rect 127222 200218 162986 200454
rect 163222 200218 198986 200454
rect 199222 200218 234986 200454
rect 235222 200218 270986 200454
rect 271222 200218 306986 200454
rect 307222 200218 342986 200454
rect 343222 200218 378986 200454
rect 379222 200218 414986 200454
rect 415222 200218 450986 200454
rect 451222 200218 486986 200454
rect 487222 200218 522986 200454
rect 523222 200218 558986 200454
rect 559222 200218 586422 200454
rect 586658 200218 586840 200454
rect -2916 200134 586840 200218
rect -2916 199898 -2734 200134
rect -2498 199898 18986 200134
rect 19222 199898 54986 200134
rect 55222 199898 90986 200134
rect 91222 199898 126986 200134
rect 127222 199898 162986 200134
rect 163222 199898 198986 200134
rect 199222 199898 234986 200134
rect 235222 199898 270986 200134
rect 271222 199898 306986 200134
rect 307222 199898 342986 200134
rect 343222 199898 378986 200134
rect 379222 199898 414986 200134
rect 415222 199898 450986 200134
rect 451222 199898 486986 200134
rect 487222 199898 522986 200134
rect 523222 199898 558986 200134
rect 559222 199898 586422 200134
rect 586658 199898 586840 200134
rect -2916 199876 586840 199898
rect -2916 199874 -2316 199876
rect 18804 199874 19404 199876
rect 54804 199874 55404 199876
rect 90804 199874 91404 199876
rect 126804 199874 127404 199876
rect 162804 199874 163404 199876
rect 198804 199874 199404 199876
rect 234804 199874 235404 199876
rect 270804 199874 271404 199876
rect 306804 199874 307404 199876
rect 342804 199874 343404 199876
rect 378804 199874 379404 199876
rect 414804 199874 415404 199876
rect 450804 199874 451404 199876
rect 486804 199874 487404 199876
rect 522804 199874 523404 199876
rect 558804 199874 559404 199876
rect 586240 199874 586840 199876
rect -7516 193276 -6916 193278
rect 11604 193276 12204 193278
rect 47604 193276 48204 193278
rect 83604 193276 84204 193278
rect 119604 193276 120204 193278
rect 155604 193276 156204 193278
rect 191604 193276 192204 193278
rect 227604 193276 228204 193278
rect 263604 193276 264204 193278
rect 299604 193276 300204 193278
rect 335604 193276 336204 193278
rect 371604 193276 372204 193278
rect 407604 193276 408204 193278
rect 443604 193276 444204 193278
rect 479604 193276 480204 193278
rect 515604 193276 516204 193278
rect 551604 193276 552204 193278
rect 590840 193276 591440 193278
rect -8436 193254 592360 193276
rect -8436 193018 -7334 193254
rect -7098 193018 11786 193254
rect 12022 193018 47786 193254
rect 48022 193018 83786 193254
rect 84022 193018 119786 193254
rect 120022 193018 155786 193254
rect 156022 193018 191786 193254
rect 192022 193018 227786 193254
rect 228022 193018 263786 193254
rect 264022 193018 299786 193254
rect 300022 193018 335786 193254
rect 336022 193018 371786 193254
rect 372022 193018 407786 193254
rect 408022 193018 443786 193254
rect 444022 193018 479786 193254
rect 480022 193018 515786 193254
rect 516022 193018 551786 193254
rect 552022 193018 591022 193254
rect 591258 193018 592360 193254
rect -8436 192934 592360 193018
rect -8436 192698 -7334 192934
rect -7098 192698 11786 192934
rect 12022 192698 47786 192934
rect 48022 192698 83786 192934
rect 84022 192698 119786 192934
rect 120022 192698 155786 192934
rect 156022 192698 191786 192934
rect 192022 192698 227786 192934
rect 228022 192698 263786 192934
rect 264022 192698 299786 192934
rect 300022 192698 335786 192934
rect 336022 192698 371786 192934
rect 372022 192698 407786 192934
rect 408022 192698 443786 192934
rect 444022 192698 479786 192934
rect 480022 192698 515786 192934
rect 516022 192698 551786 192934
rect 552022 192698 591022 192934
rect 591258 192698 592360 192934
rect -8436 192676 592360 192698
rect -7516 192674 -6916 192676
rect 11604 192674 12204 192676
rect 47604 192674 48204 192676
rect 83604 192674 84204 192676
rect 119604 192674 120204 192676
rect 155604 192674 156204 192676
rect 191604 192674 192204 192676
rect 227604 192674 228204 192676
rect 263604 192674 264204 192676
rect 299604 192674 300204 192676
rect 335604 192674 336204 192676
rect 371604 192674 372204 192676
rect 407604 192674 408204 192676
rect 443604 192674 444204 192676
rect 479604 192674 480204 192676
rect 515604 192674 516204 192676
rect 551604 192674 552204 192676
rect 590840 192674 591440 192676
rect -5676 189676 -5076 189678
rect 8004 189676 8604 189678
rect 44004 189676 44604 189678
rect 80004 189676 80604 189678
rect 116004 189676 116604 189678
rect 152004 189676 152604 189678
rect 188004 189676 188604 189678
rect 224004 189676 224604 189678
rect 260004 189676 260604 189678
rect 296004 189676 296604 189678
rect 332004 189676 332604 189678
rect 368004 189676 368604 189678
rect 404004 189676 404604 189678
rect 440004 189676 440604 189678
rect 476004 189676 476604 189678
rect 512004 189676 512604 189678
rect 548004 189676 548604 189678
rect 589000 189676 589600 189678
rect -6596 189654 590520 189676
rect -6596 189418 -5494 189654
rect -5258 189418 8186 189654
rect 8422 189418 44186 189654
rect 44422 189418 80186 189654
rect 80422 189418 116186 189654
rect 116422 189418 152186 189654
rect 152422 189418 188186 189654
rect 188422 189418 224186 189654
rect 224422 189418 260186 189654
rect 260422 189418 296186 189654
rect 296422 189418 332186 189654
rect 332422 189418 368186 189654
rect 368422 189418 404186 189654
rect 404422 189418 440186 189654
rect 440422 189418 476186 189654
rect 476422 189418 512186 189654
rect 512422 189418 548186 189654
rect 548422 189418 589182 189654
rect 589418 189418 590520 189654
rect -6596 189334 590520 189418
rect -6596 189098 -5494 189334
rect -5258 189098 8186 189334
rect 8422 189098 44186 189334
rect 44422 189098 80186 189334
rect 80422 189098 116186 189334
rect 116422 189098 152186 189334
rect 152422 189098 188186 189334
rect 188422 189098 224186 189334
rect 224422 189098 260186 189334
rect 260422 189098 296186 189334
rect 296422 189098 332186 189334
rect 332422 189098 368186 189334
rect 368422 189098 404186 189334
rect 404422 189098 440186 189334
rect 440422 189098 476186 189334
rect 476422 189098 512186 189334
rect 512422 189098 548186 189334
rect 548422 189098 589182 189334
rect 589418 189098 590520 189334
rect -6596 189076 590520 189098
rect -5676 189074 -5076 189076
rect 8004 189074 8604 189076
rect 44004 189074 44604 189076
rect 80004 189074 80604 189076
rect 116004 189074 116604 189076
rect 152004 189074 152604 189076
rect 188004 189074 188604 189076
rect 224004 189074 224604 189076
rect 260004 189074 260604 189076
rect 296004 189074 296604 189076
rect 332004 189074 332604 189076
rect 368004 189074 368604 189076
rect 404004 189074 404604 189076
rect 440004 189074 440604 189076
rect 476004 189074 476604 189076
rect 512004 189074 512604 189076
rect 548004 189074 548604 189076
rect 589000 189074 589600 189076
rect -3836 186076 -3236 186078
rect 4404 186076 5004 186078
rect 40404 186076 41004 186078
rect 76404 186076 77004 186078
rect 112404 186076 113004 186078
rect 148404 186076 149004 186078
rect 184404 186076 185004 186078
rect 220404 186076 221004 186078
rect 256404 186076 257004 186078
rect 292404 186076 293004 186078
rect 328404 186076 329004 186078
rect 364404 186076 365004 186078
rect 400404 186076 401004 186078
rect 436404 186076 437004 186078
rect 472404 186076 473004 186078
rect 508404 186076 509004 186078
rect 544404 186076 545004 186078
rect 580404 186076 581004 186078
rect 587160 186076 587760 186078
rect -4756 186054 588680 186076
rect -4756 185818 -3654 186054
rect -3418 185818 4586 186054
rect 4822 185818 40586 186054
rect 40822 185818 76586 186054
rect 76822 185818 112586 186054
rect 112822 185818 148586 186054
rect 148822 185818 184586 186054
rect 184822 185818 220586 186054
rect 220822 185818 256586 186054
rect 256822 185818 292586 186054
rect 292822 185818 328586 186054
rect 328822 185818 364586 186054
rect 364822 185818 400586 186054
rect 400822 185818 436586 186054
rect 436822 185818 472586 186054
rect 472822 185818 508586 186054
rect 508822 185818 544586 186054
rect 544822 185818 580586 186054
rect 580822 185818 587342 186054
rect 587578 185818 588680 186054
rect -4756 185734 588680 185818
rect -4756 185498 -3654 185734
rect -3418 185498 4586 185734
rect 4822 185498 40586 185734
rect 40822 185498 76586 185734
rect 76822 185498 112586 185734
rect 112822 185498 148586 185734
rect 148822 185498 184586 185734
rect 184822 185498 220586 185734
rect 220822 185498 256586 185734
rect 256822 185498 292586 185734
rect 292822 185498 328586 185734
rect 328822 185498 364586 185734
rect 364822 185498 400586 185734
rect 400822 185498 436586 185734
rect 436822 185498 472586 185734
rect 472822 185498 508586 185734
rect 508822 185498 544586 185734
rect 544822 185498 580586 185734
rect 580822 185498 587342 185734
rect 587578 185498 588680 185734
rect -4756 185476 588680 185498
rect -3836 185474 -3236 185476
rect 4404 185474 5004 185476
rect 40404 185474 41004 185476
rect 76404 185474 77004 185476
rect 112404 185474 113004 185476
rect 148404 185474 149004 185476
rect 184404 185474 185004 185476
rect 220404 185474 221004 185476
rect 256404 185474 257004 185476
rect 292404 185474 293004 185476
rect 328404 185474 329004 185476
rect 364404 185474 365004 185476
rect 400404 185474 401004 185476
rect 436404 185474 437004 185476
rect 472404 185474 473004 185476
rect 508404 185474 509004 185476
rect 544404 185474 545004 185476
rect 580404 185474 581004 185476
rect 587160 185474 587760 185476
rect -1996 182476 -1396 182478
rect 804 182476 1404 182478
rect 36804 182476 37404 182478
rect 72804 182476 73404 182478
rect 108804 182476 109404 182478
rect 144804 182476 145404 182478
rect 180804 182476 181404 182478
rect 216804 182476 217404 182478
rect 252804 182476 253404 182478
rect 288804 182476 289404 182478
rect 324804 182476 325404 182478
rect 360804 182476 361404 182478
rect 396804 182476 397404 182478
rect 432804 182476 433404 182478
rect 468804 182476 469404 182478
rect 504804 182476 505404 182478
rect 540804 182476 541404 182478
rect 576804 182476 577404 182478
rect 585320 182476 585920 182478
rect -2916 182454 586840 182476
rect -2916 182218 -1814 182454
rect -1578 182218 986 182454
rect 1222 182218 36986 182454
rect 37222 182218 72986 182454
rect 73222 182218 108986 182454
rect 109222 182218 144986 182454
rect 145222 182218 180986 182454
rect 181222 182218 216986 182454
rect 217222 182218 252986 182454
rect 253222 182218 288986 182454
rect 289222 182218 324986 182454
rect 325222 182218 360986 182454
rect 361222 182218 396986 182454
rect 397222 182218 432986 182454
rect 433222 182218 468986 182454
rect 469222 182218 504986 182454
rect 505222 182218 540986 182454
rect 541222 182218 576986 182454
rect 577222 182218 585502 182454
rect 585738 182218 586840 182454
rect -2916 182134 586840 182218
rect -2916 181898 -1814 182134
rect -1578 181898 986 182134
rect 1222 181898 36986 182134
rect 37222 181898 72986 182134
rect 73222 181898 108986 182134
rect 109222 181898 144986 182134
rect 145222 181898 180986 182134
rect 181222 181898 216986 182134
rect 217222 181898 252986 182134
rect 253222 181898 288986 182134
rect 289222 181898 324986 182134
rect 325222 181898 360986 182134
rect 361222 181898 396986 182134
rect 397222 181898 432986 182134
rect 433222 181898 468986 182134
rect 469222 181898 504986 182134
rect 505222 181898 540986 182134
rect 541222 181898 576986 182134
rect 577222 181898 585502 182134
rect 585738 181898 586840 182134
rect -2916 181876 586840 181898
rect -1996 181874 -1396 181876
rect 804 181874 1404 181876
rect 36804 181874 37404 181876
rect 72804 181874 73404 181876
rect 108804 181874 109404 181876
rect 144804 181874 145404 181876
rect 180804 181874 181404 181876
rect 216804 181874 217404 181876
rect 252804 181874 253404 181876
rect 288804 181874 289404 181876
rect 324804 181874 325404 181876
rect 360804 181874 361404 181876
rect 396804 181874 397404 181876
rect 432804 181874 433404 181876
rect 468804 181874 469404 181876
rect 504804 181874 505404 181876
rect 540804 181874 541404 181876
rect 576804 181874 577404 181876
rect 585320 181874 585920 181876
rect -8436 175276 -7836 175278
rect 29604 175276 30204 175278
rect 65604 175276 66204 175278
rect 101604 175276 102204 175278
rect 137604 175276 138204 175278
rect 173604 175276 174204 175278
rect 209604 175276 210204 175278
rect 245604 175276 246204 175278
rect 281604 175276 282204 175278
rect 317604 175276 318204 175278
rect 353604 175276 354204 175278
rect 389604 175276 390204 175278
rect 425604 175276 426204 175278
rect 461604 175276 462204 175278
rect 497604 175276 498204 175278
rect 533604 175276 534204 175278
rect 569604 175276 570204 175278
rect 591760 175276 592360 175278
rect -8436 175254 592360 175276
rect -8436 175018 -8254 175254
rect -8018 175018 29786 175254
rect 30022 175018 65786 175254
rect 66022 175018 101786 175254
rect 102022 175018 137786 175254
rect 138022 175018 173786 175254
rect 174022 175018 209786 175254
rect 210022 175018 245786 175254
rect 246022 175018 281786 175254
rect 282022 175018 317786 175254
rect 318022 175018 353786 175254
rect 354022 175018 389786 175254
rect 390022 175018 425786 175254
rect 426022 175018 461786 175254
rect 462022 175018 497786 175254
rect 498022 175018 533786 175254
rect 534022 175018 569786 175254
rect 570022 175018 591942 175254
rect 592178 175018 592360 175254
rect -8436 174934 592360 175018
rect -8436 174698 -8254 174934
rect -8018 174698 29786 174934
rect 30022 174698 65786 174934
rect 66022 174698 101786 174934
rect 102022 174698 137786 174934
rect 138022 174698 173786 174934
rect 174022 174698 209786 174934
rect 210022 174698 245786 174934
rect 246022 174698 281786 174934
rect 282022 174698 317786 174934
rect 318022 174698 353786 174934
rect 354022 174698 389786 174934
rect 390022 174698 425786 174934
rect 426022 174698 461786 174934
rect 462022 174698 497786 174934
rect 498022 174698 533786 174934
rect 534022 174698 569786 174934
rect 570022 174698 591942 174934
rect 592178 174698 592360 174934
rect -8436 174676 592360 174698
rect -8436 174674 -7836 174676
rect 29604 174674 30204 174676
rect 65604 174674 66204 174676
rect 101604 174674 102204 174676
rect 137604 174674 138204 174676
rect 173604 174674 174204 174676
rect 209604 174674 210204 174676
rect 245604 174674 246204 174676
rect 281604 174674 282204 174676
rect 317604 174674 318204 174676
rect 353604 174674 354204 174676
rect 389604 174674 390204 174676
rect 425604 174674 426204 174676
rect 461604 174674 462204 174676
rect 497604 174674 498204 174676
rect 533604 174674 534204 174676
rect 569604 174674 570204 174676
rect 591760 174674 592360 174676
rect -6596 171676 -5996 171678
rect 26004 171676 26604 171678
rect 62004 171676 62604 171678
rect 98004 171676 98604 171678
rect 134004 171676 134604 171678
rect 170004 171676 170604 171678
rect 206004 171676 206604 171678
rect 242004 171676 242604 171678
rect 278004 171676 278604 171678
rect 314004 171676 314604 171678
rect 350004 171676 350604 171678
rect 386004 171676 386604 171678
rect 422004 171676 422604 171678
rect 458004 171676 458604 171678
rect 494004 171676 494604 171678
rect 530004 171676 530604 171678
rect 566004 171676 566604 171678
rect 589920 171676 590520 171678
rect -6596 171654 590520 171676
rect -6596 171418 -6414 171654
rect -6178 171418 26186 171654
rect 26422 171418 62186 171654
rect 62422 171418 98186 171654
rect 98422 171418 134186 171654
rect 134422 171418 170186 171654
rect 170422 171418 206186 171654
rect 206422 171418 242186 171654
rect 242422 171418 278186 171654
rect 278422 171418 314186 171654
rect 314422 171418 350186 171654
rect 350422 171418 386186 171654
rect 386422 171418 422186 171654
rect 422422 171418 458186 171654
rect 458422 171418 494186 171654
rect 494422 171418 530186 171654
rect 530422 171418 566186 171654
rect 566422 171418 590102 171654
rect 590338 171418 590520 171654
rect -6596 171334 590520 171418
rect -6596 171098 -6414 171334
rect -6178 171098 26186 171334
rect 26422 171098 62186 171334
rect 62422 171098 98186 171334
rect 98422 171098 134186 171334
rect 134422 171098 170186 171334
rect 170422 171098 206186 171334
rect 206422 171098 242186 171334
rect 242422 171098 278186 171334
rect 278422 171098 314186 171334
rect 314422 171098 350186 171334
rect 350422 171098 386186 171334
rect 386422 171098 422186 171334
rect 422422 171098 458186 171334
rect 458422 171098 494186 171334
rect 494422 171098 530186 171334
rect 530422 171098 566186 171334
rect 566422 171098 590102 171334
rect 590338 171098 590520 171334
rect -6596 171076 590520 171098
rect -6596 171074 -5996 171076
rect 26004 171074 26604 171076
rect 62004 171074 62604 171076
rect 98004 171074 98604 171076
rect 134004 171074 134604 171076
rect 170004 171074 170604 171076
rect 206004 171074 206604 171076
rect 242004 171074 242604 171076
rect 278004 171074 278604 171076
rect 314004 171074 314604 171076
rect 350004 171074 350604 171076
rect 386004 171074 386604 171076
rect 422004 171074 422604 171076
rect 458004 171074 458604 171076
rect 494004 171074 494604 171076
rect 530004 171074 530604 171076
rect 566004 171074 566604 171076
rect 589920 171074 590520 171076
rect -4756 168076 -4156 168078
rect 22404 168076 23004 168078
rect 58404 168076 59004 168078
rect 94404 168076 95004 168078
rect 130404 168076 131004 168078
rect 166404 168076 167004 168078
rect 202404 168076 203004 168078
rect 238404 168076 239004 168078
rect 274404 168076 275004 168078
rect 310404 168076 311004 168078
rect 346404 168076 347004 168078
rect 382404 168076 383004 168078
rect 418404 168076 419004 168078
rect 454404 168076 455004 168078
rect 490404 168076 491004 168078
rect 526404 168076 527004 168078
rect 562404 168076 563004 168078
rect 588080 168076 588680 168078
rect -4756 168054 588680 168076
rect -4756 167818 -4574 168054
rect -4338 167818 22586 168054
rect 22822 167818 58586 168054
rect 58822 167818 94586 168054
rect 94822 167818 130586 168054
rect 130822 167818 166586 168054
rect 166822 167818 202586 168054
rect 202822 167818 238586 168054
rect 238822 167818 274586 168054
rect 274822 167818 310586 168054
rect 310822 167818 346586 168054
rect 346822 167818 382586 168054
rect 382822 167818 418586 168054
rect 418822 167818 454586 168054
rect 454822 167818 490586 168054
rect 490822 167818 526586 168054
rect 526822 167818 562586 168054
rect 562822 167818 588262 168054
rect 588498 167818 588680 168054
rect -4756 167734 588680 167818
rect -4756 167498 -4574 167734
rect -4338 167498 22586 167734
rect 22822 167498 58586 167734
rect 58822 167498 94586 167734
rect 94822 167498 130586 167734
rect 130822 167498 166586 167734
rect 166822 167498 202586 167734
rect 202822 167498 238586 167734
rect 238822 167498 274586 167734
rect 274822 167498 310586 167734
rect 310822 167498 346586 167734
rect 346822 167498 382586 167734
rect 382822 167498 418586 167734
rect 418822 167498 454586 167734
rect 454822 167498 490586 167734
rect 490822 167498 526586 167734
rect 526822 167498 562586 167734
rect 562822 167498 588262 167734
rect 588498 167498 588680 167734
rect -4756 167476 588680 167498
rect -4756 167474 -4156 167476
rect 22404 167474 23004 167476
rect 58404 167474 59004 167476
rect 94404 167474 95004 167476
rect 130404 167474 131004 167476
rect 166404 167474 167004 167476
rect 202404 167474 203004 167476
rect 238404 167474 239004 167476
rect 274404 167474 275004 167476
rect 310404 167474 311004 167476
rect 346404 167474 347004 167476
rect 382404 167474 383004 167476
rect 418404 167474 419004 167476
rect 454404 167474 455004 167476
rect 490404 167474 491004 167476
rect 526404 167474 527004 167476
rect 562404 167474 563004 167476
rect 588080 167474 588680 167476
rect -2916 164476 -2316 164478
rect 18804 164476 19404 164478
rect 54804 164476 55404 164478
rect 90804 164476 91404 164478
rect 126804 164476 127404 164478
rect 162804 164476 163404 164478
rect 198804 164476 199404 164478
rect 234804 164476 235404 164478
rect 270804 164476 271404 164478
rect 306804 164476 307404 164478
rect 342804 164476 343404 164478
rect 378804 164476 379404 164478
rect 414804 164476 415404 164478
rect 450804 164476 451404 164478
rect 486804 164476 487404 164478
rect 522804 164476 523404 164478
rect 558804 164476 559404 164478
rect 586240 164476 586840 164478
rect -2916 164454 586840 164476
rect -2916 164218 -2734 164454
rect -2498 164218 18986 164454
rect 19222 164218 54986 164454
rect 55222 164218 90986 164454
rect 91222 164218 126986 164454
rect 127222 164218 162986 164454
rect 163222 164218 198986 164454
rect 199222 164218 234986 164454
rect 235222 164218 270986 164454
rect 271222 164218 306986 164454
rect 307222 164218 342986 164454
rect 343222 164218 378986 164454
rect 379222 164218 414986 164454
rect 415222 164218 450986 164454
rect 451222 164218 486986 164454
rect 487222 164218 522986 164454
rect 523222 164218 558986 164454
rect 559222 164218 586422 164454
rect 586658 164218 586840 164454
rect -2916 164134 586840 164218
rect -2916 163898 -2734 164134
rect -2498 163898 18986 164134
rect 19222 163898 54986 164134
rect 55222 163898 90986 164134
rect 91222 163898 126986 164134
rect 127222 163898 162986 164134
rect 163222 163898 198986 164134
rect 199222 163898 234986 164134
rect 235222 163898 270986 164134
rect 271222 163898 306986 164134
rect 307222 163898 342986 164134
rect 343222 163898 378986 164134
rect 379222 163898 414986 164134
rect 415222 163898 450986 164134
rect 451222 163898 486986 164134
rect 487222 163898 522986 164134
rect 523222 163898 558986 164134
rect 559222 163898 586422 164134
rect 586658 163898 586840 164134
rect -2916 163876 586840 163898
rect -2916 163874 -2316 163876
rect 18804 163874 19404 163876
rect 54804 163874 55404 163876
rect 90804 163874 91404 163876
rect 126804 163874 127404 163876
rect 162804 163874 163404 163876
rect 198804 163874 199404 163876
rect 234804 163874 235404 163876
rect 270804 163874 271404 163876
rect 306804 163874 307404 163876
rect 342804 163874 343404 163876
rect 378804 163874 379404 163876
rect 414804 163874 415404 163876
rect 450804 163874 451404 163876
rect 486804 163874 487404 163876
rect 522804 163874 523404 163876
rect 558804 163874 559404 163876
rect 586240 163874 586840 163876
rect -7516 157276 -6916 157278
rect 11604 157276 12204 157278
rect 47604 157276 48204 157278
rect 83604 157276 84204 157278
rect 119604 157276 120204 157278
rect 155604 157276 156204 157278
rect 191604 157276 192204 157278
rect 227604 157276 228204 157278
rect 263604 157276 264204 157278
rect 299604 157276 300204 157278
rect 335604 157276 336204 157278
rect 371604 157276 372204 157278
rect 407604 157276 408204 157278
rect 443604 157276 444204 157278
rect 479604 157276 480204 157278
rect 515604 157276 516204 157278
rect 551604 157276 552204 157278
rect 590840 157276 591440 157278
rect -8436 157254 592360 157276
rect -8436 157018 -7334 157254
rect -7098 157018 11786 157254
rect 12022 157018 47786 157254
rect 48022 157018 83786 157254
rect 84022 157018 119786 157254
rect 120022 157018 155786 157254
rect 156022 157018 191786 157254
rect 192022 157018 227786 157254
rect 228022 157018 263786 157254
rect 264022 157018 299786 157254
rect 300022 157018 335786 157254
rect 336022 157018 371786 157254
rect 372022 157018 407786 157254
rect 408022 157018 443786 157254
rect 444022 157018 479786 157254
rect 480022 157018 515786 157254
rect 516022 157018 551786 157254
rect 552022 157018 591022 157254
rect 591258 157018 592360 157254
rect -8436 156934 592360 157018
rect -8436 156698 -7334 156934
rect -7098 156698 11786 156934
rect 12022 156698 47786 156934
rect 48022 156698 83786 156934
rect 84022 156698 119786 156934
rect 120022 156698 155786 156934
rect 156022 156698 191786 156934
rect 192022 156698 227786 156934
rect 228022 156698 263786 156934
rect 264022 156698 299786 156934
rect 300022 156698 335786 156934
rect 336022 156698 371786 156934
rect 372022 156698 407786 156934
rect 408022 156698 443786 156934
rect 444022 156698 479786 156934
rect 480022 156698 515786 156934
rect 516022 156698 551786 156934
rect 552022 156698 591022 156934
rect 591258 156698 592360 156934
rect -8436 156676 592360 156698
rect -7516 156674 -6916 156676
rect 11604 156674 12204 156676
rect 47604 156674 48204 156676
rect 83604 156674 84204 156676
rect 119604 156674 120204 156676
rect 155604 156674 156204 156676
rect 191604 156674 192204 156676
rect 227604 156674 228204 156676
rect 263604 156674 264204 156676
rect 299604 156674 300204 156676
rect 335604 156674 336204 156676
rect 371604 156674 372204 156676
rect 407604 156674 408204 156676
rect 443604 156674 444204 156676
rect 479604 156674 480204 156676
rect 515604 156674 516204 156676
rect 551604 156674 552204 156676
rect 590840 156674 591440 156676
rect -5676 153676 -5076 153678
rect 8004 153676 8604 153678
rect 44004 153676 44604 153678
rect 80004 153676 80604 153678
rect 116004 153676 116604 153678
rect 152004 153676 152604 153678
rect 188004 153676 188604 153678
rect 224004 153676 224604 153678
rect 260004 153676 260604 153678
rect 296004 153676 296604 153678
rect 332004 153676 332604 153678
rect 368004 153676 368604 153678
rect 404004 153676 404604 153678
rect 440004 153676 440604 153678
rect 476004 153676 476604 153678
rect 512004 153676 512604 153678
rect 548004 153676 548604 153678
rect 589000 153676 589600 153678
rect -6596 153654 590520 153676
rect -6596 153418 -5494 153654
rect -5258 153418 8186 153654
rect 8422 153418 44186 153654
rect 44422 153418 80186 153654
rect 80422 153418 116186 153654
rect 116422 153418 152186 153654
rect 152422 153418 188186 153654
rect 188422 153418 224186 153654
rect 224422 153418 260186 153654
rect 260422 153418 296186 153654
rect 296422 153418 332186 153654
rect 332422 153418 368186 153654
rect 368422 153418 404186 153654
rect 404422 153418 440186 153654
rect 440422 153418 476186 153654
rect 476422 153418 512186 153654
rect 512422 153418 548186 153654
rect 548422 153418 589182 153654
rect 589418 153418 590520 153654
rect -6596 153334 590520 153418
rect -6596 153098 -5494 153334
rect -5258 153098 8186 153334
rect 8422 153098 44186 153334
rect 44422 153098 80186 153334
rect 80422 153098 116186 153334
rect 116422 153098 152186 153334
rect 152422 153098 188186 153334
rect 188422 153098 224186 153334
rect 224422 153098 260186 153334
rect 260422 153098 296186 153334
rect 296422 153098 332186 153334
rect 332422 153098 368186 153334
rect 368422 153098 404186 153334
rect 404422 153098 440186 153334
rect 440422 153098 476186 153334
rect 476422 153098 512186 153334
rect 512422 153098 548186 153334
rect 548422 153098 589182 153334
rect 589418 153098 590520 153334
rect -6596 153076 590520 153098
rect -5676 153074 -5076 153076
rect 8004 153074 8604 153076
rect 44004 153074 44604 153076
rect 80004 153074 80604 153076
rect 116004 153074 116604 153076
rect 152004 153074 152604 153076
rect 188004 153074 188604 153076
rect 224004 153074 224604 153076
rect 260004 153074 260604 153076
rect 296004 153074 296604 153076
rect 332004 153074 332604 153076
rect 368004 153074 368604 153076
rect 404004 153074 404604 153076
rect 440004 153074 440604 153076
rect 476004 153074 476604 153076
rect 512004 153074 512604 153076
rect 548004 153074 548604 153076
rect 589000 153074 589600 153076
rect -3836 150076 -3236 150078
rect 4404 150076 5004 150078
rect 40404 150076 41004 150078
rect 76404 150076 77004 150078
rect 112404 150076 113004 150078
rect 148404 150076 149004 150078
rect 184404 150076 185004 150078
rect 220404 150076 221004 150078
rect 256404 150076 257004 150078
rect 292404 150076 293004 150078
rect 328404 150076 329004 150078
rect 364404 150076 365004 150078
rect 400404 150076 401004 150078
rect 436404 150076 437004 150078
rect 472404 150076 473004 150078
rect 508404 150076 509004 150078
rect 544404 150076 545004 150078
rect 580404 150076 581004 150078
rect 587160 150076 587760 150078
rect -4756 150054 588680 150076
rect -4756 149818 -3654 150054
rect -3418 149818 4586 150054
rect 4822 149818 40586 150054
rect 40822 149818 76586 150054
rect 76822 149818 112586 150054
rect 112822 149818 148586 150054
rect 148822 149818 184586 150054
rect 184822 149818 220586 150054
rect 220822 149818 256586 150054
rect 256822 149818 292586 150054
rect 292822 149818 328586 150054
rect 328822 149818 364586 150054
rect 364822 149818 400586 150054
rect 400822 149818 436586 150054
rect 436822 149818 472586 150054
rect 472822 149818 508586 150054
rect 508822 149818 544586 150054
rect 544822 149818 580586 150054
rect 580822 149818 587342 150054
rect 587578 149818 588680 150054
rect -4756 149734 588680 149818
rect -4756 149498 -3654 149734
rect -3418 149498 4586 149734
rect 4822 149498 40586 149734
rect 40822 149498 76586 149734
rect 76822 149498 112586 149734
rect 112822 149498 148586 149734
rect 148822 149498 184586 149734
rect 184822 149498 220586 149734
rect 220822 149498 256586 149734
rect 256822 149498 292586 149734
rect 292822 149498 328586 149734
rect 328822 149498 364586 149734
rect 364822 149498 400586 149734
rect 400822 149498 436586 149734
rect 436822 149498 472586 149734
rect 472822 149498 508586 149734
rect 508822 149498 544586 149734
rect 544822 149498 580586 149734
rect 580822 149498 587342 149734
rect 587578 149498 588680 149734
rect -4756 149476 588680 149498
rect -3836 149474 -3236 149476
rect 4404 149474 5004 149476
rect 40404 149474 41004 149476
rect 76404 149474 77004 149476
rect 112404 149474 113004 149476
rect 148404 149474 149004 149476
rect 184404 149474 185004 149476
rect 220404 149474 221004 149476
rect 256404 149474 257004 149476
rect 292404 149474 293004 149476
rect 328404 149474 329004 149476
rect 364404 149474 365004 149476
rect 400404 149474 401004 149476
rect 436404 149474 437004 149476
rect 472404 149474 473004 149476
rect 508404 149474 509004 149476
rect 544404 149474 545004 149476
rect 580404 149474 581004 149476
rect 587160 149474 587760 149476
rect -1996 146476 -1396 146478
rect 804 146476 1404 146478
rect 36804 146476 37404 146478
rect 72804 146476 73404 146478
rect 108804 146476 109404 146478
rect 144804 146476 145404 146478
rect 180804 146476 181404 146478
rect 216804 146476 217404 146478
rect 252804 146476 253404 146478
rect 288804 146476 289404 146478
rect 324804 146476 325404 146478
rect 360804 146476 361404 146478
rect 396804 146476 397404 146478
rect 432804 146476 433404 146478
rect 468804 146476 469404 146478
rect 504804 146476 505404 146478
rect 540804 146476 541404 146478
rect 576804 146476 577404 146478
rect 585320 146476 585920 146478
rect -2916 146454 586840 146476
rect -2916 146218 -1814 146454
rect -1578 146218 986 146454
rect 1222 146218 36986 146454
rect 37222 146218 72986 146454
rect 73222 146218 108986 146454
rect 109222 146218 144986 146454
rect 145222 146218 180986 146454
rect 181222 146218 216986 146454
rect 217222 146218 252986 146454
rect 253222 146218 288986 146454
rect 289222 146218 324986 146454
rect 325222 146218 360986 146454
rect 361222 146218 396986 146454
rect 397222 146218 432986 146454
rect 433222 146218 468986 146454
rect 469222 146218 504986 146454
rect 505222 146218 540986 146454
rect 541222 146218 576986 146454
rect 577222 146218 585502 146454
rect 585738 146218 586840 146454
rect -2916 146134 586840 146218
rect -2916 145898 -1814 146134
rect -1578 145898 986 146134
rect 1222 145898 36986 146134
rect 37222 145898 72986 146134
rect 73222 145898 108986 146134
rect 109222 145898 144986 146134
rect 145222 145898 180986 146134
rect 181222 145898 216986 146134
rect 217222 145898 252986 146134
rect 253222 145898 288986 146134
rect 289222 145898 324986 146134
rect 325222 145898 360986 146134
rect 361222 145898 396986 146134
rect 397222 145898 432986 146134
rect 433222 145898 468986 146134
rect 469222 145898 504986 146134
rect 505222 145898 540986 146134
rect 541222 145898 576986 146134
rect 577222 145898 585502 146134
rect 585738 145898 586840 146134
rect -2916 145876 586840 145898
rect -1996 145874 -1396 145876
rect 804 145874 1404 145876
rect 36804 145874 37404 145876
rect 72804 145874 73404 145876
rect 108804 145874 109404 145876
rect 144804 145874 145404 145876
rect 180804 145874 181404 145876
rect 216804 145874 217404 145876
rect 252804 145874 253404 145876
rect 288804 145874 289404 145876
rect 324804 145874 325404 145876
rect 360804 145874 361404 145876
rect 396804 145874 397404 145876
rect 432804 145874 433404 145876
rect 468804 145874 469404 145876
rect 504804 145874 505404 145876
rect 540804 145874 541404 145876
rect 576804 145874 577404 145876
rect 585320 145874 585920 145876
rect -8436 139276 -7836 139278
rect 29604 139276 30204 139278
rect 65604 139276 66204 139278
rect 101604 139276 102204 139278
rect 137604 139276 138204 139278
rect 173604 139276 174204 139278
rect 209604 139276 210204 139278
rect 245604 139276 246204 139278
rect 281604 139276 282204 139278
rect 317604 139276 318204 139278
rect 353604 139276 354204 139278
rect 389604 139276 390204 139278
rect 425604 139276 426204 139278
rect 461604 139276 462204 139278
rect 497604 139276 498204 139278
rect 533604 139276 534204 139278
rect 569604 139276 570204 139278
rect 591760 139276 592360 139278
rect -8436 139254 592360 139276
rect -8436 139018 -8254 139254
rect -8018 139018 29786 139254
rect 30022 139018 65786 139254
rect 66022 139018 101786 139254
rect 102022 139018 137786 139254
rect 138022 139018 173786 139254
rect 174022 139018 209786 139254
rect 210022 139018 245786 139254
rect 246022 139018 281786 139254
rect 282022 139018 317786 139254
rect 318022 139018 353786 139254
rect 354022 139018 389786 139254
rect 390022 139018 425786 139254
rect 426022 139018 461786 139254
rect 462022 139018 497786 139254
rect 498022 139018 533786 139254
rect 534022 139018 569786 139254
rect 570022 139018 591942 139254
rect 592178 139018 592360 139254
rect -8436 138934 592360 139018
rect -8436 138698 -8254 138934
rect -8018 138698 29786 138934
rect 30022 138698 65786 138934
rect 66022 138698 101786 138934
rect 102022 138698 137786 138934
rect 138022 138698 173786 138934
rect 174022 138698 209786 138934
rect 210022 138698 245786 138934
rect 246022 138698 281786 138934
rect 282022 138698 317786 138934
rect 318022 138698 353786 138934
rect 354022 138698 389786 138934
rect 390022 138698 425786 138934
rect 426022 138698 461786 138934
rect 462022 138698 497786 138934
rect 498022 138698 533786 138934
rect 534022 138698 569786 138934
rect 570022 138698 591942 138934
rect 592178 138698 592360 138934
rect -8436 138676 592360 138698
rect -8436 138674 -7836 138676
rect 29604 138674 30204 138676
rect 65604 138674 66204 138676
rect 101604 138674 102204 138676
rect 137604 138674 138204 138676
rect 173604 138674 174204 138676
rect 209604 138674 210204 138676
rect 245604 138674 246204 138676
rect 281604 138674 282204 138676
rect 317604 138674 318204 138676
rect 353604 138674 354204 138676
rect 389604 138674 390204 138676
rect 425604 138674 426204 138676
rect 461604 138674 462204 138676
rect 497604 138674 498204 138676
rect 533604 138674 534204 138676
rect 569604 138674 570204 138676
rect 591760 138674 592360 138676
rect -6596 135676 -5996 135678
rect 26004 135676 26604 135678
rect 62004 135676 62604 135678
rect 98004 135676 98604 135678
rect 134004 135676 134604 135678
rect 170004 135676 170604 135678
rect 206004 135676 206604 135678
rect 242004 135676 242604 135678
rect 278004 135676 278604 135678
rect 314004 135676 314604 135678
rect 350004 135676 350604 135678
rect 386004 135676 386604 135678
rect 422004 135676 422604 135678
rect 458004 135676 458604 135678
rect 494004 135676 494604 135678
rect 530004 135676 530604 135678
rect 566004 135676 566604 135678
rect 589920 135676 590520 135678
rect -6596 135654 590520 135676
rect -6596 135418 -6414 135654
rect -6178 135418 26186 135654
rect 26422 135418 62186 135654
rect 62422 135418 98186 135654
rect 98422 135418 134186 135654
rect 134422 135418 170186 135654
rect 170422 135418 206186 135654
rect 206422 135418 242186 135654
rect 242422 135418 278186 135654
rect 278422 135418 314186 135654
rect 314422 135418 350186 135654
rect 350422 135418 386186 135654
rect 386422 135418 422186 135654
rect 422422 135418 458186 135654
rect 458422 135418 494186 135654
rect 494422 135418 530186 135654
rect 530422 135418 566186 135654
rect 566422 135418 590102 135654
rect 590338 135418 590520 135654
rect -6596 135334 590520 135418
rect -6596 135098 -6414 135334
rect -6178 135098 26186 135334
rect 26422 135098 62186 135334
rect 62422 135098 98186 135334
rect 98422 135098 134186 135334
rect 134422 135098 170186 135334
rect 170422 135098 206186 135334
rect 206422 135098 242186 135334
rect 242422 135098 278186 135334
rect 278422 135098 314186 135334
rect 314422 135098 350186 135334
rect 350422 135098 386186 135334
rect 386422 135098 422186 135334
rect 422422 135098 458186 135334
rect 458422 135098 494186 135334
rect 494422 135098 530186 135334
rect 530422 135098 566186 135334
rect 566422 135098 590102 135334
rect 590338 135098 590520 135334
rect -6596 135076 590520 135098
rect -6596 135074 -5996 135076
rect 26004 135074 26604 135076
rect 62004 135074 62604 135076
rect 98004 135074 98604 135076
rect 134004 135074 134604 135076
rect 170004 135074 170604 135076
rect 206004 135074 206604 135076
rect 242004 135074 242604 135076
rect 278004 135074 278604 135076
rect 314004 135074 314604 135076
rect 350004 135074 350604 135076
rect 386004 135074 386604 135076
rect 422004 135074 422604 135076
rect 458004 135074 458604 135076
rect 494004 135074 494604 135076
rect 530004 135074 530604 135076
rect 566004 135074 566604 135076
rect 589920 135074 590520 135076
rect -4756 132076 -4156 132078
rect 22404 132076 23004 132078
rect 58404 132076 59004 132078
rect 94404 132076 95004 132078
rect 130404 132076 131004 132078
rect 166404 132076 167004 132078
rect 202404 132076 203004 132078
rect 238404 132076 239004 132078
rect 274404 132076 275004 132078
rect 310404 132076 311004 132078
rect 346404 132076 347004 132078
rect 382404 132076 383004 132078
rect 418404 132076 419004 132078
rect 454404 132076 455004 132078
rect 490404 132076 491004 132078
rect 526404 132076 527004 132078
rect 562404 132076 563004 132078
rect 588080 132076 588680 132078
rect -4756 132054 588680 132076
rect -4756 131818 -4574 132054
rect -4338 131818 22586 132054
rect 22822 131818 58586 132054
rect 58822 131818 94586 132054
rect 94822 131818 130586 132054
rect 130822 131818 166586 132054
rect 166822 131818 202586 132054
rect 202822 131818 238586 132054
rect 238822 131818 274586 132054
rect 274822 131818 310586 132054
rect 310822 131818 346586 132054
rect 346822 131818 382586 132054
rect 382822 131818 418586 132054
rect 418822 131818 454586 132054
rect 454822 131818 490586 132054
rect 490822 131818 526586 132054
rect 526822 131818 562586 132054
rect 562822 131818 588262 132054
rect 588498 131818 588680 132054
rect -4756 131734 588680 131818
rect -4756 131498 -4574 131734
rect -4338 131498 22586 131734
rect 22822 131498 58586 131734
rect 58822 131498 94586 131734
rect 94822 131498 130586 131734
rect 130822 131498 166586 131734
rect 166822 131498 202586 131734
rect 202822 131498 238586 131734
rect 238822 131498 274586 131734
rect 274822 131498 310586 131734
rect 310822 131498 346586 131734
rect 346822 131498 382586 131734
rect 382822 131498 418586 131734
rect 418822 131498 454586 131734
rect 454822 131498 490586 131734
rect 490822 131498 526586 131734
rect 526822 131498 562586 131734
rect 562822 131498 588262 131734
rect 588498 131498 588680 131734
rect -4756 131476 588680 131498
rect -4756 131474 -4156 131476
rect 22404 131474 23004 131476
rect 58404 131474 59004 131476
rect 94404 131474 95004 131476
rect 130404 131474 131004 131476
rect 166404 131474 167004 131476
rect 202404 131474 203004 131476
rect 238404 131474 239004 131476
rect 274404 131474 275004 131476
rect 310404 131474 311004 131476
rect 346404 131474 347004 131476
rect 382404 131474 383004 131476
rect 418404 131474 419004 131476
rect 454404 131474 455004 131476
rect 490404 131474 491004 131476
rect 526404 131474 527004 131476
rect 562404 131474 563004 131476
rect 588080 131474 588680 131476
rect -2916 128476 -2316 128478
rect 18804 128476 19404 128478
rect 54804 128476 55404 128478
rect 90804 128476 91404 128478
rect 126804 128476 127404 128478
rect 162804 128476 163404 128478
rect 198804 128476 199404 128478
rect 234804 128476 235404 128478
rect 270804 128476 271404 128478
rect 306804 128476 307404 128478
rect 342804 128476 343404 128478
rect 378804 128476 379404 128478
rect 414804 128476 415404 128478
rect 450804 128476 451404 128478
rect 486804 128476 487404 128478
rect 522804 128476 523404 128478
rect 558804 128476 559404 128478
rect 586240 128476 586840 128478
rect -2916 128454 586840 128476
rect -2916 128218 -2734 128454
rect -2498 128218 18986 128454
rect 19222 128218 54986 128454
rect 55222 128218 90986 128454
rect 91222 128218 126986 128454
rect 127222 128218 162986 128454
rect 163222 128218 198986 128454
rect 199222 128218 234986 128454
rect 235222 128218 270986 128454
rect 271222 128218 306986 128454
rect 307222 128218 342986 128454
rect 343222 128218 378986 128454
rect 379222 128218 414986 128454
rect 415222 128218 450986 128454
rect 451222 128218 486986 128454
rect 487222 128218 522986 128454
rect 523222 128218 558986 128454
rect 559222 128218 586422 128454
rect 586658 128218 586840 128454
rect -2916 128134 586840 128218
rect -2916 127898 -2734 128134
rect -2498 127898 18986 128134
rect 19222 127898 54986 128134
rect 55222 127898 90986 128134
rect 91222 127898 126986 128134
rect 127222 127898 162986 128134
rect 163222 127898 198986 128134
rect 199222 127898 234986 128134
rect 235222 127898 270986 128134
rect 271222 127898 306986 128134
rect 307222 127898 342986 128134
rect 343222 127898 378986 128134
rect 379222 127898 414986 128134
rect 415222 127898 450986 128134
rect 451222 127898 486986 128134
rect 487222 127898 522986 128134
rect 523222 127898 558986 128134
rect 559222 127898 586422 128134
rect 586658 127898 586840 128134
rect -2916 127876 586840 127898
rect -2916 127874 -2316 127876
rect 18804 127874 19404 127876
rect 54804 127874 55404 127876
rect 90804 127874 91404 127876
rect 126804 127874 127404 127876
rect 162804 127874 163404 127876
rect 198804 127874 199404 127876
rect 234804 127874 235404 127876
rect 270804 127874 271404 127876
rect 306804 127874 307404 127876
rect 342804 127874 343404 127876
rect 378804 127874 379404 127876
rect 414804 127874 415404 127876
rect 450804 127874 451404 127876
rect 486804 127874 487404 127876
rect 522804 127874 523404 127876
rect 558804 127874 559404 127876
rect 586240 127874 586840 127876
rect -7516 121276 -6916 121278
rect 11604 121276 12204 121278
rect 47604 121276 48204 121278
rect 83604 121276 84204 121278
rect 119604 121276 120204 121278
rect 155604 121276 156204 121278
rect 191604 121276 192204 121278
rect 227604 121276 228204 121278
rect 263604 121276 264204 121278
rect 299604 121276 300204 121278
rect 335604 121276 336204 121278
rect 371604 121276 372204 121278
rect 407604 121276 408204 121278
rect 443604 121276 444204 121278
rect 479604 121276 480204 121278
rect 515604 121276 516204 121278
rect 551604 121276 552204 121278
rect 590840 121276 591440 121278
rect -8436 121254 592360 121276
rect -8436 121018 -7334 121254
rect -7098 121018 11786 121254
rect 12022 121018 47786 121254
rect 48022 121018 83786 121254
rect 84022 121018 119786 121254
rect 120022 121018 155786 121254
rect 156022 121018 191786 121254
rect 192022 121018 227786 121254
rect 228022 121018 263786 121254
rect 264022 121018 299786 121254
rect 300022 121018 335786 121254
rect 336022 121018 371786 121254
rect 372022 121018 407786 121254
rect 408022 121018 443786 121254
rect 444022 121018 479786 121254
rect 480022 121018 515786 121254
rect 516022 121018 551786 121254
rect 552022 121018 591022 121254
rect 591258 121018 592360 121254
rect -8436 120934 592360 121018
rect -8436 120698 -7334 120934
rect -7098 120698 11786 120934
rect 12022 120698 47786 120934
rect 48022 120698 83786 120934
rect 84022 120698 119786 120934
rect 120022 120698 155786 120934
rect 156022 120698 191786 120934
rect 192022 120698 227786 120934
rect 228022 120698 263786 120934
rect 264022 120698 299786 120934
rect 300022 120698 335786 120934
rect 336022 120698 371786 120934
rect 372022 120698 407786 120934
rect 408022 120698 443786 120934
rect 444022 120698 479786 120934
rect 480022 120698 515786 120934
rect 516022 120698 551786 120934
rect 552022 120698 591022 120934
rect 591258 120698 592360 120934
rect -8436 120676 592360 120698
rect -7516 120674 -6916 120676
rect 11604 120674 12204 120676
rect 47604 120674 48204 120676
rect 83604 120674 84204 120676
rect 119604 120674 120204 120676
rect 155604 120674 156204 120676
rect 191604 120674 192204 120676
rect 227604 120674 228204 120676
rect 263604 120674 264204 120676
rect 299604 120674 300204 120676
rect 335604 120674 336204 120676
rect 371604 120674 372204 120676
rect 407604 120674 408204 120676
rect 443604 120674 444204 120676
rect 479604 120674 480204 120676
rect 515604 120674 516204 120676
rect 551604 120674 552204 120676
rect 590840 120674 591440 120676
rect -5676 117676 -5076 117678
rect 8004 117676 8604 117678
rect 44004 117676 44604 117678
rect 80004 117676 80604 117678
rect 116004 117676 116604 117678
rect 152004 117676 152604 117678
rect 188004 117676 188604 117678
rect 224004 117676 224604 117678
rect 260004 117676 260604 117678
rect 296004 117676 296604 117678
rect 332004 117676 332604 117678
rect 368004 117676 368604 117678
rect 404004 117676 404604 117678
rect 440004 117676 440604 117678
rect 476004 117676 476604 117678
rect 512004 117676 512604 117678
rect 548004 117676 548604 117678
rect 589000 117676 589600 117678
rect -6596 117654 590520 117676
rect -6596 117418 -5494 117654
rect -5258 117418 8186 117654
rect 8422 117418 44186 117654
rect 44422 117418 80186 117654
rect 80422 117418 116186 117654
rect 116422 117418 152186 117654
rect 152422 117418 188186 117654
rect 188422 117418 224186 117654
rect 224422 117418 260186 117654
rect 260422 117418 296186 117654
rect 296422 117418 332186 117654
rect 332422 117418 368186 117654
rect 368422 117418 404186 117654
rect 404422 117418 440186 117654
rect 440422 117418 476186 117654
rect 476422 117418 512186 117654
rect 512422 117418 548186 117654
rect 548422 117418 589182 117654
rect 589418 117418 590520 117654
rect -6596 117334 590520 117418
rect -6596 117098 -5494 117334
rect -5258 117098 8186 117334
rect 8422 117098 44186 117334
rect 44422 117098 80186 117334
rect 80422 117098 116186 117334
rect 116422 117098 152186 117334
rect 152422 117098 188186 117334
rect 188422 117098 224186 117334
rect 224422 117098 260186 117334
rect 260422 117098 296186 117334
rect 296422 117098 332186 117334
rect 332422 117098 368186 117334
rect 368422 117098 404186 117334
rect 404422 117098 440186 117334
rect 440422 117098 476186 117334
rect 476422 117098 512186 117334
rect 512422 117098 548186 117334
rect 548422 117098 589182 117334
rect 589418 117098 590520 117334
rect -6596 117076 590520 117098
rect -5676 117074 -5076 117076
rect 8004 117074 8604 117076
rect 44004 117074 44604 117076
rect 80004 117074 80604 117076
rect 116004 117074 116604 117076
rect 152004 117074 152604 117076
rect 188004 117074 188604 117076
rect 224004 117074 224604 117076
rect 260004 117074 260604 117076
rect 296004 117074 296604 117076
rect 332004 117074 332604 117076
rect 368004 117074 368604 117076
rect 404004 117074 404604 117076
rect 440004 117074 440604 117076
rect 476004 117074 476604 117076
rect 512004 117074 512604 117076
rect 548004 117074 548604 117076
rect 589000 117074 589600 117076
rect -3836 114076 -3236 114078
rect 4404 114076 5004 114078
rect 40404 114076 41004 114078
rect 76404 114076 77004 114078
rect 112404 114076 113004 114078
rect 148404 114076 149004 114078
rect 184404 114076 185004 114078
rect 220404 114076 221004 114078
rect 256404 114076 257004 114078
rect 292404 114076 293004 114078
rect 328404 114076 329004 114078
rect 364404 114076 365004 114078
rect 400404 114076 401004 114078
rect 436404 114076 437004 114078
rect 472404 114076 473004 114078
rect 508404 114076 509004 114078
rect 544404 114076 545004 114078
rect 580404 114076 581004 114078
rect 587160 114076 587760 114078
rect -4756 114054 588680 114076
rect -4756 113818 -3654 114054
rect -3418 113818 4586 114054
rect 4822 113818 40586 114054
rect 40822 113818 76586 114054
rect 76822 113818 112586 114054
rect 112822 113818 148586 114054
rect 148822 113818 184586 114054
rect 184822 113818 220586 114054
rect 220822 113818 256586 114054
rect 256822 113818 292586 114054
rect 292822 113818 328586 114054
rect 328822 113818 364586 114054
rect 364822 113818 400586 114054
rect 400822 113818 436586 114054
rect 436822 113818 472586 114054
rect 472822 113818 508586 114054
rect 508822 113818 544586 114054
rect 544822 113818 580586 114054
rect 580822 113818 587342 114054
rect 587578 113818 588680 114054
rect -4756 113734 588680 113818
rect -4756 113498 -3654 113734
rect -3418 113498 4586 113734
rect 4822 113498 40586 113734
rect 40822 113498 76586 113734
rect 76822 113498 112586 113734
rect 112822 113498 148586 113734
rect 148822 113498 184586 113734
rect 184822 113498 220586 113734
rect 220822 113498 256586 113734
rect 256822 113498 292586 113734
rect 292822 113498 328586 113734
rect 328822 113498 364586 113734
rect 364822 113498 400586 113734
rect 400822 113498 436586 113734
rect 436822 113498 472586 113734
rect 472822 113498 508586 113734
rect 508822 113498 544586 113734
rect 544822 113498 580586 113734
rect 580822 113498 587342 113734
rect 587578 113498 588680 113734
rect -4756 113476 588680 113498
rect -3836 113474 -3236 113476
rect 4404 113474 5004 113476
rect 40404 113474 41004 113476
rect 76404 113474 77004 113476
rect 112404 113474 113004 113476
rect 148404 113474 149004 113476
rect 184404 113474 185004 113476
rect 220404 113474 221004 113476
rect 256404 113474 257004 113476
rect 292404 113474 293004 113476
rect 328404 113474 329004 113476
rect 364404 113474 365004 113476
rect 400404 113474 401004 113476
rect 436404 113474 437004 113476
rect 472404 113474 473004 113476
rect 508404 113474 509004 113476
rect 544404 113474 545004 113476
rect 580404 113474 581004 113476
rect 587160 113474 587760 113476
rect -1996 110476 -1396 110478
rect 804 110476 1404 110478
rect 36804 110476 37404 110478
rect 72804 110476 73404 110478
rect 108804 110476 109404 110478
rect 144804 110476 145404 110478
rect 180804 110476 181404 110478
rect 216804 110476 217404 110478
rect 252804 110476 253404 110478
rect 288804 110476 289404 110478
rect 324804 110476 325404 110478
rect 360804 110476 361404 110478
rect 396804 110476 397404 110478
rect 432804 110476 433404 110478
rect 468804 110476 469404 110478
rect 504804 110476 505404 110478
rect 540804 110476 541404 110478
rect 576804 110476 577404 110478
rect 585320 110476 585920 110478
rect -2916 110454 586840 110476
rect -2916 110218 -1814 110454
rect -1578 110218 986 110454
rect 1222 110218 36986 110454
rect 37222 110218 72986 110454
rect 73222 110218 108986 110454
rect 109222 110218 144986 110454
rect 145222 110218 180986 110454
rect 181222 110218 216986 110454
rect 217222 110218 252986 110454
rect 253222 110218 288986 110454
rect 289222 110218 324986 110454
rect 325222 110218 360986 110454
rect 361222 110218 396986 110454
rect 397222 110218 432986 110454
rect 433222 110218 468986 110454
rect 469222 110218 504986 110454
rect 505222 110218 540986 110454
rect 541222 110218 576986 110454
rect 577222 110218 585502 110454
rect 585738 110218 586840 110454
rect -2916 110134 586840 110218
rect -2916 109898 -1814 110134
rect -1578 109898 986 110134
rect 1222 109898 36986 110134
rect 37222 109898 72986 110134
rect 73222 109898 108986 110134
rect 109222 109898 144986 110134
rect 145222 109898 180986 110134
rect 181222 109898 216986 110134
rect 217222 109898 252986 110134
rect 253222 109898 288986 110134
rect 289222 109898 324986 110134
rect 325222 109898 360986 110134
rect 361222 109898 396986 110134
rect 397222 109898 432986 110134
rect 433222 109898 468986 110134
rect 469222 109898 504986 110134
rect 505222 109898 540986 110134
rect 541222 109898 576986 110134
rect 577222 109898 585502 110134
rect 585738 109898 586840 110134
rect -2916 109876 586840 109898
rect -1996 109874 -1396 109876
rect 804 109874 1404 109876
rect 36804 109874 37404 109876
rect 72804 109874 73404 109876
rect 108804 109874 109404 109876
rect 144804 109874 145404 109876
rect 180804 109874 181404 109876
rect 216804 109874 217404 109876
rect 252804 109874 253404 109876
rect 288804 109874 289404 109876
rect 324804 109874 325404 109876
rect 360804 109874 361404 109876
rect 396804 109874 397404 109876
rect 432804 109874 433404 109876
rect 468804 109874 469404 109876
rect 504804 109874 505404 109876
rect 540804 109874 541404 109876
rect 576804 109874 577404 109876
rect 585320 109874 585920 109876
rect -8436 103276 -7836 103278
rect 29604 103276 30204 103278
rect 65604 103276 66204 103278
rect 101604 103276 102204 103278
rect 137604 103276 138204 103278
rect 173604 103276 174204 103278
rect 209604 103276 210204 103278
rect 245604 103276 246204 103278
rect 281604 103276 282204 103278
rect 317604 103276 318204 103278
rect 353604 103276 354204 103278
rect 389604 103276 390204 103278
rect 425604 103276 426204 103278
rect 461604 103276 462204 103278
rect 497604 103276 498204 103278
rect 533604 103276 534204 103278
rect 569604 103276 570204 103278
rect 591760 103276 592360 103278
rect -8436 103254 592360 103276
rect -8436 103018 -8254 103254
rect -8018 103018 29786 103254
rect 30022 103018 65786 103254
rect 66022 103018 101786 103254
rect 102022 103018 137786 103254
rect 138022 103018 173786 103254
rect 174022 103018 209786 103254
rect 210022 103018 245786 103254
rect 246022 103018 281786 103254
rect 282022 103018 317786 103254
rect 318022 103018 353786 103254
rect 354022 103018 389786 103254
rect 390022 103018 425786 103254
rect 426022 103018 461786 103254
rect 462022 103018 497786 103254
rect 498022 103018 533786 103254
rect 534022 103018 569786 103254
rect 570022 103018 591942 103254
rect 592178 103018 592360 103254
rect -8436 102934 592360 103018
rect -8436 102698 -8254 102934
rect -8018 102698 29786 102934
rect 30022 102698 65786 102934
rect 66022 102698 101786 102934
rect 102022 102698 137786 102934
rect 138022 102698 173786 102934
rect 174022 102698 209786 102934
rect 210022 102698 245786 102934
rect 246022 102698 281786 102934
rect 282022 102698 317786 102934
rect 318022 102698 353786 102934
rect 354022 102698 389786 102934
rect 390022 102698 425786 102934
rect 426022 102698 461786 102934
rect 462022 102698 497786 102934
rect 498022 102698 533786 102934
rect 534022 102698 569786 102934
rect 570022 102698 591942 102934
rect 592178 102698 592360 102934
rect -8436 102676 592360 102698
rect -8436 102674 -7836 102676
rect 29604 102674 30204 102676
rect 65604 102674 66204 102676
rect 101604 102674 102204 102676
rect 137604 102674 138204 102676
rect 173604 102674 174204 102676
rect 209604 102674 210204 102676
rect 245604 102674 246204 102676
rect 281604 102674 282204 102676
rect 317604 102674 318204 102676
rect 353604 102674 354204 102676
rect 389604 102674 390204 102676
rect 425604 102674 426204 102676
rect 461604 102674 462204 102676
rect 497604 102674 498204 102676
rect 533604 102674 534204 102676
rect 569604 102674 570204 102676
rect 591760 102674 592360 102676
rect -6596 99676 -5996 99678
rect 26004 99676 26604 99678
rect 62004 99676 62604 99678
rect 98004 99676 98604 99678
rect 134004 99676 134604 99678
rect 170004 99676 170604 99678
rect 206004 99676 206604 99678
rect 242004 99676 242604 99678
rect 278004 99676 278604 99678
rect 314004 99676 314604 99678
rect 350004 99676 350604 99678
rect 386004 99676 386604 99678
rect 422004 99676 422604 99678
rect 458004 99676 458604 99678
rect 494004 99676 494604 99678
rect 530004 99676 530604 99678
rect 566004 99676 566604 99678
rect 589920 99676 590520 99678
rect -6596 99654 590520 99676
rect -6596 99418 -6414 99654
rect -6178 99418 26186 99654
rect 26422 99418 62186 99654
rect 62422 99418 98186 99654
rect 98422 99418 134186 99654
rect 134422 99418 170186 99654
rect 170422 99418 206186 99654
rect 206422 99418 242186 99654
rect 242422 99418 278186 99654
rect 278422 99418 314186 99654
rect 314422 99418 350186 99654
rect 350422 99418 386186 99654
rect 386422 99418 422186 99654
rect 422422 99418 458186 99654
rect 458422 99418 494186 99654
rect 494422 99418 530186 99654
rect 530422 99418 566186 99654
rect 566422 99418 590102 99654
rect 590338 99418 590520 99654
rect -6596 99334 590520 99418
rect -6596 99098 -6414 99334
rect -6178 99098 26186 99334
rect 26422 99098 62186 99334
rect 62422 99098 98186 99334
rect 98422 99098 134186 99334
rect 134422 99098 170186 99334
rect 170422 99098 206186 99334
rect 206422 99098 242186 99334
rect 242422 99098 278186 99334
rect 278422 99098 314186 99334
rect 314422 99098 350186 99334
rect 350422 99098 386186 99334
rect 386422 99098 422186 99334
rect 422422 99098 458186 99334
rect 458422 99098 494186 99334
rect 494422 99098 530186 99334
rect 530422 99098 566186 99334
rect 566422 99098 590102 99334
rect 590338 99098 590520 99334
rect -6596 99076 590520 99098
rect -6596 99074 -5996 99076
rect 26004 99074 26604 99076
rect 62004 99074 62604 99076
rect 98004 99074 98604 99076
rect 134004 99074 134604 99076
rect 170004 99074 170604 99076
rect 206004 99074 206604 99076
rect 242004 99074 242604 99076
rect 278004 99074 278604 99076
rect 314004 99074 314604 99076
rect 350004 99074 350604 99076
rect 386004 99074 386604 99076
rect 422004 99074 422604 99076
rect 458004 99074 458604 99076
rect 494004 99074 494604 99076
rect 530004 99074 530604 99076
rect 566004 99074 566604 99076
rect 589920 99074 590520 99076
rect -4756 96076 -4156 96078
rect 22404 96076 23004 96078
rect 58404 96076 59004 96078
rect 94404 96076 95004 96078
rect 130404 96076 131004 96078
rect 166404 96076 167004 96078
rect 202404 96076 203004 96078
rect 238404 96076 239004 96078
rect 274404 96076 275004 96078
rect 310404 96076 311004 96078
rect 346404 96076 347004 96078
rect 382404 96076 383004 96078
rect 418404 96076 419004 96078
rect 454404 96076 455004 96078
rect 490404 96076 491004 96078
rect 526404 96076 527004 96078
rect 562404 96076 563004 96078
rect 588080 96076 588680 96078
rect -4756 96054 588680 96076
rect -4756 95818 -4574 96054
rect -4338 95818 22586 96054
rect 22822 95818 58586 96054
rect 58822 95818 94586 96054
rect 94822 95818 130586 96054
rect 130822 95818 166586 96054
rect 166822 95818 202586 96054
rect 202822 95818 238586 96054
rect 238822 95818 274586 96054
rect 274822 95818 310586 96054
rect 310822 95818 346586 96054
rect 346822 95818 382586 96054
rect 382822 95818 418586 96054
rect 418822 95818 454586 96054
rect 454822 95818 490586 96054
rect 490822 95818 526586 96054
rect 526822 95818 562586 96054
rect 562822 95818 588262 96054
rect 588498 95818 588680 96054
rect -4756 95734 588680 95818
rect -4756 95498 -4574 95734
rect -4338 95498 22586 95734
rect 22822 95498 58586 95734
rect 58822 95498 94586 95734
rect 94822 95498 130586 95734
rect 130822 95498 166586 95734
rect 166822 95498 202586 95734
rect 202822 95498 238586 95734
rect 238822 95498 274586 95734
rect 274822 95498 310586 95734
rect 310822 95498 346586 95734
rect 346822 95498 382586 95734
rect 382822 95498 418586 95734
rect 418822 95498 454586 95734
rect 454822 95498 490586 95734
rect 490822 95498 526586 95734
rect 526822 95498 562586 95734
rect 562822 95498 588262 95734
rect 588498 95498 588680 95734
rect -4756 95476 588680 95498
rect -4756 95474 -4156 95476
rect 22404 95474 23004 95476
rect 58404 95474 59004 95476
rect 94404 95474 95004 95476
rect 130404 95474 131004 95476
rect 166404 95474 167004 95476
rect 202404 95474 203004 95476
rect 238404 95474 239004 95476
rect 274404 95474 275004 95476
rect 310404 95474 311004 95476
rect 346404 95474 347004 95476
rect 382404 95474 383004 95476
rect 418404 95474 419004 95476
rect 454404 95474 455004 95476
rect 490404 95474 491004 95476
rect 526404 95474 527004 95476
rect 562404 95474 563004 95476
rect 588080 95474 588680 95476
rect -2916 92476 -2316 92478
rect 18804 92476 19404 92478
rect 54804 92476 55404 92478
rect 90804 92476 91404 92478
rect 126804 92476 127404 92478
rect 162804 92476 163404 92478
rect 198804 92476 199404 92478
rect 234804 92476 235404 92478
rect 270804 92476 271404 92478
rect 306804 92476 307404 92478
rect 342804 92476 343404 92478
rect 378804 92476 379404 92478
rect 414804 92476 415404 92478
rect 450804 92476 451404 92478
rect 486804 92476 487404 92478
rect 522804 92476 523404 92478
rect 558804 92476 559404 92478
rect 586240 92476 586840 92478
rect -2916 92454 586840 92476
rect -2916 92218 -2734 92454
rect -2498 92218 18986 92454
rect 19222 92218 54986 92454
rect 55222 92218 90986 92454
rect 91222 92218 126986 92454
rect 127222 92218 162986 92454
rect 163222 92218 198986 92454
rect 199222 92218 234986 92454
rect 235222 92218 270986 92454
rect 271222 92218 306986 92454
rect 307222 92218 342986 92454
rect 343222 92218 378986 92454
rect 379222 92218 414986 92454
rect 415222 92218 450986 92454
rect 451222 92218 486986 92454
rect 487222 92218 522986 92454
rect 523222 92218 558986 92454
rect 559222 92218 586422 92454
rect 586658 92218 586840 92454
rect -2916 92134 586840 92218
rect -2916 91898 -2734 92134
rect -2498 91898 18986 92134
rect 19222 91898 54986 92134
rect 55222 91898 90986 92134
rect 91222 91898 126986 92134
rect 127222 91898 162986 92134
rect 163222 91898 198986 92134
rect 199222 91898 234986 92134
rect 235222 91898 270986 92134
rect 271222 91898 306986 92134
rect 307222 91898 342986 92134
rect 343222 91898 378986 92134
rect 379222 91898 414986 92134
rect 415222 91898 450986 92134
rect 451222 91898 486986 92134
rect 487222 91898 522986 92134
rect 523222 91898 558986 92134
rect 559222 91898 586422 92134
rect 586658 91898 586840 92134
rect -2916 91876 586840 91898
rect -2916 91874 -2316 91876
rect 18804 91874 19404 91876
rect 54804 91874 55404 91876
rect 90804 91874 91404 91876
rect 126804 91874 127404 91876
rect 162804 91874 163404 91876
rect 198804 91874 199404 91876
rect 234804 91874 235404 91876
rect 270804 91874 271404 91876
rect 306804 91874 307404 91876
rect 342804 91874 343404 91876
rect 378804 91874 379404 91876
rect 414804 91874 415404 91876
rect 450804 91874 451404 91876
rect 486804 91874 487404 91876
rect 522804 91874 523404 91876
rect 558804 91874 559404 91876
rect 586240 91874 586840 91876
rect -7516 85276 -6916 85278
rect 11604 85276 12204 85278
rect 47604 85276 48204 85278
rect 83604 85276 84204 85278
rect 119604 85276 120204 85278
rect 155604 85276 156204 85278
rect 191604 85276 192204 85278
rect 227604 85276 228204 85278
rect 263604 85276 264204 85278
rect 299604 85276 300204 85278
rect 335604 85276 336204 85278
rect 371604 85276 372204 85278
rect 407604 85276 408204 85278
rect 443604 85276 444204 85278
rect 479604 85276 480204 85278
rect 515604 85276 516204 85278
rect 551604 85276 552204 85278
rect 590840 85276 591440 85278
rect -8436 85254 592360 85276
rect -8436 85018 -7334 85254
rect -7098 85018 11786 85254
rect 12022 85018 47786 85254
rect 48022 85018 83786 85254
rect 84022 85018 119786 85254
rect 120022 85018 155786 85254
rect 156022 85018 191786 85254
rect 192022 85018 227786 85254
rect 228022 85018 263786 85254
rect 264022 85018 299786 85254
rect 300022 85018 335786 85254
rect 336022 85018 371786 85254
rect 372022 85018 407786 85254
rect 408022 85018 443786 85254
rect 444022 85018 479786 85254
rect 480022 85018 515786 85254
rect 516022 85018 551786 85254
rect 552022 85018 591022 85254
rect 591258 85018 592360 85254
rect -8436 84934 592360 85018
rect -8436 84698 -7334 84934
rect -7098 84698 11786 84934
rect 12022 84698 47786 84934
rect 48022 84698 83786 84934
rect 84022 84698 119786 84934
rect 120022 84698 155786 84934
rect 156022 84698 191786 84934
rect 192022 84698 227786 84934
rect 228022 84698 263786 84934
rect 264022 84698 299786 84934
rect 300022 84698 335786 84934
rect 336022 84698 371786 84934
rect 372022 84698 407786 84934
rect 408022 84698 443786 84934
rect 444022 84698 479786 84934
rect 480022 84698 515786 84934
rect 516022 84698 551786 84934
rect 552022 84698 591022 84934
rect 591258 84698 592360 84934
rect -8436 84676 592360 84698
rect -7516 84674 -6916 84676
rect 11604 84674 12204 84676
rect 47604 84674 48204 84676
rect 83604 84674 84204 84676
rect 119604 84674 120204 84676
rect 155604 84674 156204 84676
rect 191604 84674 192204 84676
rect 227604 84674 228204 84676
rect 263604 84674 264204 84676
rect 299604 84674 300204 84676
rect 335604 84674 336204 84676
rect 371604 84674 372204 84676
rect 407604 84674 408204 84676
rect 443604 84674 444204 84676
rect 479604 84674 480204 84676
rect 515604 84674 516204 84676
rect 551604 84674 552204 84676
rect 590840 84674 591440 84676
rect -5676 81676 -5076 81678
rect 8004 81676 8604 81678
rect 44004 81676 44604 81678
rect 80004 81676 80604 81678
rect 116004 81676 116604 81678
rect 152004 81676 152604 81678
rect 188004 81676 188604 81678
rect 224004 81676 224604 81678
rect 260004 81676 260604 81678
rect 296004 81676 296604 81678
rect 332004 81676 332604 81678
rect 368004 81676 368604 81678
rect 404004 81676 404604 81678
rect 440004 81676 440604 81678
rect 476004 81676 476604 81678
rect 512004 81676 512604 81678
rect 548004 81676 548604 81678
rect 589000 81676 589600 81678
rect -6596 81654 590520 81676
rect -6596 81418 -5494 81654
rect -5258 81418 8186 81654
rect 8422 81418 44186 81654
rect 44422 81418 80186 81654
rect 80422 81418 116186 81654
rect 116422 81418 152186 81654
rect 152422 81418 188186 81654
rect 188422 81418 224186 81654
rect 224422 81418 260186 81654
rect 260422 81418 296186 81654
rect 296422 81418 332186 81654
rect 332422 81418 368186 81654
rect 368422 81418 404186 81654
rect 404422 81418 440186 81654
rect 440422 81418 476186 81654
rect 476422 81418 512186 81654
rect 512422 81418 548186 81654
rect 548422 81418 589182 81654
rect 589418 81418 590520 81654
rect -6596 81334 590520 81418
rect -6596 81098 -5494 81334
rect -5258 81098 8186 81334
rect 8422 81098 44186 81334
rect 44422 81098 80186 81334
rect 80422 81098 116186 81334
rect 116422 81098 152186 81334
rect 152422 81098 188186 81334
rect 188422 81098 224186 81334
rect 224422 81098 260186 81334
rect 260422 81098 296186 81334
rect 296422 81098 332186 81334
rect 332422 81098 368186 81334
rect 368422 81098 404186 81334
rect 404422 81098 440186 81334
rect 440422 81098 476186 81334
rect 476422 81098 512186 81334
rect 512422 81098 548186 81334
rect 548422 81098 589182 81334
rect 589418 81098 590520 81334
rect -6596 81076 590520 81098
rect -5676 81074 -5076 81076
rect 8004 81074 8604 81076
rect 44004 81074 44604 81076
rect 80004 81074 80604 81076
rect 116004 81074 116604 81076
rect 152004 81074 152604 81076
rect 188004 81074 188604 81076
rect 224004 81074 224604 81076
rect 260004 81074 260604 81076
rect 296004 81074 296604 81076
rect 332004 81074 332604 81076
rect 368004 81074 368604 81076
rect 404004 81074 404604 81076
rect 440004 81074 440604 81076
rect 476004 81074 476604 81076
rect 512004 81074 512604 81076
rect 548004 81074 548604 81076
rect 589000 81074 589600 81076
rect -3836 78076 -3236 78078
rect 4404 78076 5004 78078
rect 40404 78076 41004 78078
rect 76404 78076 77004 78078
rect 112404 78076 113004 78078
rect 148404 78076 149004 78078
rect 184404 78076 185004 78078
rect 220404 78076 221004 78078
rect 256404 78076 257004 78078
rect 292404 78076 293004 78078
rect 328404 78076 329004 78078
rect 364404 78076 365004 78078
rect 400404 78076 401004 78078
rect 436404 78076 437004 78078
rect 472404 78076 473004 78078
rect 508404 78076 509004 78078
rect 544404 78076 545004 78078
rect 580404 78076 581004 78078
rect 587160 78076 587760 78078
rect -4756 78054 588680 78076
rect -4756 77818 -3654 78054
rect -3418 77818 4586 78054
rect 4822 77818 40586 78054
rect 40822 77818 76586 78054
rect 76822 77818 112586 78054
rect 112822 77818 148586 78054
rect 148822 77818 184586 78054
rect 184822 77818 220586 78054
rect 220822 77818 256586 78054
rect 256822 77818 292586 78054
rect 292822 77818 328586 78054
rect 328822 77818 364586 78054
rect 364822 77818 400586 78054
rect 400822 77818 436586 78054
rect 436822 77818 472586 78054
rect 472822 77818 508586 78054
rect 508822 77818 544586 78054
rect 544822 77818 580586 78054
rect 580822 77818 587342 78054
rect 587578 77818 588680 78054
rect -4756 77734 588680 77818
rect -4756 77498 -3654 77734
rect -3418 77498 4586 77734
rect 4822 77498 40586 77734
rect 40822 77498 76586 77734
rect 76822 77498 112586 77734
rect 112822 77498 148586 77734
rect 148822 77498 184586 77734
rect 184822 77498 220586 77734
rect 220822 77498 256586 77734
rect 256822 77498 292586 77734
rect 292822 77498 328586 77734
rect 328822 77498 364586 77734
rect 364822 77498 400586 77734
rect 400822 77498 436586 77734
rect 436822 77498 472586 77734
rect 472822 77498 508586 77734
rect 508822 77498 544586 77734
rect 544822 77498 580586 77734
rect 580822 77498 587342 77734
rect 587578 77498 588680 77734
rect -4756 77476 588680 77498
rect -3836 77474 -3236 77476
rect 4404 77474 5004 77476
rect 40404 77474 41004 77476
rect 76404 77474 77004 77476
rect 112404 77474 113004 77476
rect 148404 77474 149004 77476
rect 184404 77474 185004 77476
rect 220404 77474 221004 77476
rect 256404 77474 257004 77476
rect 292404 77474 293004 77476
rect 328404 77474 329004 77476
rect 364404 77474 365004 77476
rect 400404 77474 401004 77476
rect 436404 77474 437004 77476
rect 472404 77474 473004 77476
rect 508404 77474 509004 77476
rect 544404 77474 545004 77476
rect 580404 77474 581004 77476
rect 587160 77474 587760 77476
rect -1996 74476 -1396 74478
rect 804 74476 1404 74478
rect 36804 74476 37404 74478
rect 72804 74476 73404 74478
rect 108804 74476 109404 74478
rect 144804 74476 145404 74478
rect 180804 74476 181404 74478
rect 216804 74476 217404 74478
rect 252804 74476 253404 74478
rect 288804 74476 289404 74478
rect 324804 74476 325404 74478
rect 360804 74476 361404 74478
rect 396804 74476 397404 74478
rect 432804 74476 433404 74478
rect 468804 74476 469404 74478
rect 504804 74476 505404 74478
rect 540804 74476 541404 74478
rect 576804 74476 577404 74478
rect 585320 74476 585920 74478
rect -2916 74454 586840 74476
rect -2916 74218 -1814 74454
rect -1578 74218 986 74454
rect 1222 74218 36986 74454
rect 37222 74218 72986 74454
rect 73222 74218 108986 74454
rect 109222 74218 144986 74454
rect 145222 74218 180986 74454
rect 181222 74218 216986 74454
rect 217222 74218 252986 74454
rect 253222 74218 288986 74454
rect 289222 74218 324986 74454
rect 325222 74218 360986 74454
rect 361222 74218 396986 74454
rect 397222 74218 432986 74454
rect 433222 74218 468986 74454
rect 469222 74218 504986 74454
rect 505222 74218 540986 74454
rect 541222 74218 576986 74454
rect 577222 74218 585502 74454
rect 585738 74218 586840 74454
rect -2916 74134 586840 74218
rect -2916 73898 -1814 74134
rect -1578 73898 986 74134
rect 1222 73898 36986 74134
rect 37222 73898 72986 74134
rect 73222 73898 108986 74134
rect 109222 73898 144986 74134
rect 145222 73898 180986 74134
rect 181222 73898 216986 74134
rect 217222 73898 252986 74134
rect 253222 73898 288986 74134
rect 289222 73898 324986 74134
rect 325222 73898 360986 74134
rect 361222 73898 396986 74134
rect 397222 73898 432986 74134
rect 433222 73898 468986 74134
rect 469222 73898 504986 74134
rect 505222 73898 540986 74134
rect 541222 73898 576986 74134
rect 577222 73898 585502 74134
rect 585738 73898 586840 74134
rect -2916 73876 586840 73898
rect -1996 73874 -1396 73876
rect 804 73874 1404 73876
rect 36804 73874 37404 73876
rect 72804 73874 73404 73876
rect 108804 73874 109404 73876
rect 144804 73874 145404 73876
rect 180804 73874 181404 73876
rect 216804 73874 217404 73876
rect 252804 73874 253404 73876
rect 288804 73874 289404 73876
rect 324804 73874 325404 73876
rect 360804 73874 361404 73876
rect 396804 73874 397404 73876
rect 432804 73874 433404 73876
rect 468804 73874 469404 73876
rect 504804 73874 505404 73876
rect 540804 73874 541404 73876
rect 576804 73874 577404 73876
rect 585320 73874 585920 73876
rect -8436 67276 -7836 67278
rect 29604 67276 30204 67278
rect 65604 67276 66204 67278
rect 101604 67276 102204 67278
rect 137604 67276 138204 67278
rect 173604 67276 174204 67278
rect 209604 67276 210204 67278
rect 245604 67276 246204 67278
rect 281604 67276 282204 67278
rect 317604 67276 318204 67278
rect 353604 67276 354204 67278
rect 389604 67276 390204 67278
rect 425604 67276 426204 67278
rect 461604 67276 462204 67278
rect 497604 67276 498204 67278
rect 533604 67276 534204 67278
rect 569604 67276 570204 67278
rect 591760 67276 592360 67278
rect -8436 67254 592360 67276
rect -8436 67018 -8254 67254
rect -8018 67018 29786 67254
rect 30022 67018 65786 67254
rect 66022 67018 101786 67254
rect 102022 67018 137786 67254
rect 138022 67018 173786 67254
rect 174022 67018 209786 67254
rect 210022 67018 245786 67254
rect 246022 67018 281786 67254
rect 282022 67018 317786 67254
rect 318022 67018 353786 67254
rect 354022 67018 389786 67254
rect 390022 67018 425786 67254
rect 426022 67018 461786 67254
rect 462022 67018 497786 67254
rect 498022 67018 533786 67254
rect 534022 67018 569786 67254
rect 570022 67018 591942 67254
rect 592178 67018 592360 67254
rect -8436 66934 592360 67018
rect -8436 66698 -8254 66934
rect -8018 66698 29786 66934
rect 30022 66698 65786 66934
rect 66022 66698 101786 66934
rect 102022 66698 137786 66934
rect 138022 66698 173786 66934
rect 174022 66698 209786 66934
rect 210022 66698 245786 66934
rect 246022 66698 281786 66934
rect 282022 66698 317786 66934
rect 318022 66698 353786 66934
rect 354022 66698 389786 66934
rect 390022 66698 425786 66934
rect 426022 66698 461786 66934
rect 462022 66698 497786 66934
rect 498022 66698 533786 66934
rect 534022 66698 569786 66934
rect 570022 66698 591942 66934
rect 592178 66698 592360 66934
rect -8436 66676 592360 66698
rect -8436 66674 -7836 66676
rect 29604 66674 30204 66676
rect 65604 66674 66204 66676
rect 101604 66674 102204 66676
rect 137604 66674 138204 66676
rect 173604 66674 174204 66676
rect 209604 66674 210204 66676
rect 245604 66674 246204 66676
rect 281604 66674 282204 66676
rect 317604 66674 318204 66676
rect 353604 66674 354204 66676
rect 389604 66674 390204 66676
rect 425604 66674 426204 66676
rect 461604 66674 462204 66676
rect 497604 66674 498204 66676
rect 533604 66674 534204 66676
rect 569604 66674 570204 66676
rect 591760 66674 592360 66676
rect -6596 63676 -5996 63678
rect 26004 63676 26604 63678
rect 62004 63676 62604 63678
rect 98004 63676 98604 63678
rect 134004 63676 134604 63678
rect 170004 63676 170604 63678
rect 206004 63676 206604 63678
rect 242004 63676 242604 63678
rect 278004 63676 278604 63678
rect 314004 63676 314604 63678
rect 350004 63676 350604 63678
rect 386004 63676 386604 63678
rect 422004 63676 422604 63678
rect 458004 63676 458604 63678
rect 494004 63676 494604 63678
rect 530004 63676 530604 63678
rect 566004 63676 566604 63678
rect 589920 63676 590520 63678
rect -6596 63654 590520 63676
rect -6596 63418 -6414 63654
rect -6178 63418 26186 63654
rect 26422 63418 62186 63654
rect 62422 63418 98186 63654
rect 98422 63418 134186 63654
rect 134422 63418 170186 63654
rect 170422 63418 206186 63654
rect 206422 63418 242186 63654
rect 242422 63418 278186 63654
rect 278422 63418 314186 63654
rect 314422 63418 350186 63654
rect 350422 63418 386186 63654
rect 386422 63418 422186 63654
rect 422422 63418 458186 63654
rect 458422 63418 494186 63654
rect 494422 63418 530186 63654
rect 530422 63418 566186 63654
rect 566422 63418 590102 63654
rect 590338 63418 590520 63654
rect -6596 63334 590520 63418
rect -6596 63098 -6414 63334
rect -6178 63098 26186 63334
rect 26422 63098 62186 63334
rect 62422 63098 98186 63334
rect 98422 63098 134186 63334
rect 134422 63098 170186 63334
rect 170422 63098 206186 63334
rect 206422 63098 242186 63334
rect 242422 63098 278186 63334
rect 278422 63098 314186 63334
rect 314422 63098 350186 63334
rect 350422 63098 386186 63334
rect 386422 63098 422186 63334
rect 422422 63098 458186 63334
rect 458422 63098 494186 63334
rect 494422 63098 530186 63334
rect 530422 63098 566186 63334
rect 566422 63098 590102 63334
rect 590338 63098 590520 63334
rect -6596 63076 590520 63098
rect -6596 63074 -5996 63076
rect 26004 63074 26604 63076
rect 62004 63074 62604 63076
rect 98004 63074 98604 63076
rect 134004 63074 134604 63076
rect 170004 63074 170604 63076
rect 206004 63074 206604 63076
rect 242004 63074 242604 63076
rect 278004 63074 278604 63076
rect 314004 63074 314604 63076
rect 350004 63074 350604 63076
rect 386004 63074 386604 63076
rect 422004 63074 422604 63076
rect 458004 63074 458604 63076
rect 494004 63074 494604 63076
rect 530004 63074 530604 63076
rect 566004 63074 566604 63076
rect 589920 63074 590520 63076
rect -4756 60076 -4156 60078
rect 22404 60076 23004 60078
rect 58404 60076 59004 60078
rect 94404 60076 95004 60078
rect 130404 60076 131004 60078
rect 166404 60076 167004 60078
rect 202404 60076 203004 60078
rect 238404 60076 239004 60078
rect 274404 60076 275004 60078
rect 310404 60076 311004 60078
rect 346404 60076 347004 60078
rect 382404 60076 383004 60078
rect 418404 60076 419004 60078
rect 454404 60076 455004 60078
rect 490404 60076 491004 60078
rect 526404 60076 527004 60078
rect 562404 60076 563004 60078
rect 588080 60076 588680 60078
rect -4756 60054 588680 60076
rect -4756 59818 -4574 60054
rect -4338 59818 22586 60054
rect 22822 59818 58586 60054
rect 58822 59818 94586 60054
rect 94822 59818 130586 60054
rect 130822 59818 166586 60054
rect 166822 59818 202586 60054
rect 202822 59818 238586 60054
rect 238822 59818 274586 60054
rect 274822 59818 310586 60054
rect 310822 59818 346586 60054
rect 346822 59818 382586 60054
rect 382822 59818 418586 60054
rect 418822 59818 454586 60054
rect 454822 59818 490586 60054
rect 490822 59818 526586 60054
rect 526822 59818 562586 60054
rect 562822 59818 588262 60054
rect 588498 59818 588680 60054
rect -4756 59734 588680 59818
rect -4756 59498 -4574 59734
rect -4338 59498 22586 59734
rect 22822 59498 58586 59734
rect 58822 59498 94586 59734
rect 94822 59498 130586 59734
rect 130822 59498 166586 59734
rect 166822 59498 202586 59734
rect 202822 59498 238586 59734
rect 238822 59498 274586 59734
rect 274822 59498 310586 59734
rect 310822 59498 346586 59734
rect 346822 59498 382586 59734
rect 382822 59498 418586 59734
rect 418822 59498 454586 59734
rect 454822 59498 490586 59734
rect 490822 59498 526586 59734
rect 526822 59498 562586 59734
rect 562822 59498 588262 59734
rect 588498 59498 588680 59734
rect -4756 59476 588680 59498
rect -4756 59474 -4156 59476
rect 22404 59474 23004 59476
rect 58404 59474 59004 59476
rect 94404 59474 95004 59476
rect 130404 59474 131004 59476
rect 166404 59474 167004 59476
rect 202404 59474 203004 59476
rect 238404 59474 239004 59476
rect 274404 59474 275004 59476
rect 310404 59474 311004 59476
rect 346404 59474 347004 59476
rect 382404 59474 383004 59476
rect 418404 59474 419004 59476
rect 454404 59474 455004 59476
rect 490404 59474 491004 59476
rect 526404 59474 527004 59476
rect 562404 59474 563004 59476
rect 588080 59474 588680 59476
rect -2916 56476 -2316 56478
rect 18804 56476 19404 56478
rect 54804 56476 55404 56478
rect 90804 56476 91404 56478
rect 126804 56476 127404 56478
rect 162804 56476 163404 56478
rect 198804 56476 199404 56478
rect 234804 56476 235404 56478
rect 270804 56476 271404 56478
rect 306804 56476 307404 56478
rect 342804 56476 343404 56478
rect 378804 56476 379404 56478
rect 414804 56476 415404 56478
rect 450804 56476 451404 56478
rect 486804 56476 487404 56478
rect 522804 56476 523404 56478
rect 558804 56476 559404 56478
rect 586240 56476 586840 56478
rect -2916 56454 586840 56476
rect -2916 56218 -2734 56454
rect -2498 56218 18986 56454
rect 19222 56218 54986 56454
rect 55222 56218 90986 56454
rect 91222 56218 126986 56454
rect 127222 56218 162986 56454
rect 163222 56218 198986 56454
rect 199222 56218 234986 56454
rect 235222 56218 270986 56454
rect 271222 56218 306986 56454
rect 307222 56218 342986 56454
rect 343222 56218 378986 56454
rect 379222 56218 414986 56454
rect 415222 56218 450986 56454
rect 451222 56218 486986 56454
rect 487222 56218 522986 56454
rect 523222 56218 558986 56454
rect 559222 56218 586422 56454
rect 586658 56218 586840 56454
rect -2916 56134 586840 56218
rect -2916 55898 -2734 56134
rect -2498 55898 18986 56134
rect 19222 55898 54986 56134
rect 55222 55898 90986 56134
rect 91222 55898 126986 56134
rect 127222 55898 162986 56134
rect 163222 55898 198986 56134
rect 199222 55898 234986 56134
rect 235222 55898 270986 56134
rect 271222 55898 306986 56134
rect 307222 55898 342986 56134
rect 343222 55898 378986 56134
rect 379222 55898 414986 56134
rect 415222 55898 450986 56134
rect 451222 55898 486986 56134
rect 487222 55898 522986 56134
rect 523222 55898 558986 56134
rect 559222 55898 586422 56134
rect 586658 55898 586840 56134
rect -2916 55876 586840 55898
rect -2916 55874 -2316 55876
rect 18804 55874 19404 55876
rect 54804 55874 55404 55876
rect 90804 55874 91404 55876
rect 126804 55874 127404 55876
rect 162804 55874 163404 55876
rect 198804 55874 199404 55876
rect 234804 55874 235404 55876
rect 270804 55874 271404 55876
rect 306804 55874 307404 55876
rect 342804 55874 343404 55876
rect 378804 55874 379404 55876
rect 414804 55874 415404 55876
rect 450804 55874 451404 55876
rect 486804 55874 487404 55876
rect 522804 55874 523404 55876
rect 558804 55874 559404 55876
rect 586240 55874 586840 55876
rect -7516 49276 -6916 49278
rect 11604 49276 12204 49278
rect 47604 49276 48204 49278
rect 83604 49276 84204 49278
rect 119604 49276 120204 49278
rect 155604 49276 156204 49278
rect 191604 49276 192204 49278
rect 227604 49276 228204 49278
rect 263604 49276 264204 49278
rect 299604 49276 300204 49278
rect 335604 49276 336204 49278
rect 371604 49276 372204 49278
rect 407604 49276 408204 49278
rect 443604 49276 444204 49278
rect 479604 49276 480204 49278
rect 515604 49276 516204 49278
rect 551604 49276 552204 49278
rect 590840 49276 591440 49278
rect -8436 49254 592360 49276
rect -8436 49018 -7334 49254
rect -7098 49018 11786 49254
rect 12022 49018 47786 49254
rect 48022 49018 83786 49254
rect 84022 49018 119786 49254
rect 120022 49018 155786 49254
rect 156022 49018 191786 49254
rect 192022 49018 227786 49254
rect 228022 49018 263786 49254
rect 264022 49018 299786 49254
rect 300022 49018 335786 49254
rect 336022 49018 371786 49254
rect 372022 49018 407786 49254
rect 408022 49018 443786 49254
rect 444022 49018 479786 49254
rect 480022 49018 515786 49254
rect 516022 49018 551786 49254
rect 552022 49018 591022 49254
rect 591258 49018 592360 49254
rect -8436 48934 592360 49018
rect -8436 48698 -7334 48934
rect -7098 48698 11786 48934
rect 12022 48698 47786 48934
rect 48022 48698 83786 48934
rect 84022 48698 119786 48934
rect 120022 48698 155786 48934
rect 156022 48698 191786 48934
rect 192022 48698 227786 48934
rect 228022 48698 263786 48934
rect 264022 48698 299786 48934
rect 300022 48698 335786 48934
rect 336022 48698 371786 48934
rect 372022 48698 407786 48934
rect 408022 48698 443786 48934
rect 444022 48698 479786 48934
rect 480022 48698 515786 48934
rect 516022 48698 551786 48934
rect 552022 48698 591022 48934
rect 591258 48698 592360 48934
rect -8436 48676 592360 48698
rect -7516 48674 -6916 48676
rect 11604 48674 12204 48676
rect 47604 48674 48204 48676
rect 83604 48674 84204 48676
rect 119604 48674 120204 48676
rect 155604 48674 156204 48676
rect 191604 48674 192204 48676
rect 227604 48674 228204 48676
rect 263604 48674 264204 48676
rect 299604 48674 300204 48676
rect 335604 48674 336204 48676
rect 371604 48674 372204 48676
rect 407604 48674 408204 48676
rect 443604 48674 444204 48676
rect 479604 48674 480204 48676
rect 515604 48674 516204 48676
rect 551604 48674 552204 48676
rect 590840 48674 591440 48676
rect -5676 45676 -5076 45678
rect 8004 45676 8604 45678
rect 44004 45676 44604 45678
rect 80004 45676 80604 45678
rect 116004 45676 116604 45678
rect 152004 45676 152604 45678
rect 188004 45676 188604 45678
rect 224004 45676 224604 45678
rect 260004 45676 260604 45678
rect 296004 45676 296604 45678
rect 332004 45676 332604 45678
rect 368004 45676 368604 45678
rect 404004 45676 404604 45678
rect 440004 45676 440604 45678
rect 476004 45676 476604 45678
rect 512004 45676 512604 45678
rect 548004 45676 548604 45678
rect 589000 45676 589600 45678
rect -6596 45654 590520 45676
rect -6596 45418 -5494 45654
rect -5258 45418 8186 45654
rect 8422 45418 44186 45654
rect 44422 45418 80186 45654
rect 80422 45418 116186 45654
rect 116422 45418 152186 45654
rect 152422 45418 188186 45654
rect 188422 45418 224186 45654
rect 224422 45418 260186 45654
rect 260422 45418 296186 45654
rect 296422 45418 332186 45654
rect 332422 45418 368186 45654
rect 368422 45418 404186 45654
rect 404422 45418 440186 45654
rect 440422 45418 476186 45654
rect 476422 45418 512186 45654
rect 512422 45418 548186 45654
rect 548422 45418 589182 45654
rect 589418 45418 590520 45654
rect -6596 45334 590520 45418
rect -6596 45098 -5494 45334
rect -5258 45098 8186 45334
rect 8422 45098 44186 45334
rect 44422 45098 80186 45334
rect 80422 45098 116186 45334
rect 116422 45098 152186 45334
rect 152422 45098 188186 45334
rect 188422 45098 224186 45334
rect 224422 45098 260186 45334
rect 260422 45098 296186 45334
rect 296422 45098 332186 45334
rect 332422 45098 368186 45334
rect 368422 45098 404186 45334
rect 404422 45098 440186 45334
rect 440422 45098 476186 45334
rect 476422 45098 512186 45334
rect 512422 45098 548186 45334
rect 548422 45098 589182 45334
rect 589418 45098 590520 45334
rect -6596 45076 590520 45098
rect -5676 45074 -5076 45076
rect 8004 45074 8604 45076
rect 44004 45074 44604 45076
rect 80004 45074 80604 45076
rect 116004 45074 116604 45076
rect 152004 45074 152604 45076
rect 188004 45074 188604 45076
rect 224004 45074 224604 45076
rect 260004 45074 260604 45076
rect 296004 45074 296604 45076
rect 332004 45074 332604 45076
rect 368004 45074 368604 45076
rect 404004 45074 404604 45076
rect 440004 45074 440604 45076
rect 476004 45074 476604 45076
rect 512004 45074 512604 45076
rect 548004 45074 548604 45076
rect 589000 45074 589600 45076
rect -3836 42076 -3236 42078
rect 4404 42076 5004 42078
rect 40404 42076 41004 42078
rect 76404 42076 77004 42078
rect 112404 42076 113004 42078
rect 148404 42076 149004 42078
rect 184404 42076 185004 42078
rect 220404 42076 221004 42078
rect 256404 42076 257004 42078
rect 292404 42076 293004 42078
rect 328404 42076 329004 42078
rect 364404 42076 365004 42078
rect 400404 42076 401004 42078
rect 436404 42076 437004 42078
rect 472404 42076 473004 42078
rect 508404 42076 509004 42078
rect 544404 42076 545004 42078
rect 580404 42076 581004 42078
rect 587160 42076 587760 42078
rect -4756 42054 588680 42076
rect -4756 41818 -3654 42054
rect -3418 41818 4586 42054
rect 4822 41818 40586 42054
rect 40822 41818 76586 42054
rect 76822 41818 112586 42054
rect 112822 41818 148586 42054
rect 148822 41818 184586 42054
rect 184822 41818 220586 42054
rect 220822 41818 256586 42054
rect 256822 41818 292586 42054
rect 292822 41818 328586 42054
rect 328822 41818 364586 42054
rect 364822 41818 400586 42054
rect 400822 41818 436586 42054
rect 436822 41818 472586 42054
rect 472822 41818 508586 42054
rect 508822 41818 544586 42054
rect 544822 41818 580586 42054
rect 580822 41818 587342 42054
rect 587578 41818 588680 42054
rect -4756 41734 588680 41818
rect -4756 41498 -3654 41734
rect -3418 41498 4586 41734
rect 4822 41498 40586 41734
rect 40822 41498 76586 41734
rect 76822 41498 112586 41734
rect 112822 41498 148586 41734
rect 148822 41498 184586 41734
rect 184822 41498 220586 41734
rect 220822 41498 256586 41734
rect 256822 41498 292586 41734
rect 292822 41498 328586 41734
rect 328822 41498 364586 41734
rect 364822 41498 400586 41734
rect 400822 41498 436586 41734
rect 436822 41498 472586 41734
rect 472822 41498 508586 41734
rect 508822 41498 544586 41734
rect 544822 41498 580586 41734
rect 580822 41498 587342 41734
rect 587578 41498 588680 41734
rect -4756 41476 588680 41498
rect -3836 41474 -3236 41476
rect 4404 41474 5004 41476
rect 40404 41474 41004 41476
rect 76404 41474 77004 41476
rect 112404 41474 113004 41476
rect 148404 41474 149004 41476
rect 184404 41474 185004 41476
rect 220404 41474 221004 41476
rect 256404 41474 257004 41476
rect 292404 41474 293004 41476
rect 328404 41474 329004 41476
rect 364404 41474 365004 41476
rect 400404 41474 401004 41476
rect 436404 41474 437004 41476
rect 472404 41474 473004 41476
rect 508404 41474 509004 41476
rect 544404 41474 545004 41476
rect 580404 41474 581004 41476
rect 587160 41474 587760 41476
rect -1996 38476 -1396 38478
rect 804 38476 1404 38478
rect 36804 38476 37404 38478
rect 72804 38476 73404 38478
rect 108804 38476 109404 38478
rect 144804 38476 145404 38478
rect 180804 38476 181404 38478
rect 216804 38476 217404 38478
rect 252804 38476 253404 38478
rect 288804 38476 289404 38478
rect 324804 38476 325404 38478
rect 360804 38476 361404 38478
rect 396804 38476 397404 38478
rect 432804 38476 433404 38478
rect 468804 38476 469404 38478
rect 504804 38476 505404 38478
rect 540804 38476 541404 38478
rect 576804 38476 577404 38478
rect 585320 38476 585920 38478
rect -2916 38454 586840 38476
rect -2916 38218 -1814 38454
rect -1578 38218 986 38454
rect 1222 38218 36986 38454
rect 37222 38218 72986 38454
rect 73222 38218 108986 38454
rect 109222 38218 144986 38454
rect 145222 38218 180986 38454
rect 181222 38218 216986 38454
rect 217222 38218 252986 38454
rect 253222 38218 288986 38454
rect 289222 38218 324986 38454
rect 325222 38218 360986 38454
rect 361222 38218 396986 38454
rect 397222 38218 432986 38454
rect 433222 38218 468986 38454
rect 469222 38218 504986 38454
rect 505222 38218 540986 38454
rect 541222 38218 576986 38454
rect 577222 38218 585502 38454
rect 585738 38218 586840 38454
rect -2916 38134 586840 38218
rect -2916 37898 -1814 38134
rect -1578 37898 986 38134
rect 1222 37898 36986 38134
rect 37222 37898 72986 38134
rect 73222 37898 108986 38134
rect 109222 37898 144986 38134
rect 145222 37898 180986 38134
rect 181222 37898 216986 38134
rect 217222 37898 252986 38134
rect 253222 37898 288986 38134
rect 289222 37898 324986 38134
rect 325222 37898 360986 38134
rect 361222 37898 396986 38134
rect 397222 37898 432986 38134
rect 433222 37898 468986 38134
rect 469222 37898 504986 38134
rect 505222 37898 540986 38134
rect 541222 37898 576986 38134
rect 577222 37898 585502 38134
rect 585738 37898 586840 38134
rect -2916 37876 586840 37898
rect -1996 37874 -1396 37876
rect 804 37874 1404 37876
rect 36804 37874 37404 37876
rect 72804 37874 73404 37876
rect 108804 37874 109404 37876
rect 144804 37874 145404 37876
rect 180804 37874 181404 37876
rect 216804 37874 217404 37876
rect 252804 37874 253404 37876
rect 288804 37874 289404 37876
rect 324804 37874 325404 37876
rect 360804 37874 361404 37876
rect 396804 37874 397404 37876
rect 432804 37874 433404 37876
rect 468804 37874 469404 37876
rect 504804 37874 505404 37876
rect 540804 37874 541404 37876
rect 576804 37874 577404 37876
rect 585320 37874 585920 37876
rect -8436 31276 -7836 31278
rect 29604 31276 30204 31278
rect 65604 31276 66204 31278
rect 101604 31276 102204 31278
rect 137604 31276 138204 31278
rect 173604 31276 174204 31278
rect 209604 31276 210204 31278
rect 245604 31276 246204 31278
rect 281604 31276 282204 31278
rect 317604 31276 318204 31278
rect 353604 31276 354204 31278
rect 389604 31276 390204 31278
rect 425604 31276 426204 31278
rect 461604 31276 462204 31278
rect 497604 31276 498204 31278
rect 533604 31276 534204 31278
rect 569604 31276 570204 31278
rect 591760 31276 592360 31278
rect -8436 31254 592360 31276
rect -8436 31018 -8254 31254
rect -8018 31018 29786 31254
rect 30022 31018 65786 31254
rect 66022 31018 101786 31254
rect 102022 31018 137786 31254
rect 138022 31018 173786 31254
rect 174022 31018 209786 31254
rect 210022 31018 245786 31254
rect 246022 31018 281786 31254
rect 282022 31018 317786 31254
rect 318022 31018 353786 31254
rect 354022 31018 389786 31254
rect 390022 31018 425786 31254
rect 426022 31018 461786 31254
rect 462022 31018 497786 31254
rect 498022 31018 533786 31254
rect 534022 31018 569786 31254
rect 570022 31018 591942 31254
rect 592178 31018 592360 31254
rect -8436 30934 592360 31018
rect -8436 30698 -8254 30934
rect -8018 30698 29786 30934
rect 30022 30698 65786 30934
rect 66022 30698 101786 30934
rect 102022 30698 137786 30934
rect 138022 30698 173786 30934
rect 174022 30698 209786 30934
rect 210022 30698 245786 30934
rect 246022 30698 281786 30934
rect 282022 30698 317786 30934
rect 318022 30698 353786 30934
rect 354022 30698 389786 30934
rect 390022 30698 425786 30934
rect 426022 30698 461786 30934
rect 462022 30698 497786 30934
rect 498022 30698 533786 30934
rect 534022 30698 569786 30934
rect 570022 30698 591942 30934
rect 592178 30698 592360 30934
rect -8436 30676 592360 30698
rect -8436 30674 -7836 30676
rect 29604 30674 30204 30676
rect 65604 30674 66204 30676
rect 101604 30674 102204 30676
rect 137604 30674 138204 30676
rect 173604 30674 174204 30676
rect 209604 30674 210204 30676
rect 245604 30674 246204 30676
rect 281604 30674 282204 30676
rect 317604 30674 318204 30676
rect 353604 30674 354204 30676
rect 389604 30674 390204 30676
rect 425604 30674 426204 30676
rect 461604 30674 462204 30676
rect 497604 30674 498204 30676
rect 533604 30674 534204 30676
rect 569604 30674 570204 30676
rect 591760 30674 592360 30676
rect -6596 27676 -5996 27678
rect 26004 27676 26604 27678
rect 62004 27676 62604 27678
rect 98004 27676 98604 27678
rect 134004 27676 134604 27678
rect 170004 27676 170604 27678
rect 206004 27676 206604 27678
rect 242004 27676 242604 27678
rect 278004 27676 278604 27678
rect 314004 27676 314604 27678
rect 350004 27676 350604 27678
rect 386004 27676 386604 27678
rect 422004 27676 422604 27678
rect 458004 27676 458604 27678
rect 494004 27676 494604 27678
rect 530004 27676 530604 27678
rect 566004 27676 566604 27678
rect 589920 27676 590520 27678
rect -6596 27654 590520 27676
rect -6596 27418 -6414 27654
rect -6178 27418 26186 27654
rect 26422 27418 62186 27654
rect 62422 27418 98186 27654
rect 98422 27418 134186 27654
rect 134422 27418 170186 27654
rect 170422 27418 206186 27654
rect 206422 27418 242186 27654
rect 242422 27418 278186 27654
rect 278422 27418 314186 27654
rect 314422 27418 350186 27654
rect 350422 27418 386186 27654
rect 386422 27418 422186 27654
rect 422422 27418 458186 27654
rect 458422 27418 494186 27654
rect 494422 27418 530186 27654
rect 530422 27418 566186 27654
rect 566422 27418 590102 27654
rect 590338 27418 590520 27654
rect -6596 27334 590520 27418
rect -6596 27098 -6414 27334
rect -6178 27098 26186 27334
rect 26422 27098 62186 27334
rect 62422 27098 98186 27334
rect 98422 27098 134186 27334
rect 134422 27098 170186 27334
rect 170422 27098 206186 27334
rect 206422 27098 242186 27334
rect 242422 27098 278186 27334
rect 278422 27098 314186 27334
rect 314422 27098 350186 27334
rect 350422 27098 386186 27334
rect 386422 27098 422186 27334
rect 422422 27098 458186 27334
rect 458422 27098 494186 27334
rect 494422 27098 530186 27334
rect 530422 27098 566186 27334
rect 566422 27098 590102 27334
rect 590338 27098 590520 27334
rect -6596 27076 590520 27098
rect -6596 27074 -5996 27076
rect 26004 27074 26604 27076
rect 62004 27074 62604 27076
rect 98004 27074 98604 27076
rect 134004 27074 134604 27076
rect 170004 27074 170604 27076
rect 206004 27074 206604 27076
rect 242004 27074 242604 27076
rect 278004 27074 278604 27076
rect 314004 27074 314604 27076
rect 350004 27074 350604 27076
rect 386004 27074 386604 27076
rect 422004 27074 422604 27076
rect 458004 27074 458604 27076
rect 494004 27074 494604 27076
rect 530004 27074 530604 27076
rect 566004 27074 566604 27076
rect 589920 27074 590520 27076
rect -4756 24076 -4156 24078
rect 22404 24076 23004 24078
rect 58404 24076 59004 24078
rect 94404 24076 95004 24078
rect 130404 24076 131004 24078
rect 166404 24076 167004 24078
rect 202404 24076 203004 24078
rect 238404 24076 239004 24078
rect 274404 24076 275004 24078
rect 310404 24076 311004 24078
rect 346404 24076 347004 24078
rect 382404 24076 383004 24078
rect 418404 24076 419004 24078
rect 454404 24076 455004 24078
rect 490404 24076 491004 24078
rect 526404 24076 527004 24078
rect 562404 24076 563004 24078
rect 588080 24076 588680 24078
rect -4756 24054 588680 24076
rect -4756 23818 -4574 24054
rect -4338 23818 22586 24054
rect 22822 23818 58586 24054
rect 58822 23818 94586 24054
rect 94822 23818 130586 24054
rect 130822 23818 166586 24054
rect 166822 23818 202586 24054
rect 202822 23818 238586 24054
rect 238822 23818 274586 24054
rect 274822 23818 310586 24054
rect 310822 23818 346586 24054
rect 346822 23818 382586 24054
rect 382822 23818 418586 24054
rect 418822 23818 454586 24054
rect 454822 23818 490586 24054
rect 490822 23818 526586 24054
rect 526822 23818 562586 24054
rect 562822 23818 588262 24054
rect 588498 23818 588680 24054
rect -4756 23734 588680 23818
rect -4756 23498 -4574 23734
rect -4338 23498 22586 23734
rect 22822 23498 58586 23734
rect 58822 23498 94586 23734
rect 94822 23498 130586 23734
rect 130822 23498 166586 23734
rect 166822 23498 202586 23734
rect 202822 23498 238586 23734
rect 238822 23498 274586 23734
rect 274822 23498 310586 23734
rect 310822 23498 346586 23734
rect 346822 23498 382586 23734
rect 382822 23498 418586 23734
rect 418822 23498 454586 23734
rect 454822 23498 490586 23734
rect 490822 23498 526586 23734
rect 526822 23498 562586 23734
rect 562822 23498 588262 23734
rect 588498 23498 588680 23734
rect -4756 23476 588680 23498
rect -4756 23474 -4156 23476
rect 22404 23474 23004 23476
rect 58404 23474 59004 23476
rect 94404 23474 95004 23476
rect 130404 23474 131004 23476
rect 166404 23474 167004 23476
rect 202404 23474 203004 23476
rect 238404 23474 239004 23476
rect 274404 23474 275004 23476
rect 310404 23474 311004 23476
rect 346404 23474 347004 23476
rect 382404 23474 383004 23476
rect 418404 23474 419004 23476
rect 454404 23474 455004 23476
rect 490404 23474 491004 23476
rect 526404 23474 527004 23476
rect 562404 23474 563004 23476
rect 588080 23474 588680 23476
rect -2916 20476 -2316 20478
rect 18804 20476 19404 20478
rect 54804 20476 55404 20478
rect 90804 20476 91404 20478
rect 126804 20476 127404 20478
rect 162804 20476 163404 20478
rect 198804 20476 199404 20478
rect 234804 20476 235404 20478
rect 270804 20476 271404 20478
rect 306804 20476 307404 20478
rect 342804 20476 343404 20478
rect 378804 20476 379404 20478
rect 414804 20476 415404 20478
rect 450804 20476 451404 20478
rect 486804 20476 487404 20478
rect 522804 20476 523404 20478
rect 558804 20476 559404 20478
rect 586240 20476 586840 20478
rect -2916 20454 586840 20476
rect -2916 20218 -2734 20454
rect -2498 20218 18986 20454
rect 19222 20218 54986 20454
rect 55222 20218 90986 20454
rect 91222 20218 126986 20454
rect 127222 20218 162986 20454
rect 163222 20218 198986 20454
rect 199222 20218 234986 20454
rect 235222 20218 270986 20454
rect 271222 20218 306986 20454
rect 307222 20218 342986 20454
rect 343222 20218 378986 20454
rect 379222 20218 414986 20454
rect 415222 20218 450986 20454
rect 451222 20218 486986 20454
rect 487222 20218 522986 20454
rect 523222 20218 558986 20454
rect 559222 20218 586422 20454
rect 586658 20218 586840 20454
rect -2916 20134 586840 20218
rect -2916 19898 -2734 20134
rect -2498 19898 18986 20134
rect 19222 19898 54986 20134
rect 55222 19898 90986 20134
rect 91222 19898 126986 20134
rect 127222 19898 162986 20134
rect 163222 19898 198986 20134
rect 199222 19898 234986 20134
rect 235222 19898 270986 20134
rect 271222 19898 306986 20134
rect 307222 19898 342986 20134
rect 343222 19898 378986 20134
rect 379222 19898 414986 20134
rect 415222 19898 450986 20134
rect 451222 19898 486986 20134
rect 487222 19898 522986 20134
rect 523222 19898 558986 20134
rect 559222 19898 586422 20134
rect 586658 19898 586840 20134
rect -2916 19876 586840 19898
rect -2916 19874 -2316 19876
rect 18804 19874 19404 19876
rect 54804 19874 55404 19876
rect 90804 19874 91404 19876
rect 126804 19874 127404 19876
rect 162804 19874 163404 19876
rect 198804 19874 199404 19876
rect 234804 19874 235404 19876
rect 270804 19874 271404 19876
rect 306804 19874 307404 19876
rect 342804 19874 343404 19876
rect 378804 19874 379404 19876
rect 414804 19874 415404 19876
rect 450804 19874 451404 19876
rect 486804 19874 487404 19876
rect 522804 19874 523404 19876
rect 558804 19874 559404 19876
rect 586240 19874 586840 19876
rect -7516 13276 -6916 13278
rect 11604 13276 12204 13278
rect 47604 13276 48204 13278
rect 83604 13276 84204 13278
rect 119604 13276 120204 13278
rect 155604 13276 156204 13278
rect 191604 13276 192204 13278
rect 227604 13276 228204 13278
rect 263604 13276 264204 13278
rect 299604 13276 300204 13278
rect 335604 13276 336204 13278
rect 371604 13276 372204 13278
rect 407604 13276 408204 13278
rect 443604 13276 444204 13278
rect 479604 13276 480204 13278
rect 515604 13276 516204 13278
rect 551604 13276 552204 13278
rect 590840 13276 591440 13278
rect -8436 13254 592360 13276
rect -8436 13018 -7334 13254
rect -7098 13018 11786 13254
rect 12022 13018 47786 13254
rect 48022 13018 83786 13254
rect 84022 13018 119786 13254
rect 120022 13018 155786 13254
rect 156022 13018 191786 13254
rect 192022 13018 227786 13254
rect 228022 13018 263786 13254
rect 264022 13018 299786 13254
rect 300022 13018 335786 13254
rect 336022 13018 371786 13254
rect 372022 13018 407786 13254
rect 408022 13018 443786 13254
rect 444022 13018 479786 13254
rect 480022 13018 515786 13254
rect 516022 13018 551786 13254
rect 552022 13018 591022 13254
rect 591258 13018 592360 13254
rect -8436 12934 592360 13018
rect -8436 12698 -7334 12934
rect -7098 12698 11786 12934
rect 12022 12698 47786 12934
rect 48022 12698 83786 12934
rect 84022 12698 119786 12934
rect 120022 12698 155786 12934
rect 156022 12698 191786 12934
rect 192022 12698 227786 12934
rect 228022 12698 263786 12934
rect 264022 12698 299786 12934
rect 300022 12698 335786 12934
rect 336022 12698 371786 12934
rect 372022 12698 407786 12934
rect 408022 12698 443786 12934
rect 444022 12698 479786 12934
rect 480022 12698 515786 12934
rect 516022 12698 551786 12934
rect 552022 12698 591022 12934
rect 591258 12698 592360 12934
rect -8436 12676 592360 12698
rect -7516 12674 -6916 12676
rect 11604 12674 12204 12676
rect 47604 12674 48204 12676
rect 83604 12674 84204 12676
rect 119604 12674 120204 12676
rect 155604 12674 156204 12676
rect 191604 12674 192204 12676
rect 227604 12674 228204 12676
rect 263604 12674 264204 12676
rect 299604 12674 300204 12676
rect 335604 12674 336204 12676
rect 371604 12674 372204 12676
rect 407604 12674 408204 12676
rect 443604 12674 444204 12676
rect 479604 12674 480204 12676
rect 515604 12674 516204 12676
rect 551604 12674 552204 12676
rect 590840 12674 591440 12676
rect -5676 9676 -5076 9678
rect 8004 9676 8604 9678
rect 44004 9676 44604 9678
rect 80004 9676 80604 9678
rect 116004 9676 116604 9678
rect 152004 9676 152604 9678
rect 188004 9676 188604 9678
rect 224004 9676 224604 9678
rect 260004 9676 260604 9678
rect 296004 9676 296604 9678
rect 332004 9676 332604 9678
rect 368004 9676 368604 9678
rect 404004 9676 404604 9678
rect 440004 9676 440604 9678
rect 476004 9676 476604 9678
rect 512004 9676 512604 9678
rect 548004 9676 548604 9678
rect 589000 9676 589600 9678
rect -6596 9654 590520 9676
rect -6596 9418 -5494 9654
rect -5258 9418 8186 9654
rect 8422 9418 44186 9654
rect 44422 9418 80186 9654
rect 80422 9418 116186 9654
rect 116422 9418 152186 9654
rect 152422 9418 188186 9654
rect 188422 9418 224186 9654
rect 224422 9418 260186 9654
rect 260422 9418 296186 9654
rect 296422 9418 332186 9654
rect 332422 9418 368186 9654
rect 368422 9418 404186 9654
rect 404422 9418 440186 9654
rect 440422 9418 476186 9654
rect 476422 9418 512186 9654
rect 512422 9418 548186 9654
rect 548422 9418 589182 9654
rect 589418 9418 590520 9654
rect -6596 9334 590520 9418
rect -6596 9098 -5494 9334
rect -5258 9098 8186 9334
rect 8422 9098 44186 9334
rect 44422 9098 80186 9334
rect 80422 9098 116186 9334
rect 116422 9098 152186 9334
rect 152422 9098 188186 9334
rect 188422 9098 224186 9334
rect 224422 9098 260186 9334
rect 260422 9098 296186 9334
rect 296422 9098 332186 9334
rect 332422 9098 368186 9334
rect 368422 9098 404186 9334
rect 404422 9098 440186 9334
rect 440422 9098 476186 9334
rect 476422 9098 512186 9334
rect 512422 9098 548186 9334
rect 548422 9098 589182 9334
rect 589418 9098 590520 9334
rect -6596 9076 590520 9098
rect -5676 9074 -5076 9076
rect 8004 9074 8604 9076
rect 44004 9074 44604 9076
rect 80004 9074 80604 9076
rect 116004 9074 116604 9076
rect 152004 9074 152604 9076
rect 188004 9074 188604 9076
rect 224004 9074 224604 9076
rect 260004 9074 260604 9076
rect 296004 9074 296604 9076
rect 332004 9074 332604 9076
rect 368004 9074 368604 9076
rect 404004 9074 404604 9076
rect 440004 9074 440604 9076
rect 476004 9074 476604 9076
rect 512004 9074 512604 9076
rect 548004 9074 548604 9076
rect 589000 9074 589600 9076
rect -3836 6076 -3236 6078
rect 4404 6076 5004 6078
rect 40404 6076 41004 6078
rect 76404 6076 77004 6078
rect 112404 6076 113004 6078
rect 148404 6076 149004 6078
rect 184404 6076 185004 6078
rect 220404 6076 221004 6078
rect 256404 6076 257004 6078
rect 292404 6076 293004 6078
rect 328404 6076 329004 6078
rect 364404 6076 365004 6078
rect 400404 6076 401004 6078
rect 436404 6076 437004 6078
rect 472404 6076 473004 6078
rect 508404 6076 509004 6078
rect 544404 6076 545004 6078
rect 580404 6076 581004 6078
rect 587160 6076 587760 6078
rect -4756 6054 588680 6076
rect -4756 5818 -3654 6054
rect -3418 5818 4586 6054
rect 4822 5818 40586 6054
rect 40822 5818 76586 6054
rect 76822 5818 112586 6054
rect 112822 5818 148586 6054
rect 148822 5818 184586 6054
rect 184822 5818 220586 6054
rect 220822 5818 256586 6054
rect 256822 5818 292586 6054
rect 292822 5818 328586 6054
rect 328822 5818 364586 6054
rect 364822 5818 400586 6054
rect 400822 5818 436586 6054
rect 436822 5818 472586 6054
rect 472822 5818 508586 6054
rect 508822 5818 544586 6054
rect 544822 5818 580586 6054
rect 580822 5818 587342 6054
rect 587578 5818 588680 6054
rect -4756 5734 588680 5818
rect -4756 5498 -3654 5734
rect -3418 5498 4586 5734
rect 4822 5498 40586 5734
rect 40822 5498 76586 5734
rect 76822 5498 112586 5734
rect 112822 5498 148586 5734
rect 148822 5498 184586 5734
rect 184822 5498 220586 5734
rect 220822 5498 256586 5734
rect 256822 5498 292586 5734
rect 292822 5498 328586 5734
rect 328822 5498 364586 5734
rect 364822 5498 400586 5734
rect 400822 5498 436586 5734
rect 436822 5498 472586 5734
rect 472822 5498 508586 5734
rect 508822 5498 544586 5734
rect 544822 5498 580586 5734
rect 580822 5498 587342 5734
rect 587578 5498 588680 5734
rect -4756 5476 588680 5498
rect -3836 5474 -3236 5476
rect 4404 5474 5004 5476
rect 40404 5474 41004 5476
rect 76404 5474 77004 5476
rect 112404 5474 113004 5476
rect 148404 5474 149004 5476
rect 184404 5474 185004 5476
rect 220404 5474 221004 5476
rect 256404 5474 257004 5476
rect 292404 5474 293004 5476
rect 328404 5474 329004 5476
rect 364404 5474 365004 5476
rect 400404 5474 401004 5476
rect 436404 5474 437004 5476
rect 472404 5474 473004 5476
rect 508404 5474 509004 5476
rect 544404 5474 545004 5476
rect 580404 5474 581004 5476
rect 587160 5474 587760 5476
rect -1996 2476 -1396 2478
rect 804 2476 1404 2478
rect 36804 2476 37404 2478
rect 72804 2476 73404 2478
rect 108804 2476 109404 2478
rect 144804 2476 145404 2478
rect 180804 2476 181404 2478
rect 216804 2476 217404 2478
rect 252804 2476 253404 2478
rect 288804 2476 289404 2478
rect 324804 2476 325404 2478
rect 360804 2476 361404 2478
rect 396804 2476 397404 2478
rect 432804 2476 433404 2478
rect 468804 2476 469404 2478
rect 504804 2476 505404 2478
rect 540804 2476 541404 2478
rect 576804 2476 577404 2478
rect 585320 2476 585920 2478
rect -2916 2454 586840 2476
rect -2916 2218 -1814 2454
rect -1578 2218 986 2454
rect 1222 2218 36986 2454
rect 37222 2218 72986 2454
rect 73222 2218 108986 2454
rect 109222 2218 144986 2454
rect 145222 2218 180986 2454
rect 181222 2218 216986 2454
rect 217222 2218 252986 2454
rect 253222 2218 288986 2454
rect 289222 2218 324986 2454
rect 325222 2218 360986 2454
rect 361222 2218 396986 2454
rect 397222 2218 432986 2454
rect 433222 2218 468986 2454
rect 469222 2218 504986 2454
rect 505222 2218 540986 2454
rect 541222 2218 576986 2454
rect 577222 2218 585502 2454
rect 585738 2218 586840 2454
rect -2916 2134 586840 2218
rect -2916 1898 -1814 2134
rect -1578 1898 986 2134
rect 1222 1898 36986 2134
rect 37222 1898 72986 2134
rect 73222 1898 108986 2134
rect 109222 1898 144986 2134
rect 145222 1898 180986 2134
rect 181222 1898 216986 2134
rect 217222 1898 252986 2134
rect 253222 1898 288986 2134
rect 289222 1898 324986 2134
rect 325222 1898 360986 2134
rect 361222 1898 396986 2134
rect 397222 1898 432986 2134
rect 433222 1898 468986 2134
rect 469222 1898 504986 2134
rect 505222 1898 540986 2134
rect 541222 1898 576986 2134
rect 577222 1898 585502 2134
rect 585738 1898 586840 2134
rect -2916 1876 586840 1898
rect -1996 1874 -1396 1876
rect 804 1874 1404 1876
rect 36804 1874 37404 1876
rect 72804 1874 73404 1876
rect 108804 1874 109404 1876
rect 144804 1874 145404 1876
rect 180804 1874 181404 1876
rect 216804 1874 217404 1876
rect 252804 1874 253404 1876
rect 288804 1874 289404 1876
rect 324804 1874 325404 1876
rect 360804 1874 361404 1876
rect 396804 1874 397404 1876
rect 432804 1874 433404 1876
rect 468804 1874 469404 1876
rect 504804 1874 505404 1876
rect 540804 1874 541404 1876
rect 576804 1874 577404 1876
rect 585320 1874 585920 1876
rect -1996 -324 -1396 -322
rect 804 -324 1404 -322
rect 36804 -324 37404 -322
rect 72804 -324 73404 -322
rect 108804 -324 109404 -322
rect 144804 -324 145404 -322
rect 180804 -324 181404 -322
rect 216804 -324 217404 -322
rect 252804 -324 253404 -322
rect 288804 -324 289404 -322
rect 324804 -324 325404 -322
rect 360804 -324 361404 -322
rect 396804 -324 397404 -322
rect 432804 -324 433404 -322
rect 468804 -324 469404 -322
rect 504804 -324 505404 -322
rect 540804 -324 541404 -322
rect 576804 -324 577404 -322
rect 585320 -324 585920 -322
rect -1996 -346 585920 -324
rect -1996 -582 -1814 -346
rect -1578 -582 986 -346
rect 1222 -582 36986 -346
rect 37222 -582 72986 -346
rect 73222 -582 108986 -346
rect 109222 -582 144986 -346
rect 145222 -582 180986 -346
rect 181222 -582 216986 -346
rect 217222 -582 252986 -346
rect 253222 -582 288986 -346
rect 289222 -582 324986 -346
rect 325222 -582 360986 -346
rect 361222 -582 396986 -346
rect 397222 -582 432986 -346
rect 433222 -582 468986 -346
rect 469222 -582 504986 -346
rect 505222 -582 540986 -346
rect 541222 -582 576986 -346
rect 577222 -582 585502 -346
rect 585738 -582 585920 -346
rect -1996 -666 585920 -582
rect -1996 -902 -1814 -666
rect -1578 -902 986 -666
rect 1222 -902 36986 -666
rect 37222 -902 72986 -666
rect 73222 -902 108986 -666
rect 109222 -902 144986 -666
rect 145222 -902 180986 -666
rect 181222 -902 216986 -666
rect 217222 -902 252986 -666
rect 253222 -902 288986 -666
rect 289222 -902 324986 -666
rect 325222 -902 360986 -666
rect 361222 -902 396986 -666
rect 397222 -902 432986 -666
rect 433222 -902 468986 -666
rect 469222 -902 504986 -666
rect 505222 -902 540986 -666
rect 541222 -902 576986 -666
rect 577222 -902 585502 -666
rect 585738 -902 585920 -666
rect -1996 -924 585920 -902
rect -1996 -926 -1396 -924
rect 804 -926 1404 -924
rect 36804 -926 37404 -924
rect 72804 -926 73404 -924
rect 108804 -926 109404 -924
rect 144804 -926 145404 -924
rect 180804 -926 181404 -924
rect 216804 -926 217404 -924
rect 252804 -926 253404 -924
rect 288804 -926 289404 -924
rect 324804 -926 325404 -924
rect 360804 -926 361404 -924
rect 396804 -926 397404 -924
rect 432804 -926 433404 -924
rect 468804 -926 469404 -924
rect 504804 -926 505404 -924
rect 540804 -926 541404 -924
rect 576804 -926 577404 -924
rect 585320 -926 585920 -924
rect -2916 -1244 -2316 -1242
rect 18804 -1244 19404 -1242
rect 54804 -1244 55404 -1242
rect 90804 -1244 91404 -1242
rect 126804 -1244 127404 -1242
rect 162804 -1244 163404 -1242
rect 198804 -1244 199404 -1242
rect 234804 -1244 235404 -1242
rect 270804 -1244 271404 -1242
rect 306804 -1244 307404 -1242
rect 342804 -1244 343404 -1242
rect 378804 -1244 379404 -1242
rect 414804 -1244 415404 -1242
rect 450804 -1244 451404 -1242
rect 486804 -1244 487404 -1242
rect 522804 -1244 523404 -1242
rect 558804 -1244 559404 -1242
rect 586240 -1244 586840 -1242
rect -2916 -1266 586840 -1244
rect -2916 -1502 -2734 -1266
rect -2498 -1502 18986 -1266
rect 19222 -1502 54986 -1266
rect 55222 -1502 90986 -1266
rect 91222 -1502 126986 -1266
rect 127222 -1502 162986 -1266
rect 163222 -1502 198986 -1266
rect 199222 -1502 234986 -1266
rect 235222 -1502 270986 -1266
rect 271222 -1502 306986 -1266
rect 307222 -1502 342986 -1266
rect 343222 -1502 378986 -1266
rect 379222 -1502 414986 -1266
rect 415222 -1502 450986 -1266
rect 451222 -1502 486986 -1266
rect 487222 -1502 522986 -1266
rect 523222 -1502 558986 -1266
rect 559222 -1502 586422 -1266
rect 586658 -1502 586840 -1266
rect -2916 -1586 586840 -1502
rect -2916 -1822 -2734 -1586
rect -2498 -1822 18986 -1586
rect 19222 -1822 54986 -1586
rect 55222 -1822 90986 -1586
rect 91222 -1822 126986 -1586
rect 127222 -1822 162986 -1586
rect 163222 -1822 198986 -1586
rect 199222 -1822 234986 -1586
rect 235222 -1822 270986 -1586
rect 271222 -1822 306986 -1586
rect 307222 -1822 342986 -1586
rect 343222 -1822 378986 -1586
rect 379222 -1822 414986 -1586
rect 415222 -1822 450986 -1586
rect 451222 -1822 486986 -1586
rect 487222 -1822 522986 -1586
rect 523222 -1822 558986 -1586
rect 559222 -1822 586422 -1586
rect 586658 -1822 586840 -1586
rect -2916 -1844 586840 -1822
rect -2916 -1846 -2316 -1844
rect 18804 -1846 19404 -1844
rect 54804 -1846 55404 -1844
rect 90804 -1846 91404 -1844
rect 126804 -1846 127404 -1844
rect 162804 -1846 163404 -1844
rect 198804 -1846 199404 -1844
rect 234804 -1846 235404 -1844
rect 270804 -1846 271404 -1844
rect 306804 -1846 307404 -1844
rect 342804 -1846 343404 -1844
rect 378804 -1846 379404 -1844
rect 414804 -1846 415404 -1844
rect 450804 -1846 451404 -1844
rect 486804 -1846 487404 -1844
rect 522804 -1846 523404 -1844
rect 558804 -1846 559404 -1844
rect 586240 -1846 586840 -1844
rect -3836 -2164 -3236 -2162
rect 4404 -2164 5004 -2162
rect 40404 -2164 41004 -2162
rect 76404 -2164 77004 -2162
rect 112404 -2164 113004 -2162
rect 148404 -2164 149004 -2162
rect 184404 -2164 185004 -2162
rect 220404 -2164 221004 -2162
rect 256404 -2164 257004 -2162
rect 292404 -2164 293004 -2162
rect 328404 -2164 329004 -2162
rect 364404 -2164 365004 -2162
rect 400404 -2164 401004 -2162
rect 436404 -2164 437004 -2162
rect 472404 -2164 473004 -2162
rect 508404 -2164 509004 -2162
rect 544404 -2164 545004 -2162
rect 580404 -2164 581004 -2162
rect 587160 -2164 587760 -2162
rect -3836 -2186 587760 -2164
rect -3836 -2422 -3654 -2186
rect -3418 -2422 4586 -2186
rect 4822 -2422 40586 -2186
rect 40822 -2422 76586 -2186
rect 76822 -2422 112586 -2186
rect 112822 -2422 148586 -2186
rect 148822 -2422 184586 -2186
rect 184822 -2422 220586 -2186
rect 220822 -2422 256586 -2186
rect 256822 -2422 292586 -2186
rect 292822 -2422 328586 -2186
rect 328822 -2422 364586 -2186
rect 364822 -2422 400586 -2186
rect 400822 -2422 436586 -2186
rect 436822 -2422 472586 -2186
rect 472822 -2422 508586 -2186
rect 508822 -2422 544586 -2186
rect 544822 -2422 580586 -2186
rect 580822 -2422 587342 -2186
rect 587578 -2422 587760 -2186
rect -3836 -2506 587760 -2422
rect -3836 -2742 -3654 -2506
rect -3418 -2742 4586 -2506
rect 4822 -2742 40586 -2506
rect 40822 -2742 76586 -2506
rect 76822 -2742 112586 -2506
rect 112822 -2742 148586 -2506
rect 148822 -2742 184586 -2506
rect 184822 -2742 220586 -2506
rect 220822 -2742 256586 -2506
rect 256822 -2742 292586 -2506
rect 292822 -2742 328586 -2506
rect 328822 -2742 364586 -2506
rect 364822 -2742 400586 -2506
rect 400822 -2742 436586 -2506
rect 436822 -2742 472586 -2506
rect 472822 -2742 508586 -2506
rect 508822 -2742 544586 -2506
rect 544822 -2742 580586 -2506
rect 580822 -2742 587342 -2506
rect 587578 -2742 587760 -2506
rect -3836 -2764 587760 -2742
rect -3836 -2766 -3236 -2764
rect 4404 -2766 5004 -2764
rect 40404 -2766 41004 -2764
rect 76404 -2766 77004 -2764
rect 112404 -2766 113004 -2764
rect 148404 -2766 149004 -2764
rect 184404 -2766 185004 -2764
rect 220404 -2766 221004 -2764
rect 256404 -2766 257004 -2764
rect 292404 -2766 293004 -2764
rect 328404 -2766 329004 -2764
rect 364404 -2766 365004 -2764
rect 400404 -2766 401004 -2764
rect 436404 -2766 437004 -2764
rect 472404 -2766 473004 -2764
rect 508404 -2766 509004 -2764
rect 544404 -2766 545004 -2764
rect 580404 -2766 581004 -2764
rect 587160 -2766 587760 -2764
rect -4756 -3084 -4156 -3082
rect 22404 -3084 23004 -3082
rect 58404 -3084 59004 -3082
rect 94404 -3084 95004 -3082
rect 130404 -3084 131004 -3082
rect 166404 -3084 167004 -3082
rect 202404 -3084 203004 -3082
rect 238404 -3084 239004 -3082
rect 274404 -3084 275004 -3082
rect 310404 -3084 311004 -3082
rect 346404 -3084 347004 -3082
rect 382404 -3084 383004 -3082
rect 418404 -3084 419004 -3082
rect 454404 -3084 455004 -3082
rect 490404 -3084 491004 -3082
rect 526404 -3084 527004 -3082
rect 562404 -3084 563004 -3082
rect 588080 -3084 588680 -3082
rect -4756 -3106 588680 -3084
rect -4756 -3342 -4574 -3106
rect -4338 -3342 22586 -3106
rect 22822 -3342 58586 -3106
rect 58822 -3342 94586 -3106
rect 94822 -3342 130586 -3106
rect 130822 -3342 166586 -3106
rect 166822 -3342 202586 -3106
rect 202822 -3342 238586 -3106
rect 238822 -3342 274586 -3106
rect 274822 -3342 310586 -3106
rect 310822 -3342 346586 -3106
rect 346822 -3342 382586 -3106
rect 382822 -3342 418586 -3106
rect 418822 -3342 454586 -3106
rect 454822 -3342 490586 -3106
rect 490822 -3342 526586 -3106
rect 526822 -3342 562586 -3106
rect 562822 -3342 588262 -3106
rect 588498 -3342 588680 -3106
rect -4756 -3426 588680 -3342
rect -4756 -3662 -4574 -3426
rect -4338 -3662 22586 -3426
rect 22822 -3662 58586 -3426
rect 58822 -3662 94586 -3426
rect 94822 -3662 130586 -3426
rect 130822 -3662 166586 -3426
rect 166822 -3662 202586 -3426
rect 202822 -3662 238586 -3426
rect 238822 -3662 274586 -3426
rect 274822 -3662 310586 -3426
rect 310822 -3662 346586 -3426
rect 346822 -3662 382586 -3426
rect 382822 -3662 418586 -3426
rect 418822 -3662 454586 -3426
rect 454822 -3662 490586 -3426
rect 490822 -3662 526586 -3426
rect 526822 -3662 562586 -3426
rect 562822 -3662 588262 -3426
rect 588498 -3662 588680 -3426
rect -4756 -3684 588680 -3662
rect -4756 -3686 -4156 -3684
rect 22404 -3686 23004 -3684
rect 58404 -3686 59004 -3684
rect 94404 -3686 95004 -3684
rect 130404 -3686 131004 -3684
rect 166404 -3686 167004 -3684
rect 202404 -3686 203004 -3684
rect 238404 -3686 239004 -3684
rect 274404 -3686 275004 -3684
rect 310404 -3686 311004 -3684
rect 346404 -3686 347004 -3684
rect 382404 -3686 383004 -3684
rect 418404 -3686 419004 -3684
rect 454404 -3686 455004 -3684
rect 490404 -3686 491004 -3684
rect 526404 -3686 527004 -3684
rect 562404 -3686 563004 -3684
rect 588080 -3686 588680 -3684
rect -5676 -4004 -5076 -4002
rect 8004 -4004 8604 -4002
rect 44004 -4004 44604 -4002
rect 80004 -4004 80604 -4002
rect 116004 -4004 116604 -4002
rect 152004 -4004 152604 -4002
rect 188004 -4004 188604 -4002
rect 224004 -4004 224604 -4002
rect 260004 -4004 260604 -4002
rect 296004 -4004 296604 -4002
rect 332004 -4004 332604 -4002
rect 368004 -4004 368604 -4002
rect 404004 -4004 404604 -4002
rect 440004 -4004 440604 -4002
rect 476004 -4004 476604 -4002
rect 512004 -4004 512604 -4002
rect 548004 -4004 548604 -4002
rect 589000 -4004 589600 -4002
rect -5676 -4026 589600 -4004
rect -5676 -4262 -5494 -4026
rect -5258 -4262 8186 -4026
rect 8422 -4262 44186 -4026
rect 44422 -4262 80186 -4026
rect 80422 -4262 116186 -4026
rect 116422 -4262 152186 -4026
rect 152422 -4262 188186 -4026
rect 188422 -4262 224186 -4026
rect 224422 -4262 260186 -4026
rect 260422 -4262 296186 -4026
rect 296422 -4262 332186 -4026
rect 332422 -4262 368186 -4026
rect 368422 -4262 404186 -4026
rect 404422 -4262 440186 -4026
rect 440422 -4262 476186 -4026
rect 476422 -4262 512186 -4026
rect 512422 -4262 548186 -4026
rect 548422 -4262 589182 -4026
rect 589418 -4262 589600 -4026
rect -5676 -4346 589600 -4262
rect -5676 -4582 -5494 -4346
rect -5258 -4582 8186 -4346
rect 8422 -4582 44186 -4346
rect 44422 -4582 80186 -4346
rect 80422 -4582 116186 -4346
rect 116422 -4582 152186 -4346
rect 152422 -4582 188186 -4346
rect 188422 -4582 224186 -4346
rect 224422 -4582 260186 -4346
rect 260422 -4582 296186 -4346
rect 296422 -4582 332186 -4346
rect 332422 -4582 368186 -4346
rect 368422 -4582 404186 -4346
rect 404422 -4582 440186 -4346
rect 440422 -4582 476186 -4346
rect 476422 -4582 512186 -4346
rect 512422 -4582 548186 -4346
rect 548422 -4582 589182 -4346
rect 589418 -4582 589600 -4346
rect -5676 -4604 589600 -4582
rect -5676 -4606 -5076 -4604
rect 8004 -4606 8604 -4604
rect 44004 -4606 44604 -4604
rect 80004 -4606 80604 -4604
rect 116004 -4606 116604 -4604
rect 152004 -4606 152604 -4604
rect 188004 -4606 188604 -4604
rect 224004 -4606 224604 -4604
rect 260004 -4606 260604 -4604
rect 296004 -4606 296604 -4604
rect 332004 -4606 332604 -4604
rect 368004 -4606 368604 -4604
rect 404004 -4606 404604 -4604
rect 440004 -4606 440604 -4604
rect 476004 -4606 476604 -4604
rect 512004 -4606 512604 -4604
rect 548004 -4606 548604 -4604
rect 589000 -4606 589600 -4604
rect -6596 -4924 -5996 -4922
rect 26004 -4924 26604 -4922
rect 62004 -4924 62604 -4922
rect 98004 -4924 98604 -4922
rect 134004 -4924 134604 -4922
rect 170004 -4924 170604 -4922
rect 206004 -4924 206604 -4922
rect 242004 -4924 242604 -4922
rect 278004 -4924 278604 -4922
rect 314004 -4924 314604 -4922
rect 350004 -4924 350604 -4922
rect 386004 -4924 386604 -4922
rect 422004 -4924 422604 -4922
rect 458004 -4924 458604 -4922
rect 494004 -4924 494604 -4922
rect 530004 -4924 530604 -4922
rect 566004 -4924 566604 -4922
rect 589920 -4924 590520 -4922
rect -6596 -4946 590520 -4924
rect -6596 -5182 -6414 -4946
rect -6178 -5182 26186 -4946
rect 26422 -5182 62186 -4946
rect 62422 -5182 98186 -4946
rect 98422 -5182 134186 -4946
rect 134422 -5182 170186 -4946
rect 170422 -5182 206186 -4946
rect 206422 -5182 242186 -4946
rect 242422 -5182 278186 -4946
rect 278422 -5182 314186 -4946
rect 314422 -5182 350186 -4946
rect 350422 -5182 386186 -4946
rect 386422 -5182 422186 -4946
rect 422422 -5182 458186 -4946
rect 458422 -5182 494186 -4946
rect 494422 -5182 530186 -4946
rect 530422 -5182 566186 -4946
rect 566422 -5182 590102 -4946
rect 590338 -5182 590520 -4946
rect -6596 -5266 590520 -5182
rect -6596 -5502 -6414 -5266
rect -6178 -5502 26186 -5266
rect 26422 -5502 62186 -5266
rect 62422 -5502 98186 -5266
rect 98422 -5502 134186 -5266
rect 134422 -5502 170186 -5266
rect 170422 -5502 206186 -5266
rect 206422 -5502 242186 -5266
rect 242422 -5502 278186 -5266
rect 278422 -5502 314186 -5266
rect 314422 -5502 350186 -5266
rect 350422 -5502 386186 -5266
rect 386422 -5502 422186 -5266
rect 422422 -5502 458186 -5266
rect 458422 -5502 494186 -5266
rect 494422 -5502 530186 -5266
rect 530422 -5502 566186 -5266
rect 566422 -5502 590102 -5266
rect 590338 -5502 590520 -5266
rect -6596 -5524 590520 -5502
rect -6596 -5526 -5996 -5524
rect 26004 -5526 26604 -5524
rect 62004 -5526 62604 -5524
rect 98004 -5526 98604 -5524
rect 134004 -5526 134604 -5524
rect 170004 -5526 170604 -5524
rect 206004 -5526 206604 -5524
rect 242004 -5526 242604 -5524
rect 278004 -5526 278604 -5524
rect 314004 -5526 314604 -5524
rect 350004 -5526 350604 -5524
rect 386004 -5526 386604 -5524
rect 422004 -5526 422604 -5524
rect 458004 -5526 458604 -5524
rect 494004 -5526 494604 -5524
rect 530004 -5526 530604 -5524
rect 566004 -5526 566604 -5524
rect 589920 -5526 590520 -5524
rect -7516 -5844 -6916 -5842
rect 11604 -5844 12204 -5842
rect 47604 -5844 48204 -5842
rect 83604 -5844 84204 -5842
rect 119604 -5844 120204 -5842
rect 155604 -5844 156204 -5842
rect 191604 -5844 192204 -5842
rect 227604 -5844 228204 -5842
rect 263604 -5844 264204 -5842
rect 299604 -5844 300204 -5842
rect 335604 -5844 336204 -5842
rect 371604 -5844 372204 -5842
rect 407604 -5844 408204 -5842
rect 443604 -5844 444204 -5842
rect 479604 -5844 480204 -5842
rect 515604 -5844 516204 -5842
rect 551604 -5844 552204 -5842
rect 590840 -5844 591440 -5842
rect -7516 -5866 591440 -5844
rect -7516 -6102 -7334 -5866
rect -7098 -6102 11786 -5866
rect 12022 -6102 47786 -5866
rect 48022 -6102 83786 -5866
rect 84022 -6102 119786 -5866
rect 120022 -6102 155786 -5866
rect 156022 -6102 191786 -5866
rect 192022 -6102 227786 -5866
rect 228022 -6102 263786 -5866
rect 264022 -6102 299786 -5866
rect 300022 -6102 335786 -5866
rect 336022 -6102 371786 -5866
rect 372022 -6102 407786 -5866
rect 408022 -6102 443786 -5866
rect 444022 -6102 479786 -5866
rect 480022 -6102 515786 -5866
rect 516022 -6102 551786 -5866
rect 552022 -6102 591022 -5866
rect 591258 -6102 591440 -5866
rect -7516 -6186 591440 -6102
rect -7516 -6422 -7334 -6186
rect -7098 -6422 11786 -6186
rect 12022 -6422 47786 -6186
rect 48022 -6422 83786 -6186
rect 84022 -6422 119786 -6186
rect 120022 -6422 155786 -6186
rect 156022 -6422 191786 -6186
rect 192022 -6422 227786 -6186
rect 228022 -6422 263786 -6186
rect 264022 -6422 299786 -6186
rect 300022 -6422 335786 -6186
rect 336022 -6422 371786 -6186
rect 372022 -6422 407786 -6186
rect 408022 -6422 443786 -6186
rect 444022 -6422 479786 -6186
rect 480022 -6422 515786 -6186
rect 516022 -6422 551786 -6186
rect 552022 -6422 591022 -6186
rect 591258 -6422 591440 -6186
rect -7516 -6444 591440 -6422
rect -7516 -6446 -6916 -6444
rect 11604 -6446 12204 -6444
rect 47604 -6446 48204 -6444
rect 83604 -6446 84204 -6444
rect 119604 -6446 120204 -6444
rect 155604 -6446 156204 -6444
rect 191604 -6446 192204 -6444
rect 227604 -6446 228204 -6444
rect 263604 -6446 264204 -6444
rect 299604 -6446 300204 -6444
rect 335604 -6446 336204 -6444
rect 371604 -6446 372204 -6444
rect 407604 -6446 408204 -6444
rect 443604 -6446 444204 -6444
rect 479604 -6446 480204 -6444
rect 515604 -6446 516204 -6444
rect 551604 -6446 552204 -6444
rect 590840 -6446 591440 -6444
rect -8436 -6764 -7836 -6762
rect 29604 -6764 30204 -6762
rect 65604 -6764 66204 -6762
rect 101604 -6764 102204 -6762
rect 137604 -6764 138204 -6762
rect 173604 -6764 174204 -6762
rect 209604 -6764 210204 -6762
rect 245604 -6764 246204 -6762
rect 281604 -6764 282204 -6762
rect 317604 -6764 318204 -6762
rect 353604 -6764 354204 -6762
rect 389604 -6764 390204 -6762
rect 425604 -6764 426204 -6762
rect 461604 -6764 462204 -6762
rect 497604 -6764 498204 -6762
rect 533604 -6764 534204 -6762
rect 569604 -6764 570204 -6762
rect 591760 -6764 592360 -6762
rect -8436 -6786 592360 -6764
rect -8436 -7022 -8254 -6786
rect -8018 -7022 29786 -6786
rect 30022 -7022 65786 -6786
rect 66022 -7022 101786 -6786
rect 102022 -7022 137786 -6786
rect 138022 -7022 173786 -6786
rect 174022 -7022 209786 -6786
rect 210022 -7022 245786 -6786
rect 246022 -7022 281786 -6786
rect 282022 -7022 317786 -6786
rect 318022 -7022 353786 -6786
rect 354022 -7022 389786 -6786
rect 390022 -7022 425786 -6786
rect 426022 -7022 461786 -6786
rect 462022 -7022 497786 -6786
rect 498022 -7022 533786 -6786
rect 534022 -7022 569786 -6786
rect 570022 -7022 591942 -6786
rect 592178 -7022 592360 -6786
rect -8436 -7106 592360 -7022
rect -8436 -7342 -8254 -7106
rect -8018 -7342 29786 -7106
rect 30022 -7342 65786 -7106
rect 66022 -7342 101786 -7106
rect 102022 -7342 137786 -7106
rect 138022 -7342 173786 -7106
rect 174022 -7342 209786 -7106
rect 210022 -7342 245786 -7106
rect 246022 -7342 281786 -7106
rect 282022 -7342 317786 -7106
rect 318022 -7342 353786 -7106
rect 354022 -7342 389786 -7106
rect 390022 -7342 425786 -7106
rect 426022 -7342 461786 -7106
rect 462022 -7342 497786 -7106
rect 498022 -7342 533786 -7106
rect 534022 -7342 569786 -7106
rect 570022 -7342 591942 -7106
rect 592178 -7342 592360 -7106
rect -8436 -7364 592360 -7342
rect -8436 -7366 -7836 -7364
rect 29604 -7366 30204 -7364
rect 65604 -7366 66204 -7364
rect 101604 -7366 102204 -7364
rect 137604 -7366 138204 -7364
rect 173604 -7366 174204 -7364
rect 209604 -7366 210204 -7364
rect 245604 -7366 246204 -7364
rect 281604 -7366 282204 -7364
rect 317604 -7366 318204 -7364
rect 353604 -7366 354204 -7364
rect 389604 -7366 390204 -7364
rect 425604 -7366 426204 -7364
rect 461604 -7366 462204 -7364
rect 497604 -7366 498204 -7364
rect 533604 -7366 534204 -7364
rect 569604 -7366 570204 -7364
rect 591760 -7366 592360 -7364
use user_proj_example  mprj
timestamp 1608118436
transform 1 0 230000 0 1 340000
box 0 0 59856 60000
<< labels >>
rlabel metal3 s 583520 5796 584960 6036 6 analog_io[0]
port 0 nsew default bidirectional
rlabel metal3 s 583520 474996 584960 475236 6 analog_io[10]
port 1 nsew default bidirectional
rlabel metal3 s 583520 521916 584960 522156 6 analog_io[11]
port 2 nsew default bidirectional
rlabel metal3 s 583520 568836 584960 569076 6 analog_io[12]
port 3 nsew default bidirectional
rlabel metal3 s 583520 615756 584960 615996 6 analog_io[13]
port 4 nsew default bidirectional
rlabel metal3 s 583520 662676 584960 662916 6 analog_io[14]
port 5 nsew default bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[15]
port 6 nsew default bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[16]
port 7 nsew default bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[17]
port 8 nsew default bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[18]
port 9 nsew default bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[19]
port 10 nsew default bidirectional
rlabel metal3 s 583520 52716 584960 52956 6 analog_io[1]
port 11 nsew default bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[20]
port 12 nsew default bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[21]
port 13 nsew default bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[22]
port 14 nsew default bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[23]
port 15 nsew default bidirectional
rlabel metal3 s -960 696540 480 696780 4 analog_io[24]
port 16 nsew default bidirectional
rlabel metal3 s -960 639012 480 639252 4 analog_io[25]
port 17 nsew default bidirectional
rlabel metal3 s -960 581620 480 581860 4 analog_io[26]
port 18 nsew default bidirectional
rlabel metal3 s -960 524092 480 524332 4 analog_io[27]
port 19 nsew default bidirectional
rlabel metal3 s -960 466700 480 466940 4 analog_io[28]
port 20 nsew default bidirectional
rlabel metal3 s -960 409172 480 409412 4 analog_io[29]
port 21 nsew default bidirectional
rlabel metal3 s 583520 99636 584960 99876 6 analog_io[2]
port 22 nsew default bidirectional
rlabel metal3 s -960 351780 480 352020 4 analog_io[30]
port 23 nsew default bidirectional
rlabel metal3 s 583520 146556 584960 146796 6 analog_io[3]
port 24 nsew default bidirectional
rlabel metal3 s 583520 193476 584960 193716 6 analog_io[4]
port 25 nsew default bidirectional
rlabel metal3 s 583520 240396 584960 240636 6 analog_io[5]
port 26 nsew default bidirectional
rlabel metal3 s 583520 287316 584960 287556 6 analog_io[6]
port 27 nsew default bidirectional
rlabel metal3 s 583520 334236 584960 334476 6 analog_io[7]
port 28 nsew default bidirectional
rlabel metal3 s 583520 381156 584960 381396 6 analog_io[8]
port 29 nsew default bidirectional
rlabel metal3 s 583520 428076 584960 428316 6 analog_io[9]
port 30 nsew default bidirectional
rlabel metal3 s 583520 17492 584960 17732 6 io_in[0]
port 31 nsew default input
rlabel metal3 s 583520 486692 584960 486932 6 io_in[10]
port 32 nsew default input
rlabel metal3 s 583520 533748 584960 533988 6 io_in[11]
port 33 nsew default input
rlabel metal3 s 583520 580668 584960 580908 6 io_in[12]
port 34 nsew default input
rlabel metal3 s 583520 627588 584960 627828 6 io_in[13]
port 35 nsew default input
rlabel metal3 s 583520 674508 584960 674748 6 io_in[14]
port 36 nsew default input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 37 nsew default input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 38 nsew default input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 39 nsew default input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 40 nsew default input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 41 nsew default input
rlabel metal3 s 583520 64412 584960 64652 6 io_in[1]
port 42 nsew default input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 43 nsew default input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 44 nsew default input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 45 nsew default input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 46 nsew default input
rlabel metal3 s -960 682124 480 682364 4 io_in[24]
port 47 nsew default input
rlabel metal3 s -960 624732 480 624972 4 io_in[25]
port 48 nsew default input
rlabel metal3 s -960 567204 480 567444 4 io_in[26]
port 49 nsew default input
rlabel metal3 s -960 509812 480 510052 4 io_in[27]
port 50 nsew default input
rlabel metal3 s -960 452284 480 452524 4 io_in[28]
port 51 nsew default input
rlabel metal3 s -960 394892 480 395132 4 io_in[29]
port 52 nsew default input
rlabel metal3 s 583520 111332 584960 111572 6 io_in[2]
port 53 nsew default input
rlabel metal3 s -960 337364 480 337604 4 io_in[30]
port 54 nsew default input
rlabel metal3 s -960 294252 480 294492 4 io_in[31]
port 55 nsew default input
rlabel metal3 s -960 251140 480 251380 4 io_in[32]
port 56 nsew default input
rlabel metal3 s -960 208028 480 208268 4 io_in[33]
port 57 nsew default input
rlabel metal3 s -960 164916 480 165156 4 io_in[34]
port 58 nsew default input
rlabel metal3 s -960 121940 480 122180 4 io_in[35]
port 59 nsew default input
rlabel metal3 s -960 78828 480 79068 4 io_in[36]
port 60 nsew default input
rlabel metal3 s -960 35716 480 35956 4 io_in[37]
port 61 nsew default input
rlabel metal3 s 583520 158252 584960 158492 6 io_in[3]
port 62 nsew default input
rlabel metal3 s 583520 205172 584960 205412 6 io_in[4]
port 63 nsew default input
rlabel metal3 s 583520 252092 584960 252332 6 io_in[5]
port 64 nsew default input
rlabel metal3 s 583520 299012 584960 299252 6 io_in[6]
port 65 nsew default input
rlabel metal3 s 583520 345932 584960 346172 6 io_in[7]
port 66 nsew default input
rlabel metal3 s 583520 392852 584960 393092 6 io_in[8]
port 67 nsew default input
rlabel metal3 s 583520 439772 584960 440012 6 io_in[9]
port 68 nsew default input
rlabel metal3 s 583520 40884 584960 41124 6 io_oeb[0]
port 69 nsew default tristate
rlabel metal3 s 583520 510220 584960 510460 6 io_oeb[10]
port 70 nsew default tristate
rlabel metal3 s 583520 557140 584960 557380 6 io_oeb[11]
port 71 nsew default tristate
rlabel metal3 s 583520 604060 584960 604300 6 io_oeb[12]
port 72 nsew default tristate
rlabel metal3 s 583520 650980 584960 651220 6 io_oeb[13]
port 73 nsew default tristate
rlabel metal3 s 583520 697900 584960 698140 6 io_oeb[14]
port 74 nsew default tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 75 nsew default tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 76 nsew default tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 77 nsew default tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 78 nsew default tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 79 nsew default tristate
rlabel metal3 s 583520 87804 584960 88044 6 io_oeb[1]
port 80 nsew default tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 81 nsew default tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 82 nsew default tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 83 nsew default tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 84 nsew default tristate
rlabel metal3 s -960 653428 480 653668 4 io_oeb[24]
port 85 nsew default tristate
rlabel metal3 s -960 595900 480 596140 4 io_oeb[25]
port 86 nsew default tristate
rlabel metal3 s -960 538508 480 538748 4 io_oeb[26]
port 87 nsew default tristate
rlabel metal3 s -960 480980 480 481220 4 io_oeb[27]
port 88 nsew default tristate
rlabel metal3 s -960 423588 480 423828 4 io_oeb[28]
port 89 nsew default tristate
rlabel metal3 s -960 366060 480 366300 4 io_oeb[29]
port 90 nsew default tristate
rlabel metal3 s 583520 134724 584960 134964 6 io_oeb[2]
port 91 nsew default tristate
rlabel metal3 s -960 308668 480 308908 4 io_oeb[30]
port 92 nsew default tristate
rlabel metal3 s -960 265556 480 265796 4 io_oeb[31]
port 93 nsew default tristate
rlabel metal3 s -960 222444 480 222684 4 io_oeb[32]
port 94 nsew default tristate
rlabel metal3 s -960 179332 480 179572 4 io_oeb[33]
port 95 nsew default tristate
rlabel metal3 s -960 136220 480 136460 4 io_oeb[34]
port 96 nsew default tristate
rlabel metal3 s -960 93108 480 93348 4 io_oeb[35]
port 97 nsew default tristate
rlabel metal3 s -960 49996 480 50236 4 io_oeb[36]
port 98 nsew default tristate
rlabel metal3 s -960 7020 480 7260 4 io_oeb[37]
port 99 nsew default tristate
rlabel metal3 s 583520 181780 584960 182020 6 io_oeb[3]
port 100 nsew default tristate
rlabel metal3 s 583520 228700 584960 228940 6 io_oeb[4]
port 101 nsew default tristate
rlabel metal3 s 583520 275620 584960 275860 6 io_oeb[5]
port 102 nsew default tristate
rlabel metal3 s 583520 322540 584960 322780 6 io_oeb[6]
port 103 nsew default tristate
rlabel metal3 s 583520 369460 584960 369700 6 io_oeb[7]
port 104 nsew default tristate
rlabel metal3 s 583520 416380 584960 416620 6 io_oeb[8]
port 105 nsew default tristate
rlabel metal3 s 583520 463300 584960 463540 6 io_oeb[9]
port 106 nsew default tristate
rlabel metal3 s 583520 29188 584960 29428 6 io_out[0]
port 107 nsew default tristate
rlabel metal3 s 583520 498524 584960 498764 6 io_out[10]
port 108 nsew default tristate
rlabel metal3 s 583520 545444 584960 545684 6 io_out[11]
port 109 nsew default tristate
rlabel metal3 s 583520 592364 584960 592604 6 io_out[12]
port 110 nsew default tristate
rlabel metal3 s 583520 639284 584960 639524 6 io_out[13]
port 111 nsew default tristate
rlabel metal3 s 583520 686204 584960 686444 6 io_out[14]
port 112 nsew default tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 113 nsew default tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 114 nsew default tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 115 nsew default tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 116 nsew default tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 117 nsew default tristate
rlabel metal3 s 583520 76108 584960 76348 6 io_out[1]
port 118 nsew default tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 119 nsew default tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 120 nsew default tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 121 nsew default tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 122 nsew default tristate
rlabel metal3 s -960 667844 480 668084 4 io_out[24]
port 123 nsew default tristate
rlabel metal3 s -960 610316 480 610556 4 io_out[25]
port 124 nsew default tristate
rlabel metal3 s -960 552924 480 553164 4 io_out[26]
port 125 nsew default tristate
rlabel metal3 s -960 495396 480 495636 4 io_out[27]
port 126 nsew default tristate
rlabel metal3 s -960 437868 480 438108 4 io_out[28]
port 127 nsew default tristate
rlabel metal3 s -960 380476 480 380716 4 io_out[29]
port 128 nsew default tristate
rlabel metal3 s 583520 123028 584960 123268 6 io_out[2]
port 129 nsew default tristate
rlabel metal3 s -960 322948 480 323188 4 io_out[30]
port 130 nsew default tristate
rlabel metal3 s -960 279972 480 280212 4 io_out[31]
port 131 nsew default tristate
rlabel metal3 s -960 236860 480 237100 4 io_out[32]
port 132 nsew default tristate
rlabel metal3 s -960 193748 480 193988 4 io_out[33]
port 133 nsew default tristate
rlabel metal3 s -960 150636 480 150876 4 io_out[34]
port 134 nsew default tristate
rlabel metal3 s -960 107524 480 107764 4 io_out[35]
port 135 nsew default tristate
rlabel metal3 s -960 64412 480 64652 4 io_out[36]
port 136 nsew default tristate
rlabel metal3 s -960 21300 480 21540 4 io_out[37]
port 137 nsew default tristate
rlabel metal3 s 583520 169948 584960 170188 6 io_out[3]
port 138 nsew default tristate
rlabel metal3 s 583520 216868 584960 217108 6 io_out[4]
port 139 nsew default tristate
rlabel metal3 s 583520 263788 584960 264028 6 io_out[5]
port 140 nsew default tristate
rlabel metal3 s 583520 310708 584960 310948 6 io_out[6]
port 141 nsew default tristate
rlabel metal3 s 583520 357764 584960 358004 6 io_out[7]
port 142 nsew default tristate
rlabel metal3 s 583520 404684 584960 404924 6 io_out[8]
port 143 nsew default tristate
rlabel metal3 s 583520 451604 584960 451844 6 io_out[9]
port 144 nsew default tristate
rlabel metal2 s 126582 -960 126694 480 8 la_data_in[0]
port 145 nsew default input
rlabel metal2 s 483450 -960 483562 480 8 la_data_in[100]
port 146 nsew default input
rlabel metal2 s 486946 -960 487058 480 8 la_data_in[101]
port 147 nsew default input
rlabel metal2 s 490534 -960 490646 480 8 la_data_in[102]
port 148 nsew default input
rlabel metal2 s 494122 -960 494234 480 8 la_data_in[103]
port 149 nsew default input
rlabel metal2 s 497710 -960 497822 480 8 la_data_in[104]
port 150 nsew default input
rlabel metal2 s 501206 -960 501318 480 8 la_data_in[105]
port 151 nsew default input
rlabel metal2 s 504794 -960 504906 480 8 la_data_in[106]
port 152 nsew default input
rlabel metal2 s 508382 -960 508494 480 8 la_data_in[107]
port 153 nsew default input
rlabel metal2 s 511970 -960 512082 480 8 la_data_in[108]
port 154 nsew default input
rlabel metal2 s 515558 -960 515670 480 8 la_data_in[109]
port 155 nsew default input
rlabel metal2 s 162278 -960 162390 480 8 la_data_in[10]
port 156 nsew default input
rlabel metal2 s 519054 -960 519166 480 8 la_data_in[110]
port 157 nsew default input
rlabel metal2 s 522642 -960 522754 480 8 la_data_in[111]
port 158 nsew default input
rlabel metal2 s 526230 -960 526342 480 8 la_data_in[112]
port 159 nsew default input
rlabel metal2 s 529818 -960 529930 480 8 la_data_in[113]
port 160 nsew default input
rlabel metal2 s 533406 -960 533518 480 8 la_data_in[114]
port 161 nsew default input
rlabel metal2 s 536902 -960 537014 480 8 la_data_in[115]
port 162 nsew default input
rlabel metal2 s 540490 -960 540602 480 8 la_data_in[116]
port 163 nsew default input
rlabel metal2 s 544078 -960 544190 480 8 la_data_in[117]
port 164 nsew default input
rlabel metal2 s 547666 -960 547778 480 8 la_data_in[118]
port 165 nsew default input
rlabel metal2 s 551162 -960 551274 480 8 la_data_in[119]
port 166 nsew default input
rlabel metal2 s 165866 -960 165978 480 8 la_data_in[11]
port 167 nsew default input
rlabel metal2 s 554750 -960 554862 480 8 la_data_in[120]
port 168 nsew default input
rlabel metal2 s 558338 -960 558450 480 8 la_data_in[121]
port 169 nsew default input
rlabel metal2 s 561926 -960 562038 480 8 la_data_in[122]
port 170 nsew default input
rlabel metal2 s 565514 -960 565626 480 8 la_data_in[123]
port 171 nsew default input
rlabel metal2 s 569010 -960 569122 480 8 la_data_in[124]
port 172 nsew default input
rlabel metal2 s 572598 -960 572710 480 8 la_data_in[125]
port 173 nsew default input
rlabel metal2 s 576186 -960 576298 480 8 la_data_in[126]
port 174 nsew default input
rlabel metal2 s 579774 -960 579886 480 8 la_data_in[127]
port 175 nsew default input
rlabel metal2 s 169362 -960 169474 480 8 la_data_in[12]
port 176 nsew default input
rlabel metal2 s 172950 -960 173062 480 8 la_data_in[13]
port 177 nsew default input
rlabel metal2 s 176538 -960 176650 480 8 la_data_in[14]
port 178 nsew default input
rlabel metal2 s 180126 -960 180238 480 8 la_data_in[15]
port 179 nsew default input
rlabel metal2 s 183714 -960 183826 480 8 la_data_in[16]
port 180 nsew default input
rlabel metal2 s 187210 -960 187322 480 8 la_data_in[17]
port 181 nsew default input
rlabel metal2 s 190798 -960 190910 480 8 la_data_in[18]
port 182 nsew default input
rlabel metal2 s 194386 -960 194498 480 8 la_data_in[19]
port 183 nsew default input
rlabel metal2 s 130170 -960 130282 480 8 la_data_in[1]
port 184 nsew default input
rlabel metal2 s 197974 -960 198086 480 8 la_data_in[20]
port 185 nsew default input
rlabel metal2 s 201470 -960 201582 480 8 la_data_in[21]
port 186 nsew default input
rlabel metal2 s 205058 -960 205170 480 8 la_data_in[22]
port 187 nsew default input
rlabel metal2 s 208646 -960 208758 480 8 la_data_in[23]
port 188 nsew default input
rlabel metal2 s 212234 -960 212346 480 8 la_data_in[24]
port 189 nsew default input
rlabel metal2 s 215822 -960 215934 480 8 la_data_in[25]
port 190 nsew default input
rlabel metal2 s 219318 -960 219430 480 8 la_data_in[26]
port 191 nsew default input
rlabel metal2 s 222906 -960 223018 480 8 la_data_in[27]
port 192 nsew default input
rlabel metal2 s 226494 -960 226606 480 8 la_data_in[28]
port 193 nsew default input
rlabel metal2 s 230082 -960 230194 480 8 la_data_in[29]
port 194 nsew default input
rlabel metal2 s 133758 -960 133870 480 8 la_data_in[2]
port 195 nsew default input
rlabel metal2 s 233670 -960 233782 480 8 la_data_in[30]
port 196 nsew default input
rlabel metal2 s 237166 -960 237278 480 8 la_data_in[31]
port 197 nsew default input
rlabel metal2 s 240754 -960 240866 480 8 la_data_in[32]
port 198 nsew default input
rlabel metal2 s 244342 -960 244454 480 8 la_data_in[33]
port 199 nsew default input
rlabel metal2 s 247930 -960 248042 480 8 la_data_in[34]
port 200 nsew default input
rlabel metal2 s 251426 -960 251538 480 8 la_data_in[35]
port 201 nsew default input
rlabel metal2 s 255014 -960 255126 480 8 la_data_in[36]
port 202 nsew default input
rlabel metal2 s 258602 -960 258714 480 8 la_data_in[37]
port 203 nsew default input
rlabel metal2 s 262190 -960 262302 480 8 la_data_in[38]
port 204 nsew default input
rlabel metal2 s 265778 -960 265890 480 8 la_data_in[39]
port 205 nsew default input
rlabel metal2 s 137254 -960 137366 480 8 la_data_in[3]
port 206 nsew default input
rlabel metal2 s 269274 -960 269386 480 8 la_data_in[40]
port 207 nsew default input
rlabel metal2 s 272862 -960 272974 480 8 la_data_in[41]
port 208 nsew default input
rlabel metal2 s 276450 -960 276562 480 8 la_data_in[42]
port 209 nsew default input
rlabel metal2 s 280038 -960 280150 480 8 la_data_in[43]
port 210 nsew default input
rlabel metal2 s 283626 -960 283738 480 8 la_data_in[44]
port 211 nsew default input
rlabel metal2 s 287122 -960 287234 480 8 la_data_in[45]
port 212 nsew default input
rlabel metal2 s 290710 -960 290822 480 8 la_data_in[46]
port 213 nsew default input
rlabel metal2 s 294298 -960 294410 480 8 la_data_in[47]
port 214 nsew default input
rlabel metal2 s 297886 -960 297998 480 8 la_data_in[48]
port 215 nsew default input
rlabel metal2 s 301382 -960 301494 480 8 la_data_in[49]
port 216 nsew default input
rlabel metal2 s 140842 -960 140954 480 8 la_data_in[4]
port 217 nsew default input
rlabel metal2 s 304970 -960 305082 480 8 la_data_in[50]
port 218 nsew default input
rlabel metal2 s 308558 -960 308670 480 8 la_data_in[51]
port 219 nsew default input
rlabel metal2 s 312146 -960 312258 480 8 la_data_in[52]
port 220 nsew default input
rlabel metal2 s 315734 -960 315846 480 8 la_data_in[53]
port 221 nsew default input
rlabel metal2 s 319230 -960 319342 480 8 la_data_in[54]
port 222 nsew default input
rlabel metal2 s 322818 -960 322930 480 8 la_data_in[55]
port 223 nsew default input
rlabel metal2 s 326406 -960 326518 480 8 la_data_in[56]
port 224 nsew default input
rlabel metal2 s 329994 -960 330106 480 8 la_data_in[57]
port 225 nsew default input
rlabel metal2 s 333582 -960 333694 480 8 la_data_in[58]
port 226 nsew default input
rlabel metal2 s 337078 -960 337190 480 8 la_data_in[59]
port 227 nsew default input
rlabel metal2 s 144430 -960 144542 480 8 la_data_in[5]
port 228 nsew default input
rlabel metal2 s 340666 -960 340778 480 8 la_data_in[60]
port 229 nsew default input
rlabel metal2 s 344254 -960 344366 480 8 la_data_in[61]
port 230 nsew default input
rlabel metal2 s 347842 -960 347954 480 8 la_data_in[62]
port 231 nsew default input
rlabel metal2 s 351338 -960 351450 480 8 la_data_in[63]
port 232 nsew default input
rlabel metal2 s 354926 -960 355038 480 8 la_data_in[64]
port 233 nsew default input
rlabel metal2 s 358514 -960 358626 480 8 la_data_in[65]
port 234 nsew default input
rlabel metal2 s 362102 -960 362214 480 8 la_data_in[66]
port 235 nsew default input
rlabel metal2 s 365690 -960 365802 480 8 la_data_in[67]
port 236 nsew default input
rlabel metal2 s 369186 -960 369298 480 8 la_data_in[68]
port 237 nsew default input
rlabel metal2 s 372774 -960 372886 480 8 la_data_in[69]
port 238 nsew default input
rlabel metal2 s 148018 -960 148130 480 8 la_data_in[6]
port 239 nsew default input
rlabel metal2 s 376362 -960 376474 480 8 la_data_in[70]
port 240 nsew default input
rlabel metal2 s 379950 -960 380062 480 8 la_data_in[71]
port 241 nsew default input
rlabel metal2 s 383538 -960 383650 480 8 la_data_in[72]
port 242 nsew default input
rlabel metal2 s 387034 -960 387146 480 8 la_data_in[73]
port 243 nsew default input
rlabel metal2 s 390622 -960 390734 480 8 la_data_in[74]
port 244 nsew default input
rlabel metal2 s 394210 -960 394322 480 8 la_data_in[75]
port 245 nsew default input
rlabel metal2 s 397798 -960 397910 480 8 la_data_in[76]
port 246 nsew default input
rlabel metal2 s 401294 -960 401406 480 8 la_data_in[77]
port 247 nsew default input
rlabel metal2 s 404882 -960 404994 480 8 la_data_in[78]
port 248 nsew default input
rlabel metal2 s 408470 -960 408582 480 8 la_data_in[79]
port 249 nsew default input
rlabel metal2 s 151514 -960 151626 480 8 la_data_in[7]
port 250 nsew default input
rlabel metal2 s 412058 -960 412170 480 8 la_data_in[80]
port 251 nsew default input
rlabel metal2 s 415646 -960 415758 480 8 la_data_in[81]
port 252 nsew default input
rlabel metal2 s 419142 -960 419254 480 8 la_data_in[82]
port 253 nsew default input
rlabel metal2 s 422730 -960 422842 480 8 la_data_in[83]
port 254 nsew default input
rlabel metal2 s 426318 -960 426430 480 8 la_data_in[84]
port 255 nsew default input
rlabel metal2 s 429906 -960 430018 480 8 la_data_in[85]
port 256 nsew default input
rlabel metal2 s 433494 -960 433606 480 8 la_data_in[86]
port 257 nsew default input
rlabel metal2 s 436990 -960 437102 480 8 la_data_in[87]
port 258 nsew default input
rlabel metal2 s 440578 -960 440690 480 8 la_data_in[88]
port 259 nsew default input
rlabel metal2 s 444166 -960 444278 480 8 la_data_in[89]
port 260 nsew default input
rlabel metal2 s 155102 -960 155214 480 8 la_data_in[8]
port 261 nsew default input
rlabel metal2 s 447754 -960 447866 480 8 la_data_in[90]
port 262 nsew default input
rlabel metal2 s 451250 -960 451362 480 8 la_data_in[91]
port 263 nsew default input
rlabel metal2 s 454838 -960 454950 480 8 la_data_in[92]
port 264 nsew default input
rlabel metal2 s 458426 -960 458538 480 8 la_data_in[93]
port 265 nsew default input
rlabel metal2 s 462014 -960 462126 480 8 la_data_in[94]
port 266 nsew default input
rlabel metal2 s 465602 -960 465714 480 8 la_data_in[95]
port 267 nsew default input
rlabel metal2 s 469098 -960 469210 480 8 la_data_in[96]
port 268 nsew default input
rlabel metal2 s 472686 -960 472798 480 8 la_data_in[97]
port 269 nsew default input
rlabel metal2 s 476274 -960 476386 480 8 la_data_in[98]
port 270 nsew default input
rlabel metal2 s 479862 -960 479974 480 8 la_data_in[99]
port 271 nsew default input
rlabel metal2 s 158690 -960 158802 480 8 la_data_in[9]
port 272 nsew default input
rlabel metal2 s 127778 -960 127890 480 8 la_data_out[0]
port 273 nsew default tristate
rlabel metal2 s 484554 -960 484666 480 8 la_data_out[100]
port 274 nsew default tristate
rlabel metal2 s 488142 -960 488254 480 8 la_data_out[101]
port 275 nsew default tristate
rlabel metal2 s 491730 -960 491842 480 8 la_data_out[102]
port 276 nsew default tristate
rlabel metal2 s 495318 -960 495430 480 8 la_data_out[103]
port 277 nsew default tristate
rlabel metal2 s 498906 -960 499018 480 8 la_data_out[104]
port 278 nsew default tristate
rlabel metal2 s 502402 -960 502514 480 8 la_data_out[105]
port 279 nsew default tristate
rlabel metal2 s 505990 -960 506102 480 8 la_data_out[106]
port 280 nsew default tristate
rlabel metal2 s 509578 -960 509690 480 8 la_data_out[107]
port 281 nsew default tristate
rlabel metal2 s 513166 -960 513278 480 8 la_data_out[108]
port 282 nsew default tristate
rlabel metal2 s 516754 -960 516866 480 8 la_data_out[109]
port 283 nsew default tristate
rlabel metal2 s 163474 -960 163586 480 8 la_data_out[10]
port 284 nsew default tristate
rlabel metal2 s 520250 -960 520362 480 8 la_data_out[110]
port 285 nsew default tristate
rlabel metal2 s 523838 -960 523950 480 8 la_data_out[111]
port 286 nsew default tristate
rlabel metal2 s 527426 -960 527538 480 8 la_data_out[112]
port 287 nsew default tristate
rlabel metal2 s 531014 -960 531126 480 8 la_data_out[113]
port 288 nsew default tristate
rlabel metal2 s 534510 -960 534622 480 8 la_data_out[114]
port 289 nsew default tristate
rlabel metal2 s 538098 -960 538210 480 8 la_data_out[115]
port 290 nsew default tristate
rlabel metal2 s 541686 -960 541798 480 8 la_data_out[116]
port 291 nsew default tristate
rlabel metal2 s 545274 -960 545386 480 8 la_data_out[117]
port 292 nsew default tristate
rlabel metal2 s 548862 -960 548974 480 8 la_data_out[118]
port 293 nsew default tristate
rlabel metal2 s 552358 -960 552470 480 8 la_data_out[119]
port 294 nsew default tristate
rlabel metal2 s 167062 -960 167174 480 8 la_data_out[11]
port 295 nsew default tristate
rlabel metal2 s 555946 -960 556058 480 8 la_data_out[120]
port 296 nsew default tristate
rlabel metal2 s 559534 -960 559646 480 8 la_data_out[121]
port 297 nsew default tristate
rlabel metal2 s 563122 -960 563234 480 8 la_data_out[122]
port 298 nsew default tristate
rlabel metal2 s 566710 -960 566822 480 8 la_data_out[123]
port 299 nsew default tristate
rlabel metal2 s 570206 -960 570318 480 8 la_data_out[124]
port 300 nsew default tristate
rlabel metal2 s 573794 -960 573906 480 8 la_data_out[125]
port 301 nsew default tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[126]
port 302 nsew default tristate
rlabel metal2 s 580970 -960 581082 480 8 la_data_out[127]
port 303 nsew default tristate
rlabel metal2 s 170558 -960 170670 480 8 la_data_out[12]
port 304 nsew default tristate
rlabel metal2 s 174146 -960 174258 480 8 la_data_out[13]
port 305 nsew default tristate
rlabel metal2 s 177734 -960 177846 480 8 la_data_out[14]
port 306 nsew default tristate
rlabel metal2 s 181322 -960 181434 480 8 la_data_out[15]
port 307 nsew default tristate
rlabel metal2 s 184818 -960 184930 480 8 la_data_out[16]
port 308 nsew default tristate
rlabel metal2 s 188406 -960 188518 480 8 la_data_out[17]
port 309 nsew default tristate
rlabel metal2 s 191994 -960 192106 480 8 la_data_out[18]
port 310 nsew default tristate
rlabel metal2 s 195582 -960 195694 480 8 la_data_out[19]
port 311 nsew default tristate
rlabel metal2 s 131366 -960 131478 480 8 la_data_out[1]
port 312 nsew default tristate
rlabel metal2 s 199170 -960 199282 480 8 la_data_out[20]
port 313 nsew default tristate
rlabel metal2 s 202666 -960 202778 480 8 la_data_out[21]
port 314 nsew default tristate
rlabel metal2 s 206254 -960 206366 480 8 la_data_out[22]
port 315 nsew default tristate
rlabel metal2 s 209842 -960 209954 480 8 la_data_out[23]
port 316 nsew default tristate
rlabel metal2 s 213430 -960 213542 480 8 la_data_out[24]
port 317 nsew default tristate
rlabel metal2 s 217018 -960 217130 480 8 la_data_out[25]
port 318 nsew default tristate
rlabel metal2 s 220514 -960 220626 480 8 la_data_out[26]
port 319 nsew default tristate
rlabel metal2 s 224102 -960 224214 480 8 la_data_out[27]
port 320 nsew default tristate
rlabel metal2 s 227690 -960 227802 480 8 la_data_out[28]
port 321 nsew default tristate
rlabel metal2 s 231278 -960 231390 480 8 la_data_out[29]
port 322 nsew default tristate
rlabel metal2 s 134862 -960 134974 480 8 la_data_out[2]
port 323 nsew default tristate
rlabel metal2 s 234774 -960 234886 480 8 la_data_out[30]
port 324 nsew default tristate
rlabel metal2 s 238362 -960 238474 480 8 la_data_out[31]
port 325 nsew default tristate
rlabel metal2 s 241950 -960 242062 480 8 la_data_out[32]
port 326 nsew default tristate
rlabel metal2 s 245538 -960 245650 480 8 la_data_out[33]
port 327 nsew default tristate
rlabel metal2 s 249126 -960 249238 480 8 la_data_out[34]
port 328 nsew default tristate
rlabel metal2 s 252622 -960 252734 480 8 la_data_out[35]
port 329 nsew default tristate
rlabel metal2 s 256210 -960 256322 480 8 la_data_out[36]
port 330 nsew default tristate
rlabel metal2 s 259798 -960 259910 480 8 la_data_out[37]
port 331 nsew default tristate
rlabel metal2 s 263386 -960 263498 480 8 la_data_out[38]
port 332 nsew default tristate
rlabel metal2 s 266974 -960 267086 480 8 la_data_out[39]
port 333 nsew default tristate
rlabel metal2 s 138450 -960 138562 480 8 la_data_out[3]
port 334 nsew default tristate
rlabel metal2 s 270470 -960 270582 480 8 la_data_out[40]
port 335 nsew default tristate
rlabel metal2 s 274058 -960 274170 480 8 la_data_out[41]
port 336 nsew default tristate
rlabel metal2 s 277646 -960 277758 480 8 la_data_out[42]
port 337 nsew default tristate
rlabel metal2 s 281234 -960 281346 480 8 la_data_out[43]
port 338 nsew default tristate
rlabel metal2 s 284730 -960 284842 480 8 la_data_out[44]
port 339 nsew default tristate
rlabel metal2 s 288318 -960 288430 480 8 la_data_out[45]
port 340 nsew default tristate
rlabel metal2 s 291906 -960 292018 480 8 la_data_out[46]
port 341 nsew default tristate
rlabel metal2 s 295494 -960 295606 480 8 la_data_out[47]
port 342 nsew default tristate
rlabel metal2 s 299082 -960 299194 480 8 la_data_out[48]
port 343 nsew default tristate
rlabel metal2 s 302578 -960 302690 480 8 la_data_out[49]
port 344 nsew default tristate
rlabel metal2 s 142038 -960 142150 480 8 la_data_out[4]
port 345 nsew default tristate
rlabel metal2 s 306166 -960 306278 480 8 la_data_out[50]
port 346 nsew default tristate
rlabel metal2 s 309754 -960 309866 480 8 la_data_out[51]
port 347 nsew default tristate
rlabel metal2 s 313342 -960 313454 480 8 la_data_out[52]
port 348 nsew default tristate
rlabel metal2 s 316930 -960 317042 480 8 la_data_out[53]
port 349 nsew default tristate
rlabel metal2 s 320426 -960 320538 480 8 la_data_out[54]
port 350 nsew default tristate
rlabel metal2 s 324014 -960 324126 480 8 la_data_out[55]
port 351 nsew default tristate
rlabel metal2 s 327602 -960 327714 480 8 la_data_out[56]
port 352 nsew default tristate
rlabel metal2 s 331190 -960 331302 480 8 la_data_out[57]
port 353 nsew default tristate
rlabel metal2 s 334686 -960 334798 480 8 la_data_out[58]
port 354 nsew default tristate
rlabel metal2 s 338274 -960 338386 480 8 la_data_out[59]
port 355 nsew default tristate
rlabel metal2 s 145626 -960 145738 480 8 la_data_out[5]
port 356 nsew default tristate
rlabel metal2 s 341862 -960 341974 480 8 la_data_out[60]
port 357 nsew default tristate
rlabel metal2 s 345450 -960 345562 480 8 la_data_out[61]
port 358 nsew default tristate
rlabel metal2 s 349038 -960 349150 480 8 la_data_out[62]
port 359 nsew default tristate
rlabel metal2 s 352534 -960 352646 480 8 la_data_out[63]
port 360 nsew default tristate
rlabel metal2 s 356122 -960 356234 480 8 la_data_out[64]
port 361 nsew default tristate
rlabel metal2 s 359710 -960 359822 480 8 la_data_out[65]
port 362 nsew default tristate
rlabel metal2 s 363298 -960 363410 480 8 la_data_out[66]
port 363 nsew default tristate
rlabel metal2 s 366886 -960 366998 480 8 la_data_out[67]
port 364 nsew default tristate
rlabel metal2 s 370382 -960 370494 480 8 la_data_out[68]
port 365 nsew default tristate
rlabel metal2 s 373970 -960 374082 480 8 la_data_out[69]
port 366 nsew default tristate
rlabel metal2 s 149214 -960 149326 480 8 la_data_out[6]
port 367 nsew default tristate
rlabel metal2 s 377558 -960 377670 480 8 la_data_out[70]
port 368 nsew default tristate
rlabel metal2 s 381146 -960 381258 480 8 la_data_out[71]
port 369 nsew default tristate
rlabel metal2 s 384642 -960 384754 480 8 la_data_out[72]
port 370 nsew default tristate
rlabel metal2 s 388230 -960 388342 480 8 la_data_out[73]
port 371 nsew default tristate
rlabel metal2 s 391818 -960 391930 480 8 la_data_out[74]
port 372 nsew default tristate
rlabel metal2 s 395406 -960 395518 480 8 la_data_out[75]
port 373 nsew default tristate
rlabel metal2 s 398994 -960 399106 480 8 la_data_out[76]
port 374 nsew default tristate
rlabel metal2 s 402490 -960 402602 480 8 la_data_out[77]
port 375 nsew default tristate
rlabel metal2 s 406078 -960 406190 480 8 la_data_out[78]
port 376 nsew default tristate
rlabel metal2 s 409666 -960 409778 480 8 la_data_out[79]
port 377 nsew default tristate
rlabel metal2 s 152710 -960 152822 480 8 la_data_out[7]
port 378 nsew default tristate
rlabel metal2 s 413254 -960 413366 480 8 la_data_out[80]
port 379 nsew default tristate
rlabel metal2 s 416842 -960 416954 480 8 la_data_out[81]
port 380 nsew default tristate
rlabel metal2 s 420338 -960 420450 480 8 la_data_out[82]
port 381 nsew default tristate
rlabel metal2 s 423926 -960 424038 480 8 la_data_out[83]
port 382 nsew default tristate
rlabel metal2 s 427514 -960 427626 480 8 la_data_out[84]
port 383 nsew default tristate
rlabel metal2 s 431102 -960 431214 480 8 la_data_out[85]
port 384 nsew default tristate
rlabel metal2 s 434598 -960 434710 480 8 la_data_out[86]
port 385 nsew default tristate
rlabel metal2 s 438186 -960 438298 480 8 la_data_out[87]
port 386 nsew default tristate
rlabel metal2 s 441774 -960 441886 480 8 la_data_out[88]
port 387 nsew default tristate
rlabel metal2 s 445362 -960 445474 480 8 la_data_out[89]
port 388 nsew default tristate
rlabel metal2 s 156298 -960 156410 480 8 la_data_out[8]
port 389 nsew default tristate
rlabel metal2 s 448950 -960 449062 480 8 la_data_out[90]
port 390 nsew default tristate
rlabel metal2 s 452446 -960 452558 480 8 la_data_out[91]
port 391 nsew default tristate
rlabel metal2 s 456034 -960 456146 480 8 la_data_out[92]
port 392 nsew default tristate
rlabel metal2 s 459622 -960 459734 480 8 la_data_out[93]
port 393 nsew default tristate
rlabel metal2 s 463210 -960 463322 480 8 la_data_out[94]
port 394 nsew default tristate
rlabel metal2 s 466798 -960 466910 480 8 la_data_out[95]
port 395 nsew default tristate
rlabel metal2 s 470294 -960 470406 480 8 la_data_out[96]
port 396 nsew default tristate
rlabel metal2 s 473882 -960 473994 480 8 la_data_out[97]
port 397 nsew default tristate
rlabel metal2 s 477470 -960 477582 480 8 la_data_out[98]
port 398 nsew default tristate
rlabel metal2 s 481058 -960 481170 480 8 la_data_out[99]
port 399 nsew default tristate
rlabel metal2 s 159886 -960 159998 480 8 la_data_out[9]
port 400 nsew default tristate
rlabel metal2 s 128974 -960 129086 480 8 la_oen[0]
port 401 nsew default input
rlabel metal2 s 485750 -960 485862 480 8 la_oen[100]
port 402 nsew default input
rlabel metal2 s 489338 -960 489450 480 8 la_oen[101]
port 403 nsew default input
rlabel metal2 s 492926 -960 493038 480 8 la_oen[102]
port 404 nsew default input
rlabel metal2 s 496514 -960 496626 480 8 la_oen[103]
port 405 nsew default input
rlabel metal2 s 500102 -960 500214 480 8 la_oen[104]
port 406 nsew default input
rlabel metal2 s 503598 -960 503710 480 8 la_oen[105]
port 407 nsew default input
rlabel metal2 s 507186 -960 507298 480 8 la_oen[106]
port 408 nsew default input
rlabel metal2 s 510774 -960 510886 480 8 la_oen[107]
port 409 nsew default input
rlabel metal2 s 514362 -960 514474 480 8 la_oen[108]
port 410 nsew default input
rlabel metal2 s 517858 -960 517970 480 8 la_oen[109]
port 411 nsew default input
rlabel metal2 s 164670 -960 164782 480 8 la_oen[10]
port 412 nsew default input
rlabel metal2 s 521446 -960 521558 480 8 la_oen[110]
port 413 nsew default input
rlabel metal2 s 525034 -960 525146 480 8 la_oen[111]
port 414 nsew default input
rlabel metal2 s 528622 -960 528734 480 8 la_oen[112]
port 415 nsew default input
rlabel metal2 s 532210 -960 532322 480 8 la_oen[113]
port 416 nsew default input
rlabel metal2 s 535706 -960 535818 480 8 la_oen[114]
port 417 nsew default input
rlabel metal2 s 539294 -960 539406 480 8 la_oen[115]
port 418 nsew default input
rlabel metal2 s 542882 -960 542994 480 8 la_oen[116]
port 419 nsew default input
rlabel metal2 s 546470 -960 546582 480 8 la_oen[117]
port 420 nsew default input
rlabel metal2 s 550058 -960 550170 480 8 la_oen[118]
port 421 nsew default input
rlabel metal2 s 553554 -960 553666 480 8 la_oen[119]
port 422 nsew default input
rlabel metal2 s 168166 -960 168278 480 8 la_oen[11]
port 423 nsew default input
rlabel metal2 s 557142 -960 557254 480 8 la_oen[120]
port 424 nsew default input
rlabel metal2 s 560730 -960 560842 480 8 la_oen[121]
port 425 nsew default input
rlabel metal2 s 564318 -960 564430 480 8 la_oen[122]
port 426 nsew default input
rlabel metal2 s 567814 -960 567926 480 8 la_oen[123]
port 427 nsew default input
rlabel metal2 s 571402 -960 571514 480 8 la_oen[124]
port 428 nsew default input
rlabel metal2 s 574990 -960 575102 480 8 la_oen[125]
port 429 nsew default input
rlabel metal2 s 578578 -960 578690 480 8 la_oen[126]
port 430 nsew default input
rlabel metal2 s 582166 -960 582278 480 8 la_oen[127]
port 431 nsew default input
rlabel metal2 s 171754 -960 171866 480 8 la_oen[12]
port 432 nsew default input
rlabel metal2 s 175342 -960 175454 480 8 la_oen[13]
port 433 nsew default input
rlabel metal2 s 178930 -960 179042 480 8 la_oen[14]
port 434 nsew default input
rlabel metal2 s 182518 -960 182630 480 8 la_oen[15]
port 435 nsew default input
rlabel metal2 s 186014 -960 186126 480 8 la_oen[16]
port 436 nsew default input
rlabel metal2 s 189602 -960 189714 480 8 la_oen[17]
port 437 nsew default input
rlabel metal2 s 193190 -960 193302 480 8 la_oen[18]
port 438 nsew default input
rlabel metal2 s 196778 -960 196890 480 8 la_oen[19]
port 439 nsew default input
rlabel metal2 s 132562 -960 132674 480 8 la_oen[1]
port 440 nsew default input
rlabel metal2 s 200366 -960 200478 480 8 la_oen[20]
port 441 nsew default input
rlabel metal2 s 203862 -960 203974 480 8 la_oen[21]
port 442 nsew default input
rlabel metal2 s 207450 -960 207562 480 8 la_oen[22]
port 443 nsew default input
rlabel metal2 s 211038 -960 211150 480 8 la_oen[23]
port 444 nsew default input
rlabel metal2 s 214626 -960 214738 480 8 la_oen[24]
port 445 nsew default input
rlabel metal2 s 218122 -960 218234 480 8 la_oen[25]
port 446 nsew default input
rlabel metal2 s 221710 -960 221822 480 8 la_oen[26]
port 447 nsew default input
rlabel metal2 s 225298 -960 225410 480 8 la_oen[27]
port 448 nsew default input
rlabel metal2 s 228886 -960 228998 480 8 la_oen[28]
port 449 nsew default input
rlabel metal2 s 232474 -960 232586 480 8 la_oen[29]
port 450 nsew default input
rlabel metal2 s 136058 -960 136170 480 8 la_oen[2]
port 451 nsew default input
rlabel metal2 s 235970 -960 236082 480 8 la_oen[30]
port 452 nsew default input
rlabel metal2 s 239558 -960 239670 480 8 la_oen[31]
port 453 nsew default input
rlabel metal2 s 243146 -960 243258 480 8 la_oen[32]
port 454 nsew default input
rlabel metal2 s 246734 -960 246846 480 8 la_oen[33]
port 455 nsew default input
rlabel metal2 s 250322 -960 250434 480 8 la_oen[34]
port 456 nsew default input
rlabel metal2 s 253818 -960 253930 480 8 la_oen[35]
port 457 nsew default input
rlabel metal2 s 257406 -960 257518 480 8 la_oen[36]
port 458 nsew default input
rlabel metal2 s 260994 -960 261106 480 8 la_oen[37]
port 459 nsew default input
rlabel metal2 s 264582 -960 264694 480 8 la_oen[38]
port 460 nsew default input
rlabel metal2 s 268078 -960 268190 480 8 la_oen[39]
port 461 nsew default input
rlabel metal2 s 139646 -960 139758 480 8 la_oen[3]
port 462 nsew default input
rlabel metal2 s 271666 -960 271778 480 8 la_oen[40]
port 463 nsew default input
rlabel metal2 s 275254 -960 275366 480 8 la_oen[41]
port 464 nsew default input
rlabel metal2 s 278842 -960 278954 480 8 la_oen[42]
port 465 nsew default input
rlabel metal2 s 282430 -960 282542 480 8 la_oen[43]
port 466 nsew default input
rlabel metal2 s 285926 -960 286038 480 8 la_oen[44]
port 467 nsew default input
rlabel metal2 s 289514 -960 289626 480 8 la_oen[45]
port 468 nsew default input
rlabel metal2 s 293102 -960 293214 480 8 la_oen[46]
port 469 nsew default input
rlabel metal2 s 296690 -960 296802 480 8 la_oen[47]
port 470 nsew default input
rlabel metal2 s 300278 -960 300390 480 8 la_oen[48]
port 471 nsew default input
rlabel metal2 s 303774 -960 303886 480 8 la_oen[49]
port 472 nsew default input
rlabel metal2 s 143234 -960 143346 480 8 la_oen[4]
port 473 nsew default input
rlabel metal2 s 307362 -960 307474 480 8 la_oen[50]
port 474 nsew default input
rlabel metal2 s 310950 -960 311062 480 8 la_oen[51]
port 475 nsew default input
rlabel metal2 s 314538 -960 314650 480 8 la_oen[52]
port 476 nsew default input
rlabel metal2 s 318034 -960 318146 480 8 la_oen[53]
port 477 nsew default input
rlabel metal2 s 321622 -960 321734 480 8 la_oen[54]
port 478 nsew default input
rlabel metal2 s 325210 -960 325322 480 8 la_oen[55]
port 479 nsew default input
rlabel metal2 s 328798 -960 328910 480 8 la_oen[56]
port 480 nsew default input
rlabel metal2 s 332386 -960 332498 480 8 la_oen[57]
port 481 nsew default input
rlabel metal2 s 335882 -960 335994 480 8 la_oen[58]
port 482 nsew default input
rlabel metal2 s 339470 -960 339582 480 8 la_oen[59]
port 483 nsew default input
rlabel metal2 s 146822 -960 146934 480 8 la_oen[5]
port 484 nsew default input
rlabel metal2 s 343058 -960 343170 480 8 la_oen[60]
port 485 nsew default input
rlabel metal2 s 346646 -960 346758 480 8 la_oen[61]
port 486 nsew default input
rlabel metal2 s 350234 -960 350346 480 8 la_oen[62]
port 487 nsew default input
rlabel metal2 s 353730 -960 353842 480 8 la_oen[63]
port 488 nsew default input
rlabel metal2 s 357318 -960 357430 480 8 la_oen[64]
port 489 nsew default input
rlabel metal2 s 360906 -960 361018 480 8 la_oen[65]
port 490 nsew default input
rlabel metal2 s 364494 -960 364606 480 8 la_oen[66]
port 491 nsew default input
rlabel metal2 s 367990 -960 368102 480 8 la_oen[67]
port 492 nsew default input
rlabel metal2 s 371578 -960 371690 480 8 la_oen[68]
port 493 nsew default input
rlabel metal2 s 375166 -960 375278 480 8 la_oen[69]
port 494 nsew default input
rlabel metal2 s 150410 -960 150522 480 8 la_oen[6]
port 495 nsew default input
rlabel metal2 s 378754 -960 378866 480 8 la_oen[70]
port 496 nsew default input
rlabel metal2 s 382342 -960 382454 480 8 la_oen[71]
port 497 nsew default input
rlabel metal2 s 385838 -960 385950 480 8 la_oen[72]
port 498 nsew default input
rlabel metal2 s 389426 -960 389538 480 8 la_oen[73]
port 499 nsew default input
rlabel metal2 s 393014 -960 393126 480 8 la_oen[74]
port 500 nsew default input
rlabel metal2 s 396602 -960 396714 480 8 la_oen[75]
port 501 nsew default input
rlabel metal2 s 400190 -960 400302 480 8 la_oen[76]
port 502 nsew default input
rlabel metal2 s 403686 -960 403798 480 8 la_oen[77]
port 503 nsew default input
rlabel metal2 s 407274 -960 407386 480 8 la_oen[78]
port 504 nsew default input
rlabel metal2 s 410862 -960 410974 480 8 la_oen[79]
port 505 nsew default input
rlabel metal2 s 153906 -960 154018 480 8 la_oen[7]
port 506 nsew default input
rlabel metal2 s 414450 -960 414562 480 8 la_oen[80]
port 507 nsew default input
rlabel metal2 s 417946 -960 418058 480 8 la_oen[81]
port 508 nsew default input
rlabel metal2 s 421534 -960 421646 480 8 la_oen[82]
port 509 nsew default input
rlabel metal2 s 425122 -960 425234 480 8 la_oen[83]
port 510 nsew default input
rlabel metal2 s 428710 -960 428822 480 8 la_oen[84]
port 511 nsew default input
rlabel metal2 s 432298 -960 432410 480 8 la_oen[85]
port 512 nsew default input
rlabel metal2 s 435794 -960 435906 480 8 la_oen[86]
port 513 nsew default input
rlabel metal2 s 439382 -960 439494 480 8 la_oen[87]
port 514 nsew default input
rlabel metal2 s 442970 -960 443082 480 8 la_oen[88]
port 515 nsew default input
rlabel metal2 s 446558 -960 446670 480 8 la_oen[89]
port 516 nsew default input
rlabel metal2 s 157494 -960 157606 480 8 la_oen[8]
port 517 nsew default input
rlabel metal2 s 450146 -960 450258 480 8 la_oen[90]
port 518 nsew default input
rlabel metal2 s 453642 -960 453754 480 8 la_oen[91]
port 519 nsew default input
rlabel metal2 s 457230 -960 457342 480 8 la_oen[92]
port 520 nsew default input
rlabel metal2 s 460818 -960 460930 480 8 la_oen[93]
port 521 nsew default input
rlabel metal2 s 464406 -960 464518 480 8 la_oen[94]
port 522 nsew default input
rlabel metal2 s 467902 -960 468014 480 8 la_oen[95]
port 523 nsew default input
rlabel metal2 s 471490 -960 471602 480 8 la_oen[96]
port 524 nsew default input
rlabel metal2 s 475078 -960 475190 480 8 la_oen[97]
port 525 nsew default input
rlabel metal2 s 478666 -960 478778 480 8 la_oen[98]
port 526 nsew default input
rlabel metal2 s 482254 -960 482366 480 8 la_oen[99]
port 527 nsew default input
rlabel metal2 s 161082 -960 161194 480 8 la_oen[9]
port 528 nsew default input
rlabel metal2 s 583362 -960 583474 480 8 user_clock2
port 529 nsew default input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 530 nsew default input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 531 nsew default input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 532 nsew default tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 533 nsew default input
rlabel metal2 s 48106 -960 48218 480 8 wbs_adr_i[10]
port 534 nsew default input
rlabel metal2 s 51602 -960 51714 480 8 wbs_adr_i[11]
port 535 nsew default input
rlabel metal2 s 55190 -960 55302 480 8 wbs_adr_i[12]
port 536 nsew default input
rlabel metal2 s 58778 -960 58890 480 8 wbs_adr_i[13]
port 537 nsew default input
rlabel metal2 s 62366 -960 62478 480 8 wbs_adr_i[14]
port 538 nsew default input
rlabel metal2 s 65954 -960 66066 480 8 wbs_adr_i[15]
port 539 nsew default input
rlabel metal2 s 69450 -960 69562 480 8 wbs_adr_i[16]
port 540 nsew default input
rlabel metal2 s 73038 -960 73150 480 8 wbs_adr_i[17]
port 541 nsew default input
rlabel metal2 s 76626 -960 76738 480 8 wbs_adr_i[18]
port 542 nsew default input
rlabel metal2 s 80214 -960 80326 480 8 wbs_adr_i[19]
port 543 nsew default input
rlabel metal2 s 12410 -960 12522 480 8 wbs_adr_i[1]
port 544 nsew default input
rlabel metal2 s 83802 -960 83914 480 8 wbs_adr_i[20]
port 545 nsew default input
rlabel metal2 s 87298 -960 87410 480 8 wbs_adr_i[21]
port 546 nsew default input
rlabel metal2 s 90886 -960 90998 480 8 wbs_adr_i[22]
port 547 nsew default input
rlabel metal2 s 94474 -960 94586 480 8 wbs_adr_i[23]
port 548 nsew default input
rlabel metal2 s 98062 -960 98174 480 8 wbs_adr_i[24]
port 549 nsew default input
rlabel metal2 s 101558 -960 101670 480 8 wbs_adr_i[25]
port 550 nsew default input
rlabel metal2 s 105146 -960 105258 480 8 wbs_adr_i[26]
port 551 nsew default input
rlabel metal2 s 108734 -960 108846 480 8 wbs_adr_i[27]
port 552 nsew default input
rlabel metal2 s 112322 -960 112434 480 8 wbs_adr_i[28]
port 553 nsew default input
rlabel metal2 s 115910 -960 116022 480 8 wbs_adr_i[29]
port 554 nsew default input
rlabel metal2 s 17194 -960 17306 480 8 wbs_adr_i[2]
port 555 nsew default input
rlabel metal2 s 119406 -960 119518 480 8 wbs_adr_i[30]
port 556 nsew default input
rlabel metal2 s 122994 -960 123106 480 8 wbs_adr_i[31]
port 557 nsew default input
rlabel metal2 s 21886 -960 21998 480 8 wbs_adr_i[3]
port 558 nsew default input
rlabel metal2 s 26670 -960 26782 480 8 wbs_adr_i[4]
port 559 nsew default input
rlabel metal2 s 30258 -960 30370 480 8 wbs_adr_i[5]
port 560 nsew default input
rlabel metal2 s 33846 -960 33958 480 8 wbs_adr_i[6]
port 561 nsew default input
rlabel metal2 s 37342 -960 37454 480 8 wbs_adr_i[7]
port 562 nsew default input
rlabel metal2 s 40930 -960 41042 480 8 wbs_adr_i[8]
port 563 nsew default input
rlabel metal2 s 44518 -960 44630 480 8 wbs_adr_i[9]
port 564 nsew default input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 565 nsew default input
rlabel metal2 s 8822 -960 8934 480 8 wbs_dat_i[0]
port 566 nsew default input
rlabel metal2 s 49302 -960 49414 480 8 wbs_dat_i[10]
port 567 nsew default input
rlabel metal2 s 52798 -960 52910 480 8 wbs_dat_i[11]
port 568 nsew default input
rlabel metal2 s 56386 -960 56498 480 8 wbs_dat_i[12]
port 569 nsew default input
rlabel metal2 s 59974 -960 60086 480 8 wbs_dat_i[13]
port 570 nsew default input
rlabel metal2 s 63562 -960 63674 480 8 wbs_dat_i[14]
port 571 nsew default input
rlabel metal2 s 67150 -960 67262 480 8 wbs_dat_i[15]
port 572 nsew default input
rlabel metal2 s 70646 -960 70758 480 8 wbs_dat_i[16]
port 573 nsew default input
rlabel metal2 s 74234 -960 74346 480 8 wbs_dat_i[17]
port 574 nsew default input
rlabel metal2 s 77822 -960 77934 480 8 wbs_dat_i[18]
port 575 nsew default input
rlabel metal2 s 81410 -960 81522 480 8 wbs_dat_i[19]
port 576 nsew default input
rlabel metal2 s 13606 -960 13718 480 8 wbs_dat_i[1]
port 577 nsew default input
rlabel metal2 s 84906 -960 85018 480 8 wbs_dat_i[20]
port 578 nsew default input
rlabel metal2 s 88494 -960 88606 480 8 wbs_dat_i[21]
port 579 nsew default input
rlabel metal2 s 92082 -960 92194 480 8 wbs_dat_i[22]
port 580 nsew default input
rlabel metal2 s 95670 -960 95782 480 8 wbs_dat_i[23]
port 581 nsew default input
rlabel metal2 s 99258 -960 99370 480 8 wbs_dat_i[24]
port 582 nsew default input
rlabel metal2 s 102754 -960 102866 480 8 wbs_dat_i[25]
port 583 nsew default input
rlabel metal2 s 106342 -960 106454 480 8 wbs_dat_i[26]
port 584 nsew default input
rlabel metal2 s 109930 -960 110042 480 8 wbs_dat_i[27]
port 585 nsew default input
rlabel metal2 s 113518 -960 113630 480 8 wbs_dat_i[28]
port 586 nsew default input
rlabel metal2 s 117106 -960 117218 480 8 wbs_dat_i[29]
port 587 nsew default input
rlabel metal2 s 18298 -960 18410 480 8 wbs_dat_i[2]
port 588 nsew default input
rlabel metal2 s 120602 -960 120714 480 8 wbs_dat_i[30]
port 589 nsew default input
rlabel metal2 s 124190 -960 124302 480 8 wbs_dat_i[31]
port 590 nsew default input
rlabel metal2 s 23082 -960 23194 480 8 wbs_dat_i[3]
port 591 nsew default input
rlabel metal2 s 27866 -960 27978 480 8 wbs_dat_i[4]
port 592 nsew default input
rlabel metal2 s 31454 -960 31566 480 8 wbs_dat_i[5]
port 593 nsew default input
rlabel metal2 s 34950 -960 35062 480 8 wbs_dat_i[6]
port 594 nsew default input
rlabel metal2 s 38538 -960 38650 480 8 wbs_dat_i[7]
port 595 nsew default input
rlabel metal2 s 42126 -960 42238 480 8 wbs_dat_i[8]
port 596 nsew default input
rlabel metal2 s 45714 -960 45826 480 8 wbs_dat_i[9]
port 597 nsew default input
rlabel metal2 s 10018 -960 10130 480 8 wbs_dat_o[0]
port 598 nsew default tristate
rlabel metal2 s 50498 -960 50610 480 8 wbs_dat_o[10]
port 599 nsew default tristate
rlabel metal2 s 53994 -960 54106 480 8 wbs_dat_o[11]
port 600 nsew default tristate
rlabel metal2 s 57582 -960 57694 480 8 wbs_dat_o[12]
port 601 nsew default tristate
rlabel metal2 s 61170 -960 61282 480 8 wbs_dat_o[13]
port 602 nsew default tristate
rlabel metal2 s 64758 -960 64870 480 8 wbs_dat_o[14]
port 603 nsew default tristate
rlabel metal2 s 68254 -960 68366 480 8 wbs_dat_o[15]
port 604 nsew default tristate
rlabel metal2 s 71842 -960 71954 480 8 wbs_dat_o[16]
port 605 nsew default tristate
rlabel metal2 s 75430 -960 75542 480 8 wbs_dat_o[17]
port 606 nsew default tristate
rlabel metal2 s 79018 -960 79130 480 8 wbs_dat_o[18]
port 607 nsew default tristate
rlabel metal2 s 82606 -960 82718 480 8 wbs_dat_o[19]
port 608 nsew default tristate
rlabel metal2 s 14802 -960 14914 480 8 wbs_dat_o[1]
port 609 nsew default tristate
rlabel metal2 s 86102 -960 86214 480 8 wbs_dat_o[20]
port 610 nsew default tristate
rlabel metal2 s 89690 -960 89802 480 8 wbs_dat_o[21]
port 611 nsew default tristate
rlabel metal2 s 93278 -960 93390 480 8 wbs_dat_o[22]
port 612 nsew default tristate
rlabel metal2 s 96866 -960 96978 480 8 wbs_dat_o[23]
port 613 nsew default tristate
rlabel metal2 s 100454 -960 100566 480 8 wbs_dat_o[24]
port 614 nsew default tristate
rlabel metal2 s 103950 -960 104062 480 8 wbs_dat_o[25]
port 615 nsew default tristate
rlabel metal2 s 107538 -960 107650 480 8 wbs_dat_o[26]
port 616 nsew default tristate
rlabel metal2 s 111126 -960 111238 480 8 wbs_dat_o[27]
port 617 nsew default tristate
rlabel metal2 s 114714 -960 114826 480 8 wbs_dat_o[28]
port 618 nsew default tristate
rlabel metal2 s 118210 -960 118322 480 8 wbs_dat_o[29]
port 619 nsew default tristate
rlabel metal2 s 19494 -960 19606 480 8 wbs_dat_o[2]
port 620 nsew default tristate
rlabel metal2 s 121798 -960 121910 480 8 wbs_dat_o[30]
port 621 nsew default tristate
rlabel metal2 s 125386 -960 125498 480 8 wbs_dat_o[31]
port 622 nsew default tristate
rlabel metal2 s 24278 -960 24390 480 8 wbs_dat_o[3]
port 623 nsew default tristate
rlabel metal2 s 29062 -960 29174 480 8 wbs_dat_o[4]
port 624 nsew default tristate
rlabel metal2 s 32650 -960 32762 480 8 wbs_dat_o[5]
port 625 nsew default tristate
rlabel metal2 s 36146 -960 36258 480 8 wbs_dat_o[6]
port 626 nsew default tristate
rlabel metal2 s 39734 -960 39846 480 8 wbs_dat_o[7]
port 627 nsew default tristate
rlabel metal2 s 43322 -960 43434 480 8 wbs_dat_o[8]
port 628 nsew default tristate
rlabel metal2 s 46910 -960 47022 480 8 wbs_dat_o[9]
port 629 nsew default tristate
rlabel metal2 s 11214 -960 11326 480 8 wbs_sel_i[0]
port 630 nsew default input
rlabel metal2 s 15998 -960 16110 480 8 wbs_sel_i[1]
port 631 nsew default input
rlabel metal2 s 20690 -960 20802 480 8 wbs_sel_i[2]
port 632 nsew default input
rlabel metal2 s 25474 -960 25586 480 8 wbs_sel_i[3]
port 633 nsew default input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 634 nsew default input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 635 nsew default input
rlabel metal5 s -1996 -924 585920 -324 8 vccd1
port 636 nsew default input
rlabel metal5 s -2916 -1844 586840 -1244 8 vssd1
port 637 nsew default input
rlabel metal5 s -3836 -2764 587760 -2164 8 vccd2
port 638 nsew default input
rlabel metal5 s -4756 -3684 588680 -3084 8 vssd2
port 639 nsew default input
rlabel metal5 s -5676 -4604 589600 -4004 8 vdda1
port 640 nsew default input
rlabel metal5 s -6596 -5524 590520 -4924 8 vssa1
port 641 nsew default input
rlabel metal5 s -7516 -6444 591440 -5844 8 vdda2
port 642 nsew default input
rlabel metal5 s -8436 -7364 592360 -6764 8 vssa2
port 643 nsew default input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
