magic
tech sky130A
timestamp 1607784188
<< end >>
