VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO LATCH
  CLASS CORE ;
  FOREIGN LATCH ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.440 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 6.440 2.960 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 6.440 0.240 ;
    END
  END gnd
  PIN Q
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 5.840 2.050 6.130 2.310 ;
        RECT 4.530 2.020 6.130 2.050 ;
        RECT 4.530 1.910 6.050 2.020 ;
        RECT 4.530 1.770 4.670 1.910 ;
        RECT 4.460 1.480 4.750 1.770 ;
        RECT 4.530 1.230 4.670 1.480 ;
        RECT 4.460 0.940 4.750 1.230 ;
        RECT 5.910 0.690 6.050 1.910 ;
        RECT 5.840 0.400 6.130 0.690 ;
    END
  END Q
  PIN CLK
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 3.540 1.480 3.830 1.770 ;
    END
    PORT
      LAYER met1 ;
        RECT 0.780 0.940 1.070 1.230 ;
        RECT 0.850 0.790 0.990 0.940 ;
        RECT 2.620 0.790 2.910 0.870 ;
        RECT 0.850 0.650 2.910 0.790 ;
        RECT 2.620 0.580 2.910 0.650 ;
    END
  END CLK
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 1.700 0.940 1.990 1.230 ;
    END
  END D
END LATCH
END LIBRARY

