MACRO HAX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN HAX1 0 0 ;
 SITE CORE ;
 SYMMETRY X Y R90 ;
  PIN VDD
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.00000000 2.52500000 9.20000000 2.91500000 ;
    END
  END VDD

  PIN GND
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.00000000 -0.19500000 9.20000000 0.19500000 ;
    END
  END GND

  PIN YS
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        POLYGON 8.62500000 0.60000000 8.62500000 0.83000000 8.67000000 0.83000000 8.67000000 1.90000000 8.62500000 1.90000000 8.62500000 2.13000000 8.85500000 2.13000000 8.85500000 1.90000000 8.81000000 1.90000000 8.81000000 0.83000000 8.85500000 0.83000000 8.85500000 0.60000000 ;
    END
  END YS

  PIN YC
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 1.26500000 0.60000000 1.49500000 0.83000000 ;
       LAYER metal2 ;
        RECT 1.26500000 1.90000000 1.49500000 2.13000000 ;
    END
  END YC

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        POLYGON 3.56500000 1.51000000 3.56500000 1.74000000 3.79500000 1.74000000 3.79500000 1.69500000 5.40500000 1.69500000 5.40500000 1.74000000 5.63500000 1.74000000 5.63500000 1.51000000 5.40500000 1.51000000 5.40500000 1.55500000 3.79500000 1.55500000 3.79500000 1.51000000 ;
    END
  END A

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 2.64500000 1.51000000 2.87500000 1.74000000 ;
       LAYER metal2 ;
        RECT 6.32500000 1.51000000 6.55500000 1.74000000 ;
    END
  END B


END HAX1
