MACRO NOR3X1
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN NOR3X1 0 0 ;
 SITE CORE ;
 SYMMETRY X Y R90 ;
  PIN VDD
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.00000000 2.52500000 6.44000000 2.91500000 ;
    END
  END VDD

  PIN GND
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.00000000 -0.19500000 6.44000000 0.19500000 ;
    END
  END GND

  PIN Y
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        POLYGON 1.26500000 0.60000000 1.26500000 0.83000000 1.31000000 0.83000000 1.31000000 1.42500000 0.39000000 1.42500000 0.39000000 1.90000000 0.34500000 1.90000000 0.34500000 2.13000000 0.57500000 2.13000000 0.57500000 1.90000000 0.53000000 1.90000000 0.53000000 1.56500000 1.45000000 1.56500000 1.45000000 0.83000000 1.49500000 0.83000000 1.49500000 0.60000000 ;
       LAYER metal2 ;
        RECT 3.10500000 0.60000000 3.33500000 0.83000000 ;
       LAYER metal2 ;
        RECT 5.86500000 1.90000000 6.09500000 2.13000000 ;
    END
  END Y

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        POLYGON 2.64500000 1.38000000 2.64500000 1.61000000 2.87500000 1.61000000 2.87500000 1.56500000 3.56500000 1.56500000 3.56500000 1.61000000 3.79500000 1.61000000 3.79500000 1.38000000 3.56500000 1.38000000 3.56500000 1.42500000 2.87500000 1.42500000 2.87500000 1.38000000 ;
    END
  END A

  PIN C
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.80500000 0.99000000 1.03500000 1.22000000 ;
       LAYER metal2 ;
        RECT 5.40500000 1.51000000 5.63500000 1.74000000 ;
    END
  END C

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 4.48500000 1.38000000 4.71500000 1.61000000 ;
       LAYER metal2 ;
        RECT 1.72500000 0.99000000 1.95500000 1.22000000 ;
    END
  END B


END NOR3X1
