magic
tech sky130A
timestamp 1607799982
<< end >>
