MACRO INVX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN INVX1 0 0 ;
 SIZE 2.08 BY 4.16 ;
 SYMMETRY X Y R90 ;
 SITE unithd ;
  PIN vdd
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 0.00000000 3965.00000000 2080.00000000 4355.00000000 ;
    END
  END vdd

  PIN gnd
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 0.00000000 -195.00000000 2080.00000000 195.00000000 ;
    END
  END gnd

  PIN Y
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        POLYGON 1445.00000000 730.00000000 1445.00000000 960.00000000 1490.00000000 960.00000000 1490.00000000 3200.00000000 1445.00000000 3200.00000000 1445.00000000 3430.00000000 1675.00000000 3430.00000000 1675.00000000 3200.00000000 1630.00000000 3200.00000000 1630.00000000 960.00000000 1675.00000000 960.00000000 1675.00000000 730.00000000 ;
    END
  END Y

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        POLYGON 925.00000000 1120.00000000 925.00000000 1350.00000000 970.00000000 1350.00000000 970.00000000 2810.00000000 925.00000000 2810.00000000 925.00000000 3040.00000000 1155.00000000 3040.00000000 1155.00000000 2810.00000000 1110.00000000 2810.00000000 1110.00000000 1350.00000000 1155.00000000 1350.00000000 1155.00000000 1120.00000000 ;
    END
  END A


END INVX1
