magic
tech sky130A
magscale 1 2
timestamp 1607592090
<< locali >>
rect 219081 685899 219115 695453
rect 154313 676243 154347 685797
rect 218989 666587 219023 676141
rect 299857 666587 299891 684437
rect 219265 647275 219299 656829
rect 219357 616879 219391 626501
rect 219081 608719 219115 611405
rect 219265 601579 219299 608549
rect 299673 601715 299707 608549
rect 219173 589339 219207 598893
rect 299857 589339 299891 598893
rect 154313 579751 154347 589237
rect 218897 569959 218931 579581
rect 218897 550647 218931 553401
rect 154405 521679 154439 531233
rect 154405 502367 154439 511921
rect 219081 505087 219115 510561
rect 299673 485775 299707 492609
rect 299673 466395 299707 473297
rect 154221 444431 154255 453985
rect 218989 444431 219023 453985
rect 299489 440283 299523 449837
rect 154405 427771 154439 434673
rect 299581 427771 299615 436781
rect 154313 405739 154347 415361
rect 299673 405739 299707 415361
rect 260113 402611 260147 402781
rect 261125 402475 261159 402985
rect 262229 402611 262263 402781
rect 261861 402135 261895 402577
rect 248337 401931 248371 402101
rect 262781 402067 262815 402509
rect 244841 401863 244875 401897
rect 244841 401829 245485 401863
rect 248187 401761 248337 401795
rect 248187 401625 248337 401659
rect 235457 399279 235491 399449
rect 234169 399007 234203 399245
rect 234537 399075 234571 399245
rect 242081 398871 242115 399857
rect 282469 399143 282503 399313
rect 288357 399211 288391 399313
rect 288725 398939 288759 399313
rect 237297 337807 237331 337909
rect 237665 337739 237699 338045
rect 268393 337875 268427 338045
rect 273177 337807 273211 337977
rect 235917 337331 235951 337569
rect 235825 336175 235859 336549
rect 240057 335427 240091 337093
rect 229569 328491 229603 335393
rect 233985 327131 234019 334305
rect 248797 332163 248831 335665
rect 251741 334951 251775 335937
rect 250545 328491 250579 333285
rect 254685 328491 254719 335733
rect 237021 318835 237055 328389
rect 245209 320331 245243 328389
rect 229477 310811 229511 318733
rect 229477 299523 229511 309077
rect 235273 301971 235307 317373
rect 245209 311831 245243 318733
rect 254869 316115 254903 333897
rect 255881 328491 255915 335665
rect 261769 328491 261803 337297
rect 262505 336311 262539 337569
rect 262873 336719 262907 337501
rect 265173 335359 265207 337433
rect 265633 336787 265667 337705
rect 265449 327403 265483 335665
rect 266277 327131 266311 336685
rect 266829 334883 266863 336685
rect 267473 332299 267507 337501
rect 268301 337059 268335 337569
rect 269037 327131 269071 336685
rect 272533 335495 272567 337637
rect 273269 337127 273303 337909
rect 275293 337875 275327 337977
rect 275937 337535 275971 337773
rect 271889 332231 271923 332401
rect 273177 327131 273211 336685
rect 274373 327131 274407 336685
rect 274741 336583 274775 337501
rect 277041 335427 277075 338521
rect 277317 335359 277351 338113
rect 282963 338045 283055 338079
rect 282595 337977 282779 338011
rect 277869 337331 277903 337705
rect 280537 335359 280571 337705
rect 280813 337603 280847 337909
rect 280997 335223 281031 337841
rect 282561 336855 282595 337637
rect 282745 336991 282779 337977
rect 283021 337807 283055 338045
rect 286977 337943 287011 338113
rect 287897 337875 287931 337977
rect 282837 336787 282871 337365
rect 284585 337127 284619 337297
rect 285413 336855 285447 337637
rect 278789 333727 278823 333965
rect 280111 333625 280353 333659
rect 280295 333557 280445 333591
rect 260665 314687 260699 321861
rect 267473 317475 267507 318801
rect 274373 316047 274407 325601
rect 277317 324343 277351 331245
rect 285597 329103 285631 337025
rect 287437 336923 287471 337569
rect 287529 337195 287563 337773
rect 287989 337263 288023 338113
rect 289863 337909 290105 337943
rect 289955 337773 290013 337807
rect 289587 337705 289737 337739
rect 289863 337705 290231 337739
rect 289955 337569 290105 337603
rect 289863 337501 290013 337535
rect 289955 337433 290105 337467
rect 287529 337161 287897 337195
rect 289829 336719 289863 337365
rect 290197 337331 290231 337705
rect 289829 335971 289863 336481
rect 288357 333795 288391 333965
rect 288633 329579 288667 335665
rect 290105 334747 290139 337297
rect 291485 337059 291519 337365
rect 298845 337331 298879 337841
rect 308999 337365 309091 337399
rect 309057 337331 309091 337365
rect 321569 337331 321603 337365
rect 311851 337297 312001 337331
rect 321511 337297 321603 337331
rect 328469 337195 328503 337297
rect 338129 337059 338163 337161
rect 347697 337059 347731 337297
rect 347789 337195 347823 337297
rect 352113 337195 352147 337297
rect 357449 337195 357483 337297
rect 367017 337195 367051 337297
rect 367109 337195 367143 337297
rect 371433 337195 371467 337297
rect 376769 337195 376803 337297
rect 386337 337195 386371 337297
rect 386429 337195 386463 337297
rect 390753 337195 390787 337297
rect 396089 337195 396123 337297
rect 405657 337195 405691 337297
rect 405749 337195 405783 337297
rect 410073 337195 410107 337297
rect 415409 337195 415443 337297
rect 424977 337195 425011 337297
rect 425069 337195 425103 337297
rect 429393 337195 429427 337297
rect 434729 337195 434763 337297
rect 444297 337195 444331 337297
rect 444389 337195 444423 337297
rect 448713 337195 448747 337297
rect 454049 337195 454083 337297
rect 463617 337195 463651 337297
rect 463709 337195 463743 337297
rect 468033 337195 468067 337297
rect 473369 337195 473403 337297
rect 482937 337195 482971 337365
rect 483581 336719 483615 337365
rect 298109 333727 298143 333965
rect 307677 333863 307711 333965
rect 299523 333625 299673 333659
rect 279893 326519 279927 326757
rect 309183 326553 309425 326587
rect 289863 326485 290013 326519
rect 309275 326485 309333 326519
rect 357357 326451 357391 326757
rect 280169 326043 280203 326145
rect 289737 326043 289771 326417
rect 299397 326315 299431 326417
rect 299489 326247 299523 326417
rect 308965 326247 308999 326417
rect 309149 326315 309183 326417
rect 318717 326315 318751 326417
rect 318809 326247 318843 326417
rect 328377 326247 328411 326417
rect 338129 326247 338163 326417
rect 347605 326247 347639 326417
rect 289185 318835 289219 323561
rect 237205 298163 237239 307717
rect 235365 289799 235399 298061
rect 273637 296735 273671 309077
rect 254869 285719 254903 295273
rect 255789 289119 255823 295273
rect 284585 288439 284619 298061
rect 288357 289119 288391 298061
rect 289093 288439 289127 298061
rect 229569 270555 229603 280109
rect 235181 260899 235215 273921
rect 235549 270555 235583 280109
rect 255789 264979 255823 274601
rect 229569 251243 229603 260797
rect 235181 244035 235215 259369
rect 250729 253827 250763 260797
rect 277041 256751 277075 266305
rect 277225 264979 277259 274601
rect 237113 241519 237147 251141
rect 252201 249815 252235 251277
rect 254869 249815 254903 251209
rect 238953 231863 238987 241417
rect 255789 237439 255823 255221
rect 259929 245667 259963 255221
rect 276949 249747 276983 256649
rect 277225 247027 277259 255221
rect 260573 237439 260607 246993
rect 274189 237439 274223 246993
rect 277225 237439 277259 241485
rect 262505 229075 262539 234685
rect 264253 219487 264287 237337
rect 255881 208403 255915 217957
rect 238953 191879 238987 202793
rect 252201 198747 252235 208301
rect 262689 198747 262723 217957
rect 264253 208403 264287 217957
rect 255789 191335 255823 198645
rect 245025 171139 245059 180761
rect 252109 176715 252143 186269
rect 254777 179435 254811 188989
rect 255789 184195 255823 188989
rect 260665 187731 260699 197149
rect 262689 179435 262723 188989
rect 264253 179435 264287 188989
rect 271613 186371 271647 195925
rect 277133 187731 277167 197285
rect 273821 180795 273855 184229
rect 260665 178075 260699 179401
rect 252201 168351 252235 173961
rect 235181 157403 235215 162741
rect 245025 151827 245059 161381
rect 254869 158763 254903 168317
rect 262689 160123 262723 169677
rect 264253 160123 264287 169677
rect 268853 168419 268887 177973
rect 255881 154547 255915 157369
rect 260573 149107 260607 158661
rect 268853 150467 268887 160021
rect 271613 149175 271647 160021
rect 235273 133943 235307 143497
rect 235549 135303 235583 144857
rect 245209 135167 245243 138669
rect 250545 128299 250579 140709
rect 260573 129795 260607 140709
rect 262689 131155 262723 140709
rect 264253 131155 264287 140709
rect 271613 139519 271647 149005
rect 277133 139451 277167 149005
rect 271521 129795 271555 139349
rect 235273 122859 235307 124185
rect 235549 115991 235583 125545
rect 245117 114563 245151 124117
rect 255053 113203 255087 122757
rect 257261 114563 257295 124117
rect 274097 121499 274131 131053
rect 268853 111911 268887 121397
rect 233801 95251 233835 104805
rect 250637 102187 250671 111741
rect 254869 95251 254903 104805
rect 256525 95251 256559 104805
rect 260481 102119 260515 110381
rect 262689 102255 262723 111741
rect 257261 93891 257295 95217
rect 259929 92531 259963 95217
rect 262689 91103 262723 102085
rect 264253 92531 264287 102085
rect 268853 100759 268887 111741
rect 273913 110483 273947 120037
rect 276949 102187 276983 111741
rect 277225 102255 277259 115957
rect 268853 87091 268887 92429
rect 229569 67643 229603 77197
rect 235273 75939 235307 85493
rect 237021 76007 237055 85493
rect 245209 75939 245243 85493
rect 274097 82875 274131 99297
rect 235549 57987 235583 67541
rect 237205 57987 237239 75837
rect 245117 67643 245151 70465
rect 250729 68323 250763 82773
rect 250913 72471 250947 77197
rect 251005 71723 251039 77129
rect 251097 70431 251131 77197
rect 264253 75803 264287 82773
rect 255789 63563 255823 73049
rect 256433 63563 256467 73117
rect 257169 63563 257203 68357
rect 267473 66283 267507 75837
rect 268945 71791 268979 76585
rect 273913 63563 273947 76585
rect 277133 74579 277167 84133
rect 277133 63563 277167 73049
rect 229569 48331 229603 57885
rect 245209 48331 245243 57885
rect 254961 51119 254995 60605
rect 255789 52479 255823 61965
rect 269589 53635 269623 56525
rect 229569 29019 229603 38573
rect 235181 37315 235215 46869
rect 255881 42823 255915 44217
rect 235549 19363 235583 28917
rect 250453 9707 250487 19261
rect 256617 18003 256651 44081
rect 257169 34527 257203 39321
rect 264253 35955 264287 45509
rect 276857 37315 276891 44965
rect 257261 18003 257295 27557
rect 264253 16643 264287 26197
rect 268853 16643 268887 26197
rect 271613 18003 271647 37213
rect 274281 18003 274315 27557
rect 256525 8347 256559 9673
rect 260665 9163 260699 16541
rect 262597 6987 262631 16541
rect 264253 5695 264287 6817
rect 244289 5219 244323 5389
rect 224141 4607 224175 4981
rect 224233 4811 224267 4981
rect 278053 4743 278087 4913
rect 225061 3451 225095 3553
rect 225245 3519 225279 3825
rect 229753 3723 229787 3825
rect 226165 3621 226383 3655
rect 226165 3587 226199 3621
rect 224969 3349 225153 3383
rect 224969 3315 225003 3349
rect 225061 3247 225095 3281
rect 225061 3213 225245 3247
rect 226257 2975 226291 3553
rect 226349 3043 226383 3621
rect 229845 3587 229879 3689
rect 229661 3383 229695 3485
rect 226349 3009 226441 3043
rect 229109 2771 229143 3349
rect 229753 3043 229787 3281
rect 234169 2771 234203 3553
rect 567761 3383 567795 3553
<< viali >>
rect 219081 695453 219115 695487
rect 219081 685865 219115 685899
rect 154313 685797 154347 685831
rect 154313 676209 154347 676243
rect 299857 684437 299891 684471
rect 218989 676141 219023 676175
rect 218989 666553 219023 666587
rect 299857 666553 299891 666587
rect 219265 656829 219299 656863
rect 219265 647241 219299 647275
rect 219357 626501 219391 626535
rect 219357 616845 219391 616879
rect 219081 611405 219115 611439
rect 219081 608685 219115 608719
rect 219265 608549 219299 608583
rect 299673 608549 299707 608583
rect 299673 601681 299707 601715
rect 219265 601545 219299 601579
rect 219173 598893 219207 598927
rect 219173 589305 219207 589339
rect 299857 598893 299891 598927
rect 299857 589305 299891 589339
rect 154313 589237 154347 589271
rect 154313 579717 154347 579751
rect 218897 579581 218931 579615
rect 218897 569925 218931 569959
rect 218897 553401 218931 553435
rect 218897 550613 218931 550647
rect 154405 531233 154439 531267
rect 154405 521645 154439 521679
rect 154405 511921 154439 511955
rect 219081 510561 219115 510595
rect 219081 505053 219115 505087
rect 154405 502333 154439 502367
rect 299673 492609 299707 492643
rect 299673 485741 299707 485775
rect 299673 473297 299707 473331
rect 299673 466361 299707 466395
rect 154221 453985 154255 454019
rect 154221 444397 154255 444431
rect 218989 453985 219023 454019
rect 218989 444397 219023 444431
rect 299489 449837 299523 449871
rect 299489 440249 299523 440283
rect 299581 436781 299615 436815
rect 154405 434673 154439 434707
rect 154405 427737 154439 427771
rect 299581 427737 299615 427771
rect 154313 415361 154347 415395
rect 154313 405705 154347 405739
rect 299673 415361 299707 415395
rect 299673 405705 299707 405739
rect 261125 402985 261159 403019
rect 260113 402781 260147 402815
rect 260113 402577 260147 402611
rect 262229 402781 262263 402815
rect 261125 402441 261159 402475
rect 261861 402577 261895 402611
rect 262229 402577 262263 402611
rect 248337 402101 248371 402135
rect 261861 402101 261895 402135
rect 262781 402509 262815 402543
rect 262781 402033 262815 402067
rect 244841 401897 244875 401931
rect 248337 401897 248371 401931
rect 245485 401829 245519 401863
rect 248153 401761 248187 401795
rect 248337 401761 248371 401795
rect 248153 401625 248187 401659
rect 248337 401625 248371 401659
rect 242081 399857 242115 399891
rect 235457 399449 235491 399483
rect 234169 399245 234203 399279
rect 234537 399245 234571 399279
rect 235457 399245 235491 399279
rect 234537 399041 234571 399075
rect 234169 398973 234203 399007
rect 282469 399313 282503 399347
rect 288357 399313 288391 399347
rect 288357 399177 288391 399211
rect 288725 399313 288759 399347
rect 282469 399109 282503 399143
rect 288725 398905 288759 398939
rect 242081 398837 242115 398871
rect 277041 338521 277075 338555
rect 237665 338045 237699 338079
rect 237297 337909 237331 337943
rect 237297 337773 237331 337807
rect 268393 338045 268427 338079
rect 268393 337841 268427 337875
rect 273177 337977 273211 338011
rect 275293 337977 275327 338011
rect 273177 337773 273211 337807
rect 273269 337909 273303 337943
rect 237665 337705 237699 337739
rect 265633 337705 265667 337739
rect 235917 337569 235951 337603
rect 262505 337569 262539 337603
rect 235917 337297 235951 337331
rect 261769 337297 261803 337331
rect 240057 337093 240091 337127
rect 235825 336549 235859 336583
rect 235825 336141 235859 336175
rect 251741 335937 251775 335971
rect 229569 335393 229603 335427
rect 240057 335393 240091 335427
rect 248797 335665 248831 335699
rect 229569 328457 229603 328491
rect 233985 334305 234019 334339
rect 251741 334917 251775 334951
rect 254685 335733 254719 335767
rect 248797 332129 248831 332163
rect 250545 333285 250579 333319
rect 250545 328457 250579 328491
rect 255881 335665 255915 335699
rect 254685 328457 254719 328491
rect 254869 333897 254903 333931
rect 233985 327097 234019 327131
rect 237021 328389 237055 328423
rect 245209 328389 245243 328423
rect 245209 320297 245243 320331
rect 237021 318801 237055 318835
rect 229477 318733 229511 318767
rect 245209 318733 245243 318767
rect 229477 310777 229511 310811
rect 235273 317373 235307 317407
rect 229477 309077 229511 309111
rect 255881 328457 255915 328491
rect 262873 337501 262907 337535
rect 262873 336685 262907 336719
rect 265173 337433 265207 337467
rect 262505 336277 262539 336311
rect 272533 337637 272567 337671
rect 268301 337569 268335 337603
rect 265633 336753 265667 336787
rect 267473 337501 267507 337535
rect 266277 336685 266311 336719
rect 265173 335325 265207 335359
rect 265449 335665 265483 335699
rect 261769 328457 261803 328491
rect 265449 327369 265483 327403
rect 266829 336685 266863 336719
rect 266829 334849 266863 334883
rect 268301 337025 268335 337059
rect 267473 332265 267507 332299
rect 269037 336685 269071 336719
rect 266277 327097 266311 327131
rect 275293 337841 275327 337875
rect 275937 337773 275971 337807
rect 273269 337093 273303 337127
rect 274741 337501 274775 337535
rect 275937 337501 275971 337535
rect 272533 335461 272567 335495
rect 273177 336685 273211 336719
rect 271889 332401 271923 332435
rect 271889 332197 271923 332231
rect 269037 327097 269071 327131
rect 273177 327097 273211 327131
rect 274373 336685 274407 336719
rect 274741 336549 274775 336583
rect 277041 335393 277075 335427
rect 277317 338113 277351 338147
rect 286977 338113 287011 338147
rect 282929 338045 282963 338079
rect 282561 337977 282595 338011
rect 280813 337909 280847 337943
rect 277869 337705 277903 337739
rect 277869 337297 277903 337331
rect 280537 337705 280571 337739
rect 277317 335325 277351 335359
rect 280813 337569 280847 337603
rect 280997 337841 281031 337875
rect 280537 335325 280571 335359
rect 282561 337637 282595 337671
rect 287989 338113 288023 338147
rect 286977 337909 287011 337943
rect 287897 337977 287931 338011
rect 287897 337841 287931 337875
rect 283021 337773 283055 337807
rect 287529 337773 287563 337807
rect 285413 337637 285447 337671
rect 282745 336957 282779 336991
rect 282837 337365 282871 337399
rect 282561 336821 282595 336855
rect 284585 337297 284619 337331
rect 284585 337093 284619 337127
rect 287437 337569 287471 337603
rect 285413 336821 285447 336855
rect 285597 337025 285631 337059
rect 282837 336753 282871 336787
rect 280997 335189 281031 335223
rect 278789 333965 278823 333999
rect 278789 333693 278823 333727
rect 280077 333625 280111 333659
rect 280353 333625 280387 333659
rect 280261 333557 280295 333591
rect 280445 333557 280479 333591
rect 274373 327097 274407 327131
rect 277317 331245 277351 331279
rect 274373 325601 274407 325635
rect 254869 316081 254903 316115
rect 260665 321861 260699 321895
rect 267473 318801 267507 318835
rect 267473 317441 267507 317475
rect 289829 337909 289863 337943
rect 290105 337909 290139 337943
rect 298845 337841 298879 337875
rect 289921 337773 289955 337807
rect 290013 337773 290047 337807
rect 289553 337705 289587 337739
rect 289737 337705 289771 337739
rect 289829 337705 289863 337739
rect 289921 337569 289955 337603
rect 290105 337569 290139 337603
rect 289829 337501 289863 337535
rect 290013 337501 290047 337535
rect 289921 337433 289955 337467
rect 290105 337433 290139 337467
rect 287989 337229 288023 337263
rect 289829 337365 289863 337399
rect 287897 337161 287931 337195
rect 287437 336889 287471 336923
rect 289829 336685 289863 336719
rect 290105 337297 290139 337331
rect 290197 337297 290231 337331
rect 291485 337365 291519 337399
rect 289829 336481 289863 336515
rect 289829 335937 289863 335971
rect 288633 335665 288667 335699
rect 288357 333965 288391 333999
rect 288357 333761 288391 333795
rect 308965 337365 308999 337399
rect 298845 337297 298879 337331
rect 321569 337365 321603 337399
rect 482937 337365 482971 337399
rect 309057 337297 309091 337331
rect 311817 337297 311851 337331
rect 312001 337297 312035 337331
rect 321477 337297 321511 337331
rect 328469 337297 328503 337331
rect 347697 337297 347731 337331
rect 328469 337161 328503 337195
rect 338129 337161 338163 337195
rect 291485 337025 291519 337059
rect 338129 337025 338163 337059
rect 347789 337297 347823 337331
rect 347789 337161 347823 337195
rect 352113 337297 352147 337331
rect 352113 337161 352147 337195
rect 357449 337297 357483 337331
rect 357449 337161 357483 337195
rect 367017 337297 367051 337331
rect 367017 337161 367051 337195
rect 367109 337297 367143 337331
rect 367109 337161 367143 337195
rect 371433 337297 371467 337331
rect 371433 337161 371467 337195
rect 376769 337297 376803 337331
rect 376769 337161 376803 337195
rect 386337 337297 386371 337331
rect 386337 337161 386371 337195
rect 386429 337297 386463 337331
rect 386429 337161 386463 337195
rect 390753 337297 390787 337331
rect 390753 337161 390787 337195
rect 396089 337297 396123 337331
rect 396089 337161 396123 337195
rect 405657 337297 405691 337331
rect 405657 337161 405691 337195
rect 405749 337297 405783 337331
rect 405749 337161 405783 337195
rect 410073 337297 410107 337331
rect 410073 337161 410107 337195
rect 415409 337297 415443 337331
rect 415409 337161 415443 337195
rect 424977 337297 425011 337331
rect 424977 337161 425011 337195
rect 425069 337297 425103 337331
rect 425069 337161 425103 337195
rect 429393 337297 429427 337331
rect 429393 337161 429427 337195
rect 434729 337297 434763 337331
rect 434729 337161 434763 337195
rect 444297 337297 444331 337331
rect 444297 337161 444331 337195
rect 444389 337297 444423 337331
rect 444389 337161 444423 337195
rect 448713 337297 448747 337331
rect 448713 337161 448747 337195
rect 454049 337297 454083 337331
rect 454049 337161 454083 337195
rect 463617 337297 463651 337331
rect 463617 337161 463651 337195
rect 463709 337297 463743 337331
rect 463709 337161 463743 337195
rect 468033 337297 468067 337331
rect 468033 337161 468067 337195
rect 473369 337297 473403 337331
rect 473369 337161 473403 337195
rect 482937 337161 482971 337195
rect 483581 337365 483615 337399
rect 347697 337025 347731 337059
rect 483581 336685 483615 336719
rect 290105 334713 290139 334747
rect 298109 333965 298143 333999
rect 307677 333965 307711 333999
rect 307677 333829 307711 333863
rect 298109 333693 298143 333727
rect 299489 333625 299523 333659
rect 299673 333625 299707 333659
rect 288633 329545 288667 329579
rect 285597 329069 285631 329103
rect 279893 326757 279927 326791
rect 357357 326757 357391 326791
rect 309149 326553 309183 326587
rect 309425 326553 309459 326587
rect 279893 326485 279927 326519
rect 289829 326485 289863 326519
rect 290013 326485 290047 326519
rect 309241 326485 309275 326519
rect 309333 326485 309367 326519
rect 289737 326417 289771 326451
rect 280169 326145 280203 326179
rect 280169 326009 280203 326043
rect 299397 326417 299431 326451
rect 299397 326281 299431 326315
rect 299489 326417 299523 326451
rect 299489 326213 299523 326247
rect 308965 326417 308999 326451
rect 309149 326417 309183 326451
rect 309149 326281 309183 326315
rect 318717 326417 318751 326451
rect 318717 326281 318751 326315
rect 318809 326417 318843 326451
rect 308965 326213 308999 326247
rect 318809 326213 318843 326247
rect 328377 326417 328411 326451
rect 328377 326213 328411 326247
rect 338129 326417 338163 326451
rect 338129 326213 338163 326247
rect 347605 326417 347639 326451
rect 357357 326417 357391 326451
rect 347605 326213 347639 326247
rect 289737 326009 289771 326043
rect 277317 324309 277351 324343
rect 289185 323561 289219 323595
rect 289185 318801 289219 318835
rect 274373 316013 274407 316047
rect 260665 314653 260699 314687
rect 245209 311797 245243 311831
rect 273637 309077 273671 309111
rect 235273 301937 235307 301971
rect 237205 307717 237239 307751
rect 229477 299489 229511 299523
rect 237205 298129 237239 298163
rect 235365 298061 235399 298095
rect 273637 296701 273671 296735
rect 284585 298061 284619 298095
rect 235365 289765 235399 289799
rect 254869 295273 254903 295307
rect 255789 295273 255823 295307
rect 255789 289085 255823 289119
rect 288357 298061 288391 298095
rect 288357 289085 288391 289119
rect 289093 298061 289127 298095
rect 284585 288405 284619 288439
rect 289093 288405 289127 288439
rect 254869 285685 254903 285719
rect 229569 280109 229603 280143
rect 235549 280109 235583 280143
rect 229569 270521 229603 270555
rect 235181 273921 235215 273955
rect 235549 270521 235583 270555
rect 255789 274601 255823 274635
rect 277225 274601 277259 274635
rect 255789 264945 255823 264979
rect 277041 266305 277075 266339
rect 235181 260865 235215 260899
rect 229569 260797 229603 260831
rect 250729 260797 250763 260831
rect 229569 251209 229603 251243
rect 235181 259369 235215 259403
rect 277225 264945 277259 264979
rect 277041 256717 277075 256751
rect 276949 256649 276983 256683
rect 250729 253793 250763 253827
rect 255789 255221 255823 255255
rect 252201 251277 252235 251311
rect 235181 244001 235215 244035
rect 237113 251141 237147 251175
rect 252201 249781 252235 249815
rect 254869 251209 254903 251243
rect 254869 249781 254903 249815
rect 237113 241485 237147 241519
rect 238953 241417 238987 241451
rect 259929 255221 259963 255255
rect 276949 249713 276983 249747
rect 277225 255221 277259 255255
rect 259929 245633 259963 245667
rect 260573 246993 260607 247027
rect 255789 237405 255823 237439
rect 260573 237405 260607 237439
rect 274189 246993 274223 247027
rect 277225 246993 277259 247027
rect 274189 237405 274223 237439
rect 277225 241485 277259 241519
rect 277225 237405 277259 237439
rect 264253 237337 264287 237371
rect 238953 231829 238987 231863
rect 262505 234685 262539 234719
rect 262505 229041 262539 229075
rect 264253 219453 264287 219487
rect 255881 217957 255915 217991
rect 255881 208369 255915 208403
rect 262689 217957 262723 217991
rect 252201 208301 252235 208335
rect 238953 202793 238987 202827
rect 252201 198713 252235 198747
rect 264253 217957 264287 217991
rect 264253 208369 264287 208403
rect 262689 198713 262723 198747
rect 238953 191845 238987 191879
rect 255789 198645 255823 198679
rect 277133 197285 277167 197319
rect 255789 191301 255823 191335
rect 260665 197149 260699 197183
rect 254777 188989 254811 189023
rect 252109 186269 252143 186303
rect 245025 180761 245059 180795
rect 255789 188989 255823 189023
rect 271613 195925 271647 195959
rect 260665 187697 260699 187731
rect 262689 188989 262723 189023
rect 255789 184161 255823 184195
rect 254777 179401 254811 179435
rect 260665 179401 260699 179435
rect 262689 179401 262723 179435
rect 264253 188989 264287 189023
rect 277133 187697 277167 187731
rect 271613 186337 271647 186371
rect 273821 184229 273855 184263
rect 273821 180761 273855 180795
rect 264253 179401 264287 179435
rect 260665 178041 260699 178075
rect 252109 176681 252143 176715
rect 268853 177973 268887 178007
rect 245025 171105 245059 171139
rect 252201 173961 252235 173995
rect 262689 169677 262723 169711
rect 252201 168317 252235 168351
rect 254869 168317 254903 168351
rect 235181 162741 235215 162775
rect 235181 157369 235215 157403
rect 245025 161381 245059 161415
rect 262689 160089 262723 160123
rect 264253 169677 264287 169711
rect 268853 168385 268887 168419
rect 264253 160089 264287 160123
rect 254869 158729 254903 158763
rect 268853 160021 268887 160055
rect 260573 158661 260607 158695
rect 255881 157369 255915 157403
rect 255881 154513 255915 154547
rect 245025 151793 245059 151827
rect 268853 150433 268887 150467
rect 271613 160021 271647 160055
rect 271613 149141 271647 149175
rect 260573 149073 260607 149107
rect 271613 149005 271647 149039
rect 235549 144857 235583 144891
rect 235273 143497 235307 143531
rect 250545 140709 250579 140743
rect 235549 135269 235583 135303
rect 245209 138669 245243 138703
rect 245209 135133 245243 135167
rect 235273 133909 235307 133943
rect 260573 140709 260607 140743
rect 262689 140709 262723 140743
rect 262689 131121 262723 131155
rect 264253 140709 264287 140743
rect 271613 139485 271647 139519
rect 277133 149005 277167 149039
rect 277133 139417 277167 139451
rect 264253 131121 264287 131155
rect 271521 139349 271555 139383
rect 260573 129761 260607 129795
rect 271521 129761 271555 129795
rect 274097 131053 274131 131087
rect 250545 128265 250579 128299
rect 235549 125545 235583 125579
rect 235273 124185 235307 124219
rect 235273 122825 235307 122859
rect 235549 115957 235583 115991
rect 245117 124117 245151 124151
rect 257261 124117 257295 124151
rect 245117 114529 245151 114563
rect 255053 122757 255087 122791
rect 274097 121465 274131 121499
rect 257261 114529 257295 114563
rect 268853 121397 268887 121431
rect 255053 113169 255087 113203
rect 268853 111877 268887 111911
rect 273913 120037 273947 120071
rect 250637 111741 250671 111775
rect 233801 104805 233835 104839
rect 262689 111741 262723 111775
rect 260481 110381 260515 110415
rect 250637 102153 250671 102187
rect 254869 104805 254903 104839
rect 233801 95217 233835 95251
rect 254869 95217 254903 95251
rect 256525 104805 256559 104839
rect 262689 102221 262723 102255
rect 268853 111741 268887 111775
rect 260481 102085 260515 102119
rect 262689 102085 262723 102119
rect 256525 95217 256559 95251
rect 257261 95217 257295 95251
rect 257261 93857 257295 93891
rect 259929 95217 259963 95251
rect 259929 92497 259963 92531
rect 264253 102085 264287 102119
rect 277225 115957 277259 115991
rect 273913 110449 273947 110483
rect 276949 111741 276983 111775
rect 277225 102221 277259 102255
rect 276949 102153 276983 102187
rect 268853 100725 268887 100759
rect 264253 92497 264287 92531
rect 274097 99297 274131 99331
rect 262689 91069 262723 91103
rect 268853 92429 268887 92463
rect 268853 87057 268887 87091
rect 235273 85493 235307 85527
rect 229569 77197 229603 77231
rect 237021 85493 237055 85527
rect 237021 75973 237055 76007
rect 245209 85493 245243 85527
rect 235273 75905 235307 75939
rect 274097 82841 274131 82875
rect 277133 84133 277167 84167
rect 245209 75905 245243 75939
rect 250729 82773 250763 82807
rect 229569 67609 229603 67643
rect 237205 75837 237239 75871
rect 235549 67541 235583 67575
rect 235549 57953 235583 57987
rect 245117 70465 245151 70499
rect 264253 82773 264287 82807
rect 250913 77197 250947 77231
rect 251097 77197 251131 77231
rect 250913 72437 250947 72471
rect 251005 77129 251039 77163
rect 251005 71689 251039 71723
rect 268945 76585 268979 76619
rect 264253 75769 264287 75803
rect 267473 75837 267507 75871
rect 256433 73117 256467 73151
rect 251097 70397 251131 70431
rect 255789 73049 255823 73083
rect 250729 68289 250763 68323
rect 245117 67609 245151 67643
rect 255789 63529 255823 63563
rect 256433 63529 256467 63563
rect 257169 68357 257203 68391
rect 268945 71757 268979 71791
rect 273913 76585 273947 76619
rect 267473 66249 267507 66283
rect 257169 63529 257203 63563
rect 277133 74545 277167 74579
rect 273913 63529 273947 63563
rect 277133 73049 277167 73083
rect 277133 63529 277167 63563
rect 255789 61965 255823 61999
rect 237205 57953 237239 57987
rect 254961 60605 254995 60639
rect 229569 57885 229603 57919
rect 229569 48297 229603 48331
rect 245209 57885 245243 57919
rect 269589 56525 269623 56559
rect 269589 53601 269623 53635
rect 255789 52445 255823 52479
rect 254961 51085 254995 51119
rect 245209 48297 245243 48331
rect 235181 46869 235215 46903
rect 229569 38573 229603 38607
rect 264253 45509 264287 45543
rect 255881 44217 255915 44251
rect 255881 42789 255915 42823
rect 256617 44081 256651 44115
rect 235181 37281 235215 37315
rect 229569 28985 229603 29019
rect 235549 28917 235583 28951
rect 235549 19329 235583 19363
rect 250453 19261 250487 19295
rect 257169 39321 257203 39355
rect 276857 44965 276891 44999
rect 276857 37281 276891 37315
rect 264253 35921 264287 35955
rect 271613 37213 271647 37247
rect 257169 34493 257203 34527
rect 256617 17969 256651 18003
rect 257261 27557 257295 27591
rect 257261 17969 257295 18003
rect 264253 26197 264287 26231
rect 264253 16609 264287 16643
rect 268853 26197 268887 26231
rect 271613 17969 271647 18003
rect 274281 27557 274315 27591
rect 274281 17969 274315 18003
rect 268853 16609 268887 16643
rect 260665 16541 260699 16575
rect 250453 9673 250487 9707
rect 256525 9673 256559 9707
rect 260665 9129 260699 9163
rect 262597 16541 262631 16575
rect 256525 8313 256559 8347
rect 262597 6953 262631 6987
rect 264253 6817 264287 6851
rect 264253 5661 264287 5695
rect 244289 5389 244323 5423
rect 244289 5185 244323 5219
rect 224141 4981 224175 5015
rect 224233 4981 224267 5015
rect 224233 4777 224267 4811
rect 278053 4913 278087 4947
rect 278053 4709 278087 4743
rect 224141 4573 224175 4607
rect 225245 3825 225279 3859
rect 225061 3553 225095 3587
rect 229753 3825 229787 3859
rect 229753 3689 229787 3723
rect 229845 3689 229879 3723
rect 226165 3553 226199 3587
rect 226257 3553 226291 3587
rect 225245 3485 225279 3519
rect 225061 3417 225095 3451
rect 225153 3349 225187 3383
rect 224969 3281 225003 3315
rect 225061 3281 225095 3315
rect 225245 3213 225279 3247
rect 229845 3553 229879 3587
rect 234169 3553 234203 3587
rect 229661 3485 229695 3519
rect 229109 3349 229143 3383
rect 229661 3349 229695 3383
rect 226441 3009 226475 3043
rect 226257 2941 226291 2975
rect 229753 3281 229787 3315
rect 229753 3009 229787 3043
rect 229109 2737 229143 2771
rect 567761 3553 567795 3587
rect 567761 3349 567795 3383
rect 234169 2737 234203 2771
<< metal1 >>
rect 257890 700952 257896 701004
rect 257948 700992 257954 701004
rect 397454 700992 397460 701004
rect 257948 700964 397460 700992
rect 257948 700952 257954 700964
rect 397454 700952 397460 700964
rect 397512 700952 397518 701004
rect 259270 700884 259276 700936
rect 259328 700924 259334 700936
rect 413646 700924 413652 700936
rect 259328 700896 413652 700924
rect 259328 700884 259334 700896
rect 413646 700884 413652 700896
rect 413704 700884 413710 700936
rect 257982 700816 257988 700868
rect 258040 700856 258046 700868
rect 429838 700856 429844 700868
rect 258040 700828 429844 700856
rect 258040 700816 258046 700828
rect 429838 700816 429844 700828
rect 429896 700816 429902 700868
rect 72970 700748 72976 700800
rect 73028 700788 73034 700800
rect 265066 700788 265072 700800
rect 73028 700760 265072 700788
rect 73028 700748 73034 700760
rect 265066 700748 265072 700760
rect 265124 700748 265130 700800
rect 256418 700680 256424 700732
rect 256476 700720 256482 700732
rect 462314 700720 462320 700732
rect 256476 700692 462320 700720
rect 256476 700680 256482 700692
rect 462314 700680 462320 700692
rect 462372 700680 462378 700732
rect 256510 700612 256516 700664
rect 256568 700652 256574 700664
rect 478506 700652 478512 700664
rect 256568 700624 478512 700652
rect 256568 700612 256574 700624
rect 478506 700612 478512 700624
rect 478564 700612 478570 700664
rect 256602 700544 256608 700596
rect 256660 700584 256666 700596
rect 494790 700584 494796 700596
rect 256660 700556 494796 700584
rect 256660 700544 256666 700556
rect 494790 700544 494796 700556
rect 494848 700544 494854 700596
rect 8110 700476 8116 700528
rect 8168 700516 8174 700528
rect 266538 700516 266544 700528
rect 8168 700488 266544 700516
rect 8168 700476 8174 700488
rect 266538 700476 266544 700488
rect 266596 700476 266602 700528
rect 255222 700408 255228 700460
rect 255280 700448 255286 700460
rect 527174 700448 527180 700460
rect 255280 700420 527180 700448
rect 255280 700408 255286 700420
rect 527174 700408 527180 700420
rect 527232 700408 527238 700460
rect 40494 700340 40500 700392
rect 40552 700380 40558 700392
rect 41322 700380 41328 700392
rect 40552 700352 41328 700380
rect 40552 700340 40558 700352
rect 41322 700340 41328 700352
rect 41380 700340 41386 700392
rect 255130 700340 255136 700392
rect 255188 700380 255194 700392
rect 543458 700380 543464 700392
rect 255188 700352 543464 700380
rect 255188 700340 255194 700352
rect 543458 700340 543464 700352
rect 543516 700340 543522 700392
rect 253842 700272 253848 700324
rect 253900 700312 253906 700324
rect 559650 700312 559656 700324
rect 253900 700284 559656 700312
rect 253900 700272 253906 700284
rect 559650 700272 559656 700284
rect 559708 700272 559714 700324
rect 137830 700204 137836 700256
rect 137888 700244 137894 700256
rect 263778 700244 263784 700256
rect 137888 700216 263784 700244
rect 137888 700204 137894 700216
rect 263778 700204 263784 700216
rect 263836 700204 263842 700256
rect 259362 700136 259368 700188
rect 259420 700176 259426 700188
rect 364978 700176 364984 700188
rect 259420 700148 364984 700176
rect 259420 700136 259426 700148
rect 364978 700136 364984 700148
rect 365036 700136 365042 700188
rect 260650 700068 260656 700120
rect 260708 700108 260714 700120
rect 348786 700108 348792 700120
rect 260708 700080 348792 700108
rect 260708 700068 260714 700080
rect 348786 700068 348792 700080
rect 348844 700068 348850 700120
rect 259178 700000 259184 700052
rect 259236 700040 259242 700052
rect 332502 700040 332508 700052
rect 259236 700012 332508 700040
rect 259236 700000 259242 700012
rect 332502 700000 332508 700012
rect 332560 700000 332566 700052
rect 202782 699932 202788 699984
rect 202840 699972 202846 699984
rect 262214 699972 262220 699984
rect 202840 699944 262220 699972
rect 202840 699932 202846 699944
rect 262214 699932 262220 699944
rect 262272 699932 262278 699984
rect 262122 699864 262128 699916
rect 262180 699904 262186 699916
rect 283834 699904 283840 699916
rect 262180 699876 283840 699904
rect 262180 699864 262186 699876
rect 283834 699864 283840 699876
rect 283892 699864 283898 699916
rect 24302 699660 24308 699712
rect 24360 699700 24366 699712
rect 24762 699700 24768 699712
rect 24360 699672 24768 699700
rect 24360 699660 24366 699672
rect 24762 699660 24768 699672
rect 24820 699660 24826 699712
rect 89162 699660 89168 699712
rect 89220 699700 89226 699712
rect 89622 699700 89628 699712
rect 89220 699672 89628 699700
rect 89220 699660 89226 699672
rect 89622 699660 89628 699672
rect 89680 699660 89686 699712
rect 105446 699660 105452 699712
rect 105504 699700 105510 699712
rect 106182 699700 106188 699712
rect 105504 699672 106188 699700
rect 105504 699660 105510 699672
rect 106182 699660 106188 699672
rect 106240 699660 106246 699712
rect 170306 699660 170312 699712
rect 170364 699700 170370 699712
rect 171042 699700 171048 699712
rect 170364 699672 171048 699700
rect 170364 699660 170370 699672
rect 171042 699660 171048 699672
rect 171100 699660 171106 699712
rect 235166 699660 235172 699712
rect 235224 699700 235230 699712
rect 235902 699700 235908 699712
rect 235224 699672 235908 699700
rect 235224 699660 235230 699672
rect 235902 699660 235908 699672
rect 235960 699660 235966 699712
rect 260742 699660 260748 699712
rect 260800 699700 260806 699712
rect 267642 699700 267648 699712
rect 260800 699672 267648 699700
rect 260800 699660 260806 699672
rect 267642 699660 267648 699672
rect 267700 699660 267706 699712
rect 253750 696940 253756 696992
rect 253808 696980 253814 696992
rect 580166 696980 580172 696992
rect 253808 696952 580172 696980
rect 253808 696940 253814 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 154114 695512 154120 695564
rect 154172 695552 154178 695564
rect 154206 695552 154212 695564
rect 154172 695524 154212 695552
rect 154172 695512 154178 695524
rect 154206 695512 154212 695524
rect 154264 695512 154270 695564
rect 219069 695487 219127 695493
rect 219069 695453 219081 695487
rect 219115 695484 219127 695487
rect 219158 695484 219164 695496
rect 219115 695456 219164 695484
rect 219115 695453 219127 695456
rect 219069 695447 219127 695453
rect 219158 695444 219164 695456
rect 219216 695444 219222 695496
rect 154206 688576 154212 688628
rect 154264 688616 154270 688628
rect 154390 688616 154396 688628
rect 154264 688588 154396 688616
rect 154264 688576 154270 688588
rect 154390 688576 154396 688588
rect 154448 688576 154454 688628
rect 299658 688576 299664 688628
rect 299716 688616 299722 688628
rect 300118 688616 300124 688628
rect 299716 688588 300124 688616
rect 299716 688576 299722 688588
rect 300118 688576 300124 688588
rect 300176 688576 300182 688628
rect 299492 685936 301268 685964
rect 219066 685896 219072 685908
rect 219027 685868 219072 685896
rect 219066 685856 219072 685868
rect 219124 685856 219130 685908
rect 253658 685856 253664 685908
rect 253716 685896 253722 685908
rect 299492 685896 299520 685936
rect 253716 685868 299520 685896
rect 301240 685896 301268 685936
rect 580166 685896 580172 685908
rect 301240 685868 580172 685896
rect 253716 685856 253722 685868
rect 580166 685856 580172 685868
rect 580224 685856 580230 685908
rect 154301 685831 154359 685837
rect 154301 685797 154313 685831
rect 154347 685828 154359 685831
rect 154390 685828 154396 685840
rect 154347 685800 154396 685828
rect 154347 685797 154359 685800
rect 154301 685791 154359 685797
rect 154390 685788 154396 685800
rect 154448 685788 154454 685840
rect 299566 684428 299572 684480
rect 299624 684468 299630 684480
rect 299845 684471 299903 684477
rect 299845 684468 299857 684471
rect 299624 684440 299857 684468
rect 299624 684428 299630 684440
rect 299845 684437 299857 684440
rect 299891 684437 299903 684471
rect 299845 684431 299903 684437
rect 154298 676240 154304 676252
rect 154259 676212 154304 676240
rect 154298 676200 154304 676212
rect 154356 676200 154362 676252
rect 218974 676172 218980 676184
rect 218935 676144 218980 676172
rect 218974 676132 218980 676144
rect 219032 676132 219038 676184
rect 154298 673480 154304 673532
rect 154356 673520 154362 673532
rect 154482 673520 154488 673532
rect 154356 673492 154488 673520
rect 154356 673480 154362 673492
rect 154482 673480 154488 673492
rect 154540 673480 154546 673532
rect 252462 673480 252468 673532
rect 252520 673520 252526 673532
rect 580166 673520 580172 673532
rect 252520 673492 580172 673520
rect 252520 673480 252526 673492
rect 580166 673480 580172 673492
rect 580224 673480 580230 673532
rect 3510 667904 3516 667956
rect 3568 667944 3574 667956
rect 262858 667944 262864 667956
rect 3568 667916 262864 667944
rect 3568 667904 3574 667916
rect 262858 667904 262864 667916
rect 262916 667904 262922 667956
rect 218977 666587 219035 666593
rect 218977 666553 218989 666587
rect 219023 666584 219035 666587
rect 219066 666584 219072 666596
rect 219023 666556 219072 666584
rect 219023 666553 219035 666556
rect 218977 666547 219035 666553
rect 219066 666544 219072 666556
rect 219124 666544 219130 666596
rect 299845 666587 299903 666593
rect 299845 666553 299857 666587
rect 299891 666584 299903 666587
rect 299934 666584 299940 666596
rect 299891 666556 299940 666584
rect 299891 666553 299903 666556
rect 299845 666547 299903 666553
rect 299934 666544 299940 666556
rect 299992 666544 299998 666596
rect 219158 659608 219164 659660
rect 219216 659648 219222 659660
rect 219342 659648 219348 659660
rect 219216 659620 219348 659648
rect 219216 659608 219222 659620
rect 219342 659608 219348 659620
rect 219400 659608 219406 659660
rect 219253 656863 219311 656869
rect 219253 656829 219265 656863
rect 219299 656860 219311 656863
rect 219342 656860 219348 656872
rect 219299 656832 219348 656860
rect 219299 656829 219311 656832
rect 219253 656823 219311 656829
rect 219342 656820 219348 656832
rect 219400 656820 219406 656872
rect 154298 654100 154304 654152
rect 154356 654140 154362 654152
rect 154482 654140 154488 654152
rect 154356 654112 154488 654140
rect 154356 654100 154362 654112
rect 154482 654100 154488 654112
rect 154540 654100 154546 654152
rect 3050 652740 3056 652792
rect 3108 652780 3114 652792
rect 267826 652780 267832 652792
rect 3108 652752 267832 652780
rect 3108 652740 3114 652752
rect 267826 652740 267832 652752
rect 267884 652740 267890 652792
rect 252370 650020 252376 650072
rect 252428 650060 252434 650072
rect 580166 650060 580172 650072
rect 252428 650032 580172 650060
rect 252428 650020 252434 650032
rect 580166 650020 580172 650032
rect 580224 650020 580230 650072
rect 219250 647272 219256 647284
rect 219211 647244 219256 647272
rect 219250 647232 219256 647244
rect 219308 647232 219314 647284
rect 299658 647232 299664 647284
rect 299716 647272 299722 647284
rect 299750 647272 299756 647284
rect 299716 647244 299756 647272
rect 299716 647232 299722 647244
rect 299750 647232 299756 647244
rect 299808 647232 299814 647284
rect 219250 640404 219256 640416
rect 219084 640376 219256 640404
rect 219084 640280 219112 640376
rect 219250 640364 219256 640376
rect 219308 640364 219314 640416
rect 299658 640364 299664 640416
rect 299716 640404 299722 640416
rect 299750 640404 299756 640416
rect 299716 640376 299756 640404
rect 299716 640364 299722 640376
rect 299750 640364 299756 640376
rect 299808 640364 299814 640416
rect 219066 640228 219072 640280
rect 219124 640228 219130 640280
rect 252278 638936 252284 638988
rect 252336 638976 252342 638988
rect 580166 638976 580172 638988
rect 252336 638948 580172 638976
rect 252336 638936 252342 638948
rect 580166 638936 580172 638948
rect 580224 638936 580230 638988
rect 219066 637508 219072 637560
rect 219124 637548 219130 637560
rect 219158 637548 219164 637560
rect 219124 637520 219164 637548
rect 219124 637508 219130 637520
rect 219158 637508 219164 637520
rect 219216 637508 219222 637560
rect 154298 634788 154304 634840
rect 154356 634828 154362 634840
rect 154482 634828 154488 634840
rect 154356 634800 154488 634828
rect 154356 634788 154362 634800
rect 154482 634788 154488 634800
rect 154540 634788 154546 634840
rect 299566 630640 299572 630692
rect 299624 630680 299630 630692
rect 299750 630680 299756 630692
rect 299624 630652 299756 630680
rect 299624 630640 299630 630652
rect 299750 630640 299756 630652
rect 299808 630640 299814 630692
rect 251082 626560 251088 626612
rect 251140 626600 251146 626612
rect 580166 626600 580172 626612
rect 251140 626572 580172 626600
rect 251140 626560 251146 626572
rect 580166 626560 580172 626572
rect 580224 626560 580230 626612
rect 219342 626532 219348 626544
rect 219303 626504 219348 626532
rect 219342 626492 219348 626504
rect 219400 626492 219406 626544
rect 219342 616876 219348 616888
rect 219303 616848 219348 616876
rect 219342 616836 219348 616848
rect 219400 616836 219406 616888
rect 154298 615476 154304 615528
rect 154356 615516 154362 615528
rect 154482 615516 154488 615528
rect 154356 615488 154488 615516
rect 154356 615476 154362 615488
rect 154482 615476 154488 615488
rect 154540 615476 154546 615528
rect 219069 611439 219127 611445
rect 219069 611405 219081 611439
rect 219115 611436 219127 611439
rect 219342 611436 219348 611448
rect 219115 611408 219348 611436
rect 219115 611405 219127 611408
rect 219069 611399 219127 611405
rect 219342 611396 219348 611408
rect 219400 611396 219406 611448
rect 299566 611328 299572 611380
rect 299624 611368 299630 611380
rect 299750 611368 299756 611380
rect 299624 611340 299756 611368
rect 299624 611328 299630 611340
rect 299750 611328 299756 611340
rect 299808 611328 299814 611380
rect 3602 609968 3608 610020
rect 3660 610008 3666 610020
rect 264238 610008 264244 610020
rect 3660 609980 264244 610008
rect 3660 609968 3666 609980
rect 264238 609968 264244 609980
rect 264296 609968 264302 610020
rect 219066 608716 219072 608728
rect 219027 608688 219072 608716
rect 219066 608676 219072 608688
rect 219124 608676 219130 608728
rect 219066 608540 219072 608592
rect 219124 608580 219130 608592
rect 219253 608583 219311 608589
rect 219253 608580 219265 608583
rect 219124 608552 219265 608580
rect 219124 608540 219130 608552
rect 219253 608549 219265 608552
rect 219299 608549 219311 608583
rect 299658 608580 299664 608592
rect 299619 608552 299664 608580
rect 219253 608543 219311 608549
rect 299658 608540 299664 608552
rect 299716 608540 299722 608592
rect 249702 603100 249708 603152
rect 249760 603140 249766 603152
rect 580166 603140 580172 603152
rect 249760 603112 580172 603140
rect 249760 603100 249766 603112
rect 580166 603100 580172 603112
rect 580224 603100 580230 603152
rect 299661 601715 299719 601721
rect 299661 601681 299673 601715
rect 299707 601712 299719 601715
rect 299842 601712 299848 601724
rect 299707 601684 299848 601712
rect 299707 601681 299719 601684
rect 299661 601675 299719 601681
rect 299842 601672 299848 601684
rect 299900 601672 299906 601724
rect 219250 601576 219256 601588
rect 219211 601548 219256 601576
rect 219250 601536 219256 601548
rect 219308 601536 219314 601588
rect 219161 598927 219219 598933
rect 219161 598893 219173 598927
rect 219207 598924 219219 598927
rect 219250 598924 219256 598936
rect 219207 598896 219256 598924
rect 219207 598893 219219 598896
rect 219161 598887 219219 598893
rect 219250 598884 219256 598896
rect 219308 598884 219314 598936
rect 299842 598924 299848 598936
rect 299803 598896 299848 598924
rect 299842 598884 299848 598896
rect 299900 598884 299906 598936
rect 154298 596164 154304 596216
rect 154356 596204 154362 596216
rect 154482 596204 154488 596216
rect 154356 596176 154488 596204
rect 154356 596164 154362 596176
rect 154482 596164 154488 596176
rect 154540 596164 154546 596216
rect 3326 594804 3332 594856
rect 3384 594844 3390 594856
rect 269298 594844 269304 594856
rect 3384 594816 269304 594844
rect 3384 594804 3390 594816
rect 269298 594804 269304 594816
rect 269356 594804 269362 594856
rect 250990 592016 250996 592068
rect 251048 592056 251054 592068
rect 580166 592056 580172 592068
rect 251048 592028 580172 592056
rect 251048 592016 251054 592028
rect 580166 592016 580172 592028
rect 580224 592016 580230 592068
rect 219158 589336 219164 589348
rect 219119 589308 219164 589336
rect 219158 589296 219164 589308
rect 219216 589296 219222 589348
rect 299845 589339 299903 589345
rect 299845 589305 299857 589339
rect 299891 589336 299903 589339
rect 299934 589336 299940 589348
rect 299891 589308 299940 589336
rect 299891 589305 299903 589308
rect 299845 589299 299903 589305
rect 299934 589296 299940 589308
rect 299992 589296 299998 589348
rect 154298 589268 154304 589280
rect 154259 589240 154304 589268
rect 154298 589228 154304 589240
rect 154356 589228 154362 589280
rect 299934 582468 299940 582480
rect 299860 582440 299940 582468
rect 218974 582360 218980 582412
rect 219032 582400 219038 582412
rect 219158 582400 219164 582412
rect 219032 582372 219164 582400
rect 219032 582360 219038 582372
rect 219158 582360 219164 582372
rect 219216 582360 219222 582412
rect 299860 582344 299888 582440
rect 299934 582428 299940 582440
rect 299992 582428 299998 582480
rect 299842 582292 299848 582344
rect 299900 582292 299906 582344
rect 154298 579748 154304 579760
rect 154259 579720 154304 579748
rect 154298 579708 154304 579720
rect 154356 579708 154362 579760
rect 249610 579640 249616 579692
rect 249668 579680 249674 579692
rect 580166 579680 580172 579692
rect 249668 579652 580172 579680
rect 249668 579640 249674 579652
rect 580166 579640 580172 579652
rect 580224 579640 580230 579692
rect 154206 579572 154212 579624
rect 154264 579612 154270 579624
rect 154390 579612 154396 579624
rect 154264 579584 154396 579612
rect 154264 579572 154270 579584
rect 154390 579572 154396 579584
rect 154448 579572 154454 579624
rect 218885 579615 218943 579621
rect 218885 579581 218897 579615
rect 218931 579612 218943 579615
rect 218974 579612 218980 579624
rect 218931 579584 218980 579612
rect 218931 579581 218943 579584
rect 218885 579575 218943 579581
rect 218974 579572 218980 579584
rect 219032 579572 219038 579624
rect 218882 569956 218888 569968
rect 218843 569928 218888 569956
rect 218882 569916 218888 569928
rect 218940 569916 218946 569968
rect 299566 563116 299572 563168
rect 299624 563116 299630 563168
rect 218882 563048 218888 563100
rect 218940 563048 218946 563100
rect 154206 562912 154212 562964
rect 154264 562952 154270 562964
rect 154390 562952 154396 562964
rect 154264 562924 154396 562952
rect 154264 562912 154270 562924
rect 154390 562912 154396 562924
rect 154448 562912 154454 562964
rect 218900 562952 218928 563048
rect 299584 563032 299612 563116
rect 299566 562980 299572 563032
rect 299624 562980 299630 563032
rect 218974 562952 218980 562964
rect 218900 562924 218980 562952
rect 218974 562912 218980 562924
rect 219032 562912 219038 562964
rect 248322 556180 248328 556232
rect 248380 556220 248386 556232
rect 580166 556220 580172 556232
rect 248380 556192 580172 556220
rect 248380 556180 248386 556192
rect 580166 556180 580172 556192
rect 580224 556180 580230 556232
rect 299566 553500 299572 553512
rect 299492 553472 299572 553500
rect 218882 553432 218888 553444
rect 218843 553404 218888 553432
rect 218882 553392 218888 553404
rect 218940 553392 218946 553444
rect 299492 553376 299520 553472
rect 299566 553460 299572 553472
rect 299624 553460 299630 553512
rect 299474 553324 299480 553376
rect 299532 553324 299538 553376
rect 3326 552032 3332 552084
rect 3384 552072 3390 552084
rect 265618 552072 265624 552084
rect 3384 552044 265624 552072
rect 3384 552032 3390 552044
rect 265618 552032 265624 552044
rect 265676 552032 265682 552084
rect 218882 550644 218888 550656
rect 218843 550616 218888 550644
rect 218882 550604 218888 550616
rect 218940 550604 218946 550656
rect 249518 545096 249524 545148
rect 249576 545136 249582 545148
rect 580166 545136 580172 545148
rect 249576 545108 580172 545136
rect 249576 545096 249582 545108
rect 580166 545096 580172 545108
rect 580224 545096 580230 545148
rect 218882 543736 218888 543788
rect 218940 543736 218946 543788
rect 218900 543640 218928 543736
rect 299290 543668 299296 543720
rect 299348 543708 299354 543720
rect 299474 543708 299480 543720
rect 299348 543680 299480 543708
rect 299348 543668 299354 543680
rect 299474 543668 299480 543680
rect 299532 543668 299538 543720
rect 218974 543640 218980 543652
rect 218900 543612 218980 543640
rect 218974 543600 218980 543612
rect 219032 543600 219038 543652
rect 3234 538228 3240 538280
rect 3292 538268 3298 538280
rect 270770 538268 270776 538280
rect 3292 538240 270776 538268
rect 3292 538228 3298 538240
rect 270770 538228 270776 538240
rect 270828 538228 270834 538280
rect 248230 532720 248236 532772
rect 248288 532760 248294 532772
rect 580166 532760 580172 532772
rect 248288 532732 580172 532760
rect 248288 532720 248294 532732
rect 580166 532720 580172 532732
rect 580224 532720 580230 532772
rect 299566 531292 299572 531344
rect 299624 531332 299630 531344
rect 299750 531332 299756 531344
rect 299624 531304 299756 531332
rect 299624 531292 299630 531304
rect 299750 531292 299756 531304
rect 299808 531292 299814 531344
rect 154390 531264 154396 531276
rect 154351 531236 154396 531264
rect 154390 531224 154396 531236
rect 154448 531224 154454 531276
rect 299750 524424 299756 524476
rect 299808 524424 299814 524476
rect 299768 524396 299796 524424
rect 299842 524396 299848 524408
rect 299768 524368 299848 524396
rect 299842 524356 299848 524368
rect 299900 524356 299906 524408
rect 218974 524288 218980 524340
rect 219032 524328 219038 524340
rect 219158 524328 219164 524340
rect 219032 524300 219164 524328
rect 219032 524288 219038 524300
rect 219158 524288 219164 524300
rect 219216 524288 219222 524340
rect 154393 521679 154451 521685
rect 154393 521645 154405 521679
rect 154439 521676 154451 521679
rect 154482 521676 154488 521688
rect 154439 521648 154488 521676
rect 154439 521645 154451 521648
rect 154393 521639 154451 521645
rect 154482 521636 154488 521648
rect 154540 521636 154546 521688
rect 218790 514632 218796 514684
rect 218848 514672 218854 514684
rect 219066 514672 219072 514684
rect 218848 514644 219072 514672
rect 218848 514632 218854 514644
rect 219066 514632 219072 514644
rect 219124 514632 219130 514684
rect 299658 511980 299664 512032
rect 299716 512020 299722 512032
rect 299934 512020 299940 512032
rect 299716 511992 299940 512020
rect 299716 511980 299722 511992
rect 299934 511980 299940 511992
rect 299992 511980 299998 512032
rect 154390 511952 154396 511964
rect 154351 511924 154396 511952
rect 154390 511912 154396 511924
rect 154448 511912 154454 511964
rect 219066 510592 219072 510604
rect 219027 510564 219072 510592
rect 219066 510552 219072 510564
rect 219124 510552 219130 510604
rect 246942 509260 246948 509312
rect 247000 509300 247006 509312
rect 580166 509300 580172 509312
rect 247000 509272 580172 509300
rect 247000 509260 247006 509272
rect 580166 509260 580172 509272
rect 580224 509260 580230 509312
rect 219066 505084 219072 505096
rect 219027 505056 219072 505084
rect 219066 505044 219072 505056
rect 219124 505044 219130 505096
rect 154393 502367 154451 502373
rect 154393 502333 154405 502367
rect 154439 502364 154451 502367
rect 154482 502364 154488 502376
rect 154439 502336 154488 502364
rect 154439 502333 154451 502336
rect 154393 502327 154451 502333
rect 154482 502324 154488 502336
rect 154540 502324 154546 502376
rect 299750 502324 299756 502376
rect 299808 502364 299814 502376
rect 299934 502364 299940 502376
rect 299808 502336 299940 502364
rect 299808 502324 299814 502336
rect 299934 502324 299940 502336
rect 299992 502324 299998 502376
rect 248138 498176 248144 498228
rect 248196 498216 248202 498228
rect 580166 498216 580172 498228
rect 248196 498188 580172 498216
rect 248196 498176 248202 498188
rect 580166 498176 580172 498188
rect 580224 498176 580230 498228
rect 3326 495456 3332 495508
rect 3384 495496 3390 495508
rect 266998 495496 267004 495508
rect 3384 495468 267004 495496
rect 3384 495456 3390 495468
rect 266998 495456 267004 495468
rect 267056 495456 267062 495508
rect 219066 492668 219072 492720
rect 219124 492708 219130 492720
rect 219158 492708 219164 492720
rect 219124 492680 219164 492708
rect 219124 492668 219130 492680
rect 219158 492668 219164 492680
rect 219216 492668 219222 492720
rect 154206 492600 154212 492652
rect 154264 492640 154270 492652
rect 154390 492640 154396 492652
rect 154264 492612 154396 492640
rect 154264 492600 154270 492612
rect 154390 492600 154396 492612
rect 154448 492600 154454 492652
rect 299658 492640 299664 492652
rect 299619 492612 299664 492640
rect 299658 492600 299664 492612
rect 299716 492600 299722 492652
rect 219158 485800 219164 485852
rect 219216 485800 219222 485852
rect 246850 485800 246856 485852
rect 246908 485840 246914 485852
rect 580166 485840 580172 485852
rect 246908 485812 580172 485840
rect 246908 485800 246914 485812
rect 580166 485800 580172 485812
rect 580224 485800 580230 485852
rect 219176 485704 219204 485800
rect 299658 485772 299664 485784
rect 299619 485744 299664 485772
rect 299658 485732 299664 485744
rect 299716 485732 299722 485784
rect 219250 485704 219256 485716
rect 219176 485676 219256 485704
rect 219250 485664 219256 485676
rect 219308 485664 219314 485716
rect 2958 480224 2964 480276
rect 3016 480264 3022 480276
rect 272518 480264 272524 480276
rect 3016 480236 272524 480264
rect 3016 480224 3022 480236
rect 272518 480224 272524 480236
rect 272576 480224 272582 480276
rect 299566 476076 299572 476128
rect 299624 476116 299630 476128
rect 299750 476116 299756 476128
rect 299624 476088 299756 476116
rect 299624 476076 299630 476088
rect 299750 476076 299756 476088
rect 299808 476076 299814 476128
rect 299658 473328 299664 473340
rect 299619 473300 299664 473328
rect 299658 473288 299664 473300
rect 299716 473288 299722 473340
rect 154298 466420 154304 466472
rect 154356 466460 154362 466472
rect 154482 466460 154488 466472
rect 154356 466432 154488 466460
rect 154356 466420 154362 466432
rect 154482 466420 154488 466432
rect 154540 466420 154546 466472
rect 218974 466420 218980 466472
rect 219032 466420 219038 466472
rect 218992 466324 219020 466420
rect 299658 466392 299664 466404
rect 299619 466364 299664 466392
rect 299658 466352 299664 466364
rect 299716 466352 299722 466404
rect 219342 466324 219348 466336
rect 218992 466296 219348 466324
rect 219342 466284 219348 466296
rect 219400 466284 219406 466336
rect 245562 462340 245568 462392
rect 245620 462380 245626 462392
rect 580166 462380 580172 462392
rect 245620 462352 580172 462380
rect 245620 462340 245626 462352
rect 580166 462340 580172 462352
rect 580224 462340 580230 462392
rect 299382 460844 299388 460896
rect 299440 460884 299446 460896
rect 299750 460884 299756 460896
rect 299440 460856 299756 460884
rect 299440 460844 299446 460856
rect 299750 460844 299756 460856
rect 299808 460844 299814 460896
rect 154209 454019 154267 454025
rect 154209 453985 154221 454019
rect 154255 454016 154267 454019
rect 154298 454016 154304 454028
rect 154255 453988 154304 454016
rect 154255 453985 154267 453988
rect 154209 453979 154267 453985
rect 154298 453976 154304 453988
rect 154356 453976 154362 454028
rect 218977 454019 219035 454025
rect 218977 453985 218989 454019
rect 219023 454016 219035 454019
rect 219066 454016 219072 454028
rect 219023 453988 219072 454016
rect 219023 453985 219035 453988
rect 218977 453979 219035 453985
rect 219066 453976 219072 453988
rect 219124 453976 219130 454028
rect 299400 451336 299888 451364
rect 245470 451256 245476 451308
rect 245528 451296 245534 451308
rect 299400 451296 299428 451336
rect 245528 451268 299428 451296
rect 299860 451296 299888 451336
rect 580166 451296 580172 451308
rect 299860 451268 580172 451296
rect 245528 451256 245534 451268
rect 580166 451256 580172 451268
rect 580224 451256 580230 451308
rect 299474 449868 299480 449880
rect 299435 449840 299480 449868
rect 299474 449828 299480 449840
rect 299532 449828 299538 449880
rect 154206 444428 154212 444440
rect 154167 444400 154212 444428
rect 154206 444388 154212 444400
rect 154264 444388 154270 444440
rect 218974 444428 218980 444440
rect 218935 444400 218980 444428
rect 218974 444388 218980 444400
rect 219032 444388 219038 444440
rect 299477 440283 299535 440289
rect 299477 440249 299489 440283
rect 299523 440280 299535 440283
rect 299566 440280 299572 440292
rect 299523 440252 299572 440280
rect 299523 440249 299535 440252
rect 299477 440243 299535 440249
rect 299566 440240 299572 440252
rect 299624 440240 299630 440292
rect 245378 438880 245384 438932
rect 245436 438920 245442 438932
rect 580166 438920 580172 438932
rect 245436 438892 580172 438920
rect 245436 438880 245442 438892
rect 580166 438880 580172 438892
rect 580224 438880 580230 438932
rect 3326 437452 3332 437504
rect 3384 437492 3390 437504
rect 269758 437492 269764 437504
rect 3384 437464 269764 437492
rect 3384 437452 3390 437464
rect 269758 437452 269764 437464
rect 269816 437452 269822 437504
rect 299566 436812 299572 436824
rect 299527 436784 299572 436812
rect 299566 436772 299572 436784
rect 299624 436772 299630 436824
rect 154390 434704 154396 434716
rect 154351 434676 154396 434704
rect 154390 434664 154396 434676
rect 154448 434664 154454 434716
rect 218974 434664 218980 434716
rect 219032 434704 219038 434716
rect 219066 434704 219072 434716
rect 219032 434676 219072 434704
rect 219032 434664 219038 434676
rect 219066 434664 219072 434676
rect 219124 434664 219130 434716
rect 154390 427768 154396 427780
rect 154351 427740 154396 427768
rect 154390 427728 154396 427740
rect 154448 427728 154454 427780
rect 299566 427768 299572 427780
rect 299527 427740 299572 427768
rect 299566 427728 299572 427740
rect 299624 427728 299630 427780
rect 3326 423648 3332 423700
rect 3384 423688 3390 423700
rect 273898 423688 273904 423700
rect 3384 423660 273904 423688
rect 3384 423648 3390 423660
rect 273898 423648 273904 423660
rect 273956 423648 273962 423700
rect 244182 415420 244188 415472
rect 244240 415460 244246 415472
rect 580166 415460 580172 415472
rect 244240 415432 580172 415460
rect 244240 415420 244246 415432
rect 580166 415420 580172 415432
rect 580224 415420 580230 415472
rect 154298 415392 154304 415404
rect 154259 415364 154304 415392
rect 154298 415352 154304 415364
rect 154356 415352 154362 415404
rect 299661 415395 299719 415401
rect 299661 415361 299673 415395
rect 299707 415392 299719 415395
rect 299750 415392 299756 415404
rect 299707 415364 299756 415392
rect 299707 415361 299719 415364
rect 299661 415355 299719 415361
rect 299750 415352 299756 415364
rect 299808 415352 299814 415404
rect 258442 407736 258448 407788
rect 258500 407776 258506 407788
rect 259270 407776 259276 407788
rect 258500 407748 259276 407776
rect 258500 407736 258506 407748
rect 259270 407736 259276 407748
rect 259328 407736 259334 407788
rect 154301 405739 154359 405745
rect 154301 405705 154313 405739
rect 154347 405736 154359 405739
rect 154390 405736 154396 405748
rect 154347 405708 154396 405736
rect 154347 405705 154359 405708
rect 154301 405699 154359 405705
rect 154390 405696 154396 405708
rect 154448 405696 154454 405748
rect 299658 405736 299664 405748
rect 299619 405708 299664 405736
rect 299658 405696 299664 405708
rect 299716 405696 299722 405748
rect 243814 404336 243820 404388
rect 243872 404376 243878 404388
rect 580166 404376 580172 404388
rect 243872 404348 580172 404376
rect 243872 404336 243878 404348
rect 580166 404336 580172 404348
rect 580224 404336 580230 404388
rect 261113 403019 261171 403025
rect 261113 402985 261125 403019
rect 261159 403016 261171 403019
rect 261159 402988 263456 403016
rect 261159 402985 261171 402988
rect 261113 402979 261171 402985
rect 171042 402908 171048 402960
rect 171100 402948 171106 402960
rect 263318 402948 263324 402960
rect 171100 402920 263324 402948
rect 171100 402908 171106 402920
rect 263318 402908 263324 402920
rect 263376 402908 263382 402960
rect 263428 402948 263456 402988
rect 269206 402948 269212 402960
rect 263428 402920 269212 402948
rect 269206 402908 269212 402920
rect 269264 402908 269270 402960
rect 154390 402840 154396 402892
rect 154448 402880 154454 402892
rect 264330 402880 264336 402892
rect 154448 402852 264336 402880
rect 154448 402840 154454 402852
rect 264330 402840 264336 402852
rect 264388 402840 264394 402892
rect 106182 402772 106188 402824
rect 106240 402812 106246 402824
rect 260101 402815 260159 402821
rect 106240 402784 258396 402812
rect 106240 402772 106246 402784
rect 89622 402704 89628 402756
rect 89680 402744 89686 402756
rect 258368 402744 258396 402784
rect 260101 402781 260113 402815
rect 260147 402812 260159 402815
rect 262217 402815 262275 402821
rect 262217 402812 262229 402815
rect 260147 402784 262229 402812
rect 260147 402781 260159 402784
rect 260101 402775 260159 402781
rect 262217 402781 262229 402784
rect 262263 402781 262275 402815
rect 262217 402775 262275 402781
rect 264238 402772 264244 402824
rect 264296 402812 264302 402824
rect 270678 402812 270684 402824
rect 264296 402784 270684 402812
rect 264296 402772 264302 402784
rect 270678 402772 270684 402784
rect 270736 402772 270742 402824
rect 264882 402744 264888 402756
rect 89680 402716 258304 402744
rect 258368 402716 264888 402744
rect 89680 402704 89686 402716
rect 41322 402636 41328 402688
rect 41380 402676 41386 402688
rect 258276 402676 258304 402716
rect 264882 402704 264888 402716
rect 264940 402704 264946 402756
rect 265618 402704 265624 402756
rect 265676 402744 265682 402756
rect 272242 402744 272248 402756
rect 265676 402716 272248 402744
rect 265676 402704 265682 402716
rect 272242 402704 272248 402716
rect 272300 402704 272306 402756
rect 265894 402676 265900 402688
rect 41380 402648 258212 402676
rect 258276 402648 265900 402676
rect 41380 402636 41386 402648
rect 24762 402568 24768 402620
rect 24820 402608 24826 402620
rect 258074 402608 258080 402620
rect 24820 402580 258080 402608
rect 24820 402568 24826 402580
rect 258074 402568 258080 402580
rect 258132 402568 258138 402620
rect 258184 402608 258212 402648
rect 265894 402636 265900 402648
rect 265952 402636 265958 402688
rect 260101 402611 260159 402617
rect 260101 402608 260113 402611
rect 258184 402580 260113 402608
rect 260101 402577 260113 402580
rect 260147 402577 260159 402611
rect 260101 402571 260159 402577
rect 260190 402568 260196 402620
rect 260248 402608 260254 402620
rect 261849 402611 261907 402617
rect 261849 402608 261861 402611
rect 260248 402580 261861 402608
rect 260248 402568 260254 402580
rect 261849 402577 261861 402580
rect 261895 402577 261907 402611
rect 261849 402571 261907 402577
rect 262217 402611 262275 402617
rect 262217 402577 262229 402611
rect 262263 402608 262275 402611
rect 266446 402608 266452 402620
rect 262263 402580 266452 402608
rect 262263 402577 262275 402580
rect 262217 402571 262275 402577
rect 266446 402568 266452 402580
rect 266504 402568 266510 402620
rect 266998 402568 267004 402620
rect 267056 402608 267062 402620
rect 273806 402608 273812 402620
rect 267056 402580 273812 402608
rect 267056 402568 267062 402580
rect 273806 402568 273812 402580
rect 273864 402568 273870 402620
rect 3418 402500 3424 402552
rect 3476 402540 3482 402552
rect 262769 402543 262827 402549
rect 262769 402540 262781 402543
rect 3476 402512 262781 402540
rect 3476 402500 3482 402512
rect 262769 402509 262781 402512
rect 262815 402509 262827 402543
rect 267550 402540 267556 402552
rect 262769 402503 262827 402509
rect 262876 402512 267556 402540
rect 3510 402432 3516 402484
rect 3568 402472 3574 402484
rect 261113 402475 261171 402481
rect 261113 402472 261125 402475
rect 3568 402444 261125 402472
rect 3568 402432 3574 402444
rect 261113 402441 261125 402444
rect 261159 402441 261171 402475
rect 261113 402435 261171 402441
rect 261202 402432 261208 402484
rect 261260 402472 261266 402484
rect 262876 402472 262904 402512
rect 267550 402500 267556 402512
rect 267608 402500 267614 402552
rect 261260 402444 262904 402472
rect 261260 402432 261266 402444
rect 262950 402432 262956 402484
rect 263008 402472 263014 402484
rect 269114 402472 269120 402484
rect 263008 402444 269120 402472
rect 263008 402432 263014 402444
rect 269114 402432 269120 402444
rect 269172 402432 269178 402484
rect 3694 402364 3700 402416
rect 3752 402404 3758 402416
rect 271230 402404 271236 402416
rect 3752 402376 271236 402404
rect 3752 402364 3758 402376
rect 271230 402364 271236 402376
rect 271288 402364 271294 402416
rect 3878 402296 3884 402348
rect 3936 402336 3942 402348
rect 272794 402336 272800 402348
rect 3936 402308 272800 402336
rect 3936 402296 3942 402308
rect 272794 402296 272800 402308
rect 272852 402296 272858 402348
rect 4062 402228 4068 402280
rect 4120 402268 4126 402280
rect 274358 402268 274364 402280
rect 4120 402240 274364 402268
rect 4120 402228 4126 402240
rect 274358 402228 274364 402240
rect 274416 402228 274422 402280
rect 219342 402160 219348 402212
rect 219400 402200 219406 402212
rect 262766 402200 262772 402212
rect 219400 402172 262772 402200
rect 219400 402160 219406 402172
rect 262766 402160 262772 402172
rect 262824 402160 262830 402212
rect 269758 402160 269764 402212
rect 269816 402200 269822 402212
rect 275370 402200 275376 402212
rect 269816 402172 275376 402200
rect 269816 402160 269822 402172
rect 275370 402160 275376 402172
rect 275428 402160 275434 402212
rect 240686 402092 240692 402144
rect 240744 402132 240750 402144
rect 248325 402135 248383 402141
rect 248325 402132 248337 402135
rect 240744 402104 248337 402132
rect 240744 402092 240750 402104
rect 248325 402101 248337 402104
rect 248371 402101 248383 402135
rect 248325 402095 248383 402101
rect 248598 402092 248604 402144
rect 248656 402132 248662 402144
rect 249518 402132 249524 402144
rect 248656 402104 249524 402132
rect 248656 402092 248662 402104
rect 249518 402092 249524 402104
rect 249576 402092 249582 402144
rect 250162 402092 250168 402144
rect 250220 402132 250226 402144
rect 250990 402132 250996 402144
rect 250220 402104 250996 402132
rect 250220 402092 250226 402104
rect 250990 402092 250996 402104
rect 251048 402092 251054 402144
rect 251174 402092 251180 402144
rect 251232 402132 251238 402144
rect 252370 402132 252376 402144
rect 251232 402104 252376 402132
rect 251232 402092 251238 402104
rect 252370 402092 252376 402104
rect 252428 402092 252434 402144
rect 252738 402092 252744 402144
rect 252796 402132 252802 402144
rect 253750 402132 253756 402144
rect 252796 402104 253756 402132
rect 252796 402092 252802 402104
rect 253750 402092 253756 402104
rect 253808 402092 253814 402144
rect 254394 402092 254400 402144
rect 254452 402132 254458 402144
rect 255222 402132 255228 402144
rect 254452 402104 255228 402132
rect 254452 402092 254458 402104
rect 255222 402092 255228 402104
rect 255280 402092 255286 402144
rect 255406 402092 255412 402144
rect 255464 402132 255470 402144
rect 256602 402132 256608 402144
rect 255464 402104 256608 402132
rect 255464 402092 255470 402104
rect 256602 402092 256608 402104
rect 256660 402092 256666 402144
rect 256970 402092 256976 402144
rect 257028 402132 257034 402144
rect 257982 402132 257988 402144
rect 257028 402104 257988 402132
rect 257028 402092 257034 402104
rect 257982 402092 257988 402104
rect 258040 402092 258046 402144
rect 261754 402132 261760 402144
rect 258460 402104 261760 402132
rect 235902 402024 235908 402076
rect 235960 402064 235966 402076
rect 258460 402064 258488 402104
rect 261754 402092 261760 402104
rect 261812 402092 261818 402144
rect 261849 402135 261907 402141
rect 261849 402101 261861 402135
rect 261895 402132 261907 402135
rect 299658 402132 299664 402144
rect 261895 402104 299664 402132
rect 261895 402101 261907 402104
rect 261849 402095 261907 402101
rect 299658 402092 299664 402104
rect 299716 402092 299722 402144
rect 235960 402036 258488 402064
rect 235960 402024 235966 402036
rect 258534 402024 258540 402076
rect 258592 402064 258598 402076
rect 259362 402064 259368 402076
rect 258592 402036 259368 402064
rect 258592 402024 258598 402036
rect 259362 402024 259368 402036
rect 259420 402024 259426 402076
rect 259638 402024 259644 402076
rect 259696 402064 259702 402076
rect 260650 402064 260656 402076
rect 259696 402036 260656 402064
rect 259696 402024 259702 402036
rect 260650 402024 260656 402036
rect 260708 402024 260714 402076
rect 261202 402024 261208 402076
rect 261260 402064 261266 402076
rect 262122 402064 262128 402076
rect 261260 402036 262128 402064
rect 261260 402024 261266 402036
rect 262122 402024 262128 402036
rect 262180 402024 262186 402076
rect 262769 402067 262827 402073
rect 262769 402033 262781 402067
rect 262815 402064 262827 402067
rect 268010 402064 268016 402076
rect 262815 402036 268016 402064
rect 262815 402033 262827 402036
rect 262769 402027 262827 402033
rect 268010 402024 268016 402036
rect 268068 402024 268074 402076
rect 272518 402024 272524 402076
rect 272576 402064 272582 402076
rect 273254 402064 273260 402076
rect 272576 402036 273260 402064
rect 272576 402024 272582 402036
rect 273254 402024 273260 402036
rect 273312 402024 273318 402076
rect 273898 402024 273904 402076
rect 273956 402064 273962 402076
rect 274910 402064 274916 402076
rect 273956 402036 274916 402064
rect 273956 402024 273962 402036
rect 274910 402024 274916 402036
rect 274968 402024 274974 402076
rect 493318 401996 493324 402008
rect 235920 401968 493324 401996
rect 235920 401940 235948 401968
rect 493318 401956 493324 401968
rect 493376 401956 493382 402008
rect 235902 401888 235908 401940
rect 235960 401888 235966 401940
rect 239122 401888 239128 401940
rect 239180 401928 239186 401940
rect 244829 401931 244887 401937
rect 244829 401928 244841 401931
rect 239180 401900 244841 401928
rect 239180 401888 239186 401900
rect 244829 401897 244841 401900
rect 244875 401897 244887 401931
rect 244829 401891 244887 401897
rect 244918 401888 244924 401940
rect 244976 401928 244982 401940
rect 245562 401928 245568 401940
rect 244976 401900 245568 401928
rect 244976 401888 244982 401900
rect 245562 401888 245568 401900
rect 245620 401888 245626 401940
rect 245672 401900 246988 401928
rect 243262 401820 243268 401872
rect 243320 401860 243326 401872
rect 244182 401860 244188 401872
rect 243320 401832 244188 401860
rect 243320 401820 243326 401832
rect 244182 401820 244188 401832
rect 244240 401820 244246 401872
rect 244366 401820 244372 401872
rect 244424 401860 244430 401872
rect 245378 401860 245384 401872
rect 244424 401832 245384 401860
rect 244424 401820 244430 401832
rect 245378 401820 245384 401832
rect 245436 401820 245442 401872
rect 245473 401863 245531 401869
rect 245473 401829 245485 401863
rect 245519 401860 245531 401863
rect 245672 401860 245700 401900
rect 245519 401832 245700 401860
rect 245519 401829 245531 401832
rect 245473 401823 245531 401829
rect 245930 401820 245936 401872
rect 245988 401860 245994 401872
rect 246850 401860 246856 401872
rect 245988 401832 246856 401860
rect 245988 401820 245994 401832
rect 246850 401820 246856 401832
rect 246908 401820 246914 401872
rect 246960 401860 246988 401900
rect 247034 401888 247040 401940
rect 247092 401928 247098 401940
rect 248138 401928 248144 401940
rect 247092 401900 248144 401928
rect 247092 401888 247098 401900
rect 248138 401888 248144 401900
rect 248196 401888 248202 401940
rect 248325 401931 248383 401937
rect 248325 401897 248337 401931
rect 248371 401928 248383 401931
rect 500218 401928 500224 401940
rect 248371 401900 500224 401928
rect 248371 401897 248383 401900
rect 248325 401891 248383 401897
rect 500218 401888 500224 401900
rect 500276 401888 500282 401940
rect 498838 401860 498844 401872
rect 246960 401832 498844 401860
rect 498838 401820 498844 401832
rect 498896 401820 498902 401872
rect 3970 401752 3976 401804
rect 4028 401792 4034 401804
rect 248141 401795 248199 401801
rect 248141 401792 248153 401795
rect 4028 401764 248153 401792
rect 4028 401752 4034 401764
rect 248141 401761 248153 401764
rect 248187 401761 248199 401795
rect 248141 401755 248199 401761
rect 248325 401795 248383 401801
rect 248325 401761 248337 401795
rect 248371 401792 248383 401795
rect 278590 401792 278596 401804
rect 248371 401764 278596 401792
rect 248371 401761 248383 401764
rect 248325 401755 248383 401761
rect 278590 401752 278596 401764
rect 278648 401752 278654 401804
rect 3786 401684 3792 401736
rect 3844 401724 3850 401736
rect 280154 401724 280160 401736
rect 3844 401696 280160 401724
rect 3844 401684 3850 401696
rect 280154 401684 280160 401696
rect 280212 401684 280218 401736
rect 3602 401616 3608 401668
rect 3660 401656 3666 401668
rect 248141 401659 248199 401665
rect 248141 401656 248153 401659
rect 3660 401628 248153 401656
rect 3660 401616 3666 401628
rect 248141 401625 248153 401628
rect 248187 401625 248199 401659
rect 248141 401619 248199 401625
rect 248325 401659 248383 401665
rect 248325 401625 248337 401659
rect 248371 401656 248383 401659
rect 281718 401656 281724 401668
rect 248371 401628 281724 401656
rect 248371 401625 248383 401628
rect 248325 401619 248383 401625
rect 281718 401616 281724 401628
rect 281776 401616 281782 401668
rect 13078 401276 13084 401328
rect 13136 401316 13142 401328
rect 277486 401316 277492 401328
rect 13136 401288 277492 401316
rect 13136 401276 13142 401288
rect 277486 401276 277492 401288
rect 277544 401276 277550 401328
rect 226978 401208 226984 401260
rect 227036 401248 227042 401260
rect 276474 401248 276480 401260
rect 227036 401220 276480 401248
rect 227036 401208 227042 401220
rect 276474 401208 276480 401220
rect 276532 401208 276538 401260
rect 241238 401140 241244 401192
rect 241296 401180 241302 401192
rect 290458 401180 290464 401192
rect 241296 401152 290464 401180
rect 241296 401140 241302 401152
rect 290458 401140 290464 401152
rect 290516 401140 290522 401192
rect 225782 401072 225788 401124
rect 225840 401112 225846 401124
rect 280706 401112 280712 401124
rect 225840 401084 280712 401112
rect 225840 401072 225846 401084
rect 280706 401072 280712 401084
rect 280764 401072 280770 401124
rect 227070 401004 227076 401056
rect 227128 401044 227134 401056
rect 284846 401044 284852 401056
rect 227128 401016 284852 401044
rect 227128 401004 227134 401016
rect 284846 401004 284852 401016
rect 284904 401004 284910 401056
rect 234890 400936 234896 400988
rect 234948 400976 234954 400988
rect 297450 400976 297456 400988
rect 234948 400948 297456 400976
rect 234948 400936 234954 400948
rect 297450 400936 297456 400948
rect 297508 400936 297514 400988
rect 231762 400868 231768 400920
rect 231820 400908 231826 400920
rect 294598 400908 294604 400920
rect 231820 400880 294604 400908
rect 231820 400868 231826 400880
rect 294598 400868 294604 400880
rect 294656 400868 294662 400920
rect 238018 400800 238024 400852
rect 238076 400840 238082 400852
rect 301590 400840 301596 400852
rect 238076 400812 301596 400840
rect 238076 400800 238082 400812
rect 301590 400800 301596 400812
rect 301648 400800 301654 400852
rect 218698 400732 218704 400784
rect 218756 400772 218762 400784
rect 283834 400772 283840 400784
rect 218756 400744 283840 400772
rect 218756 400732 218762 400744
rect 283834 400732 283840 400744
rect 283892 400732 283898 400784
rect 211798 400664 211804 400716
rect 211856 400704 211862 400716
rect 278038 400704 278044 400716
rect 211856 400676 278044 400704
rect 211856 400664 211862 400676
rect 278038 400664 278044 400676
rect 278096 400664 278102 400716
rect 214558 400596 214564 400648
rect 214616 400636 214622 400648
rect 286962 400636 286968 400648
rect 214616 400608 286968 400636
rect 214616 400596 214622 400608
rect 286962 400596 286968 400608
rect 287020 400596 287026 400648
rect 207658 400528 207664 400580
rect 207716 400568 207722 400580
rect 281166 400568 281172 400580
rect 207716 400540 281172 400568
rect 207716 400528 207722 400540
rect 281166 400528 281172 400540
rect 281224 400528 281230 400580
rect 230658 400460 230664 400512
rect 230716 400500 230722 400512
rect 304258 400500 304264 400512
rect 230716 400472 304264 400500
rect 230716 400460 230722 400472
rect 304258 400460 304264 400472
rect 304316 400460 304322 400512
rect 235442 400392 235448 400444
rect 235500 400432 235506 400444
rect 308398 400432 308404 400444
rect 235500 400404 308404 400432
rect 235500 400392 235506 400404
rect 308398 400392 308404 400404
rect 308456 400392 308462 400444
rect 203518 400324 203524 400376
rect 203576 400364 203582 400376
rect 285950 400364 285956 400376
rect 203576 400336 285956 400364
rect 203576 400324 203582 400336
rect 285950 400324 285956 400336
rect 286008 400324 286014 400376
rect 237558 400256 237564 400308
rect 237616 400296 237622 400308
rect 413278 400296 413284 400308
rect 237616 400268 413284 400296
rect 237616 400256 237622 400268
rect 413278 400256 413284 400268
rect 413336 400256 413342 400308
rect 240134 400188 240140 400240
rect 240192 400228 240198 400240
rect 290550 400228 290556 400240
rect 240192 400200 290556 400228
rect 240192 400188 240198 400200
rect 290550 400188 290556 400200
rect 290608 400188 290614 400240
rect 10962 399916 10968 399968
rect 11020 399956 11026 399968
rect 275646 399956 275652 399968
rect 11020 399928 275652 399956
rect 11020 399916 11026 399928
rect 275646 399916 275652 399928
rect 275704 399916 275710 399968
rect 242066 399888 242072 399900
rect 242027 399860 242072 399888
rect 242066 399848 242072 399860
rect 242124 399848 242130 399900
rect 242894 399848 242900 399900
rect 242952 399888 242958 399900
rect 290642 399888 290648 399900
rect 242952 399860 290648 399888
rect 242952 399848 242958 399860
rect 290642 399848 290648 399860
rect 290700 399848 290706 399900
rect 227162 399780 227168 399832
rect 227220 399820 227226 399832
rect 278774 399820 278780 399832
rect 227220 399792 278780 399820
rect 227220 399780 227226 399792
rect 278774 399780 278780 399792
rect 278832 399780 278838 399832
rect 222930 399712 222936 399764
rect 222988 399752 222994 399764
rect 281902 399752 281908 399764
rect 222988 399724 281908 399752
rect 222988 399712 222994 399724
rect 281902 399712 281908 399724
rect 281960 399712 281966 399764
rect 233602 399644 233608 399696
rect 233660 399684 233666 399696
rect 291930 399684 291936 399696
rect 233660 399656 291936 399684
rect 233660 399644 233666 399656
rect 291930 399644 291936 399656
rect 291988 399644 291994 399696
rect 236730 399576 236736 399628
rect 236788 399616 236794 399628
rect 298830 399616 298836 399628
rect 236788 399588 298836 399616
rect 236788 399576 236794 399588
rect 298830 399576 298836 399588
rect 298888 399576 298894 399628
rect 225598 399508 225604 399560
rect 225656 399548 225662 399560
rect 289262 399548 289268 399560
rect 225656 399520 289268 399548
rect 225656 399508 225662 399520
rect 289262 399508 289268 399520
rect 289320 399508 289326 399560
rect 232498 399440 232504 399492
rect 232556 399480 232562 399492
rect 235445 399483 235503 399489
rect 235445 399480 235457 399483
rect 232556 399452 235457 399480
rect 232556 399440 232562 399452
rect 235445 399449 235457 399452
rect 235491 399449 235503 399483
rect 235445 399443 235503 399449
rect 239858 399440 239864 399492
rect 239916 399480 239922 399492
rect 302970 399480 302976 399492
rect 239916 399452 302976 399480
rect 239916 399440 239922 399452
rect 302970 399440 302976 399452
rect 303028 399440 303034 399492
rect 215938 399372 215944 399424
rect 215996 399412 216002 399424
rect 285030 399412 285036 399424
rect 215996 399384 285036 399412
rect 215996 399372 216002 399384
rect 285030 399372 285036 399384
rect 285088 399372 285094 399424
rect 209038 399304 209044 399356
rect 209096 399344 209102 399356
rect 279326 399344 279332 399356
rect 209096 399316 279332 399344
rect 209096 399304 209102 399316
rect 279326 399304 279332 399316
rect 279384 399304 279390 399356
rect 282454 399344 282460 399356
rect 282415 399316 282460 399344
rect 282454 399304 282460 399316
rect 282512 399304 282518 399356
rect 288342 399344 288348 399356
rect 288303 399316 288348 399344
rect 288342 399304 288348 399316
rect 288400 399304 288406 399356
rect 288710 399344 288716 399356
rect 288671 399316 288716 399344
rect 288710 399304 288716 399316
rect 288768 399304 288774 399356
rect 234154 399276 234160 399288
rect 234115 399248 234160 399276
rect 234154 399236 234160 399248
rect 234212 399236 234218 399288
rect 234522 399276 234528 399288
rect 234483 399248 234528 399276
rect 234522 399236 234528 399248
rect 234580 399236 234586 399288
rect 235445 399279 235503 399285
rect 235445 399245 235457 399279
rect 235491 399276 235503 399279
rect 305638 399276 305644 399288
rect 235491 399248 305644 399276
rect 235491 399245 235503 399248
rect 235445 399239 235503 399245
rect 305638 399236 305644 399248
rect 305696 399236 305702 399288
rect 213178 399168 213184 399220
rect 213236 399208 213242 399220
rect 288345 399211 288403 399217
rect 288345 399208 288357 399211
rect 213236 399180 288357 399208
rect 213236 399168 213242 399180
rect 288345 399177 288357 399180
rect 288391 399177 288403 399211
rect 288345 399171 288403 399177
rect 204898 399100 204904 399152
rect 204956 399140 204962 399152
rect 282457 399143 282515 399149
rect 282457 399140 282469 399143
rect 204956 399112 282469 399140
rect 204956 399100 204962 399112
rect 282457 399109 282469 399112
rect 282503 399109 282515 399143
rect 282457 399103 282515 399109
rect 234525 399075 234583 399081
rect 234525 399041 234537 399075
rect 234571 399072 234583 399075
rect 312538 399072 312544 399084
rect 234571 399044 312544 399072
rect 234571 399041 234583 399044
rect 234525 399035 234583 399041
rect 312538 399032 312544 399044
rect 312596 399032 312602 399084
rect 234157 399007 234215 399013
rect 234157 398973 234169 399007
rect 234203 399004 234215 399007
rect 319438 399004 319444 399016
rect 234203 398976 319444 399004
rect 234203 398973 234215 398976
rect 234157 398967 234215 398973
rect 319438 398964 319444 398976
rect 319496 398964 319502 399016
rect 135898 398896 135904 398948
rect 135956 398936 135962 398948
rect 288713 398939 288771 398945
rect 288713 398936 288725 398939
rect 135956 398908 288725 398936
rect 135956 398896 135962 398908
rect 288713 398905 288725 398908
rect 288759 398905 288771 398939
rect 288713 398899 288771 398905
rect 242069 398871 242127 398877
rect 242069 398837 242081 398871
rect 242115 398868 242127 398871
rect 291838 398868 291844 398880
rect 242115 398840 291844 398868
rect 242115 398837 242127 398840
rect 242069 398831 242127 398837
rect 291838 398828 291844 398840
rect 291896 398828 291902 398880
rect 3142 395972 3148 396024
rect 3200 396012 3206 396024
rect 10962 396012 10968 396024
rect 3200 395984 10968 396012
rect 3200 395972 3206 395984
rect 10962 395972 10968 395984
rect 11020 395972 11026 396024
rect 290642 393252 290648 393304
rect 290700 393292 290706 393304
rect 579798 393292 579804 393304
rect 290700 393264 579804 393292
rect 290700 393252 290706 393264
rect 579798 393252 579804 393264
rect 579856 393252 579862 393304
rect 3418 380808 3424 380860
rect 3476 380848 3482 380860
rect 225690 380848 225696 380860
rect 3476 380820 225696 380848
rect 3476 380808 3482 380820
rect 225690 380808 225696 380820
rect 225748 380808 225754 380860
rect 291838 369792 291844 369844
rect 291896 369832 291902 369844
rect 580166 369832 580172 369844
rect 291896 369804 580172 369832
rect 291896 369792 291902 369804
rect 580166 369792 580172 369804
rect 580224 369792 580230 369844
rect 2958 367004 2964 367056
rect 3016 367044 3022 367056
rect 226978 367044 226984 367056
rect 3016 367016 226984 367044
rect 3016 367004 3022 367016
rect 226978 367004 226984 367016
rect 227036 367004 227042 367056
rect 326338 358708 326344 358760
rect 326396 358748 326402 358760
rect 580074 358748 580080 358760
rect 326396 358720 580080 358748
rect 326396 358708 326402 358720
rect 580074 358708 580080 358720
rect 580132 358708 580138 358760
rect 290458 346332 290464 346384
rect 290516 346372 290522 346384
rect 579798 346372 579804 346384
rect 290516 346344 579804 346372
rect 290516 346332 290522 346344
rect 579798 346332 579804 346344
rect 579856 346332 579862 346384
rect 277026 338552 277032 338564
rect 276987 338524 277032 338552
rect 277026 338512 277032 338524
rect 277084 338512 277090 338564
rect 263594 338376 263600 338428
rect 263652 338416 263658 338428
rect 265894 338416 265900 338428
rect 263652 338388 265900 338416
rect 263652 338376 263658 338388
rect 265894 338376 265900 338388
rect 265952 338376 265958 338428
rect 247402 338172 247408 338224
rect 247460 338212 247466 338224
rect 247678 338212 247684 338224
rect 247460 338184 247684 338212
rect 247460 338172 247466 338184
rect 247678 338172 247684 338184
rect 247736 338172 247742 338224
rect 282196 338184 283052 338212
rect 253014 338104 253020 338156
rect 253072 338144 253078 338156
rect 253198 338144 253204 338156
rect 253072 338116 253204 338144
rect 253072 338104 253078 338116
rect 253198 338104 253204 338116
rect 253256 338104 253262 338156
rect 270862 338104 270868 338156
rect 270920 338144 270926 338156
rect 277305 338147 277363 338153
rect 277305 338144 277317 338147
rect 270920 338116 277317 338144
rect 270920 338104 270926 338116
rect 277305 338113 277317 338116
rect 277351 338113 277363 338147
rect 277305 338107 277363 338113
rect 3418 338036 3424 338088
rect 3476 338076 3482 338088
rect 13078 338076 13084 338088
rect 3476 338048 13084 338076
rect 3476 338036 3482 338048
rect 13078 338036 13084 338048
rect 13136 338036 13142 338088
rect 125502 338036 125508 338088
rect 125560 338076 125566 338088
rect 237653 338079 237711 338085
rect 237653 338076 237665 338079
rect 125560 338048 237665 338076
rect 125560 338036 125566 338048
rect 237653 338045 237665 338048
rect 237699 338045 237711 338079
rect 240962 338076 240968 338088
rect 237653 338039 237711 338045
rect 237760 338048 240968 338076
rect 107562 337968 107568 338020
rect 107620 338008 107626 338020
rect 237760 338008 237788 338048
rect 240962 338036 240968 338048
rect 241020 338036 241026 338088
rect 247678 338036 247684 338088
rect 247736 338076 247742 338088
rect 255038 338076 255044 338088
rect 247736 338048 255044 338076
rect 247736 338036 247742 338048
rect 255038 338036 255044 338048
rect 255096 338036 255102 338088
rect 261294 338036 261300 338088
rect 261352 338076 261358 338088
rect 268381 338079 268439 338085
rect 268381 338076 268393 338079
rect 261352 338048 268393 338076
rect 261352 338036 261358 338048
rect 268381 338045 268393 338048
rect 268427 338045 268439 338079
rect 268381 338039 268439 338045
rect 271966 338036 271972 338088
rect 272024 338076 272030 338088
rect 272024 338048 273208 338076
rect 272024 338036 272030 338048
rect 107620 337980 237788 338008
rect 107620 337968 107626 337980
rect 240226 337968 240232 338020
rect 240284 337968 240290 338020
rect 262766 337968 262772 338020
rect 262824 338008 262830 338020
rect 273180 338017 273208 338048
rect 279694 338036 279700 338088
rect 279752 338076 279758 338088
rect 282196 338076 282224 338184
rect 279752 338048 282224 338076
rect 279752 338036 279758 338048
rect 282270 338036 282276 338088
rect 282328 338076 282334 338088
rect 282917 338079 282975 338085
rect 282917 338076 282929 338079
rect 282328 338048 282929 338076
rect 282328 338036 282334 338048
rect 282917 338045 282929 338048
rect 282963 338045 282975 338079
rect 283024 338076 283052 338184
rect 286965 338147 287023 338153
rect 286965 338113 286977 338147
rect 287011 338144 287023 338147
rect 287977 338147 288035 338153
rect 287977 338144 287989 338147
rect 287011 338116 287989 338144
rect 287011 338113 287023 338116
rect 286965 338107 287023 338113
rect 287977 338113 287989 338116
rect 288023 338113 288035 338147
rect 287977 338107 288035 338113
rect 291194 338076 291200 338088
rect 283024 338048 291200 338076
rect 282917 338039 282975 338045
rect 291194 338036 291200 338048
rect 291252 338036 291258 338088
rect 273165 338011 273223 338017
rect 262824 337980 273024 338008
rect 262824 337968 262830 337980
rect 115842 337900 115848 337952
rect 115900 337940 115906 337952
rect 237285 337943 237343 337949
rect 237285 337940 237297 337943
rect 115900 337912 237297 337940
rect 115900 337900 115906 337912
rect 237285 337909 237297 337912
rect 237331 337909 237343 337943
rect 240244 337940 240272 337968
rect 237285 337903 237343 337909
rect 237392 337912 240272 337940
rect 100662 337832 100668 337884
rect 100720 337872 100726 337884
rect 237392 337872 237420 337912
rect 253198 337900 253204 337952
rect 253256 337940 253262 337952
rect 254210 337940 254216 337952
rect 253256 337912 254216 337940
rect 253256 337900 253262 337912
rect 254210 337900 254216 337912
rect 254268 337900 254274 337952
rect 263962 337900 263968 337952
rect 264020 337940 264026 337952
rect 268102 337940 268108 337952
rect 264020 337912 268108 337940
rect 264020 337900 264026 337912
rect 268102 337900 268108 337912
rect 268160 337900 268166 337952
rect 100720 337844 237420 337872
rect 100720 337832 100726 337844
rect 240226 337832 240232 337884
rect 240284 337872 240290 337884
rect 246574 337872 246580 337884
rect 240284 337844 246580 337872
rect 240284 337832 240290 337844
rect 246574 337832 246580 337844
rect 246632 337832 246638 337884
rect 268381 337875 268439 337881
rect 268381 337841 268393 337875
rect 268427 337872 268439 337875
rect 272996 337872 273024 337980
rect 273165 337977 273177 338011
rect 273211 337977 273223 338011
rect 273165 337971 273223 337977
rect 275281 338011 275339 338017
rect 275281 337977 275293 338011
rect 275327 338008 275339 338011
rect 280706 338008 280712 338020
rect 275327 337980 280712 338008
rect 275327 337977 275339 337980
rect 275281 337971 275339 337977
rect 280706 337968 280712 337980
rect 280764 337968 280770 338020
rect 281166 337968 281172 338020
rect 281224 338008 281230 338020
rect 282549 338011 282607 338017
rect 282549 338008 282561 338011
rect 281224 337980 282561 338008
rect 281224 337968 281230 337980
rect 282549 337977 282561 337980
rect 282595 337977 282607 338011
rect 282549 337971 282607 337977
rect 287054 337968 287060 338020
rect 287112 338008 287118 338020
rect 287885 338011 287943 338017
rect 287112 337980 287836 338008
rect 287112 337968 287118 337980
rect 273257 337943 273315 337949
rect 273257 337909 273269 337943
rect 273303 337940 273315 337943
rect 280801 337943 280859 337949
rect 280801 337940 280813 337943
rect 273303 337912 280813 337940
rect 273303 337909 273315 337912
rect 273257 337903 273315 337909
rect 280801 337909 280813 337912
rect 280847 337909 280859 337943
rect 280801 337903 280859 337909
rect 283006 337900 283012 337952
rect 283064 337940 283070 337952
rect 286965 337943 287023 337949
rect 286965 337940 286977 337943
rect 283064 337912 286977 337940
rect 283064 337900 283070 337912
rect 286965 337909 286977 337912
rect 287011 337909 287023 337943
rect 287808 337940 287836 337980
rect 287885 337977 287897 338011
rect 287931 338008 287943 338011
rect 297358 338008 297364 338020
rect 287931 337980 297364 338008
rect 287931 337977 287943 337980
rect 287885 337971 287943 337977
rect 297358 337968 297364 337980
rect 297416 337968 297422 338020
rect 289817 337943 289875 337949
rect 289817 337940 289829 337943
rect 287808 337912 289829 337940
rect 286965 337903 287023 337909
rect 289817 337909 289829 337912
rect 289863 337909 289875 337943
rect 289817 337903 289875 337909
rect 290093 337943 290151 337949
rect 290093 337909 290105 337943
rect 290139 337940 290151 337943
rect 290826 337940 290832 337952
rect 290139 337912 290832 337940
rect 290139 337909 290151 337912
rect 290093 337903 290151 337909
rect 290826 337900 290832 337912
rect 290884 337900 290890 337952
rect 275281 337875 275339 337881
rect 275281 337872 275293 337875
rect 268427 337844 272748 337872
rect 272996 337844 275293 337872
rect 268427 337841 268439 337844
rect 268381 337835 268439 337841
rect 35158 337764 35164 337816
rect 35216 337804 35222 337816
rect 232866 337804 232872 337816
rect 35216 337776 232872 337804
rect 35216 337764 35222 337776
rect 232866 337764 232872 337776
rect 232924 337764 232930 337816
rect 237285 337807 237343 337813
rect 237285 337773 237297 337807
rect 237331 337804 237343 337807
rect 241698 337804 241704 337816
rect 237331 337776 241704 337804
rect 237331 337773 237343 337776
rect 237285 337767 237343 337773
rect 241698 337764 241704 337776
rect 241756 337764 241762 337816
rect 264146 337764 264152 337816
rect 264204 337804 264210 337816
rect 264204 337776 272656 337804
rect 264204 337764 264210 337776
rect 39298 337696 39304 337748
rect 39356 337736 39362 337748
rect 233602 337736 233608 337748
rect 39356 337708 233608 337736
rect 39356 337696 39362 337708
rect 233602 337696 233608 337708
rect 233660 337696 233666 337748
rect 237653 337739 237711 337745
rect 237653 337705 237665 337739
rect 237699 337736 237711 337739
rect 242802 337736 242808 337748
rect 237699 337708 242808 337736
rect 237699 337705 237711 337708
rect 237653 337699 237711 337705
rect 242802 337696 242808 337708
rect 242860 337696 242866 337748
rect 265250 337696 265256 337748
rect 265308 337736 265314 337748
rect 265621 337739 265679 337745
rect 265621 337736 265633 337739
rect 265308 337708 265633 337736
rect 265308 337696 265314 337708
rect 265621 337705 265633 337708
rect 265667 337705 265679 337739
rect 265621 337699 265679 337705
rect 32398 337628 32404 337680
rect 32456 337668 32462 337680
rect 231946 337668 231952 337680
rect 32456 337640 231952 337668
rect 32456 337628 32462 337640
rect 231946 337628 231952 337640
rect 232004 337628 232010 337680
rect 258258 337628 258264 337680
rect 258316 337668 258322 337680
rect 272521 337671 272579 337677
rect 272521 337668 272533 337671
rect 258316 337640 272533 337668
rect 258316 337628 258322 337640
rect 272521 337637 272533 337640
rect 272567 337637 272579 337671
rect 272628 337668 272656 337776
rect 272720 337736 272748 337844
rect 275281 337841 275293 337844
rect 275327 337841 275339 337875
rect 275281 337835 275339 337841
rect 277486 337832 277492 337884
rect 277544 337872 277550 337884
rect 280985 337875 281043 337881
rect 280985 337872 280997 337875
rect 277544 337844 280997 337872
rect 277544 337832 277550 337844
rect 280985 337841 280997 337844
rect 281031 337841 281043 337875
rect 280985 337835 281043 337841
rect 284110 337832 284116 337884
rect 284168 337872 284174 337884
rect 287885 337875 287943 337881
rect 287885 337872 287897 337875
rect 284168 337844 287897 337872
rect 284168 337832 284174 337844
rect 287885 337841 287897 337844
rect 287931 337841 287943 337875
rect 287885 337835 287943 337841
rect 288066 337832 288072 337884
rect 288124 337872 288130 337884
rect 298738 337872 298744 337884
rect 288124 337844 298744 337872
rect 288124 337832 288130 337844
rect 298738 337832 298744 337844
rect 298796 337832 298802 337884
rect 298833 337875 298891 337881
rect 298833 337841 298845 337875
rect 298879 337872 298891 337875
rect 302878 337872 302884 337884
rect 298879 337844 302884 337872
rect 298879 337841 298891 337844
rect 298833 337835 298891 337841
rect 302878 337832 302884 337844
rect 302936 337832 302942 337884
rect 273165 337807 273223 337813
rect 273165 337773 273177 337807
rect 273211 337804 273223 337807
rect 275925 337807 275983 337813
rect 275925 337804 275937 337807
rect 273211 337776 275937 337804
rect 273211 337773 273223 337776
rect 273165 337767 273223 337773
rect 275925 337773 275937 337776
rect 275971 337773 275983 337807
rect 275925 337767 275983 337773
rect 276014 337764 276020 337816
rect 276072 337804 276078 337816
rect 276072 337776 280016 337804
rect 276072 337764 276078 337776
rect 277857 337739 277915 337745
rect 277857 337736 277869 337739
rect 272720 337708 277869 337736
rect 277857 337705 277869 337708
rect 277903 337705 277915 337739
rect 279988 337736 280016 337776
rect 280062 337764 280068 337816
rect 280120 337804 280126 337816
rect 283009 337807 283067 337813
rect 280120 337776 282776 337804
rect 280120 337764 280126 337776
rect 280525 337739 280583 337745
rect 280525 337736 280537 337739
rect 279988 337708 280537 337736
rect 277857 337699 277915 337705
rect 280525 337705 280537 337708
rect 280571 337705 280583 337739
rect 280525 337699 280583 337705
rect 282549 337671 282607 337677
rect 282549 337668 282561 337671
rect 272628 337640 282561 337668
rect 272521 337631 272579 337637
rect 282549 337637 282561 337640
rect 282595 337637 282607 337671
rect 282549 337631 282607 337637
rect 28258 337560 28264 337612
rect 28316 337600 28322 337612
rect 232038 337600 232044 337612
rect 28316 337572 232044 337600
rect 28316 337560 28322 337572
rect 232038 337560 232044 337572
rect 232096 337560 232102 337612
rect 233602 337560 233608 337612
rect 233660 337600 233666 337612
rect 234890 337600 234896 337612
rect 233660 337572 234896 337600
rect 233660 337560 233666 337572
rect 234890 337560 234896 337572
rect 234948 337560 234954 337612
rect 235905 337603 235963 337609
rect 235905 337569 235917 337603
rect 235951 337600 235963 337603
rect 246942 337600 246948 337612
rect 235951 337572 246948 337600
rect 235951 337569 235963 337572
rect 235905 337563 235963 337569
rect 246942 337560 246948 337572
rect 247000 337560 247006 337612
rect 257154 337560 257160 337612
rect 257212 337600 257218 337612
rect 262493 337603 262551 337609
rect 262493 337600 262505 337603
rect 257212 337572 262505 337600
rect 257212 337560 257218 337572
rect 262493 337569 262505 337572
rect 262539 337569 262551 337603
rect 268289 337603 268347 337609
rect 262493 337563 262551 337569
rect 265544 337572 267596 337600
rect 14458 337492 14464 337544
rect 14516 337532 14522 337544
rect 230934 337532 230940 337544
rect 14516 337504 230940 337532
rect 14516 337492 14522 337504
rect 230934 337492 230940 337504
rect 230992 337492 230998 337544
rect 240318 337492 240324 337544
rect 240376 337532 240382 337544
rect 242986 337532 242992 337544
rect 240376 337504 242992 337532
rect 240376 337492 240382 337504
rect 242986 337492 242992 337504
rect 243044 337492 243050 337544
rect 257522 337492 257528 337544
rect 257580 337532 257586 337544
rect 262861 337535 262919 337541
rect 262861 337532 262873 337535
rect 257580 337504 262873 337532
rect 257580 337492 257586 337504
rect 262861 337501 262873 337504
rect 262907 337501 262919 337535
rect 262861 337495 262919 337501
rect 15838 337424 15844 337476
rect 15896 337464 15902 337476
rect 231026 337464 231032 337476
rect 15896 337436 231032 337464
rect 15896 337424 15902 337436
rect 231026 337424 231032 337436
rect 231084 337424 231090 337476
rect 231854 337424 231860 337476
rect 231912 337464 231918 337476
rect 235258 337464 235264 337476
rect 231912 337436 235264 337464
rect 231912 337424 231918 337436
rect 235258 337424 235264 337436
rect 235316 337424 235322 337476
rect 242894 337424 242900 337476
rect 242952 337464 242958 337476
rect 251358 337464 251364 337476
rect 242952 337436 251364 337464
rect 242952 337424 242958 337436
rect 251358 337424 251364 337436
rect 251416 337424 251422 337476
rect 257246 337424 257252 337476
rect 257304 337464 257310 337476
rect 265161 337467 265219 337473
rect 265161 337464 265173 337467
rect 257304 337436 265173 337464
rect 257304 337424 257310 337436
rect 265161 337433 265173 337436
rect 265207 337433 265219 337467
rect 265161 337427 265219 337433
rect 10318 337356 10324 337408
rect 10376 337396 10382 337408
rect 230474 337396 230480 337408
rect 10376 337368 230480 337396
rect 10376 337356 10382 337368
rect 230474 337356 230480 337368
rect 230532 337356 230538 337408
rect 231946 337356 231952 337408
rect 232004 337396 232010 337408
rect 253014 337396 253020 337408
rect 232004 337368 253020 337396
rect 232004 337356 232010 337368
rect 253014 337356 253020 337368
rect 253072 337356 253078 337408
rect 260558 337356 260564 337408
rect 260616 337396 260622 337408
rect 265544 337396 265572 337572
rect 266354 337492 266360 337544
rect 266412 337532 266418 337544
rect 266630 337532 266636 337544
rect 266412 337504 266636 337532
rect 266412 337492 266418 337504
rect 266630 337492 266636 337504
rect 266688 337492 266694 337544
rect 266722 337492 266728 337544
rect 266780 337532 266786 337544
rect 267461 337535 267519 337541
rect 267461 337532 267473 337535
rect 266780 337504 267473 337532
rect 266780 337492 266786 337504
rect 267461 337501 267473 337504
rect 267507 337501 267519 337535
rect 267568 337532 267596 337572
rect 268289 337569 268301 337603
rect 268335 337600 268347 337603
rect 280338 337600 280344 337612
rect 268335 337572 280344 337600
rect 268335 337569 268347 337572
rect 268289 337563 268347 337569
rect 280338 337560 280344 337572
rect 280396 337560 280402 337612
rect 280798 337600 280804 337612
rect 280759 337572 280804 337600
rect 280798 337560 280804 337572
rect 280856 337560 280862 337612
rect 282748 337600 282776 337776
rect 283009 337773 283021 337807
rect 283055 337804 283067 337807
rect 287517 337807 287575 337813
rect 287517 337804 287529 337807
rect 283055 337776 287529 337804
rect 283055 337773 283067 337776
rect 283009 337767 283067 337773
rect 287517 337773 287529 337776
rect 287563 337773 287575 337807
rect 287517 337767 287575 337773
rect 287698 337764 287704 337816
rect 287756 337804 287762 337816
rect 289909 337807 289967 337813
rect 289909 337804 289921 337807
rect 287756 337776 289921 337804
rect 287756 337764 287762 337776
rect 289909 337773 289921 337776
rect 289955 337773 289967 337807
rect 289909 337767 289967 337773
rect 290001 337807 290059 337813
rect 290001 337773 290013 337807
rect 290047 337804 290059 337807
rect 301498 337804 301504 337816
rect 290047 337776 301504 337804
rect 290047 337773 290059 337776
rect 290001 337767 290059 337773
rect 301498 337764 301504 337776
rect 301556 337764 301562 337816
rect 289538 337696 289544 337748
rect 289596 337736 289602 337748
rect 289725 337739 289783 337745
rect 289596 337708 289641 337736
rect 289596 337696 289602 337708
rect 289725 337705 289737 337739
rect 289771 337736 289783 337739
rect 289817 337739 289875 337745
rect 289817 337736 289829 337739
rect 289771 337708 289829 337736
rect 289771 337705 289783 337708
rect 289725 337699 289783 337705
rect 289817 337705 289829 337708
rect 289863 337705 289875 337739
rect 289817 337699 289875 337705
rect 284478 337628 284484 337680
rect 284536 337668 284542 337680
rect 285401 337671 285459 337677
rect 285401 337668 285413 337671
rect 284536 337640 285413 337668
rect 284536 337628 284542 337640
rect 285401 337637 285413 337640
rect 285447 337637 285459 337671
rect 285401 337631 285459 337637
rect 287790 337628 287796 337680
rect 287848 337668 287854 337680
rect 320818 337668 320824 337680
rect 287848 337640 320824 337668
rect 287848 337628 287854 337640
rect 320818 337628 320824 337640
rect 320876 337628 320882 337680
rect 282748 337572 284340 337600
rect 274729 337535 274787 337541
rect 274729 337532 274741 337535
rect 267568 337504 274741 337532
rect 267461 337495 267519 337501
rect 274729 337501 274741 337504
rect 274775 337501 274787 337535
rect 274729 337495 274787 337501
rect 275925 337535 275983 337541
rect 275925 337501 275937 337535
rect 275971 337532 275983 337535
rect 283006 337532 283012 337544
rect 275971 337504 283012 337532
rect 275971 337501 275983 337504
rect 275925 337495 275983 337501
rect 283006 337492 283012 337504
rect 283064 337492 283070 337544
rect 283742 337492 283748 337544
rect 283800 337532 283806 337544
rect 284110 337532 284116 337544
rect 283800 337504 284116 337532
rect 283800 337492 283806 337504
rect 284110 337492 284116 337504
rect 284168 337492 284174 337544
rect 284312 337532 284340 337572
rect 284846 337560 284852 337612
rect 284904 337600 284910 337612
rect 285490 337600 285496 337612
rect 284904 337572 285496 337600
rect 284904 337560 284910 337572
rect 285490 337560 285496 337572
rect 285548 337560 285554 337612
rect 287425 337603 287483 337609
rect 287425 337569 287437 337603
rect 287471 337600 287483 337603
rect 289909 337603 289967 337609
rect 289909 337600 289921 337603
rect 287471 337572 289921 337600
rect 287471 337569 287483 337572
rect 287425 337563 287483 337569
rect 289909 337569 289921 337572
rect 289955 337569 289967 337603
rect 289909 337563 289967 337569
rect 290093 337603 290151 337609
rect 290093 337569 290105 337603
rect 290139 337600 290151 337603
rect 316678 337600 316684 337612
rect 290139 337572 316684 337600
rect 290139 337569 290151 337572
rect 290093 337563 290151 337569
rect 316678 337560 316684 337572
rect 316736 337560 316742 337612
rect 289817 337535 289875 337541
rect 289817 337532 289829 337535
rect 284312 337504 289829 337532
rect 289817 337501 289829 337504
rect 289863 337501 289875 337535
rect 289817 337495 289875 337501
rect 290001 337535 290059 337541
rect 290001 337501 290013 337535
rect 290047 337532 290059 337535
rect 315298 337532 315304 337544
rect 290047 337504 315304 337532
rect 290047 337501 290059 337504
rect 290001 337495 290059 337501
rect 315298 337492 315304 337504
rect 315356 337492 315362 337544
rect 265618 337424 265624 337476
rect 265676 337464 265682 337476
rect 289909 337467 289967 337473
rect 289909 337464 289921 337467
rect 265676 337436 289921 337464
rect 265676 337424 265682 337436
rect 289909 337433 289921 337436
rect 289955 337433 289967 337467
rect 289909 337427 289967 337433
rect 290093 337467 290151 337473
rect 290093 337433 290105 337467
rect 290139 337464 290151 337467
rect 346394 337464 346400 337476
rect 290139 337436 346400 337464
rect 290139 337433 290151 337436
rect 290093 337427 290151 337433
rect 346394 337424 346400 337436
rect 346452 337424 346458 337476
rect 260616 337368 265572 337396
rect 260616 337356 260622 337368
rect 273254 337356 273260 337408
rect 273312 337396 273318 337408
rect 273438 337396 273444 337408
rect 273312 337368 273444 337396
rect 273312 337356 273318 337368
rect 273438 337356 273444 337368
rect 273496 337356 273502 337408
rect 276934 337356 276940 337408
rect 276992 337396 276998 337408
rect 277210 337396 277216 337408
rect 276992 337368 277216 337396
rect 276992 337356 276998 337368
rect 277210 337356 277216 337368
rect 277268 337356 277274 337408
rect 280430 337356 280436 337408
rect 280488 337396 280494 337408
rect 282825 337399 282883 337405
rect 282825 337396 282837 337399
rect 280488 337368 282837 337396
rect 280488 337356 280494 337368
rect 282825 337365 282837 337368
rect 282871 337365 282883 337399
rect 282825 337359 282883 337365
rect 285950 337356 285956 337408
rect 286008 337396 286014 337408
rect 289817 337399 289875 337405
rect 289817 337396 289829 337399
rect 286008 337368 289829 337396
rect 286008 337356 286014 337368
rect 289817 337365 289829 337368
rect 289863 337365 289875 337399
rect 289817 337359 289875 337365
rect 291473 337399 291531 337405
rect 291473 337365 291485 337399
rect 291519 337396 291531 337399
rect 308953 337399 309011 337405
rect 308953 337396 308965 337399
rect 291519 337368 308965 337396
rect 291519 337365 291531 337368
rect 291473 337359 291531 337365
rect 308953 337365 308965 337368
rect 308999 337365 309011 337399
rect 308953 337359 309011 337365
rect 321557 337399 321615 337405
rect 321557 337365 321569 337399
rect 321603 337396 321615 337399
rect 482925 337399 482983 337405
rect 321603 337368 328500 337396
rect 321603 337365 321615 337368
rect 321557 337359 321615 337365
rect 226978 337288 226984 337340
rect 227036 337328 227042 337340
rect 235905 337331 235963 337337
rect 235905 337328 235917 337331
rect 227036 337300 235917 337328
rect 227036 337288 227042 337300
rect 235905 337297 235917 337300
rect 235951 337297 235963 337331
rect 235905 337291 235963 337297
rect 258626 337288 258632 337340
rect 258684 337328 258690 337340
rect 261757 337331 261815 337337
rect 261757 337328 261769 337331
rect 258684 337300 261769 337328
rect 258684 337288 258690 337300
rect 261757 337297 261769 337300
rect 261803 337297 261815 337331
rect 261757 337291 261815 337297
rect 264330 337288 264336 337340
rect 264388 337328 264394 337340
rect 264790 337328 264796 337340
rect 264388 337300 264796 337328
rect 264388 337288 264394 337300
rect 264790 337288 264796 337300
rect 264848 337288 264854 337340
rect 268010 337288 268016 337340
rect 268068 337328 268074 337340
rect 269022 337328 269028 337340
rect 268068 337300 269028 337328
rect 268068 337288 268074 337300
rect 269022 337288 269028 337300
rect 269080 337288 269086 337340
rect 277857 337331 277915 337337
rect 277857 337297 277869 337331
rect 277903 337328 277915 337331
rect 281074 337328 281080 337340
rect 277903 337300 281080 337328
rect 277903 337297 277915 337300
rect 277857 337291 277915 337297
rect 281074 337288 281080 337300
rect 281132 337288 281138 337340
rect 328472 337337 328500 337368
rect 347700 337368 347820 337396
rect 347700 337337 347728 337368
rect 347792 337337 347820 337368
rect 367020 337368 367140 337396
rect 367020 337337 367048 337368
rect 367112 337337 367140 337368
rect 386340 337368 386460 337396
rect 386340 337337 386368 337368
rect 386432 337337 386460 337368
rect 405660 337368 405780 337396
rect 405660 337337 405688 337368
rect 405752 337337 405780 337368
rect 424980 337368 425100 337396
rect 424980 337337 425008 337368
rect 425072 337337 425100 337368
rect 444300 337368 444420 337396
rect 444300 337337 444328 337368
rect 444392 337337 444420 337368
rect 463620 337368 463740 337396
rect 463620 337337 463648 337368
rect 463712 337337 463740 337368
rect 482925 337365 482937 337399
rect 482971 337396 482983 337399
rect 483569 337399 483627 337405
rect 483569 337396 483581 337399
rect 482971 337368 483581 337396
rect 482971 337365 482983 337368
rect 482925 337359 482983 337365
rect 483569 337365 483581 337368
rect 483615 337365 483627 337399
rect 483569 337359 483627 337365
rect 284573 337331 284631 337337
rect 284573 337297 284585 337331
rect 284619 337328 284631 337331
rect 290093 337331 290151 337337
rect 290093 337328 290105 337331
rect 284619 337300 290105 337328
rect 284619 337297 284631 337300
rect 284573 337291 284631 337297
rect 290093 337297 290105 337300
rect 290139 337297 290151 337331
rect 290093 337291 290151 337297
rect 290185 337331 290243 337337
rect 290185 337297 290197 337331
rect 290231 337328 290243 337331
rect 298833 337331 298891 337337
rect 298833 337328 298845 337331
rect 290231 337300 298845 337328
rect 290231 337297 290243 337300
rect 290185 337291 290243 337297
rect 298833 337297 298845 337300
rect 298879 337297 298891 337331
rect 298833 337291 298891 337297
rect 309045 337331 309103 337337
rect 309045 337297 309057 337331
rect 309091 337328 309103 337331
rect 311805 337331 311863 337337
rect 311805 337328 311817 337331
rect 309091 337300 311817 337328
rect 309091 337297 309103 337300
rect 309045 337291 309103 337297
rect 311805 337297 311817 337300
rect 311851 337297 311863 337331
rect 311805 337291 311863 337297
rect 311989 337331 312047 337337
rect 311989 337297 312001 337331
rect 312035 337328 312047 337331
rect 321465 337331 321523 337337
rect 321465 337328 321477 337331
rect 312035 337300 321477 337328
rect 312035 337297 312047 337300
rect 311989 337291 312047 337297
rect 321465 337297 321477 337300
rect 321511 337297 321523 337331
rect 321465 337291 321523 337297
rect 328457 337331 328515 337337
rect 328457 337297 328469 337331
rect 328503 337297 328515 337331
rect 328457 337291 328515 337297
rect 347685 337331 347743 337337
rect 347685 337297 347697 337331
rect 347731 337297 347743 337331
rect 347685 337291 347743 337297
rect 347777 337331 347835 337337
rect 347777 337297 347789 337331
rect 347823 337297 347835 337331
rect 347777 337291 347835 337297
rect 352101 337331 352159 337337
rect 352101 337297 352113 337331
rect 352147 337328 352159 337331
rect 357437 337331 357495 337337
rect 357437 337328 357449 337331
rect 352147 337300 357449 337328
rect 352147 337297 352159 337300
rect 352101 337291 352159 337297
rect 357437 337297 357449 337300
rect 357483 337297 357495 337331
rect 357437 337291 357495 337297
rect 367005 337331 367063 337337
rect 367005 337297 367017 337331
rect 367051 337297 367063 337331
rect 367005 337291 367063 337297
rect 367097 337331 367155 337337
rect 367097 337297 367109 337331
rect 367143 337297 367155 337331
rect 367097 337291 367155 337297
rect 371421 337331 371479 337337
rect 371421 337297 371433 337331
rect 371467 337328 371479 337331
rect 376757 337331 376815 337337
rect 376757 337328 376769 337331
rect 371467 337300 376769 337328
rect 371467 337297 371479 337300
rect 371421 337291 371479 337297
rect 376757 337297 376769 337300
rect 376803 337297 376815 337331
rect 376757 337291 376815 337297
rect 386325 337331 386383 337337
rect 386325 337297 386337 337331
rect 386371 337297 386383 337331
rect 386325 337291 386383 337297
rect 386417 337331 386475 337337
rect 386417 337297 386429 337331
rect 386463 337297 386475 337331
rect 386417 337291 386475 337297
rect 390741 337331 390799 337337
rect 390741 337297 390753 337331
rect 390787 337328 390799 337331
rect 396077 337331 396135 337337
rect 396077 337328 396089 337331
rect 390787 337300 396089 337328
rect 390787 337297 390799 337300
rect 390741 337291 390799 337297
rect 396077 337297 396089 337300
rect 396123 337297 396135 337331
rect 396077 337291 396135 337297
rect 405645 337331 405703 337337
rect 405645 337297 405657 337331
rect 405691 337297 405703 337331
rect 405645 337291 405703 337297
rect 405737 337331 405795 337337
rect 405737 337297 405749 337331
rect 405783 337297 405795 337331
rect 405737 337291 405795 337297
rect 410061 337331 410119 337337
rect 410061 337297 410073 337331
rect 410107 337328 410119 337331
rect 415397 337331 415455 337337
rect 415397 337328 415409 337331
rect 410107 337300 415409 337328
rect 410107 337297 410119 337300
rect 410061 337291 410119 337297
rect 415397 337297 415409 337300
rect 415443 337297 415455 337331
rect 415397 337291 415455 337297
rect 424965 337331 425023 337337
rect 424965 337297 424977 337331
rect 425011 337297 425023 337331
rect 424965 337291 425023 337297
rect 425057 337331 425115 337337
rect 425057 337297 425069 337331
rect 425103 337297 425115 337331
rect 425057 337291 425115 337297
rect 429381 337331 429439 337337
rect 429381 337297 429393 337331
rect 429427 337328 429439 337331
rect 434717 337331 434775 337337
rect 434717 337328 434729 337331
rect 429427 337300 434729 337328
rect 429427 337297 429439 337300
rect 429381 337291 429439 337297
rect 434717 337297 434729 337300
rect 434763 337297 434775 337331
rect 434717 337291 434775 337297
rect 444285 337331 444343 337337
rect 444285 337297 444297 337331
rect 444331 337297 444343 337331
rect 444285 337291 444343 337297
rect 444377 337331 444435 337337
rect 444377 337297 444389 337331
rect 444423 337297 444435 337331
rect 444377 337291 444435 337297
rect 448701 337331 448759 337337
rect 448701 337297 448713 337331
rect 448747 337328 448759 337331
rect 454037 337331 454095 337337
rect 454037 337328 454049 337331
rect 448747 337300 454049 337328
rect 448747 337297 448759 337300
rect 448701 337291 448759 337297
rect 454037 337297 454049 337300
rect 454083 337297 454095 337331
rect 454037 337291 454095 337297
rect 463605 337331 463663 337337
rect 463605 337297 463617 337331
rect 463651 337297 463663 337331
rect 463605 337291 463663 337297
rect 463697 337331 463755 337337
rect 463697 337297 463709 337331
rect 463743 337297 463755 337331
rect 463697 337291 463755 337297
rect 468021 337331 468079 337337
rect 468021 337297 468033 337331
rect 468067 337328 468079 337331
rect 473357 337331 473415 337337
rect 473357 337328 473369 337331
rect 468067 337300 473369 337328
rect 468067 337297 468079 337300
rect 468021 337291 468079 337297
rect 473357 337297 473369 337300
rect 473403 337297 473415 337331
rect 473357 337291 473415 337297
rect 222838 337220 222844 337272
rect 222896 337260 222902 337272
rect 241974 337260 241980 337272
rect 222896 337232 241980 337260
rect 222896 337220 222902 337232
rect 241974 337220 241980 337232
rect 242032 337220 242038 337272
rect 242986 337220 242992 337272
rect 243044 337260 243050 337272
rect 246206 337260 246212 337272
rect 243044 337232 246212 337260
rect 243044 337220 243050 337232
rect 246206 337220 246212 337232
rect 246264 337220 246270 337272
rect 259638 337220 259644 337272
rect 259696 337260 259702 337272
rect 262214 337260 262220 337272
rect 259696 337232 262220 337260
rect 259696 337220 259702 337232
rect 262214 337220 262220 337232
rect 262272 337220 262278 337272
rect 266722 337220 266728 337272
rect 266780 337260 266786 337272
rect 267550 337260 267556 337272
rect 266780 337232 267556 337260
rect 266780 337220 266786 337232
rect 267550 337220 267556 337232
rect 267608 337220 267614 337272
rect 277026 337220 277032 337272
rect 277084 337260 277090 337272
rect 277394 337260 277400 337272
rect 277084 337232 277400 337260
rect 277084 337220 277090 337232
rect 277394 337220 277400 337232
rect 277452 337220 277458 337272
rect 287977 337263 288035 337269
rect 287977 337229 287989 337263
rect 288023 337260 288035 337263
rect 290458 337260 290464 337272
rect 288023 337232 290464 337260
rect 288023 337229 288035 337232
rect 287977 337223 288035 337229
rect 290458 337220 290464 337232
rect 290516 337220 290522 337272
rect 225690 337152 225696 337204
rect 225748 337192 225754 337204
rect 245102 337192 245108 337204
rect 225748 337164 245108 337192
rect 225748 337152 225754 337164
rect 245102 337152 245108 337164
rect 245160 337152 245166 337204
rect 260098 337152 260104 337204
rect 260156 337192 260162 337204
rect 260742 337192 260748 337204
rect 260156 337164 260748 337192
rect 260156 337152 260162 337164
rect 260742 337152 260748 337164
rect 260800 337152 260806 337204
rect 262490 337152 262496 337204
rect 262548 337192 262554 337204
rect 262950 337192 262956 337204
rect 262548 337164 262956 337192
rect 262548 337152 262554 337164
rect 262950 337152 262956 337164
rect 263008 337152 263014 337204
rect 268010 337152 268016 337204
rect 268068 337192 268074 337204
rect 268654 337192 268660 337204
rect 268068 337164 268660 337192
rect 268068 337152 268074 337164
rect 268654 337152 268660 337164
rect 268712 337152 268718 337204
rect 277854 337152 277860 337204
rect 277912 337192 277918 337204
rect 279234 337192 279240 337204
rect 277912 337164 279240 337192
rect 277912 337152 277918 337164
rect 279234 337152 279240 337164
rect 279292 337152 279298 337204
rect 280706 337152 280712 337204
rect 280764 337192 280770 337204
rect 281166 337192 281172 337204
rect 280764 337164 281172 337192
rect 280764 337152 280770 337164
rect 281166 337152 281172 337164
rect 281224 337152 281230 337204
rect 281534 337152 281540 337204
rect 281592 337192 281598 337204
rect 281592 337164 282592 337192
rect 281592 337152 281598 337164
rect 228358 337084 228364 337136
rect 228416 337124 228422 337136
rect 240045 337127 240103 337133
rect 228416 337096 239444 337124
rect 228416 337084 228422 337096
rect 239416 337056 239444 337096
rect 240045 337093 240057 337127
rect 240091 337124 240103 337127
rect 254578 337124 254584 337136
rect 240091 337096 254584 337124
rect 240091 337093 240103 337096
rect 240045 337087 240103 337093
rect 254578 337084 254584 337096
rect 254636 337084 254642 337136
rect 257430 337084 257436 337136
rect 257488 337124 257494 337136
rect 257488 337096 259684 337124
rect 257488 337084 257494 337096
rect 246758 337056 246764 337068
rect 239416 337028 246764 337056
rect 246758 337016 246764 337028
rect 246816 337016 246822 337068
rect 246942 337016 246948 337068
rect 247000 337056 247006 337068
rect 252922 337056 252928 337068
rect 247000 337028 252928 337056
rect 247000 337016 247006 337028
rect 252922 337016 252928 337028
rect 252980 337016 252986 337068
rect 256694 337016 256700 337068
rect 256752 337056 256758 337068
rect 258534 337056 258540 337068
rect 256752 337028 258540 337056
rect 256752 337016 256758 337028
rect 258534 337016 258540 337028
rect 258592 337016 258598 337068
rect 248506 336948 248512 337000
rect 248564 336988 248570 337000
rect 251266 336988 251272 337000
rect 248564 336960 251272 336988
rect 248564 336948 248570 336960
rect 251266 336948 251272 336960
rect 251324 336948 251330 337000
rect 252186 336948 252192 337000
rect 252244 336988 252250 337000
rect 252554 336988 252560 337000
rect 252244 336960 252560 336988
rect 252244 336948 252250 336960
rect 252554 336948 252560 336960
rect 252612 336948 252618 337000
rect 256786 336880 256792 336932
rect 256844 336920 256850 336932
rect 257706 336920 257712 336932
rect 256844 336892 257712 336920
rect 256844 336880 256850 336892
rect 257706 336880 257712 336892
rect 257764 336880 257770 336932
rect 258258 336880 258264 336932
rect 258316 336920 258322 336932
rect 259086 336920 259092 336932
rect 258316 336892 259092 336920
rect 258316 336880 258322 336892
rect 259086 336880 259092 336892
rect 259144 336880 259150 336932
rect 251266 336812 251272 336864
rect 251324 336852 251330 336864
rect 253750 336852 253756 336864
rect 251324 336824 253756 336852
rect 251324 336812 251330 336824
rect 253750 336812 253756 336824
rect 253808 336812 253814 336864
rect 256510 336812 256516 336864
rect 256568 336852 256574 336864
rect 257338 336852 257344 336864
rect 256568 336824 257344 336852
rect 256568 336812 256574 336824
rect 257338 336812 257344 336824
rect 257396 336812 257402 336864
rect 258902 336812 258908 336864
rect 258960 336852 258966 336864
rect 259270 336852 259276 336864
rect 258960 336824 259276 336852
rect 258960 336812 258966 336824
rect 259270 336812 259276 336824
rect 259328 336812 259334 336864
rect 259656 336852 259684 337096
rect 259730 337084 259736 337136
rect 259788 337124 259794 337136
rect 263686 337124 263692 337136
rect 259788 337096 263692 337124
rect 259788 337084 259794 337096
rect 263686 337084 263692 337096
rect 263744 337084 263750 337136
rect 263962 337084 263968 337136
rect 264020 337124 264026 337136
rect 264882 337124 264888 337136
rect 264020 337096 264888 337124
rect 264020 337084 264026 337096
rect 264882 337084 264888 337096
rect 264940 337084 264946 337136
rect 267734 337084 267740 337136
rect 267792 337124 267798 337136
rect 273257 337127 273315 337133
rect 273257 337124 273269 337127
rect 267792 337096 273269 337124
rect 267792 337084 267798 337096
rect 273257 337093 273269 337096
rect 273303 337093 273315 337127
rect 273257 337087 273315 337093
rect 277394 337084 277400 337136
rect 277452 337124 277458 337136
rect 278590 337124 278596 337136
rect 277452 337096 278596 337124
rect 277452 337084 277458 337096
rect 278590 337084 278596 337096
rect 278648 337084 278654 337136
rect 282564 337124 282592 337164
rect 282914 337152 282920 337204
rect 282972 337192 282978 337204
rect 283282 337192 283288 337204
rect 282972 337164 283288 337192
rect 282972 337152 282978 337164
rect 283282 337152 283288 337164
rect 283340 337152 283346 337204
rect 283374 337152 283380 337204
rect 283432 337192 283438 337204
rect 284018 337192 284024 337204
rect 283432 337164 284024 337192
rect 283432 337152 283438 337164
rect 284018 337152 284024 337164
rect 284076 337152 284082 337204
rect 284386 337152 284392 337204
rect 284444 337192 284450 337204
rect 285398 337192 285404 337204
rect 284444 337164 285404 337192
rect 284444 337152 284450 337164
rect 285398 337152 285404 337164
rect 285456 337152 285462 337204
rect 287422 337152 287428 337204
rect 287480 337192 287486 337204
rect 287790 337192 287796 337204
rect 287480 337164 287796 337192
rect 287480 337152 287486 337164
rect 287790 337152 287796 337164
rect 287848 337152 287854 337204
rect 287885 337195 287943 337201
rect 287885 337161 287897 337195
rect 287931 337192 287943 337195
rect 291838 337192 291844 337204
rect 287931 337164 291844 337192
rect 287931 337161 287943 337164
rect 287885 337155 287943 337161
rect 291838 337152 291844 337164
rect 291896 337152 291902 337204
rect 328457 337195 328515 337201
rect 328457 337161 328469 337195
rect 328503 337192 328515 337195
rect 338117 337195 338175 337201
rect 338117 337192 338129 337195
rect 328503 337164 338129 337192
rect 328503 337161 328515 337164
rect 328457 337155 328515 337161
rect 338117 337161 338129 337164
rect 338163 337161 338175 337195
rect 338117 337155 338175 337161
rect 347777 337195 347835 337201
rect 347777 337161 347789 337195
rect 347823 337192 347835 337195
rect 352101 337195 352159 337201
rect 352101 337192 352113 337195
rect 347823 337164 352113 337192
rect 347823 337161 347835 337164
rect 347777 337155 347835 337161
rect 352101 337161 352113 337164
rect 352147 337161 352159 337195
rect 352101 337155 352159 337161
rect 357437 337195 357495 337201
rect 357437 337161 357449 337195
rect 357483 337192 357495 337195
rect 367005 337195 367063 337201
rect 367005 337192 367017 337195
rect 357483 337164 367017 337192
rect 357483 337161 357495 337164
rect 357437 337155 357495 337161
rect 367005 337161 367017 337164
rect 367051 337161 367063 337195
rect 367005 337155 367063 337161
rect 367097 337195 367155 337201
rect 367097 337161 367109 337195
rect 367143 337192 367155 337195
rect 371421 337195 371479 337201
rect 371421 337192 371433 337195
rect 367143 337164 371433 337192
rect 367143 337161 367155 337164
rect 367097 337155 367155 337161
rect 371421 337161 371433 337164
rect 371467 337161 371479 337195
rect 371421 337155 371479 337161
rect 376757 337195 376815 337201
rect 376757 337161 376769 337195
rect 376803 337192 376815 337195
rect 386325 337195 386383 337201
rect 386325 337192 386337 337195
rect 376803 337164 386337 337192
rect 376803 337161 376815 337164
rect 376757 337155 376815 337161
rect 386325 337161 386337 337164
rect 386371 337161 386383 337195
rect 386325 337155 386383 337161
rect 386417 337195 386475 337201
rect 386417 337161 386429 337195
rect 386463 337192 386475 337195
rect 390741 337195 390799 337201
rect 390741 337192 390753 337195
rect 386463 337164 390753 337192
rect 386463 337161 386475 337164
rect 386417 337155 386475 337161
rect 390741 337161 390753 337164
rect 390787 337161 390799 337195
rect 390741 337155 390799 337161
rect 396077 337195 396135 337201
rect 396077 337161 396089 337195
rect 396123 337192 396135 337195
rect 405645 337195 405703 337201
rect 405645 337192 405657 337195
rect 396123 337164 405657 337192
rect 396123 337161 396135 337164
rect 396077 337155 396135 337161
rect 405645 337161 405657 337164
rect 405691 337161 405703 337195
rect 405645 337155 405703 337161
rect 405737 337195 405795 337201
rect 405737 337161 405749 337195
rect 405783 337192 405795 337195
rect 410061 337195 410119 337201
rect 410061 337192 410073 337195
rect 405783 337164 410073 337192
rect 405783 337161 405795 337164
rect 405737 337155 405795 337161
rect 410061 337161 410073 337164
rect 410107 337161 410119 337195
rect 410061 337155 410119 337161
rect 415397 337195 415455 337201
rect 415397 337161 415409 337195
rect 415443 337192 415455 337195
rect 424965 337195 425023 337201
rect 424965 337192 424977 337195
rect 415443 337164 424977 337192
rect 415443 337161 415455 337164
rect 415397 337155 415455 337161
rect 424965 337161 424977 337164
rect 425011 337161 425023 337195
rect 424965 337155 425023 337161
rect 425057 337195 425115 337201
rect 425057 337161 425069 337195
rect 425103 337192 425115 337195
rect 429381 337195 429439 337201
rect 429381 337192 429393 337195
rect 425103 337164 429393 337192
rect 425103 337161 425115 337164
rect 425057 337155 425115 337161
rect 429381 337161 429393 337164
rect 429427 337161 429439 337195
rect 429381 337155 429439 337161
rect 434717 337195 434775 337201
rect 434717 337161 434729 337195
rect 434763 337192 434775 337195
rect 444285 337195 444343 337201
rect 444285 337192 444297 337195
rect 434763 337164 444297 337192
rect 434763 337161 434775 337164
rect 434717 337155 434775 337161
rect 444285 337161 444297 337164
rect 444331 337161 444343 337195
rect 444285 337155 444343 337161
rect 444377 337195 444435 337201
rect 444377 337161 444389 337195
rect 444423 337192 444435 337195
rect 448701 337195 448759 337201
rect 448701 337192 448713 337195
rect 444423 337164 448713 337192
rect 444423 337161 444435 337164
rect 444377 337155 444435 337161
rect 448701 337161 448713 337164
rect 448747 337161 448759 337195
rect 448701 337155 448759 337161
rect 454037 337195 454095 337201
rect 454037 337161 454049 337195
rect 454083 337192 454095 337195
rect 463605 337195 463663 337201
rect 463605 337192 463617 337195
rect 454083 337164 463617 337192
rect 454083 337161 454095 337164
rect 454037 337155 454095 337161
rect 463605 337161 463617 337164
rect 463651 337161 463663 337195
rect 463605 337155 463663 337161
rect 463697 337195 463755 337201
rect 463697 337161 463709 337195
rect 463743 337192 463755 337195
rect 468021 337195 468079 337201
rect 468021 337192 468033 337195
rect 463743 337164 468033 337192
rect 463743 337161 463755 337164
rect 463697 337155 463755 337161
rect 468021 337161 468033 337164
rect 468067 337161 468079 337195
rect 468021 337155 468079 337161
rect 473357 337195 473415 337201
rect 473357 337161 473369 337195
rect 473403 337192 473415 337195
rect 482925 337195 482983 337201
rect 482925 337192 482937 337195
rect 473403 337164 482937 337192
rect 473403 337161 473415 337164
rect 473357 337155 473415 337161
rect 482925 337161 482937 337164
rect 482971 337161 482983 337195
rect 482925 337155 482983 337161
rect 284573 337127 284631 337133
rect 284573 337124 284585 337127
rect 282564 337096 284585 337124
rect 284573 337093 284585 337096
rect 284619 337093 284631 337127
rect 284573 337087 284631 337093
rect 289262 337084 289268 337136
rect 289320 337124 289326 337136
rect 289538 337124 289544 337136
rect 289320 337096 289544 337124
rect 289320 337084 289326 337096
rect 289538 337084 289544 337096
rect 289596 337084 289602 337136
rect 260190 337016 260196 337068
rect 260248 337056 260254 337068
rect 268289 337059 268347 337065
rect 268289 337056 268301 337059
rect 260248 337028 268301 337056
rect 260248 337016 260254 337028
rect 268289 337025 268301 337028
rect 268335 337025 268347 337059
rect 268289 337019 268347 337025
rect 269114 337016 269120 337068
rect 269172 337056 269178 337068
rect 269850 337056 269856 337068
rect 269172 337028 269856 337056
rect 269172 337016 269178 337028
rect 269850 337016 269856 337028
rect 269908 337016 269914 337068
rect 273346 337016 273352 337068
rect 273404 337056 273410 337068
rect 274358 337056 274364 337068
rect 273404 337028 274364 337056
rect 273404 337016 273410 337028
rect 274358 337016 274364 337028
rect 274416 337016 274422 337068
rect 274910 337016 274916 337068
rect 274968 337056 274974 337068
rect 274968 337028 277440 337056
rect 274968 337016 274974 337028
rect 263778 336948 263784 337000
rect 263836 336988 263842 337000
rect 264422 336988 264428 337000
rect 263836 336960 264428 336988
rect 263836 336948 263842 336960
rect 264422 336948 264428 336960
rect 264480 336948 264486 337000
rect 266354 336948 266360 337000
rect 266412 336988 266418 337000
rect 267182 336988 267188 337000
rect 266412 336960 267188 336988
rect 266412 336948 266418 336960
rect 267182 336948 267188 336960
rect 267240 336948 267246 337000
rect 269390 336948 269396 337000
rect 269448 336988 269454 337000
rect 269448 336960 270264 336988
rect 269448 336948 269454 336960
rect 261202 336880 261208 336932
rect 261260 336920 261266 336932
rect 261846 336920 261852 336932
rect 261260 336892 261852 336920
rect 261260 336880 261266 336892
rect 261846 336880 261852 336892
rect 261904 336880 261910 336932
rect 269482 336880 269488 336932
rect 269540 336920 269546 336932
rect 270034 336920 270040 336932
rect 269540 336892 270040 336920
rect 269540 336880 269546 336892
rect 270034 336880 270040 336892
rect 270092 336880 270098 336932
rect 259656 336824 260972 336852
rect 230382 336744 230388 336796
rect 230440 336784 230446 336796
rect 231302 336784 231308 336796
rect 230440 336756 231308 336784
rect 230440 336744 230446 336756
rect 231302 336744 231308 336756
rect 231360 336744 231366 336796
rect 237098 336744 237104 336796
rect 237156 336784 237162 336796
rect 239030 336784 239036 336796
rect 237156 336756 239036 336784
rect 237156 336744 237162 336756
rect 239030 336744 239036 336756
rect 239088 336744 239094 336796
rect 240962 336744 240968 336796
rect 241020 336784 241026 336796
rect 241606 336784 241612 336796
rect 241020 336756 241612 336784
rect 241020 336744 241026 336756
rect 241606 336744 241612 336756
rect 241664 336744 241670 336796
rect 244274 336744 244280 336796
rect 244332 336784 244338 336796
rect 245838 336784 245844 336796
rect 244332 336756 245844 336784
rect 244332 336744 244338 336756
rect 245838 336744 245844 336756
rect 245896 336744 245902 336796
rect 254578 336744 254584 336796
rect 254636 336784 254642 336796
rect 255406 336784 255412 336796
rect 254636 336756 255412 336784
rect 254636 336744 254642 336756
rect 255406 336744 255412 336756
rect 255464 336744 255470 336796
rect 257430 336744 257436 336796
rect 257488 336784 257494 336796
rect 257890 336784 257896 336796
rect 257488 336756 257896 336784
rect 257488 336744 257494 336756
rect 257890 336744 257896 336756
rect 257948 336744 257954 336796
rect 258166 336744 258172 336796
rect 258224 336784 258230 336796
rect 258626 336784 258632 336796
rect 258224 336756 258632 336784
rect 258224 336744 258230 336756
rect 258626 336744 258632 336756
rect 258684 336744 258690 336796
rect 258718 336744 258724 336796
rect 258776 336784 258782 336796
rect 259086 336784 259092 336796
rect 258776 336756 259092 336784
rect 258776 336744 258782 336756
rect 259086 336744 259092 336756
rect 259144 336744 259150 336796
rect 259454 336744 259460 336796
rect 259512 336784 259518 336796
rect 260374 336784 260380 336796
rect 259512 336756 260380 336784
rect 259512 336744 259518 336756
rect 260374 336744 260380 336756
rect 260432 336744 260438 336796
rect 233786 336608 233792 336660
rect 233844 336648 233850 336660
rect 236822 336648 236828 336660
rect 233844 336620 236828 336648
rect 233844 336608 233850 336620
rect 236822 336608 236828 336620
rect 236880 336608 236886 336660
rect 260944 336648 260972 336824
rect 262858 336812 262864 336864
rect 262916 336852 262922 336864
rect 263226 336852 263232 336864
rect 262916 336824 263232 336852
rect 262916 336812 262922 336824
rect 263226 336812 263232 336824
rect 263284 336812 263290 336864
rect 264146 336812 264152 336864
rect 264204 336852 264210 336864
rect 264606 336852 264612 336864
rect 264204 336824 264612 336852
rect 264204 336812 264210 336824
rect 264606 336812 264612 336824
rect 264664 336812 264670 336864
rect 265342 336812 265348 336864
rect 265400 336852 265406 336864
rect 266262 336852 266268 336864
rect 265400 336824 266268 336852
rect 265400 336812 265406 336824
rect 266262 336812 266268 336824
rect 266320 336812 266326 336864
rect 267090 336812 267096 336864
rect 267148 336852 267154 336864
rect 267458 336852 267464 336864
rect 267148 336824 267464 336852
rect 267148 336812 267154 336824
rect 267458 336812 267464 336824
rect 267516 336812 267522 336864
rect 267826 336812 267832 336864
rect 267884 336852 267890 336864
rect 268378 336852 268384 336864
rect 267884 336824 268384 336852
rect 267884 336812 267890 336824
rect 268378 336812 268384 336824
rect 268436 336812 268442 336864
rect 269574 336812 269580 336864
rect 269632 336852 269638 336864
rect 270126 336852 270132 336864
rect 269632 336824 270132 336852
rect 269632 336812 269638 336824
rect 270126 336812 270132 336824
rect 270184 336812 270190 336864
rect 261018 336744 261024 336796
rect 261076 336784 261082 336796
rect 261478 336784 261484 336796
rect 261076 336756 261484 336784
rect 261076 336744 261082 336756
rect 261478 336744 261484 336756
rect 261536 336744 261542 336796
rect 262766 336744 262772 336796
rect 262824 336784 262830 336796
rect 263134 336784 263140 336796
rect 262824 336756 263140 336784
rect 262824 336744 262830 336756
rect 263134 336744 263140 336756
rect 263192 336744 263198 336796
rect 265618 336744 265624 336796
rect 265676 336784 265682 336796
rect 265676 336756 265721 336784
rect 265676 336744 265682 336756
rect 266630 336744 266636 336796
rect 266688 336784 266694 336796
rect 266688 336756 266860 336784
rect 266688 336744 266694 336756
rect 262858 336716 262864 336728
rect 262819 336688 262864 336716
rect 262858 336676 262864 336688
rect 262916 336676 262922 336728
rect 266262 336716 266268 336728
rect 266223 336688 266268 336716
rect 266262 336676 266268 336688
rect 266320 336676 266326 336728
rect 266832 336725 266860 336756
rect 266906 336744 266912 336796
rect 266964 336784 266970 336796
rect 267366 336784 267372 336796
rect 266964 336756 267372 336784
rect 266964 336744 266970 336756
rect 267366 336744 267372 336756
rect 267424 336744 267430 336796
rect 267734 336744 267740 336796
rect 267792 336784 267798 336796
rect 268286 336784 268292 336796
rect 267792 336756 268292 336784
rect 267792 336744 267798 336756
rect 268286 336744 268292 336756
rect 268344 336744 268350 336796
rect 268930 336784 268936 336796
rect 268396 336756 268936 336784
rect 266817 336719 266875 336725
rect 266817 336685 266829 336719
rect 266863 336716 266875 336719
rect 266863 336688 266897 336716
rect 266863 336685 266875 336688
rect 266817 336679 266875 336685
rect 267826 336676 267832 336728
rect 267884 336716 267890 336728
rect 268396 336716 268424 336756
rect 268930 336744 268936 336756
rect 268988 336744 268994 336796
rect 269390 336744 269396 336796
rect 269448 336784 269454 336796
rect 269758 336784 269764 336796
rect 269448 336756 269764 336784
rect 269448 336744 269454 336756
rect 269758 336744 269764 336756
rect 269816 336744 269822 336796
rect 270236 336784 270264 336960
rect 273530 336948 273536 337000
rect 273588 336988 273594 337000
rect 274082 336988 274088 337000
rect 273588 336960 274088 336988
rect 273588 336948 273594 336960
rect 274082 336948 274088 336960
rect 274140 336948 274146 337000
rect 275278 336948 275284 337000
rect 275336 336988 275342 337000
rect 275554 336988 275560 337000
rect 275336 336960 275560 336988
rect 275336 336948 275342 336960
rect 275554 336948 275560 336960
rect 275612 336948 275618 337000
rect 276014 336948 276020 337000
rect 276072 336988 276078 337000
rect 276842 336988 276848 337000
rect 276072 336960 276848 336988
rect 276072 336948 276078 336960
rect 276842 336948 276848 336960
rect 276900 336948 276906 337000
rect 273346 336880 273352 336932
rect 273404 336920 273410 336932
rect 273806 336920 273812 336932
rect 273404 336892 273812 336920
rect 273404 336880 273410 336892
rect 273806 336880 273812 336892
rect 273864 336880 273870 336932
rect 273622 336812 273628 336864
rect 273680 336852 273686 336864
rect 274174 336852 274180 336864
rect 273680 336824 274180 336852
rect 273680 336812 273686 336824
rect 274174 336812 274180 336824
rect 274232 336812 274238 336864
rect 276198 336812 276204 336864
rect 276256 336852 276262 336864
rect 277118 336852 277124 336864
rect 276256 336824 277124 336852
rect 276256 336812 276262 336824
rect 277118 336812 277124 336824
rect 277176 336812 277182 336864
rect 270144 336756 270264 336784
rect 270144 336728 270172 336756
rect 271966 336744 271972 336796
rect 272024 336784 272030 336796
rect 272242 336784 272248 336796
rect 272024 336756 272248 336784
rect 272024 336744 272030 336756
rect 272242 336744 272248 336756
rect 272300 336744 272306 336796
rect 272334 336744 272340 336796
rect 272392 336784 272398 336796
rect 272610 336784 272616 336796
rect 272392 336756 272616 336784
rect 272392 336744 272398 336756
rect 272610 336744 272616 336756
rect 272668 336744 272674 336796
rect 272702 336744 272708 336796
rect 272760 336784 272766 336796
rect 272760 336756 272840 336784
rect 272760 336744 272766 336756
rect 269022 336716 269028 336728
rect 267884 336688 268424 336716
rect 268983 336688 269028 336716
rect 267884 336676 267890 336688
rect 269022 336676 269028 336688
rect 269080 336676 269086 336728
rect 270126 336676 270132 336728
rect 270184 336676 270190 336728
rect 261018 336648 261024 336660
rect 260944 336620 261024 336648
rect 261018 336608 261024 336620
rect 261076 336608 261082 336660
rect 272812 336648 272840 336756
rect 272886 336744 272892 336796
rect 272944 336784 272950 336796
rect 273070 336784 273076 336796
rect 272944 336756 273076 336784
rect 272944 336744 272950 336756
rect 273070 336744 273076 336756
rect 273128 336744 273134 336796
rect 273438 336744 273444 336796
rect 273496 336784 273502 336796
rect 273898 336784 273904 336796
rect 273496 336756 273904 336784
rect 273496 336744 273502 336756
rect 273898 336744 273904 336756
rect 273956 336744 273962 336796
rect 274450 336784 274456 336796
rect 274008 336756 274456 336784
rect 273162 336716 273168 336728
rect 273123 336688 273168 336716
rect 273162 336676 273168 336688
rect 273220 336676 273226 336728
rect 273530 336676 273536 336728
rect 273588 336716 273594 336728
rect 274008 336716 274036 336756
rect 274450 336744 274456 336756
rect 274508 336744 274514 336796
rect 275002 336744 275008 336796
rect 275060 336784 275066 336796
rect 275186 336784 275192 336796
rect 275060 336756 275192 336784
rect 275060 336744 275066 336756
rect 275186 336744 275192 336756
rect 275244 336744 275250 336796
rect 275278 336744 275284 336796
rect 275336 336784 275342 336796
rect 275462 336784 275468 336796
rect 275336 336756 275468 336784
rect 275336 336744 275342 336756
rect 275462 336744 275468 336756
rect 275520 336744 275526 336796
rect 276474 336744 276480 336796
rect 276532 336784 276538 336796
rect 276842 336784 276848 336796
rect 276532 336756 276848 336784
rect 276532 336744 276538 336756
rect 276842 336744 276848 336756
rect 276900 336744 276906 336796
rect 277412 336784 277440 337028
rect 277854 337016 277860 337068
rect 277912 337056 277918 337068
rect 278682 337056 278688 337068
rect 277912 337028 278688 337056
rect 277912 337016 277918 337028
rect 278682 337016 278688 337028
rect 278740 337016 278746 337068
rect 281810 337016 281816 337068
rect 281868 337056 281874 337068
rect 282362 337056 282368 337068
rect 281868 337028 282368 337056
rect 281868 337016 281874 337028
rect 282362 337016 282368 337028
rect 282420 337016 282426 337068
rect 284478 337016 284484 337068
rect 284536 337056 284542 337068
rect 285306 337056 285312 337068
rect 284536 337028 285312 337056
rect 284536 337016 284542 337028
rect 285306 337016 285312 337028
rect 285364 337016 285370 337068
rect 285582 337056 285588 337068
rect 285543 337028 285588 337056
rect 285582 337016 285588 337028
rect 285640 337016 285646 337068
rect 286318 337016 286324 337068
rect 286376 337056 286382 337068
rect 286962 337056 286968 337068
rect 286376 337028 286968 337056
rect 286376 337016 286382 337028
rect 286962 337016 286968 337028
rect 287020 337016 287026 337068
rect 291473 337059 291531 337065
rect 291473 337056 291485 337059
rect 287716 337028 291485 337056
rect 277578 336948 277584 337000
rect 277636 336988 277642 337000
rect 278590 336988 278596 337000
rect 277636 336960 278596 336988
rect 277636 336948 277642 336960
rect 278590 336948 278596 336960
rect 278648 336948 278654 337000
rect 280706 336948 280712 337000
rect 280764 336988 280770 337000
rect 281350 336988 281356 337000
rect 280764 336960 281356 336988
rect 280764 336948 280770 336960
rect 281350 336948 281356 336960
rect 281408 336948 281414 337000
rect 282086 336948 282092 337000
rect 282144 336988 282150 337000
rect 282638 336988 282644 337000
rect 282144 336960 282644 336988
rect 282144 336948 282150 336960
rect 282638 336948 282644 336960
rect 282696 336948 282702 337000
rect 282733 336991 282791 336997
rect 282733 336957 282745 336991
rect 282779 336988 282791 336991
rect 287716 336988 287744 337028
rect 291473 337025 291485 337028
rect 291519 337025 291531 337059
rect 291473 337019 291531 337025
rect 338117 337059 338175 337065
rect 338117 337025 338129 337059
rect 338163 337056 338175 337059
rect 347685 337059 347743 337065
rect 347685 337056 347697 337059
rect 338163 337028 347697 337056
rect 338163 337025 338175 337028
rect 338117 337019 338175 337025
rect 347685 337025 347697 337028
rect 347731 337025 347743 337059
rect 347685 337019 347743 337025
rect 282779 336960 287744 336988
rect 282779 336957 282791 336960
rect 282733 336951 282791 336957
rect 288526 336948 288532 337000
rect 288584 336988 288590 337000
rect 290734 336988 290740 337000
rect 288584 336960 290740 336988
rect 288584 336948 288590 336960
rect 290734 336948 290740 336960
rect 290792 336948 290798 337000
rect 282270 336880 282276 336932
rect 282328 336920 282334 336932
rect 282822 336920 282828 336932
rect 282328 336892 282828 336920
rect 282328 336880 282334 336892
rect 282822 336880 282828 336892
rect 282880 336880 282886 336932
rect 287425 336923 287483 336929
rect 287425 336920 287437 336923
rect 283024 336892 287437 336920
rect 277486 336812 277492 336864
rect 277544 336852 277550 336864
rect 278314 336852 278320 336864
rect 277544 336824 278320 336852
rect 277544 336812 277550 336824
rect 278314 336812 278320 336824
rect 278372 336812 278378 336864
rect 279142 336812 279148 336864
rect 279200 336852 279206 336864
rect 280062 336852 280068 336864
rect 279200 336824 280068 336852
rect 279200 336812 279206 336824
rect 280062 336812 280068 336824
rect 280120 336812 280126 336864
rect 280614 336812 280620 336864
rect 280672 336852 280678 336864
rect 281350 336852 281356 336864
rect 280672 336824 281356 336852
rect 280672 336812 280678 336824
rect 281350 336812 281356 336824
rect 281408 336812 281414 336864
rect 281902 336812 281908 336864
rect 281960 336852 281966 336864
rect 282454 336852 282460 336864
rect 281960 336824 282460 336852
rect 281960 336812 281966 336824
rect 282454 336812 282460 336824
rect 282512 336812 282518 336864
rect 282549 336855 282607 336861
rect 282549 336821 282561 336855
rect 282595 336852 282607 336855
rect 282914 336852 282920 336864
rect 282595 336824 282920 336852
rect 282595 336821 282607 336824
rect 282549 336815 282607 336821
rect 282914 336812 282920 336824
rect 282972 336812 282978 336864
rect 277412 336756 277532 336784
rect 274358 336716 274364 336728
rect 273588 336688 274036 336716
rect 274319 336688 274364 336716
rect 273588 336676 273594 336688
rect 274358 336676 274364 336688
rect 274416 336676 274422 336728
rect 277504 336716 277532 336756
rect 277578 336744 277584 336796
rect 277636 336784 277642 336796
rect 277854 336784 277860 336796
rect 277636 336756 277860 336784
rect 277636 336744 277642 336756
rect 277854 336744 277860 336756
rect 277912 336744 277918 336796
rect 277946 336744 277952 336796
rect 278004 336784 278010 336796
rect 278406 336784 278412 336796
rect 278004 336756 278412 336784
rect 278004 336744 278010 336756
rect 278406 336744 278412 336756
rect 278464 336744 278470 336796
rect 279510 336744 279516 336796
rect 279568 336784 279574 336796
rect 279970 336784 279976 336796
rect 279568 336756 279976 336784
rect 279568 336744 279574 336756
rect 279970 336744 279976 336756
rect 280028 336744 280034 336796
rect 280154 336744 280160 336796
rect 280212 336784 280218 336796
rect 280430 336784 280436 336796
rect 280212 336756 280436 336784
rect 280212 336744 280218 336756
rect 280430 336744 280436 336756
rect 280488 336744 280494 336796
rect 280982 336744 280988 336796
rect 281040 336784 281046 336796
rect 281442 336784 281448 336796
rect 281040 336756 281448 336784
rect 281040 336744 281046 336756
rect 281442 336744 281448 336756
rect 281500 336744 281506 336796
rect 282178 336744 282184 336796
rect 282236 336784 282242 336796
rect 282730 336784 282736 336796
rect 282236 336756 282736 336784
rect 282236 336744 282242 336756
rect 282730 336744 282736 336756
rect 282788 336744 282794 336796
rect 282825 336787 282883 336793
rect 282825 336753 282837 336787
rect 282871 336784 282883 336787
rect 283024 336784 283052 336892
rect 287425 336889 287437 336892
rect 287471 336889 287483 336923
rect 287425 336883 287483 336889
rect 288986 336880 288992 336932
rect 289044 336920 289050 336932
rect 292022 336920 292028 336932
rect 289044 336892 292028 336920
rect 289044 336880 289050 336892
rect 292022 336880 292028 336892
rect 292080 336880 292086 336932
rect 283282 336812 283288 336864
rect 283340 336852 283346 336864
rect 283926 336852 283932 336864
rect 283340 336824 283932 336852
rect 283340 336812 283346 336824
rect 283926 336812 283932 336824
rect 283984 336812 283990 336864
rect 284570 336812 284576 336864
rect 284628 336852 284634 336864
rect 285122 336852 285128 336864
rect 284628 336824 285128 336852
rect 284628 336812 284634 336824
rect 285122 336812 285128 336824
rect 285180 336812 285186 336864
rect 285398 336852 285404 336864
rect 285359 336824 285404 336852
rect 285398 336812 285404 336824
rect 285456 336812 285462 336864
rect 286226 336812 286232 336864
rect 286284 336852 286290 336864
rect 286502 336852 286508 336864
rect 286284 336824 286508 336852
rect 286284 336812 286290 336824
rect 286502 336812 286508 336824
rect 286560 336812 286566 336864
rect 287330 336812 287336 336864
rect 287388 336852 287394 336864
rect 287974 336852 287980 336864
rect 287388 336824 287980 336852
rect 287388 336812 287394 336824
rect 287974 336812 287980 336824
rect 288032 336812 288038 336864
rect 288894 336812 288900 336864
rect 288952 336852 288958 336864
rect 290642 336852 290648 336864
rect 288952 336824 290648 336852
rect 288952 336812 288958 336824
rect 290642 336812 290648 336824
rect 290700 336812 290706 336864
rect 282871 336756 283052 336784
rect 282871 336753 282883 336756
rect 282825 336747 282883 336753
rect 283098 336744 283104 336796
rect 283156 336784 283162 336796
rect 283650 336784 283656 336796
rect 283156 336756 283656 336784
rect 283156 336744 283162 336756
rect 283650 336744 283656 336756
rect 283708 336744 283714 336796
rect 284294 336744 284300 336796
rect 284352 336784 284358 336796
rect 284352 336756 284892 336784
rect 284352 336744 284358 336756
rect 278682 336716 278688 336728
rect 277504 336688 278688 336716
rect 278682 336676 278688 336688
rect 278740 336676 278746 336728
rect 284864 336716 284892 336756
rect 284938 336744 284944 336796
rect 284996 336784 285002 336796
rect 285214 336784 285220 336796
rect 284996 336756 285220 336784
rect 284996 336744 285002 336756
rect 285214 336744 285220 336756
rect 285272 336744 285278 336796
rect 287238 336744 287244 336796
rect 287296 336784 287302 336796
rect 287606 336784 287612 336796
rect 287296 336756 287612 336784
rect 287296 336744 287302 336756
rect 287606 336744 287612 336756
rect 287664 336744 287670 336796
rect 285306 336716 285312 336728
rect 284864 336688 285312 336716
rect 285306 336676 285312 336688
rect 285364 336676 285370 336728
rect 289817 336719 289875 336725
rect 289817 336685 289829 336719
rect 289863 336716 289875 336719
rect 294690 336716 294696 336728
rect 289863 336688 294696 336716
rect 289863 336685 289875 336688
rect 289817 336679 289875 336685
rect 294690 336676 294696 336688
rect 294748 336676 294754 336728
rect 483569 336719 483627 336725
rect 483569 336685 483581 336719
rect 483615 336716 483627 336719
rect 489178 336716 489184 336728
rect 483615 336688 489184 336716
rect 483615 336685 483627 336688
rect 483569 336679 483627 336685
rect 489178 336676 489184 336688
rect 489236 336676 489242 336728
rect 273070 336648 273076 336660
rect 272812 336620 273076 336648
rect 273070 336608 273076 336620
rect 273128 336608 273134 336660
rect 280338 336608 280344 336660
rect 280396 336648 280402 336660
rect 293954 336648 293960 336660
rect 280396 336620 293960 336648
rect 280396 336608 280402 336620
rect 293954 336608 293960 336620
rect 294012 336608 294018 336660
rect 235813 336583 235871 336589
rect 235813 336549 235825 336583
rect 235859 336580 235871 336583
rect 240318 336580 240324 336592
rect 235859 336552 240324 336580
rect 235859 336549 235871 336552
rect 235813 336543 235871 336549
rect 240318 336540 240324 336552
rect 240376 336540 240382 336592
rect 274729 336583 274787 336589
rect 274729 336549 274741 336583
rect 274775 336580 274787 336583
rect 296714 336580 296720 336592
rect 274775 336552 296720 336580
rect 274775 336549 274787 336552
rect 274729 336543 274787 336549
rect 296714 336540 296720 336552
rect 296772 336540 296778 336592
rect 230474 336472 230480 336524
rect 230532 336512 230538 336524
rect 253566 336512 253572 336524
rect 230532 336484 253572 336512
rect 230532 336472 230538 336484
rect 253566 336472 253572 336484
rect 253624 336472 253630 336524
rect 260926 336472 260932 336524
rect 260984 336512 260990 336524
rect 289817 336515 289875 336521
rect 289817 336512 289829 336515
rect 260984 336484 289829 336512
rect 260984 336472 260990 336484
rect 289817 336481 289829 336484
rect 289863 336481 289875 336515
rect 289817 336475 289875 336481
rect 219342 336404 219348 336456
rect 219400 336444 219406 336456
rect 252462 336444 252468 336456
rect 219400 336416 252468 336444
rect 219400 336404 219406 336416
rect 252462 336404 252468 336416
rect 252520 336404 252526 336456
rect 262490 336404 262496 336456
rect 262548 336444 262554 336456
rect 314654 336444 314660 336456
rect 262548 336416 314660 336444
rect 262548 336404 262554 336416
rect 314654 336404 314660 336416
rect 314712 336404 314718 336456
rect 209682 336336 209688 336388
rect 209740 336376 209746 336388
rect 242894 336376 242900 336388
rect 209740 336348 242900 336376
rect 209740 336336 209746 336348
rect 242894 336336 242900 336348
rect 242952 336336 242958 336388
rect 268102 336336 268108 336388
rect 268160 336376 268166 336388
rect 331214 336376 331220 336388
rect 268160 336348 331220 336376
rect 268160 336336 268166 336348
rect 331214 336336 331220 336348
rect 331272 336336 331278 336388
rect 180702 336268 180708 336320
rect 180760 336308 180766 336320
rect 248414 336308 248420 336320
rect 180760 336280 248420 336308
rect 180760 336268 180766 336280
rect 248414 336268 248420 336280
rect 248472 336268 248478 336320
rect 262490 336308 262496 336320
rect 262451 336280 262496 336308
rect 262490 336268 262496 336280
rect 262548 336268 262554 336320
rect 265986 336268 265992 336320
rect 266044 336308 266050 336320
rect 349154 336308 349160 336320
rect 266044 336280 349160 336308
rect 266044 336268 266050 336280
rect 349154 336268 349160 336280
rect 349212 336268 349218 336320
rect 169662 336200 169668 336252
rect 169720 336240 169726 336252
rect 247310 336240 247316 336252
rect 169720 336212 247316 336240
rect 169720 336200 169726 336212
rect 247310 336200 247316 336212
rect 247368 336200 247374 336252
rect 275646 336200 275652 336252
rect 275704 336240 275710 336252
rect 443086 336240 443092 336252
rect 275704 336212 443092 336240
rect 275704 336200 275710 336212
rect 443086 336200 443092 336212
rect 443144 336200 443150 336252
rect 126882 336132 126888 336184
rect 126940 336172 126946 336184
rect 235813 336175 235871 336181
rect 235813 336172 235825 336175
rect 126940 336144 235825 336172
rect 126940 336132 126946 336144
rect 235813 336141 235825 336144
rect 235859 336141 235871 336175
rect 237190 336172 237196 336184
rect 235813 336135 235871 336141
rect 235920 336144 237196 336172
rect 71682 336064 71688 336116
rect 71740 336104 71746 336116
rect 235920 336104 235948 336144
rect 237190 336132 237196 336144
rect 237248 336132 237254 336184
rect 291194 336132 291200 336184
rect 291252 336172 291258 336184
rect 483014 336172 483020 336184
rect 291252 336144 483020 336172
rect 291252 336132 291258 336144
rect 483014 336132 483020 336144
rect 483072 336132 483078 336184
rect 71740 336076 235948 336104
rect 71740 336064 71746 336076
rect 236546 336064 236552 336116
rect 236604 336104 236610 336116
rect 236914 336104 236920 336116
rect 236604 336076 236920 336104
rect 236604 336064 236610 336076
rect 236914 336064 236920 336076
rect 236972 336064 236978 336116
rect 284110 336064 284116 336116
rect 284168 336104 284174 336116
rect 521654 336104 521660 336116
rect 284168 336076 521660 336104
rect 284168 336064 284174 336076
rect 521654 336064 521660 336076
rect 521712 336064 521718 336116
rect 48222 335996 48228 336048
rect 48280 336036 48286 336048
rect 233602 336036 233608 336048
rect 48280 336008 233608 336036
rect 48280 335996 48286 336008
rect 233602 335996 233608 336008
rect 233660 335996 233666 336048
rect 287790 335996 287796 336048
rect 287848 336036 287854 336048
rect 557534 336036 557540 336048
rect 287848 336008 557540 336036
rect 287848 335996 287854 336008
rect 557534 335996 557540 336008
rect 557592 335996 557598 336048
rect 233234 335928 233240 335980
rect 233292 335968 233298 335980
rect 234154 335968 234160 335980
rect 233292 335940 234160 335968
rect 233292 335928 233298 335940
rect 234154 335928 234160 335940
rect 234212 335928 234218 335980
rect 251726 335968 251732 335980
rect 251687 335940 251732 335968
rect 251726 335928 251732 335940
rect 251784 335928 251790 335980
rect 289817 335971 289875 335977
rect 289817 335937 289829 335971
rect 289863 335968 289875 335971
rect 300854 335968 300860 335980
rect 289863 335940 300860 335968
rect 289863 335937 289875 335940
rect 289817 335931 289875 335937
rect 300854 335928 300860 335940
rect 300912 335928 300918 335980
rect 232222 335860 232228 335912
rect 232280 335900 232286 335912
rect 232682 335900 232688 335912
rect 232280 335872 232688 335900
rect 232280 335860 232286 335872
rect 232682 335860 232688 335872
rect 232740 335860 232746 335912
rect 232038 335792 232044 335844
rect 232096 335832 232102 335844
rect 232774 335832 232780 335844
rect 232096 335804 232780 335832
rect 232096 335792 232102 335804
rect 232774 335792 232780 335804
rect 232832 335792 232838 335844
rect 233418 335792 233424 335844
rect 233476 335832 233482 335844
rect 234154 335832 234160 335844
rect 233476 335804 234160 335832
rect 233476 335792 233482 335804
rect 234154 335792 234160 335804
rect 234212 335792 234218 335844
rect 236454 335792 236460 335844
rect 236512 335832 236518 335844
rect 236638 335832 236644 335844
rect 236512 335804 236644 335832
rect 236512 335792 236518 335804
rect 236638 335792 236644 335804
rect 236696 335792 236702 335844
rect 242894 335792 242900 335844
rect 242952 335832 242958 335844
rect 243170 335832 243176 335844
rect 242952 335804 243176 335832
rect 242952 335792 242958 335804
rect 243170 335792 243176 335804
rect 243228 335792 243234 335844
rect 254118 335792 254124 335844
rect 254176 335832 254182 335844
rect 254486 335832 254492 335844
rect 254176 335804 254492 335832
rect 254176 335792 254182 335804
rect 254486 335792 254492 335804
rect 254544 335792 254550 335844
rect 232498 335724 232504 335776
rect 232556 335764 232562 335776
rect 232958 335764 232964 335776
rect 232556 335736 232964 335764
rect 232556 335724 232562 335736
rect 232958 335724 232964 335736
rect 233016 335724 233022 335776
rect 248874 335724 248880 335776
rect 248932 335724 248938 335776
rect 254673 335767 254731 335773
rect 254673 335733 254685 335767
rect 254719 335764 254731 335767
rect 255774 335764 255780 335776
rect 254719 335736 255780 335764
rect 254719 335733 254731 335736
rect 254673 335727 254731 335733
rect 255774 335724 255780 335736
rect 255832 335724 255838 335776
rect 258350 335724 258356 335776
rect 258408 335764 258414 335776
rect 258902 335764 258908 335776
rect 258408 335736 258908 335764
rect 258408 335724 258414 335736
rect 258902 335724 258908 335736
rect 258960 335724 258966 335776
rect 262582 335724 262588 335776
rect 262640 335764 262646 335776
rect 263410 335764 263416 335776
rect 262640 335736 263416 335764
rect 262640 335724 262646 335736
rect 263410 335724 263416 335736
rect 263468 335724 263474 335776
rect 232222 335656 232228 335708
rect 232280 335696 232286 335708
rect 232590 335696 232596 335708
rect 232280 335668 232596 335696
rect 232280 335656 232286 335668
rect 232590 335656 232596 335668
rect 232648 335656 232654 335708
rect 233418 335656 233424 335708
rect 233476 335696 233482 335708
rect 233694 335696 233700 335708
rect 233476 335668 233700 335696
rect 233476 335656 233482 335668
rect 233694 335656 233700 335668
rect 233752 335656 233758 335708
rect 234062 335656 234068 335708
rect 234120 335696 234126 335708
rect 234430 335696 234436 335708
rect 234120 335668 234436 335696
rect 234120 335656 234126 335668
rect 234430 335656 234436 335668
rect 234488 335656 234494 335708
rect 236086 335656 236092 335708
rect 236144 335656 236150 335708
rect 236362 335656 236368 335708
rect 236420 335696 236426 335708
rect 236420 335668 236592 335696
rect 236420 335656 236426 335668
rect 229186 335588 229192 335640
rect 229244 335628 229250 335640
rect 230198 335628 230204 335640
rect 229244 335600 230204 335628
rect 229244 335588 229250 335600
rect 230198 335588 230204 335600
rect 230256 335588 230262 335640
rect 230658 335588 230664 335640
rect 230716 335628 230722 335640
rect 231118 335628 231124 335640
rect 230716 335600 231124 335628
rect 230716 335588 230722 335600
rect 231118 335588 231124 335600
rect 231176 335588 231182 335640
rect 232314 335588 232320 335640
rect 232372 335628 232378 335640
rect 232774 335628 232780 335640
rect 232372 335600 232780 335628
rect 232372 335588 232378 335600
rect 232774 335588 232780 335600
rect 232832 335588 232838 335640
rect 234614 335588 234620 335640
rect 234672 335628 234678 335640
rect 235902 335628 235908 335640
rect 234672 335600 235908 335628
rect 234672 335588 234678 335600
rect 235902 335588 235908 335600
rect 235960 335588 235966 335640
rect 230566 335452 230572 335504
rect 230624 335492 230630 335504
rect 231118 335492 231124 335504
rect 230624 335464 231124 335492
rect 230624 335452 230630 335464
rect 231118 335452 231124 335464
rect 231176 335452 231182 335504
rect 229557 335427 229615 335433
rect 229557 335393 229569 335427
rect 229603 335424 229615 335427
rect 230290 335424 230296 335436
rect 229603 335396 230296 335424
rect 229603 335393 229615 335396
rect 229557 335387 229615 335393
rect 230290 335384 230296 335396
rect 230348 335384 230354 335436
rect 227622 335316 227628 335368
rect 227680 335356 227686 335368
rect 231946 335356 231952 335368
rect 227680 335328 231952 335356
rect 227680 335316 227686 335328
rect 231946 335316 231952 335328
rect 232004 335316 232010 335368
rect 236104 335220 236132 335656
rect 236564 335640 236592 335668
rect 237650 335656 237656 335708
rect 237708 335696 237714 335708
rect 238478 335696 238484 335708
rect 237708 335668 238484 335696
rect 237708 335656 237714 335668
rect 238478 335656 238484 335668
rect 238536 335656 238542 335708
rect 239122 335656 239128 335708
rect 239180 335696 239186 335708
rect 239950 335696 239956 335708
rect 239180 335668 239956 335696
rect 239180 335656 239186 335668
rect 239950 335656 239956 335668
rect 240008 335656 240014 335708
rect 240318 335656 240324 335708
rect 240376 335696 240382 335708
rect 240778 335696 240784 335708
rect 240376 335668 240784 335696
rect 240376 335656 240382 335668
rect 240778 335656 240784 335668
rect 240836 335656 240842 335708
rect 243170 335656 243176 335708
rect 243228 335696 243234 335708
rect 243814 335696 243820 335708
rect 243228 335668 243820 335696
rect 243228 335656 243234 335668
rect 243814 335656 243820 335668
rect 243872 335656 243878 335708
rect 244826 335656 244832 335708
rect 244884 335696 244890 335708
rect 245102 335696 245108 335708
rect 244884 335668 245108 335696
rect 244884 335656 244890 335668
rect 245102 335656 245108 335668
rect 245160 335656 245166 335708
rect 248782 335696 248788 335708
rect 248743 335668 248788 335696
rect 248782 335656 248788 335668
rect 248840 335656 248846 335708
rect 248892 335640 248920 335724
rect 255869 335699 255927 335705
rect 255869 335665 255881 335699
rect 255915 335696 255927 335699
rect 256050 335696 256056 335708
rect 255915 335668 256056 335696
rect 255915 335665 255927 335668
rect 255869 335659 255927 335665
rect 256050 335656 256056 335668
rect 256108 335656 256114 335708
rect 265437 335699 265495 335705
rect 265437 335665 265449 335699
rect 265483 335696 265495 335699
rect 266078 335696 266084 335708
rect 265483 335668 266084 335696
rect 265483 335665 265495 335668
rect 265437 335659 265495 335665
rect 266078 335656 266084 335668
rect 266136 335656 266142 335708
rect 266538 335656 266544 335708
rect 266596 335696 266602 335708
rect 267458 335696 267464 335708
rect 266596 335668 267464 335696
rect 266596 335656 266602 335668
rect 267458 335656 267464 335668
rect 267516 335656 267522 335708
rect 268010 335656 268016 335708
rect 268068 335656 268074 335708
rect 268562 335656 268568 335708
rect 268620 335696 268626 335708
rect 268930 335696 268936 335708
rect 268620 335668 268936 335696
rect 268620 335656 268626 335668
rect 268930 335656 268936 335668
rect 268988 335656 268994 335708
rect 276382 335656 276388 335708
rect 276440 335696 276446 335708
rect 277210 335696 277216 335708
rect 276440 335668 277216 335696
rect 276440 335656 276446 335668
rect 277210 335656 277216 335668
rect 277268 335656 277274 335708
rect 280338 335656 280344 335708
rect 280396 335696 280402 335708
rect 280706 335696 280712 335708
rect 280396 335668 280712 335696
rect 280396 335656 280402 335668
rect 280706 335656 280712 335668
rect 280764 335656 280770 335708
rect 280798 335656 280804 335708
rect 280856 335656 280862 335708
rect 284018 335656 284024 335708
rect 284076 335656 284082 335708
rect 286042 335656 286048 335708
rect 286100 335696 286106 335708
rect 286318 335696 286324 335708
rect 286100 335668 286324 335696
rect 286100 335656 286106 335668
rect 286318 335656 286324 335668
rect 286376 335656 286382 335708
rect 288621 335699 288679 335705
rect 288621 335665 288633 335699
rect 288667 335696 288679 335699
rect 289354 335696 289360 335708
rect 288667 335668 289360 335696
rect 288667 335665 288679 335668
rect 288621 335659 288679 335665
rect 289354 335656 289360 335668
rect 289412 335656 289418 335708
rect 236546 335588 236552 335640
rect 236604 335588 236610 335640
rect 236638 335588 236644 335640
rect 236696 335628 236702 335640
rect 237006 335628 237012 335640
rect 236696 335600 237012 335628
rect 236696 335588 236702 335600
rect 237006 335588 237012 335600
rect 237064 335588 237070 335640
rect 238110 335588 238116 335640
rect 238168 335628 238174 335640
rect 238386 335628 238392 335640
rect 238168 335600 238392 335628
rect 238168 335588 238174 335600
rect 238386 335588 238392 335600
rect 238444 335588 238450 335640
rect 239582 335588 239588 335640
rect 239640 335628 239646 335640
rect 239858 335628 239864 335640
rect 239640 335600 239864 335628
rect 239640 335588 239646 335600
rect 239858 335588 239864 335600
rect 239916 335588 239922 335640
rect 240686 335588 240692 335640
rect 240744 335628 240750 335640
rect 241054 335628 241060 335640
rect 240744 335600 241060 335628
rect 240744 335588 240750 335600
rect 241054 335588 241060 335600
rect 241112 335588 241118 335640
rect 242158 335588 242164 335640
rect 242216 335628 242222 335640
rect 242434 335628 242440 335640
rect 242216 335600 242440 335628
rect 242216 335588 242222 335600
rect 242434 335588 242440 335600
rect 242492 335588 242498 335640
rect 242526 335588 242532 335640
rect 242584 335628 242590 335640
rect 242710 335628 242716 335640
rect 242584 335600 242716 335628
rect 242584 335588 242590 335600
rect 242710 335588 242716 335600
rect 242768 335588 242774 335640
rect 243262 335588 243268 335640
rect 243320 335628 243326 335640
rect 243446 335628 243452 335640
rect 243320 335600 243452 335628
rect 243320 335588 243326 335600
rect 243446 335588 243452 335600
rect 243504 335588 243510 335640
rect 244918 335588 244924 335640
rect 244976 335628 244982 335640
rect 245562 335628 245568 335640
rect 244976 335600 245568 335628
rect 244976 335588 244982 335600
rect 245562 335588 245568 335600
rect 245620 335588 245626 335640
rect 245930 335588 245936 335640
rect 245988 335628 245994 335640
rect 246850 335628 246856 335640
rect 245988 335600 246856 335628
rect 245988 335588 245994 335600
rect 246850 335588 246856 335600
rect 246908 335588 246914 335640
rect 247586 335588 247592 335640
rect 247644 335628 247650 335640
rect 247862 335628 247868 335640
rect 247644 335600 247868 335628
rect 247644 335588 247650 335600
rect 247862 335588 247868 335600
rect 247920 335588 247926 335640
rect 248874 335588 248880 335640
rect 248932 335588 248938 335640
rect 249242 335588 249248 335640
rect 249300 335628 249306 335640
rect 249610 335628 249616 335640
rect 249300 335600 249616 335628
rect 249300 335588 249306 335600
rect 249610 335588 249616 335600
rect 249668 335588 249674 335640
rect 250714 335588 250720 335640
rect 250772 335628 250778 335640
rect 251082 335628 251088 335640
rect 250772 335600 251088 335628
rect 250772 335588 250778 335600
rect 251082 335588 251088 335600
rect 251140 335588 251146 335640
rect 251174 335588 251180 335640
rect 251232 335628 251238 335640
rect 251542 335628 251548 335640
rect 251232 335600 251548 335628
rect 251232 335588 251238 335600
rect 251542 335588 251548 335600
rect 251600 335588 251606 335640
rect 252922 335588 252928 335640
rect 252980 335628 252986 335640
rect 253842 335628 253848 335640
rect 252980 335600 253848 335628
rect 252980 335588 252986 335600
rect 253842 335588 253848 335600
rect 253900 335588 253906 335640
rect 254302 335588 254308 335640
rect 254360 335628 254366 335640
rect 254670 335628 254676 335640
rect 254360 335600 254676 335628
rect 254360 335588 254366 335600
rect 254670 335588 254676 335600
rect 254728 335588 254734 335640
rect 239122 335520 239128 335572
rect 239180 335560 239186 335572
rect 240042 335560 240048 335572
rect 239180 335532 240048 335560
rect 239180 335520 239186 335532
rect 240042 335520 240048 335532
rect 240100 335520 240106 335572
rect 255866 335520 255872 335572
rect 255924 335520 255930 335572
rect 236270 335452 236276 335504
rect 236328 335492 236334 335504
rect 237282 335492 237288 335504
rect 236328 335464 237288 335492
rect 236328 335452 236334 335464
rect 237282 335452 237288 335464
rect 237340 335452 237346 335504
rect 248690 335452 248696 335504
rect 248748 335492 248754 335504
rect 249058 335492 249064 335504
rect 248748 335464 249064 335492
rect 248748 335452 248754 335464
rect 249058 335452 249064 335464
rect 249116 335452 249122 335504
rect 249794 335452 249800 335504
rect 249852 335492 249858 335504
rect 250254 335492 250260 335504
rect 249852 335464 250260 335492
rect 249852 335452 249858 335464
rect 250254 335452 250260 335464
rect 250312 335452 250318 335504
rect 251450 335452 251456 335504
rect 251508 335492 251514 335504
rect 251726 335492 251732 335504
rect 251508 335464 251732 335492
rect 251508 335452 251514 335464
rect 251726 335452 251732 335464
rect 251784 335452 251790 335504
rect 240042 335424 240048 335436
rect 240003 335396 240048 335424
rect 240042 335384 240048 335396
rect 240100 335384 240106 335436
rect 236178 335316 236184 335368
rect 236236 335356 236242 335368
rect 236822 335356 236828 335368
rect 236236 335328 236828 335356
rect 236236 335316 236242 335328
rect 236822 335316 236828 335328
rect 236880 335316 236886 335368
rect 251634 335248 251640 335300
rect 251692 335248 251698 335300
rect 236822 335220 236828 335232
rect 236104 335192 236828 335220
rect 236822 335180 236828 335192
rect 236880 335180 236886 335232
rect 235994 335112 236000 335164
rect 236052 335152 236058 335164
rect 236362 335152 236368 335164
rect 236052 335124 236368 335152
rect 236052 335112 236058 335124
rect 236362 335112 236368 335124
rect 236420 335112 236426 335164
rect 224862 335044 224868 335096
rect 224920 335084 224926 335096
rect 246942 335084 246948 335096
rect 224920 335056 246948 335084
rect 224920 335044 224926 335056
rect 246942 335044 246948 335056
rect 247000 335044 247006 335096
rect 251652 335084 251680 335248
rect 251726 335084 251732 335096
rect 251652 335056 251732 335084
rect 251726 335044 251732 335056
rect 251784 335044 251790 335096
rect 255498 335044 255504 335096
rect 255556 335084 255562 335096
rect 255884 335084 255912 335520
rect 268028 335504 268056 335656
rect 269482 335588 269488 335640
rect 269540 335628 269546 335640
rect 270310 335628 270316 335640
rect 269540 335600 270316 335628
rect 269540 335588 269546 335600
rect 270310 335588 270316 335600
rect 270368 335588 270374 335640
rect 272334 335588 272340 335640
rect 272392 335628 272398 335640
rect 272518 335628 272524 335640
rect 272392 335600 272524 335628
rect 272392 335588 272398 335600
rect 272518 335588 272524 335600
rect 272576 335588 272582 335640
rect 280816 335628 280844 335656
rect 280724 335600 280844 335628
rect 280724 335504 280752 335600
rect 284036 335560 284064 335656
rect 284036 335532 284248 335560
rect 284220 335504 284248 335532
rect 265710 335452 265716 335504
rect 265768 335492 265774 335504
rect 266078 335492 266084 335504
rect 265768 335464 266084 335492
rect 265768 335452 265774 335464
rect 266078 335452 266084 335464
rect 266136 335452 266142 335504
rect 268010 335452 268016 335504
rect 268068 335452 268074 335504
rect 268562 335452 268568 335504
rect 268620 335492 268626 335504
rect 268838 335492 268844 335504
rect 268620 335464 268844 335492
rect 268620 335452 268626 335464
rect 268838 335452 268844 335464
rect 268896 335452 268902 335504
rect 272518 335492 272524 335504
rect 272479 335464 272524 335492
rect 272518 335452 272524 335464
rect 272576 335452 272582 335504
rect 279050 335452 279056 335504
rect 279108 335492 279114 335504
rect 279602 335492 279608 335504
rect 279108 335464 279608 335492
rect 279108 335452 279114 335464
rect 279602 335452 279608 335464
rect 279660 335452 279666 335504
rect 280706 335452 280712 335504
rect 280764 335452 280770 335504
rect 283466 335452 283472 335504
rect 283524 335492 283530 335504
rect 284018 335492 284024 335504
rect 283524 335464 284024 335492
rect 283524 335452 283530 335464
rect 284018 335452 284024 335464
rect 284076 335452 284082 335504
rect 284202 335452 284208 335504
rect 284260 335452 284266 335504
rect 288618 335452 288624 335504
rect 288676 335492 288682 335504
rect 289262 335492 289268 335504
rect 288676 335464 289268 335492
rect 288676 335452 288682 335464
rect 289262 335452 289268 335464
rect 289320 335452 289326 335504
rect 277026 335424 277032 335436
rect 276987 335396 277032 335424
rect 277026 335384 277032 335396
rect 277084 335384 277090 335436
rect 278958 335384 278964 335436
rect 279016 335424 279022 335436
rect 279510 335424 279516 335436
rect 279016 335396 279516 335424
rect 279016 335384 279022 335396
rect 279510 335384 279516 335396
rect 279568 335384 279574 335436
rect 283558 335384 283564 335436
rect 283616 335424 283622 335436
rect 284110 335424 284116 335436
rect 283616 335396 284116 335424
rect 283616 335384 283622 335396
rect 284110 335384 284116 335396
rect 284168 335384 284174 335436
rect 265158 335356 265164 335368
rect 265119 335328 265164 335356
rect 265158 335316 265164 335328
rect 265216 335316 265222 335368
rect 265434 335316 265440 335368
rect 265492 335356 265498 335368
rect 265526 335356 265532 335368
rect 265492 335328 265532 335356
rect 265492 335316 265498 335328
rect 265526 335316 265532 335328
rect 265584 335316 265590 335368
rect 266354 335316 266360 335368
rect 266412 335356 266418 335368
rect 266998 335356 267004 335368
rect 266412 335328 267004 335356
rect 266412 335316 266418 335328
rect 266998 335316 267004 335328
rect 267056 335316 267062 335368
rect 277305 335359 277363 335365
rect 277305 335325 277317 335359
rect 277351 335356 277363 335359
rect 280338 335356 280344 335368
rect 277351 335328 280344 335356
rect 277351 335325 277363 335328
rect 277305 335319 277363 335325
rect 280338 335316 280344 335328
rect 280396 335316 280402 335368
rect 280522 335356 280528 335368
rect 280483 335328 280528 335356
rect 280522 335316 280528 335328
rect 280580 335316 280586 335368
rect 282914 335316 282920 335368
rect 282972 335356 282978 335368
rect 283282 335356 283288 335368
rect 282972 335328 283288 335356
rect 282972 335316 282978 335328
rect 283282 335316 283288 335328
rect 283340 335316 283346 335368
rect 286134 335316 286140 335368
rect 286192 335356 286198 335368
rect 286870 335356 286876 335368
rect 286192 335328 286876 335356
rect 286192 335316 286198 335328
rect 286870 335316 286876 335328
rect 286928 335316 286934 335368
rect 278774 335180 278780 335232
rect 278832 335220 278838 335232
rect 279142 335220 279148 335232
rect 278832 335192 279148 335220
rect 278832 335180 278838 335192
rect 279142 335180 279148 335192
rect 279200 335180 279206 335232
rect 280985 335223 281043 335229
rect 280985 335189 280997 335223
rect 281031 335220 281043 335223
rect 283466 335220 283472 335232
rect 281031 335192 283472 335220
rect 281031 335189 281043 335192
rect 280985 335183 281043 335189
rect 283466 335180 283472 335192
rect 283524 335180 283530 335232
rect 281074 335112 281080 335164
rect 281132 335152 281138 335164
rect 304994 335152 305000 335164
rect 281132 335124 305000 335152
rect 281132 335112 281138 335124
rect 304994 335112 305000 335124
rect 305052 335112 305058 335164
rect 255556 335056 255912 335084
rect 255556 335044 255562 335056
rect 260742 335044 260748 335096
rect 260800 335084 260806 335096
rect 292574 335084 292580 335096
rect 260800 335056 292580 335084
rect 260800 335044 260806 335056
rect 292574 335044 292580 335056
rect 292632 335044 292638 335096
rect 223482 334976 223488 335028
rect 223540 335016 223546 335028
rect 252830 335016 252836 335028
rect 223540 334988 252836 335016
rect 223540 334976 223546 334988
rect 252830 334976 252836 334988
rect 252888 334976 252894 335028
rect 262030 334976 262036 335028
rect 262088 335016 262094 335028
rect 311894 335016 311900 335028
rect 262088 334988 311900 335016
rect 262088 334976 262094 334988
rect 311894 334976 311900 334988
rect 311952 334976 311958 335028
rect 212442 334908 212448 334960
rect 212500 334948 212506 334960
rect 251729 334951 251787 334957
rect 251729 334948 251741 334951
rect 212500 334920 251741 334948
rect 212500 334908 212506 334920
rect 251729 334917 251741 334920
rect 251775 334917 251787 334951
rect 251729 334911 251787 334917
rect 265894 334908 265900 334960
rect 265952 334948 265958 334960
rect 327074 334948 327080 334960
rect 265952 334920 327080 334948
rect 265952 334908 265958 334920
rect 327074 334908 327080 334920
rect 327132 334908 327138 334960
rect 176562 334840 176568 334892
rect 176620 334880 176626 334892
rect 248046 334880 248052 334892
rect 176620 334852 248052 334880
rect 176620 334840 176626 334852
rect 248046 334840 248052 334852
rect 248104 334840 248110 334892
rect 266817 334883 266875 334889
rect 266817 334849 266829 334883
rect 266863 334880 266875 334883
rect 353294 334880 353300 334892
rect 266863 334852 353300 334880
rect 266863 334849 266875 334852
rect 266817 334843 266875 334849
rect 353294 334840 353300 334852
rect 353352 334840 353358 334892
rect 162762 334772 162768 334824
rect 162820 334812 162826 334824
rect 240226 334812 240232 334824
rect 162820 334784 240232 334812
rect 162820 334772 162826 334784
rect 240226 334772 240232 334784
rect 240284 334772 240290 334824
rect 273254 334772 273260 334824
rect 273312 334812 273318 334824
rect 422294 334812 422300 334824
rect 273312 334784 422300 334812
rect 273312 334772 273318 334784
rect 422294 334772 422300 334784
rect 422352 334772 422358 334824
rect 160002 334704 160008 334756
rect 160060 334744 160066 334756
rect 242986 334744 242992 334756
rect 160060 334716 242992 334744
rect 160060 334704 160066 334716
rect 242986 334704 242992 334716
rect 243044 334704 243050 334756
rect 290093 334747 290151 334753
rect 290093 334713 290105 334747
rect 290139 334744 290151 334747
rect 500954 334744 500960 334756
rect 290139 334716 500960 334744
rect 290139 334713 290151 334716
rect 290093 334707 290151 334713
rect 500954 334704 500960 334716
rect 501012 334704 501018 334756
rect 74442 334636 74448 334688
rect 74500 334676 74506 334688
rect 237558 334676 237564 334688
rect 74500 334648 237564 334676
rect 74500 334636 74506 334648
rect 237558 334636 237564 334648
rect 237616 334636 237622 334688
rect 256878 334636 256884 334688
rect 256936 334676 256942 334688
rect 257154 334676 257160 334688
rect 256936 334648 257160 334676
rect 256936 334636 256942 334648
rect 257154 334636 257160 334648
rect 257212 334636 257218 334688
rect 285490 334636 285496 334688
rect 285548 334676 285554 334688
rect 532694 334676 532700 334688
rect 285548 334648 532700 334676
rect 285548 334636 285554 334648
rect 532694 334636 532700 334648
rect 532752 334636 532758 334688
rect 52362 334568 52368 334620
rect 52420 334608 52426 334620
rect 231854 334608 231860 334620
rect 52420 334580 231860 334608
rect 52420 334568 52426 334580
rect 231854 334568 231860 334580
rect 231912 334568 231918 334620
rect 240226 334568 240232 334620
rect 240284 334608 240290 334620
rect 240502 334608 240508 334620
rect 240284 334580 240508 334608
rect 240284 334568 240290 334580
rect 240502 334568 240508 334580
rect 240560 334568 240566 334620
rect 262214 334568 262220 334620
rect 262272 334608 262278 334620
rect 287054 334608 287060 334620
rect 262272 334580 287060 334608
rect 262272 334568 262278 334580
rect 287054 334568 287060 334580
rect 287112 334568 287118 334620
rect 289630 334568 289636 334620
rect 289688 334608 289694 334620
rect 573358 334608 573364 334620
rect 289688 334580 573364 334608
rect 289688 334568 289694 334580
rect 573358 334568 573364 334580
rect 573416 334568 573422 334620
rect 240686 334364 240692 334416
rect 240744 334404 240750 334416
rect 241238 334404 241244 334416
rect 240744 334376 241244 334404
rect 240744 334364 240750 334376
rect 241238 334364 241244 334376
rect 241296 334364 241302 334416
rect 233326 334296 233332 334348
rect 233384 334336 233390 334348
rect 233973 334339 234031 334345
rect 233973 334336 233985 334339
rect 233384 334308 233985 334336
rect 233384 334296 233390 334308
rect 233973 334305 233985 334308
rect 234019 334305 234031 334339
rect 233973 334299 234031 334305
rect 245746 334092 245752 334144
rect 245804 334132 245810 334144
rect 246206 334132 246212 334144
rect 245804 334104 246212 334132
rect 245804 334092 245810 334104
rect 246206 334092 246212 334104
rect 246264 334092 246270 334144
rect 270770 334092 270776 334144
rect 270828 334132 270834 334144
rect 271782 334132 271788 334144
rect 270828 334104 271788 334132
rect 270828 334092 270834 334104
rect 271782 334092 271788 334104
rect 271840 334092 271846 334144
rect 276290 334092 276296 334144
rect 276348 334132 276354 334144
rect 276474 334132 276480 334144
rect 276348 334104 276480 334132
rect 276348 334092 276354 334104
rect 276474 334092 276480 334104
rect 276532 334092 276538 334144
rect 251910 333956 251916 334008
rect 251968 333996 251974 334008
rect 252370 333996 252376 334008
rect 251968 333968 252376 333996
rect 251968 333956 251974 333968
rect 252370 333956 252376 333968
rect 252428 333956 252434 334008
rect 278777 333999 278835 334005
rect 278777 333965 278789 333999
rect 278823 333996 278835 333999
rect 288345 333999 288403 334005
rect 288345 333996 288357 333999
rect 278823 333968 288357 333996
rect 278823 333965 278835 333968
rect 278777 333959 278835 333965
rect 288345 333965 288357 333968
rect 288391 333965 288403 333999
rect 288345 333959 288403 333965
rect 298097 333999 298155 334005
rect 298097 333965 298109 333999
rect 298143 333996 298155 333999
rect 307665 333999 307723 334005
rect 307665 333996 307677 333999
rect 298143 333968 307677 333996
rect 298143 333965 298155 333968
rect 298097 333959 298155 333965
rect 307665 333965 307677 333968
rect 307711 333965 307723 333999
rect 307665 333959 307723 333965
rect 254857 333931 254915 333937
rect 254857 333897 254869 333931
rect 254903 333928 254915 333931
rect 254946 333928 254952 333940
rect 254903 333900 254952 333928
rect 254903 333897 254915 333900
rect 254857 333891 254915 333897
rect 254946 333888 254952 333900
rect 255004 333888 255010 333940
rect 233602 333820 233608 333872
rect 233660 333860 233666 333872
rect 234062 333860 234068 333872
rect 233660 333832 234068 333860
rect 233660 333820 233666 333832
rect 234062 333820 234068 333832
rect 234120 333820 234126 333872
rect 307665 333863 307723 333869
rect 307665 333829 307677 333863
rect 307711 333829 307723 333863
rect 307665 333823 307723 333829
rect 241514 333752 241520 333804
rect 241572 333792 241578 333804
rect 241882 333792 241888 333804
rect 241572 333764 241888 333792
rect 241572 333752 241578 333764
rect 241882 333752 241888 333764
rect 241940 333752 241946 333804
rect 252646 333792 252652 333804
rect 247236 333764 252652 333792
rect 220722 333616 220728 333668
rect 220780 333656 220786 333668
rect 247236 333656 247264 333764
rect 252646 333752 252652 333764
rect 252704 333752 252710 333804
rect 261662 333752 261668 333804
rect 261720 333752 261726 333804
rect 288345 333795 288403 333801
rect 288345 333761 288357 333795
rect 288391 333761 288403 333795
rect 307680 333792 307708 333823
rect 307754 333792 307760 333804
rect 307680 333764 307760 333792
rect 288345 333755 288403 333761
rect 252462 333724 252468 333736
rect 220780 333628 247264 333656
rect 247328 333696 252468 333724
rect 220780 333616 220786 333628
rect 216582 333548 216588 333600
rect 216640 333588 216646 333600
rect 247328 333588 247356 333696
rect 252462 333684 252468 333696
rect 252520 333684 252526 333736
rect 261680 333724 261708 333752
rect 278777 333727 278835 333733
rect 278777 333724 278789 333727
rect 261680 333696 278789 333724
rect 278777 333693 278789 333696
rect 278823 333693 278835 333727
rect 288360 333724 288388 333755
rect 307754 333752 307760 333764
rect 307812 333752 307818 333804
rect 298097 333727 298155 333733
rect 298097 333724 298109 333727
rect 288360 333696 298109 333724
rect 278777 333687 278835 333693
rect 298097 333693 298109 333696
rect 298143 333693 298155 333727
rect 298097 333687 298155 333693
rect 247402 333616 247408 333668
rect 247460 333616 247466 333668
rect 262950 333616 262956 333668
rect 263008 333656 263014 333668
rect 280065 333659 280123 333665
rect 280065 333656 280077 333659
rect 263008 333628 280077 333656
rect 263008 333616 263014 333628
rect 280065 333625 280077 333628
rect 280111 333625 280123 333659
rect 280065 333619 280123 333625
rect 280341 333659 280399 333665
rect 280341 333625 280353 333659
rect 280387 333656 280399 333659
rect 299477 333659 299535 333665
rect 299477 333656 299489 333659
rect 280387 333628 299489 333656
rect 280387 333625 280399 333628
rect 280341 333619 280399 333625
rect 299477 333625 299489 333628
rect 299523 333625 299535 333659
rect 299477 333619 299535 333625
rect 299661 333659 299719 333665
rect 299661 333625 299673 333659
rect 299707 333656 299719 333659
rect 316034 333656 316040 333668
rect 299707 333628 316040 333656
rect 299707 333625 299719 333628
rect 299661 333619 299719 333625
rect 316034 333616 316040 333628
rect 316092 333616 316098 333668
rect 216640 333560 247356 333588
rect 216640 333548 216646 333560
rect 173802 333480 173808 333532
rect 173860 333520 173866 333532
rect 247420 333520 247448 333616
rect 261018 333548 261024 333600
rect 261076 333588 261082 333600
rect 261570 333588 261576 333600
rect 261076 333560 261576 333588
rect 261076 333548 261082 333560
rect 261570 333548 261576 333560
rect 261628 333548 261634 333600
rect 264698 333548 264704 333600
rect 264756 333588 264762 333600
rect 280249 333591 280307 333597
rect 280249 333588 280261 333591
rect 264756 333560 280261 333588
rect 264756 333548 264762 333560
rect 280249 333557 280261 333560
rect 280295 333557 280307 333591
rect 280249 333551 280307 333557
rect 280433 333591 280491 333597
rect 280433 333557 280445 333591
rect 280479 333588 280491 333591
rect 338114 333588 338120 333600
rect 280479 333560 338120 333588
rect 280479 333557 280491 333560
rect 280433 333551 280491 333557
rect 338114 333548 338120 333560
rect 338172 333548 338178 333600
rect 173860 333492 247448 333520
rect 173860 333480 173866 333492
rect 254026 333480 254032 333532
rect 254084 333520 254090 333532
rect 254210 333520 254216 333532
rect 254084 333492 254216 333520
rect 254084 333480 254090 333492
rect 254210 333480 254216 333492
rect 254268 333480 254274 333532
rect 268930 333480 268936 333532
rect 268988 333520 268994 333532
rect 373994 333520 374000 333532
rect 268988 333492 374000 333520
rect 268988 333480 268994 333492
rect 373994 333480 374000 333492
rect 374052 333480 374058 333532
rect 142062 333412 142068 333464
rect 142120 333452 142126 333464
rect 244458 333452 244464 333464
rect 142120 333424 244464 333452
rect 142120 333412 142126 333424
rect 244458 333412 244464 333424
rect 244516 333412 244522 333464
rect 247310 333412 247316 333464
rect 247368 333452 247374 333464
rect 247954 333452 247960 333464
rect 247368 333424 247960 333452
rect 247368 333412 247374 333424
rect 247954 333412 247960 333424
rect 248012 333412 248018 333464
rect 262490 333412 262496 333464
rect 262548 333452 262554 333464
rect 262858 333452 262864 333464
rect 262548 333424 262864 333452
rect 262548 333412 262554 333424
rect 262858 333412 262864 333424
rect 262916 333412 262922 333464
rect 271230 333412 271236 333464
rect 271288 333452 271294 333464
rect 400306 333452 400312 333464
rect 271288 333424 400312 333452
rect 271288 333412 271294 333424
rect 400306 333412 400312 333424
rect 400364 333412 400370 333464
rect 129642 333344 129648 333396
rect 129700 333384 129706 333396
rect 242894 333384 242900 333396
rect 129700 333356 242900 333384
rect 129700 333344 129706 333356
rect 242894 333344 242900 333356
rect 242952 333344 242958 333396
rect 247402 333344 247408 333396
rect 247460 333384 247466 333396
rect 248322 333384 248328 333396
rect 247460 333356 248328 333384
rect 247460 333344 247466 333356
rect 248322 333344 248328 333356
rect 248380 333344 248386 333396
rect 259822 333344 259828 333396
rect 259880 333384 259886 333396
rect 260190 333384 260196 333396
rect 259880 333356 260196 333384
rect 259880 333344 259886 333356
rect 260190 333344 260196 333356
rect 260248 333344 260254 333396
rect 275554 333344 275560 333396
rect 275612 333384 275618 333396
rect 440234 333384 440240 333396
rect 275612 333356 440240 333384
rect 275612 333344 275618 333356
rect 440234 333344 440240 333356
rect 440292 333344 440298 333396
rect 92382 333276 92388 333328
rect 92440 333316 92446 333328
rect 239398 333316 239404 333328
rect 92440 333288 239404 333316
rect 92440 333276 92446 333288
rect 239398 333276 239404 333288
rect 239456 333276 239462 333328
rect 250530 333316 250536 333328
rect 250491 333288 250536 333316
rect 250530 333276 250536 333288
rect 250588 333276 250594 333328
rect 261294 333276 261300 333328
rect 261352 333316 261358 333328
rect 261754 333316 261760 333328
rect 261352 333288 261760 333316
rect 261352 333276 261358 333288
rect 261754 333276 261760 333288
rect 261812 333276 261818 333328
rect 271874 333276 271880 333328
rect 271932 333316 271938 333328
rect 272242 333316 272248 333328
rect 271932 333288 272248 333316
rect 271932 333276 271938 333288
rect 272242 333276 272248 333288
rect 272300 333276 272306 333328
rect 276106 333276 276112 333328
rect 276164 333316 276170 333328
rect 276566 333316 276572 333328
rect 276164 333288 276572 333316
rect 276164 333276 276170 333288
rect 276566 333276 276572 333288
rect 276624 333276 276630 333328
rect 277854 333276 277860 333328
rect 277912 333316 277918 333328
rect 278498 333316 278504 333328
rect 277912 333288 278504 333316
rect 277912 333276 277918 333288
rect 278498 333276 278504 333288
rect 278556 333276 278562 333328
rect 284202 333276 284208 333328
rect 284260 333316 284266 333328
rect 518894 333316 518900 333328
rect 284260 333288 518900 333316
rect 284260 333276 284266 333288
rect 518894 333276 518900 333288
rect 518952 333276 518958 333328
rect 56502 333208 56508 333260
rect 56560 333248 56566 333260
rect 235626 333248 235632 333260
rect 56560 333220 235632 333248
rect 56560 333208 56566 333220
rect 235626 333208 235632 333220
rect 235684 333208 235690 333260
rect 286962 333208 286968 333260
rect 287020 333248 287026 333260
rect 546494 333248 546500 333260
rect 287020 333220 546500 333248
rect 287020 333208 287026 333220
rect 546494 333208 546500 333220
rect 546552 333208 546558 333260
rect 274818 333004 274824 333056
rect 274876 333044 274882 333056
rect 275738 333044 275744 333056
rect 274876 333016 275744 333044
rect 274876 333004 274882 333016
rect 275738 333004 275744 333016
rect 275796 333004 275802 333056
rect 261202 332936 261208 332988
rect 261260 332976 261266 332988
rect 261386 332976 261392 332988
rect 261260 332948 261392 332976
rect 261260 332936 261266 332948
rect 261386 332936 261392 332948
rect 261444 332936 261450 332988
rect 231486 332596 231492 332648
rect 231544 332636 231550 332648
rect 231762 332636 231768 332648
rect 231544 332608 231768 332636
rect 231544 332596 231550 332608
rect 231762 332596 231768 332608
rect 231820 332596 231826 332648
rect 244366 332596 244372 332648
rect 244424 332636 244430 332648
rect 245470 332636 245476 332648
rect 244424 332608 245476 332636
rect 244424 332596 244430 332608
rect 245470 332596 245476 332608
rect 245528 332596 245534 332648
rect 264790 332392 264796 332444
rect 264848 332432 264854 332444
rect 271877 332435 271935 332441
rect 271877 332432 271889 332435
rect 264848 332404 271889 332432
rect 264848 332392 264854 332404
rect 271877 332401 271889 332404
rect 271923 332401 271935 332435
rect 271877 332395 271935 332401
rect 260466 332324 260472 332376
rect 260524 332364 260530 332376
rect 296806 332364 296812 332376
rect 260524 332336 296812 332364
rect 260524 332324 260530 332336
rect 296806 332324 296812 332336
rect 296864 332324 296870 332376
rect 267461 332299 267519 332305
rect 267461 332265 267473 332299
rect 267507 332296 267519 332299
rect 267507 332268 271828 332296
rect 267507 332265 267519 332268
rect 267461 332259 267519 332265
rect 211062 332188 211068 332240
rect 211120 332228 211126 332240
rect 251358 332228 251364 332240
rect 211120 332200 251364 332228
rect 211120 332188 211126 332200
rect 251358 332188 251364 332200
rect 251416 332188 251422 332240
rect 270862 332188 270868 332240
rect 270920 332228 270926 332240
rect 271322 332228 271328 332240
rect 270920 332200 271328 332228
rect 270920 332188 270926 332200
rect 271322 332188 271328 332200
rect 271380 332188 271386 332240
rect 184842 332120 184848 332172
rect 184900 332160 184906 332172
rect 248785 332163 248843 332169
rect 248785 332160 248797 332163
rect 184900 332132 248797 332160
rect 184900 332120 184906 332132
rect 248785 332129 248797 332132
rect 248831 332129 248843 332163
rect 248785 332123 248843 332129
rect 270954 332120 270960 332172
rect 271012 332160 271018 332172
rect 271690 332160 271696 332172
rect 271012 332132 271696 332160
rect 271012 332120 271018 332132
rect 271690 332120 271696 332132
rect 271748 332120 271754 332172
rect 271800 332160 271828 332268
rect 281166 332256 281172 332308
rect 281224 332296 281230 332308
rect 318794 332296 318800 332308
rect 281224 332268 318800 332296
rect 281224 332256 281230 332268
rect 318794 332256 318800 332268
rect 318852 332256 318858 332308
rect 271877 332231 271935 332237
rect 271877 332197 271889 332231
rect 271923 332228 271935 332231
rect 333974 332228 333980 332240
rect 271923 332200 333980 332228
rect 271923 332197 271935 332200
rect 271877 332191 271935 332197
rect 333974 332188 333980 332200
rect 334032 332188 334038 332240
rect 356054 332160 356060 332172
rect 271800 332132 356060 332160
rect 356054 332120 356060 332132
rect 356112 332120 356118 332172
rect 153102 332052 153108 332104
rect 153160 332092 153166 332104
rect 245654 332092 245660 332104
rect 153160 332064 245660 332092
rect 153160 332052 153166 332064
rect 245654 332052 245660 332064
rect 245712 332052 245718 332104
rect 271598 332052 271604 332104
rect 271656 332092 271662 332104
rect 404354 332092 404360 332104
rect 271656 332064 404360 332092
rect 271656 332052 271662 332064
rect 404354 332052 404360 332064
rect 404412 332052 404418 332104
rect 144822 331984 144828 332036
rect 144880 332024 144886 332036
rect 245102 332024 245108 332036
rect 144880 331996 245108 332024
rect 144880 331984 144886 331996
rect 245102 331984 245108 331996
rect 245160 331984 245166 332036
rect 266446 331984 266452 332036
rect 266504 332024 266510 332036
rect 266722 332024 266728 332036
rect 266504 331996 266728 332024
rect 266504 331984 266510 331996
rect 266722 331984 266728 331996
rect 266780 331984 266786 332036
rect 278222 331984 278228 332036
rect 278280 332024 278286 332036
rect 467834 332024 467840 332036
rect 278280 331996 467840 332024
rect 278280 331984 278286 331996
rect 467834 331984 467840 331996
rect 467892 331984 467898 332036
rect 89622 331916 89628 331968
rect 89680 331956 89686 331968
rect 237098 331956 237104 331968
rect 89680 331928 237104 331956
rect 89680 331916 89686 331928
rect 237098 331916 237104 331928
rect 237156 331916 237162 331968
rect 285398 331916 285404 331968
rect 285456 331956 285462 331968
rect 528554 331956 528560 331968
rect 285456 331928 528560 331956
rect 285456 331916 285462 331928
rect 528554 331916 528560 331928
rect 528612 331916 528618 331968
rect 49602 331848 49608 331900
rect 49660 331888 49666 331900
rect 234982 331888 234988 331900
rect 49660 331860 234988 331888
rect 49660 331848 49666 331860
rect 234982 331848 234988 331860
rect 235040 331848 235046 331900
rect 289538 331848 289544 331900
rect 289596 331888 289602 331900
rect 574738 331888 574744 331900
rect 289596 331860 574744 331888
rect 289596 331848 289602 331860
rect 574738 331848 574744 331860
rect 574796 331848 574802 331900
rect 234062 331780 234068 331832
rect 234120 331820 234126 331832
rect 234338 331820 234344 331832
rect 234120 331792 234344 331820
rect 234120 331780 234126 331792
rect 234338 331780 234344 331792
rect 234396 331780 234402 331832
rect 234798 331644 234804 331696
rect 234856 331684 234862 331696
rect 235074 331684 235080 331696
rect 234856 331656 235080 331684
rect 234856 331644 234862 331656
rect 235074 331644 235080 331656
rect 235132 331644 235138 331696
rect 235534 331576 235540 331628
rect 235592 331616 235598 331628
rect 235810 331616 235816 331628
rect 235592 331588 235816 331616
rect 235592 331576 235598 331588
rect 235810 331576 235816 331588
rect 235868 331576 235874 331628
rect 262674 331304 262680 331356
rect 262732 331344 262738 331356
rect 275830 331344 275836 331356
rect 262732 331316 263272 331344
rect 262732 331304 262738 331316
rect 263244 331288 263272 331316
rect 275020 331316 275836 331344
rect 235718 331236 235724 331288
rect 235776 331236 235782 331288
rect 261938 331276 261944 331288
rect 260852 331248 261944 331276
rect 233510 331168 233516 331220
rect 233568 331208 233574 331220
rect 233694 331208 233700 331220
rect 233568 331180 233700 331208
rect 233568 331168 233574 331180
rect 233694 331168 233700 331180
rect 233752 331168 233758 331220
rect 235736 331152 235764 331236
rect 260852 331220 260880 331248
rect 261938 331236 261944 331248
rect 261996 331236 262002 331288
rect 263226 331236 263232 331288
rect 263284 331236 263290 331288
rect 275020 331220 275048 331316
rect 275830 331304 275836 331316
rect 275888 331304 275894 331356
rect 281718 331304 281724 331356
rect 281776 331304 281782 331356
rect 277302 331276 277308 331288
rect 277263 331248 277308 331276
rect 277302 331236 277308 331248
rect 277360 331236 277366 331288
rect 258258 331168 258264 331220
rect 258316 331208 258322 331220
rect 259362 331208 259368 331220
rect 258316 331180 259368 331208
rect 258316 331168 258322 331180
rect 259362 331168 259368 331180
rect 259420 331168 259426 331220
rect 260834 331168 260840 331220
rect 260892 331168 260898 331220
rect 275002 331168 275008 331220
rect 275060 331168 275066 331220
rect 235718 331100 235724 331152
rect 235776 331100 235782 331152
rect 281736 331140 281764 331304
rect 287422 331236 287428 331288
rect 287480 331276 287486 331288
rect 287480 331248 288020 331276
rect 287480 331236 287486 331248
rect 287992 331220 288020 331248
rect 287974 331168 287980 331220
rect 288032 331168 288038 331220
rect 284938 331140 284944 331152
rect 281736 331112 284944 331140
rect 284938 331100 284944 331112
rect 284996 331100 285002 331152
rect 287146 331100 287152 331152
rect 287204 331140 287210 331152
rect 287698 331140 287704 331152
rect 287204 331112 287704 331140
rect 287204 331100 287210 331112
rect 287698 331100 287704 331112
rect 287756 331100 287762 331152
rect 229002 330828 229008 330880
rect 229060 330868 229066 330880
rect 253290 330868 253296 330880
rect 229060 330840 253296 330868
rect 229060 330828 229066 330840
rect 253290 330828 253296 330840
rect 253348 330828 253354 330880
rect 262122 330828 262128 330880
rect 262180 330868 262186 330880
rect 313274 330868 313280 330880
rect 262180 330840 313280 330868
rect 262180 330828 262186 330840
rect 313274 330828 313280 330840
rect 313332 330828 313338 330880
rect 208302 330760 208308 330812
rect 208360 330800 208366 330812
rect 248414 330800 248420 330812
rect 208360 330772 248420 330800
rect 208360 330760 208366 330772
rect 248414 330760 248420 330772
rect 248472 330760 248478 330812
rect 270494 330760 270500 330812
rect 270552 330800 270558 330812
rect 393314 330800 393320 330812
rect 270552 330772 393320 330800
rect 270552 330760 270558 330772
rect 393314 330760 393320 330772
rect 393372 330760 393378 330812
rect 151722 330692 151728 330744
rect 151780 330732 151786 330744
rect 244366 330732 244372 330744
rect 151780 330704 244372 330732
rect 151780 330692 151786 330704
rect 244366 330692 244372 330704
rect 244424 330692 244430 330744
rect 272610 330692 272616 330744
rect 272668 330732 272674 330744
rect 411254 330732 411260 330744
rect 272668 330704 411260 330732
rect 272668 330692 272674 330704
rect 411254 330692 411260 330704
rect 411312 330692 411318 330744
rect 128262 330624 128268 330676
rect 128320 330664 128326 330676
rect 243078 330664 243084 330676
rect 128320 330636 243084 330664
rect 128320 330624 128326 330636
rect 243078 330624 243084 330636
rect 243136 330624 243142 330676
rect 277210 330624 277216 330676
rect 277268 330664 277274 330676
rect 451274 330664 451280 330676
rect 277268 330636 451280 330664
rect 277268 330624 277274 330636
rect 451274 330624 451280 330636
rect 451332 330624 451338 330676
rect 78582 330556 78588 330608
rect 78640 330596 78646 330608
rect 237926 330596 237932 330608
rect 78640 330568 237932 330596
rect 78640 330556 78646 330568
rect 237926 330556 237932 330568
rect 237984 330556 237990 330608
rect 278590 330556 278596 330608
rect 278648 330596 278654 330608
rect 462314 330596 462320 330608
rect 278648 330568 462320 330596
rect 278648 330556 278654 330568
rect 462314 330556 462320 330568
rect 462372 330556 462378 330608
rect 34422 330488 34428 330540
rect 34480 330528 34486 330540
rect 234154 330528 234160 330540
rect 34480 330500 234160 330528
rect 34480 330488 34486 330500
rect 234154 330488 234160 330500
rect 234212 330488 234218 330540
rect 285582 330488 285588 330540
rect 285640 330528 285646 330540
rect 536834 330528 536840 330540
rect 285640 330500 536840 330528
rect 285640 330488 285646 330500
rect 536834 330488 536840 330500
rect 536892 330488 536898 330540
rect 288618 329576 288624 329588
rect 288579 329548 288624 329576
rect 288618 329536 288624 329548
rect 288676 329536 288682 329588
rect 263502 329400 263508 329452
rect 263560 329440 263566 329452
rect 322934 329440 322940 329452
rect 263560 329412 322940 329440
rect 263560 329400 263566 329412
rect 322934 329400 322940 329412
rect 322992 329400 322998 329452
rect 206922 329332 206928 329384
rect 206980 329372 206986 329384
rect 251542 329372 251548 329384
rect 206980 329344 251548 329372
rect 206980 329332 206986 329344
rect 251542 329332 251548 329344
rect 251600 329332 251606 329384
rect 265618 329332 265624 329384
rect 265676 329372 265682 329384
rect 342254 329372 342260 329384
rect 265676 329344 342260 329372
rect 265676 329332 265682 329344
rect 342254 329332 342260 329344
rect 342312 329332 342318 329384
rect 157242 329264 157248 329316
rect 157300 329304 157306 329316
rect 246022 329304 246028 329316
rect 157300 329276 246028 329304
rect 157300 329264 157306 329276
rect 246022 329264 246028 329276
rect 246080 329264 246086 329316
rect 280338 329264 280344 329316
rect 280396 329304 280402 329316
rect 397454 329304 397460 329316
rect 280396 329276 397460 329304
rect 280396 329264 280402 329276
rect 397454 329264 397460 329276
rect 397512 329264 397518 329316
rect 155862 329196 155868 329248
rect 155920 329236 155926 329248
rect 244274 329236 244280 329248
rect 155920 329208 244280 329236
rect 155920 329196 155926 329208
rect 244274 329196 244280 329208
rect 244332 329196 244338 329248
rect 273346 329196 273352 329248
rect 273404 329236 273410 329248
rect 425146 329236 425152 329248
rect 273404 329208 425152 329236
rect 273404 329196 273410 329208
rect 425146 329196 425152 329208
rect 425204 329196 425210 329248
rect 85482 329128 85488 329180
rect 85540 329168 85546 329180
rect 238662 329168 238668 329180
rect 85540 329140 238668 329168
rect 85540 329128 85546 329140
rect 238662 329128 238668 329140
rect 238720 329128 238726 329180
rect 277394 329128 277400 329180
rect 277452 329168 277458 329180
rect 471974 329168 471980 329180
rect 277452 329140 471980 329168
rect 277452 329128 277458 329140
rect 471974 329128 471980 329140
rect 472032 329128 472038 329180
rect 38562 329060 38568 329112
rect 38620 329100 38626 329112
rect 233418 329100 233424 329112
rect 38620 329072 233424 329100
rect 38620 329060 38626 329072
rect 233418 329060 233424 329072
rect 233476 329060 233482 329112
rect 285585 329103 285643 329109
rect 285585 329069 285597 329103
rect 285631 329100 285643 329103
rect 539594 329100 539600 329112
rect 285631 329072 539600 329100
rect 285631 329069 285643 329072
rect 285585 329063 285643 329069
rect 539594 329060 539600 329072
rect 539652 329060 539658 329112
rect 251818 328992 251824 329044
rect 251876 329032 251882 329044
rect 254854 329032 254860 329044
rect 251876 329004 254860 329032
rect 251876 328992 251882 329004
rect 254854 328992 254860 329004
rect 254912 328992 254918 329044
rect 229554 328488 229560 328500
rect 229515 328460 229560 328488
rect 229554 328448 229560 328460
rect 229612 328448 229618 328500
rect 250533 328491 250591 328497
rect 250533 328457 250545 328491
rect 250579 328488 250591 328491
rect 250622 328488 250628 328500
rect 250579 328460 250628 328488
rect 250579 328457 250591 328460
rect 250533 328451 250591 328457
rect 250622 328448 250628 328460
rect 250680 328448 250686 328500
rect 252002 328448 252008 328500
rect 252060 328488 252066 328500
rect 253474 328488 253480 328500
rect 252060 328460 253480 328488
rect 252060 328448 252066 328460
rect 253474 328448 253480 328460
rect 253532 328448 253538 328500
rect 254670 328488 254676 328500
rect 254631 328460 254676 328488
rect 254670 328448 254676 328460
rect 254728 328448 254734 328500
rect 255866 328488 255872 328500
rect 255827 328460 255872 328488
rect 255866 328448 255872 328460
rect 255924 328448 255930 328500
rect 261754 328488 261760 328500
rect 261715 328460 261760 328488
rect 261754 328448 261760 328460
rect 261812 328448 261818 328500
rect 237006 328420 237012 328432
rect 236967 328392 237012 328420
rect 237006 328380 237012 328392
rect 237064 328380 237070 328432
rect 245197 328423 245255 328429
rect 245197 328389 245209 328423
rect 245243 328420 245255 328423
rect 245378 328420 245384 328432
rect 245243 328392 245384 328420
rect 245243 328389 245255 328392
rect 245197 328383 245255 328389
rect 245378 328380 245384 328392
rect 245436 328380 245442 328432
rect 257154 328380 257160 328432
rect 257212 328420 257218 328432
rect 257246 328420 257252 328432
rect 257212 328392 257252 328420
rect 257212 328380 257218 328392
rect 257246 328380 257252 328392
rect 257304 328380 257310 328432
rect 256418 328108 256424 328160
rect 256476 328148 256482 328160
rect 256694 328148 256700 328160
rect 256476 328120 256700 328148
rect 256476 328108 256482 328120
rect 256694 328108 256700 328120
rect 256752 328108 256758 328160
rect 260926 328108 260932 328160
rect 260984 328148 260990 328160
rect 299474 328148 299480 328160
rect 260984 328120 299480 328148
rect 260984 328108 260990 328120
rect 299474 328108 299480 328120
rect 299532 328108 299538 328160
rect 264422 328040 264428 328092
rect 264480 328080 264486 328092
rect 328454 328080 328460 328092
rect 264480 328052 328460 328080
rect 264480 328040 264486 328052
rect 328454 328040 328460 328052
rect 328512 328040 328518 328092
rect 215202 327972 215208 328024
rect 215260 328012 215266 328024
rect 251634 328012 251640 328024
rect 215260 327984 251640 328012
rect 215260 327972 215266 327984
rect 251634 327972 251640 327984
rect 251692 327972 251698 328024
rect 269298 327972 269304 328024
rect 269356 328012 269362 328024
rect 382274 328012 382280 328024
rect 269356 327984 382280 328012
rect 269356 327972 269362 327984
rect 382274 327972 382280 327984
rect 382332 327972 382338 328024
rect 168282 327904 168288 327956
rect 168340 327944 168346 327956
rect 247126 327944 247132 327956
rect 168340 327916 247132 327944
rect 168340 327904 168346 327916
rect 247126 327904 247132 327916
rect 247184 327904 247190 327956
rect 283282 327904 283288 327956
rect 283340 327944 283346 327956
rect 408494 327944 408500 327956
rect 283340 327916 408500 327944
rect 283340 327904 283346 327916
rect 408494 327904 408500 327916
rect 408552 327904 408558 327956
rect 139302 327836 139308 327888
rect 139360 327876 139366 327888
rect 244182 327876 244188 327888
rect 139360 327848 244188 327876
rect 139360 327836 139366 327848
rect 244182 327836 244188 327848
rect 244240 327836 244246 327888
rect 273622 327836 273628 327888
rect 273680 327876 273686 327888
rect 429194 327876 429200 327888
rect 273680 327848 429200 327876
rect 273680 327836 273686 327848
rect 429194 327836 429200 327848
rect 429252 327836 429258 327888
rect 96522 327768 96528 327820
rect 96580 327808 96586 327820
rect 239766 327808 239772 327820
rect 96580 327780 239772 327808
rect 96580 327768 96586 327780
rect 239766 327768 239772 327780
rect 239824 327768 239830 327820
rect 281902 327768 281908 327820
rect 281960 327808 281966 327820
rect 509234 327808 509240 327820
rect 281960 327780 509240 327808
rect 281960 327768 281966 327780
rect 509234 327768 509240 327780
rect 509292 327768 509298 327820
rect 53742 327700 53748 327752
rect 53800 327740 53806 327752
rect 235350 327740 235356 327752
rect 53800 327712 235356 327740
rect 53800 327700 53806 327712
rect 235350 327700 235356 327712
rect 235408 327700 235414 327752
rect 258994 327700 259000 327752
rect 259052 327740 259058 327752
rect 281534 327740 281540 327752
rect 259052 327712 281540 327740
rect 259052 327700 259058 327712
rect 281534 327700 281540 327712
rect 281592 327700 281598 327752
rect 286686 327700 286692 327752
rect 286744 327740 286750 327752
rect 550634 327740 550640 327752
rect 286744 327712 550640 327740
rect 286744 327700 286750 327712
rect 550634 327700 550640 327712
rect 550692 327700 550698 327752
rect 265434 327400 265440 327412
rect 265395 327372 265440 327400
rect 265434 327360 265440 327372
rect 265492 327360 265498 327412
rect 233970 327128 233976 327140
rect 233931 327100 233976 327128
rect 233970 327088 233976 327100
rect 234028 327088 234034 327140
rect 266262 327128 266268 327140
rect 266223 327100 266268 327128
rect 266262 327088 266268 327100
rect 266320 327088 266326 327140
rect 269022 327128 269028 327140
rect 268983 327100 269028 327128
rect 269022 327088 269028 327100
rect 269080 327088 269086 327140
rect 273162 327128 273168 327140
rect 273123 327100 273168 327128
rect 273162 327088 273168 327100
rect 273220 327088 273226 327140
rect 274358 327128 274364 327140
rect 274319 327100 274364 327128
rect 274358 327088 274364 327100
rect 274416 327088 274422 327140
rect 265158 327020 265164 327072
rect 265216 327060 265222 327072
rect 265250 327060 265256 327072
rect 265216 327032 265256 327060
rect 265216 327020 265222 327032
rect 265250 327020 265256 327032
rect 265308 327020 265314 327072
rect 265526 327020 265532 327072
rect 265584 327060 265590 327072
rect 265618 327060 265624 327072
rect 265584 327032 265624 327060
rect 265584 327020 265590 327032
rect 265618 327020 265624 327032
rect 265676 327020 265682 327072
rect 277026 327020 277032 327072
rect 277084 327060 277090 327072
rect 277118 327060 277124 327072
rect 277084 327032 277124 327060
rect 277084 327020 277090 327032
rect 277118 327020 277124 327032
rect 277176 327020 277182 327072
rect 263870 326952 263876 327004
rect 263928 326992 263934 327004
rect 264330 326992 264336 327004
rect 263928 326964 264336 326992
rect 263928 326952 263934 326964
rect 264330 326952 264336 326964
rect 264388 326952 264394 327004
rect 269574 326952 269580 327004
rect 269632 326952 269638 327004
rect 269482 326748 269488 326800
rect 269540 326788 269546 326800
rect 269592 326788 269620 326952
rect 269540 326760 269620 326788
rect 269540 326748 269546 326760
rect 274726 326748 274732 326800
rect 274784 326788 274790 326800
rect 279881 326791 279939 326797
rect 279881 326788 279893 326791
rect 274784 326760 279893 326788
rect 274784 326748 274790 326760
rect 279881 326757 279893 326760
rect 279927 326757 279939 326791
rect 279881 326751 279939 326757
rect 347774 326748 347780 326800
rect 347832 326788 347838 326800
rect 357345 326791 357403 326797
rect 357345 326788 357357 326791
rect 347832 326760 357357 326788
rect 347832 326748 347838 326760
rect 357345 326757 357357 326760
rect 357391 326757 357403 326791
rect 357345 326751 357403 326757
rect 263318 326680 263324 326732
rect 263376 326720 263382 326732
rect 320174 326720 320180 326732
rect 263376 326692 320180 326720
rect 263376 326680 263382 326692
rect 320174 326680 320180 326692
rect 320232 326680 320238 326732
rect 222102 326612 222108 326664
rect 222160 326652 222166 326664
rect 252738 326652 252744 326664
rect 222160 326624 252744 326652
rect 222160 326612 222166 326624
rect 252738 326612 252744 326624
rect 252796 326612 252802 326664
rect 266354 326612 266360 326664
rect 266412 326652 266418 326664
rect 360194 326652 360200 326664
rect 266412 326624 360200 326652
rect 266412 326612 266418 326624
rect 360194 326612 360200 326624
rect 360252 326612 360258 326664
rect 171042 326544 171048 326596
rect 171100 326584 171106 326596
rect 247586 326584 247592 326596
rect 171100 326556 247592 326584
rect 171100 326544 171106 326556
rect 247586 326544 247592 326556
rect 247644 326544 247650 326596
rect 273070 326544 273076 326596
rect 273128 326584 273134 326596
rect 309137 326587 309195 326593
rect 309137 326584 309149 326587
rect 273128 326556 309149 326584
rect 273128 326544 273134 326556
rect 309137 326553 309149 326556
rect 309183 326553 309195 326587
rect 309137 326547 309195 326553
rect 309413 326587 309471 326593
rect 309413 326553 309425 326587
rect 309459 326584 309471 326587
rect 415394 326584 415400 326596
rect 309459 326556 415400 326584
rect 309459 326553 309471 326556
rect 309413 326547 309471 326553
rect 415394 326544 415400 326556
rect 415452 326544 415458 326596
rect 159910 326476 159916 326528
rect 159968 326516 159974 326528
rect 246390 326516 246396 326528
rect 159968 326488 246396 326516
rect 159968 326476 159974 326488
rect 246390 326476 246396 326488
rect 246448 326476 246454 326528
rect 279786 326476 279792 326528
rect 279844 326476 279850 326528
rect 279881 326519 279939 326525
rect 279881 326485 279893 326519
rect 279927 326516 279939 326519
rect 289817 326519 289875 326525
rect 289817 326516 289829 326519
rect 279927 326488 289829 326516
rect 279927 326485 279939 326488
rect 279881 326479 279939 326485
rect 289817 326485 289829 326488
rect 289863 326485 289875 326519
rect 289817 326479 289875 326485
rect 290001 326519 290059 326525
rect 290001 326485 290013 326519
rect 290047 326516 290059 326519
rect 309229 326519 309287 326525
rect 309229 326516 309241 326519
rect 290047 326488 309241 326516
rect 290047 326485 290059 326488
rect 290001 326479 290059 326485
rect 309229 326485 309241 326488
rect 309275 326485 309287 326519
rect 309229 326479 309287 326485
rect 309321 326519 309379 326525
rect 309321 326485 309333 326519
rect 309367 326516 309379 326519
rect 433334 326516 433340 326528
rect 309367 326488 433340 326516
rect 309367 326485 309379 326488
rect 309321 326479 309379 326485
rect 433334 326476 433340 326488
rect 433392 326476 433398 326528
rect 56410 326408 56416 326460
rect 56468 326448 56474 326460
rect 235718 326448 235724 326460
rect 56468 326420 235724 326448
rect 56468 326408 56474 326420
rect 235718 326408 235724 326420
rect 235776 326408 235782 326460
rect 19978 326340 19984 326392
rect 20036 326380 20042 326392
rect 231486 326380 231492 326392
rect 20036 326352 231492 326380
rect 20036 326340 20042 326352
rect 231486 326340 231492 326352
rect 231544 326340 231550 326392
rect 251910 326340 251916 326392
rect 251968 326380 251974 326392
rect 252094 326380 252100 326392
rect 251968 326352 252100 326380
rect 251968 326340 251974 326352
rect 252094 326340 252100 326352
rect 252152 326340 252158 326392
rect 264054 326340 264060 326392
rect 264112 326380 264118 326392
rect 264238 326380 264244 326392
rect 264112 326352 264244 326380
rect 264112 326340 264118 326352
rect 264238 326340 264244 326352
rect 264296 326340 264302 326392
rect 266630 326340 266636 326392
rect 266688 326380 266694 326392
rect 266814 326380 266820 326392
rect 266688 326352 266820 326380
rect 266688 326340 266694 326352
rect 266814 326340 266820 326352
rect 266872 326340 266878 326392
rect 267366 326340 267372 326392
rect 267424 326380 267430 326392
rect 267642 326380 267648 326392
rect 267424 326352 267648 326380
rect 267424 326340 267430 326352
rect 267642 326340 267648 326352
rect 267700 326340 267706 326392
rect 267734 326340 267740 326392
rect 267792 326380 267798 326392
rect 267918 326380 267924 326392
rect 267792 326352 267924 326380
rect 267792 326340 267798 326352
rect 267918 326340 267924 326352
rect 267976 326340 267982 326392
rect 272150 326340 272156 326392
rect 272208 326380 272214 326392
rect 272978 326380 272984 326392
rect 272208 326352 272984 326380
rect 272208 326340 272214 326352
rect 272978 326340 272984 326352
rect 273036 326340 273042 326392
rect 279326 326340 279332 326392
rect 279384 326380 279390 326392
rect 279510 326380 279516 326392
rect 279384 326352 279516 326380
rect 279384 326340 279390 326352
rect 279510 326340 279516 326352
rect 279568 326340 279574 326392
rect 261662 326272 261668 326324
rect 261720 326272 261726 326324
rect 261680 326120 261708 326272
rect 279510 326204 279516 326256
rect 279568 326244 279574 326256
rect 279804 326244 279832 326476
rect 289725 326451 289783 326457
rect 289725 326417 289737 326451
rect 289771 326448 289783 326451
rect 299385 326451 299443 326457
rect 289771 326420 289860 326448
rect 289771 326417 289783 326420
rect 289725 326411 289783 326417
rect 282086 326340 282092 326392
rect 282144 326380 282150 326392
rect 282362 326380 282368 326392
rect 282144 326352 282368 326380
rect 282144 326340 282150 326352
rect 282362 326340 282368 326352
rect 282420 326340 282426 326392
rect 284754 326340 284760 326392
rect 284812 326380 284818 326392
rect 285030 326380 285036 326392
rect 284812 326352 285036 326380
rect 284812 326340 284818 326352
rect 285030 326340 285036 326352
rect 285088 326340 285094 326392
rect 287422 326340 287428 326392
rect 287480 326380 287486 326392
rect 287790 326380 287796 326392
rect 287480 326352 287796 326380
rect 287480 326340 287486 326352
rect 287790 326340 287796 326352
rect 287848 326340 287854 326392
rect 284386 326272 284392 326324
rect 284444 326312 284450 326324
rect 284846 326312 284852 326324
rect 284444 326284 284852 326312
rect 284444 326272 284450 326284
rect 284846 326272 284852 326284
rect 284904 326272 284910 326324
rect 287606 326272 287612 326324
rect 287664 326312 287670 326324
rect 288342 326312 288348 326324
rect 287664 326284 288348 326312
rect 287664 326272 287670 326284
rect 288342 326272 288348 326284
rect 288400 326272 288406 326324
rect 289832 326312 289860 326420
rect 299385 326417 299397 326451
rect 299431 326448 299443 326451
rect 299477 326451 299535 326457
rect 299477 326448 299489 326451
rect 299431 326420 299489 326448
rect 299431 326417 299443 326420
rect 299385 326411 299443 326417
rect 299477 326417 299489 326420
rect 299523 326417 299535 326451
rect 299477 326411 299535 326417
rect 308953 326451 309011 326457
rect 308953 326417 308965 326451
rect 308999 326448 309011 326451
rect 309137 326451 309195 326457
rect 309137 326448 309149 326451
rect 308999 326420 309149 326448
rect 308999 326417 309011 326420
rect 308953 326411 309011 326417
rect 309137 326417 309149 326420
rect 309183 326417 309195 326451
rect 309137 326411 309195 326417
rect 318705 326451 318763 326457
rect 318705 326417 318717 326451
rect 318751 326448 318763 326451
rect 318797 326451 318855 326457
rect 318797 326448 318809 326451
rect 318751 326420 318809 326448
rect 318751 326417 318763 326420
rect 318705 326411 318763 326417
rect 318797 326417 318809 326420
rect 318843 326417 318855 326451
rect 318797 326411 318855 326417
rect 328365 326451 328423 326457
rect 328365 326417 328377 326451
rect 328411 326448 328423 326451
rect 338117 326451 338175 326457
rect 338117 326448 338129 326451
rect 328411 326420 338129 326448
rect 328411 326417 328423 326420
rect 328365 326411 328423 326417
rect 338117 326417 338129 326420
rect 338163 326417 338175 326451
rect 338117 326411 338175 326417
rect 347593 326451 347651 326457
rect 347593 326417 347605 326451
rect 347639 326448 347651 326451
rect 347774 326448 347780 326460
rect 347639 326420 347780 326448
rect 347639 326417 347651 326420
rect 347593 326411 347651 326417
rect 347774 326408 347780 326420
rect 347832 326408 347838 326460
rect 357345 326451 357403 326457
rect 357345 326417 357357 326451
rect 357391 326448 357403 326451
rect 465074 326448 465080 326460
rect 357391 326420 465080 326448
rect 357391 326417 357403 326420
rect 357345 326411 357403 326417
rect 465074 326408 465080 326420
rect 465132 326408 465138 326460
rect 290826 326340 290832 326392
rect 290884 326380 290890 326392
rect 554774 326380 554780 326392
rect 290884 326352 554780 326380
rect 290884 326340 290890 326352
rect 554774 326340 554780 326352
rect 554832 326340 554838 326392
rect 299385 326315 299443 326321
rect 299385 326312 299397 326315
rect 289832 326284 299397 326312
rect 299385 326281 299397 326284
rect 299431 326281 299443 326315
rect 299385 326275 299443 326281
rect 309137 326315 309195 326321
rect 309137 326281 309149 326315
rect 309183 326312 309195 326315
rect 318705 326315 318763 326321
rect 318705 326312 318717 326315
rect 309183 326284 318717 326312
rect 309183 326281 309195 326284
rect 309137 326275 309195 326281
rect 318705 326281 318717 326284
rect 318751 326281 318763 326315
rect 318705 326275 318763 326281
rect 279568 326216 279832 326244
rect 299477 326247 299535 326253
rect 279568 326204 279574 326216
rect 299477 326213 299489 326247
rect 299523 326244 299535 326247
rect 308953 326247 309011 326253
rect 308953 326244 308965 326247
rect 299523 326216 308965 326244
rect 299523 326213 299535 326216
rect 299477 326207 299535 326213
rect 308953 326213 308965 326216
rect 308999 326213 309011 326247
rect 308953 326207 309011 326213
rect 318797 326247 318855 326253
rect 318797 326213 318809 326247
rect 318843 326244 318855 326247
rect 328365 326247 328423 326253
rect 328365 326244 328377 326247
rect 318843 326216 328377 326244
rect 318843 326213 318855 326216
rect 318797 326207 318855 326213
rect 328365 326213 328377 326216
rect 328411 326213 328423 326247
rect 328365 326207 328423 326213
rect 338117 326247 338175 326253
rect 338117 326213 338129 326247
rect 338163 326244 338175 326247
rect 347593 326247 347651 326253
rect 347593 326244 347605 326247
rect 338163 326216 347605 326244
rect 338163 326213 338175 326216
rect 338117 326207 338175 326213
rect 347593 326213 347605 326216
rect 347639 326213 347651 326247
rect 347593 326207 347651 326213
rect 279234 326136 279240 326188
rect 279292 326176 279298 326188
rect 280157 326179 280215 326185
rect 280157 326176 280169 326179
rect 279292 326148 280169 326176
rect 279292 326136 279298 326148
rect 280157 326145 280169 326148
rect 280203 326145 280215 326179
rect 280157 326139 280215 326145
rect 261662 326068 261668 326120
rect 261720 326068 261726 326120
rect 278958 326068 278964 326120
rect 279016 326108 279022 326120
rect 279970 326108 279976 326120
rect 279016 326080 279976 326108
rect 279016 326068 279022 326080
rect 279970 326068 279976 326080
rect 280028 326068 280034 326120
rect 280246 326068 280252 326120
rect 280304 326108 280310 326120
rect 281442 326108 281448 326120
rect 280304 326080 281448 326108
rect 280304 326068 280310 326080
rect 281442 326068 281448 326080
rect 281500 326068 281506 326120
rect 280157 326043 280215 326049
rect 280157 326009 280169 326043
rect 280203 326040 280215 326043
rect 289725 326043 289783 326049
rect 289725 326040 289737 326043
rect 280203 326012 289737 326040
rect 280203 326009 280215 326012
rect 280157 326003 280215 326009
rect 289725 326009 289737 326012
rect 289771 326009 289783 326043
rect 289725 326003 289783 326009
rect 274358 325632 274364 325644
rect 274319 325604 274364 325632
rect 274358 325592 274364 325604
rect 274416 325592 274422 325644
rect 261846 325252 261852 325304
rect 261904 325292 261910 325304
rect 303614 325292 303620 325304
rect 261904 325264 303620 325292
rect 261904 325252 261910 325264
rect 303614 325252 303620 325264
rect 303672 325252 303678 325304
rect 268378 325184 268384 325236
rect 268436 325224 268442 325236
rect 367094 325224 367100 325236
rect 268436 325196 367100 325224
rect 268436 325184 268442 325196
rect 367094 325184 367100 325196
rect 367152 325184 367158 325236
rect 213822 325116 213828 325168
rect 213880 325156 213886 325168
rect 251450 325156 251456 325168
rect 213880 325128 251456 325156
rect 213880 325116 213886 325128
rect 251450 325116 251456 325128
rect 251508 325116 251514 325168
rect 270770 325116 270776 325168
rect 270828 325156 270834 325168
rect 398834 325156 398840 325168
rect 270828 325128 398840 325156
rect 270828 325116 270834 325128
rect 398834 325116 398840 325128
rect 398892 325116 398898 325168
rect 141970 325048 141976 325100
rect 142028 325088 142034 325100
rect 244734 325088 244740 325100
rect 142028 325060 244740 325088
rect 142028 325048 142034 325060
rect 244734 325048 244740 325060
rect 244792 325048 244798 325100
rect 272886 325048 272892 325100
rect 272944 325088 272950 325100
rect 418154 325088 418160 325100
rect 272944 325060 418160 325088
rect 272944 325048 272950 325060
rect 418154 325048 418160 325060
rect 418212 325048 418218 325100
rect 103422 324980 103428 325032
rect 103480 325020 103486 325032
rect 240226 325020 240232 325032
rect 103480 324992 240232 325020
rect 103480 324980 103486 324992
rect 240226 324980 240232 324992
rect 240284 324980 240290 325032
rect 281810 324980 281816 325032
rect 281868 325020 281874 325032
rect 502334 325020 502340 325032
rect 281868 324992 502340 325020
rect 281868 324980 281874 324992
rect 502334 324980 502340 324992
rect 502392 324980 502398 325032
rect 42058 324912 42064 324964
rect 42116 324952 42122 324964
rect 233326 324952 233332 324964
rect 42116 324924 233332 324952
rect 42116 324912 42122 324924
rect 233326 324912 233332 324924
rect 233384 324912 233390 324964
rect 288158 324912 288164 324964
rect 288216 324952 288222 324964
rect 564434 324952 564440 324964
rect 288216 324924 564440 324952
rect 288216 324912 288222 324924
rect 564434 324912 564440 324924
rect 564492 324912 564498 324964
rect 260374 324300 260380 324352
rect 260432 324340 260438 324352
rect 260650 324340 260656 324352
rect 260432 324312 260656 324340
rect 260432 324300 260438 324312
rect 260650 324300 260656 324312
rect 260708 324300 260714 324352
rect 262674 324300 262680 324352
rect 262732 324340 262738 324352
rect 263594 324340 263600 324352
rect 262732 324312 263600 324340
rect 262732 324300 262738 324312
rect 263594 324300 263600 324312
rect 263652 324300 263658 324352
rect 277305 324343 277363 324349
rect 277305 324309 277317 324343
rect 277351 324340 277363 324343
rect 277394 324340 277400 324352
rect 277351 324312 277400 324340
rect 277351 324309 277363 324312
rect 277305 324303 277363 324309
rect 277394 324300 277400 324312
rect 277452 324300 277458 324352
rect 262306 323892 262312 323944
rect 262364 323932 262370 323944
rect 313366 323932 313372 323944
rect 262364 323904 313372 323932
rect 262364 323892 262370 323904
rect 313366 323892 313372 323904
rect 313424 323892 313430 323944
rect 269758 323824 269764 323876
rect 269816 323864 269822 323876
rect 385034 323864 385040 323876
rect 269816 323836 385040 323864
rect 269816 323824 269822 323836
rect 385034 323824 385040 323836
rect 385092 323824 385098 323876
rect 217962 323756 217968 323808
rect 218020 323796 218026 323808
rect 252370 323796 252376 323808
rect 218020 323768 252376 323796
rect 218020 323756 218026 323768
rect 252370 323756 252376 323768
rect 252428 323756 252434 323808
rect 279142 323756 279148 323808
rect 279200 323796 279206 323808
rect 436094 323796 436100 323808
rect 279200 323768 436100 323796
rect 279200 323756 279206 323768
rect 436094 323756 436100 323768
rect 436152 323756 436158 323808
rect 165522 323688 165528 323740
rect 165580 323728 165586 323740
rect 245930 323728 245936 323740
rect 165580 323700 245936 323728
rect 165580 323688 165586 323700
rect 245930 323688 245936 323700
rect 245988 323688 245994 323740
rect 275186 323688 275192 323740
rect 275244 323728 275250 323740
rect 437474 323728 437480 323740
rect 275244 323700 437480 323728
rect 275244 323688 275250 323700
rect 437474 323688 437480 323700
rect 437532 323688 437538 323740
rect 114462 323620 114468 323672
rect 114520 323660 114526 323672
rect 240778 323660 240784 323672
rect 114520 323632 240784 323660
rect 114520 323620 114526 323632
rect 240778 323620 240784 323632
rect 240836 323620 240842 323672
rect 285674 323620 285680 323672
rect 285732 323660 285738 323672
rect 540974 323660 540980 323672
rect 285732 323632 540980 323660
rect 285732 323620 285738 323632
rect 540974 323620 540980 323632
rect 541032 323620 541038 323672
rect 46198 323552 46204 323604
rect 46256 323592 46262 323604
rect 234522 323592 234528 323604
rect 46256 323564 234528 323592
rect 46256 323552 46262 323564
rect 234522 323552 234528 323564
rect 234580 323552 234586 323604
rect 289170 323592 289176 323604
rect 289131 323564 289176 323592
rect 289170 323552 289176 323564
rect 289228 323552 289234 323604
rect 290734 323552 290740 323604
rect 290792 323592 290798 323604
rect 568574 323592 568580 323604
rect 290792 323564 568580 323592
rect 290792 323552 290798 323564
rect 568574 323552 568580 323564
rect 568632 323552 568638 323604
rect 287974 322872 287980 322924
rect 288032 322912 288038 322924
rect 288250 322912 288256 322924
rect 288032 322884 288256 322912
rect 288032 322872 288038 322884
rect 288250 322872 288256 322884
rect 288308 322872 288314 322924
rect 290550 322872 290556 322924
rect 290608 322912 290614 322924
rect 580166 322912 580172 322924
rect 290608 322884 580172 322912
rect 290608 322872 290614 322884
rect 580166 322872 580172 322884
rect 580224 322872 580230 322924
rect 226242 322396 226248 322448
rect 226300 322436 226306 322448
rect 253106 322436 253112 322448
rect 226300 322408 253112 322436
rect 226300 322396 226306 322408
rect 253106 322396 253112 322408
rect 253164 322396 253170 322448
rect 263042 322396 263048 322448
rect 263100 322436 263106 322448
rect 321554 322436 321560 322448
rect 263100 322408 321560 322436
rect 263100 322396 263106 322408
rect 321554 322396 321560 322408
rect 321612 322396 321618 322448
rect 146202 322328 146208 322380
rect 146260 322368 146266 322380
rect 245562 322368 245568 322380
rect 146260 322340 245568 322368
rect 146260 322328 146266 322340
rect 245562 322328 245568 322340
rect 245620 322328 245626 322380
rect 276750 322328 276756 322380
rect 276808 322368 276814 322380
rect 454034 322368 454040 322380
rect 276808 322340 454040 322368
rect 276808 322328 276814 322340
rect 454034 322328 454040 322340
rect 454092 322328 454098 322380
rect 121362 322260 121368 322312
rect 121420 322300 121426 322312
rect 242342 322300 242348 322312
rect 121420 322272 242348 322300
rect 121420 322260 121426 322272
rect 242342 322260 242348 322272
rect 242400 322260 242406 322312
rect 277486 322260 277492 322312
rect 277544 322300 277550 322312
rect 469214 322300 469220 322312
rect 277544 322272 469220 322300
rect 277544 322260 277550 322272
rect 469214 322260 469220 322272
rect 469272 322260 469278 322312
rect 67542 322192 67548 322244
rect 67600 322232 67606 322244
rect 233878 322232 233884 322244
rect 67600 322204 233884 322232
rect 67600 322192 67606 322204
rect 233878 322192 233884 322204
rect 233936 322192 233942 322244
rect 289262 322192 289268 322244
rect 289320 322232 289326 322244
rect 567838 322232 567844 322244
rect 289320 322204 567844 322232
rect 289320 322192 289326 322204
rect 567838 322192 567844 322204
rect 567896 322192 567902 322244
rect 260650 321892 260656 321904
rect 260611 321864 260656 321892
rect 260650 321852 260656 321864
rect 260708 321852 260714 321904
rect 289078 321688 289084 321700
rect 289004 321660 289084 321688
rect 233510 321580 233516 321632
rect 233568 321620 233574 321632
rect 233694 321620 233700 321632
rect 233568 321592 233700 321620
rect 233568 321580 233574 321592
rect 233694 321580 233700 321592
rect 233752 321580 233758 321632
rect 289004 321564 289032 321660
rect 289078 321648 289084 321660
rect 289136 321648 289142 321700
rect 288986 321512 288992 321564
rect 289044 321512 289050 321564
rect 270586 321036 270592 321088
rect 270644 321076 270650 321088
rect 394694 321076 394700 321088
rect 270644 321048 394700 321076
rect 270644 321036 270650 321048
rect 394694 321036 394700 321048
rect 394752 321036 394758 321088
rect 150342 320968 150348 321020
rect 150400 321008 150406 321020
rect 245194 321008 245200 321020
rect 150400 320980 245200 321008
rect 150400 320968 150406 320980
rect 245194 320968 245200 320980
rect 245252 320968 245258 321020
rect 276566 320968 276572 321020
rect 276624 321008 276630 321020
rect 448514 321008 448520 321020
rect 276624 320980 448520 321008
rect 276624 320968 276630 320980
rect 448514 320968 448520 320980
rect 448572 320968 448578 321020
rect 125410 320900 125416 320952
rect 125468 320940 125474 320952
rect 242526 320940 242532 320952
rect 125468 320912 242532 320940
rect 125468 320900 125474 320912
rect 242526 320900 242532 320912
rect 242584 320900 242590 320952
rect 279326 320900 279332 320952
rect 279384 320940 279390 320952
rect 476114 320940 476120 320952
rect 279384 320912 476120 320940
rect 279384 320900 279390 320912
rect 476114 320900 476120 320912
rect 476172 320900 476178 320952
rect 82722 320832 82728 320884
rect 82780 320872 82786 320884
rect 238294 320872 238300 320884
rect 82780 320844 238300 320872
rect 82780 320832 82786 320844
rect 238294 320832 238300 320844
rect 238352 320832 238358 320884
rect 290642 320832 290648 320884
rect 290700 320872 290706 320884
rect 571426 320872 571432 320884
rect 290700 320844 571432 320872
rect 290700 320832 290706 320844
rect 571426 320832 571432 320844
rect 571484 320832 571490 320884
rect 245194 320328 245200 320340
rect 245155 320300 245200 320328
rect 245194 320288 245200 320300
rect 245252 320288 245258 320340
rect 261662 319676 261668 319728
rect 261720 319716 261726 319728
rect 306374 319716 306380 319728
rect 261720 319688 306380 319716
rect 261720 319676 261726 319688
rect 306374 319676 306380 319688
rect 306432 319676 306438 319728
rect 267090 319608 267096 319660
rect 267148 319648 267154 319660
rect 364334 319648 364340 319660
rect 267148 319620 364340 319648
rect 267148 319608 267154 319620
rect 364334 319608 364340 319620
rect 364392 319608 364398 319660
rect 210970 319540 210976 319592
rect 211028 319580 211034 319592
rect 251726 319580 251732 319592
rect 211028 319552 251732 319580
rect 211028 319540 211034 319552
rect 251726 319540 251732 319552
rect 251784 319540 251790 319592
rect 274542 319540 274548 319592
rect 274600 319580 274606 319592
rect 433426 319580 433432 319592
rect 274600 319552 433432 319580
rect 274600 319540 274606 319552
rect 433426 319540 433432 319552
rect 433484 319540 433490 319592
rect 154482 319472 154488 319524
rect 154540 319512 154546 319524
rect 246206 319512 246212 319524
rect 154540 319484 246212 319512
rect 154540 319472 154546 319484
rect 246206 319472 246212 319484
rect 246264 319472 246270 319524
rect 280706 319472 280712 319524
rect 280764 319512 280770 319524
rect 487154 319512 487160 319524
rect 280764 319484 487160 319512
rect 280764 319472 280770 319484
rect 487154 319472 487160 319484
rect 487212 319472 487218 319524
rect 13722 319404 13728 319456
rect 13780 319444 13786 319456
rect 229738 319444 229744 319456
rect 13780 319416 229744 319444
rect 13780 319404 13786 319416
rect 229738 319404 229744 319416
rect 229796 319404 229802 319456
rect 287698 319404 287704 319456
rect 287756 319444 287762 319456
rect 554866 319444 554872 319456
rect 287756 319416 554872 319444
rect 287756 319404 287762 319416
rect 554866 319404 554872 319416
rect 554924 319404 554930 319456
rect 233970 318860 233976 318912
rect 234028 318860 234034 318912
rect 233988 318776 234016 318860
rect 237009 318835 237067 318841
rect 237009 318801 237021 318835
rect 237055 318832 237067 318835
rect 237098 318832 237104 318844
rect 237055 318804 237104 318832
rect 237055 318801 237067 318804
rect 237009 318795 237067 318801
rect 237098 318792 237104 318804
rect 237156 318792 237162 318844
rect 267458 318832 267464 318844
rect 267419 318804 267464 318832
rect 267458 318792 267464 318804
rect 267516 318792 267522 318844
rect 289173 318835 289231 318841
rect 289173 318801 289185 318835
rect 289219 318832 289231 318835
rect 289262 318832 289268 318844
rect 289219 318804 289268 318832
rect 289219 318801 289231 318804
rect 289173 318795 289231 318801
rect 289262 318792 289268 318804
rect 289320 318792 289326 318844
rect 229465 318767 229523 318773
rect 229465 318733 229477 318767
rect 229511 318764 229523 318767
rect 229554 318764 229560 318776
rect 229511 318736 229560 318764
rect 229511 318733 229523 318736
rect 229465 318727 229523 318733
rect 229554 318724 229560 318736
rect 229612 318724 229618 318776
rect 233970 318724 233976 318776
rect 234028 318724 234034 318776
rect 245194 318764 245200 318776
rect 245155 318736 245200 318764
rect 245194 318724 245200 318736
rect 245252 318724 245258 318776
rect 264514 318248 264520 318300
rect 264572 318288 264578 318300
rect 335354 318288 335360 318300
rect 264572 318260 335360 318288
rect 264572 318248 264578 318260
rect 335354 318248 335360 318260
rect 335412 318248 335418 318300
rect 136542 318180 136548 318232
rect 136600 318220 136606 318232
rect 243906 318220 243912 318232
rect 136600 318192 243912 318220
rect 136600 318180 136606 318192
rect 243906 318180 243912 318192
rect 243964 318180 243970 318232
rect 270862 318180 270868 318232
rect 270920 318220 270926 318232
rect 401594 318220 401600 318232
rect 270920 318192 401600 318220
rect 270920 318180 270926 318192
rect 401594 318180 401600 318192
rect 401652 318180 401658 318232
rect 99282 318112 99288 318164
rect 99340 318152 99346 318164
rect 240134 318152 240140 318164
rect 99340 318124 240140 318152
rect 99340 318112 99346 318124
rect 240134 318112 240140 318124
rect 240192 318112 240198 318164
rect 280522 318112 280528 318164
rect 280580 318152 280586 318164
rect 447134 318152 447140 318164
rect 280580 318124 447140 318152
rect 280580 318112 280586 318124
rect 447134 318112 447140 318124
rect 447192 318112 447198 318164
rect 50982 318044 50988 318096
rect 51040 318084 51046 318096
rect 234890 318084 234896 318096
rect 51040 318056 234896 318084
rect 51040 318044 51046 318056
rect 234890 318044 234896 318056
rect 234948 318044 234954 318096
rect 257430 318044 257436 318096
rect 257488 318084 257494 318096
rect 270494 318084 270500 318096
rect 257488 318056 270500 318084
rect 257488 318044 257494 318056
rect 270494 318044 270500 318056
rect 270552 318044 270558 318096
rect 282362 318044 282368 318096
rect 282420 318084 282426 318096
rect 505094 318084 505100 318096
rect 282420 318056 505100 318084
rect 282420 318044 282426 318056
rect 505094 318044 505100 318056
rect 505152 318044 505158 318096
rect 267458 317472 267464 317484
rect 267419 317444 267464 317472
rect 267458 317432 267464 317444
rect 267516 317432 267522 317484
rect 235166 317364 235172 317416
rect 235224 317404 235230 317416
rect 235261 317407 235319 317413
rect 235261 317404 235273 317407
rect 235224 317376 235273 317404
rect 235224 317364 235230 317376
rect 235261 317373 235273 317376
rect 235307 317373 235319 317407
rect 235261 317367 235319 317373
rect 268286 316888 268292 316940
rect 268344 316928 268350 316940
rect 371234 316928 371240 316940
rect 268344 316900 371240 316928
rect 268344 316888 268350 316900
rect 371234 316888 371240 316900
rect 371292 316888 371298 316940
rect 272058 316820 272064 316872
rect 272116 316860 272122 316872
rect 408586 316860 408592 316872
rect 272116 316832 408592 316860
rect 272116 316820 272122 316832
rect 408586 316820 408592 316832
rect 408644 316820 408650 316872
rect 140682 316752 140688 316804
rect 140740 316792 140746 316804
rect 244550 316792 244556 316804
rect 140740 316764 244556 316792
rect 140740 316752 140746 316764
rect 244550 316752 244556 316764
rect 244608 316752 244614 316804
rect 276290 316752 276296 316804
rect 276348 316792 276354 316804
rect 458174 316792 458180 316804
rect 276348 316764 458180 316792
rect 276348 316752 276354 316764
rect 458174 316752 458180 316764
rect 458232 316752 458238 316804
rect 110322 316684 110328 316736
rect 110380 316724 110386 316736
rect 240686 316724 240692 316736
rect 110380 316696 240692 316724
rect 110380 316684 110386 316696
rect 240686 316684 240692 316696
rect 240744 316684 240750 316736
rect 279326 316684 279332 316736
rect 279384 316724 279390 316736
rect 279786 316724 279792 316736
rect 279384 316696 279792 316724
rect 279384 316684 279390 316696
rect 279786 316684 279792 316696
rect 279844 316684 279850 316736
rect 283650 316684 283656 316736
rect 283708 316724 283714 316736
rect 516134 316724 516140 316736
rect 283708 316696 516140 316724
rect 283708 316684 283714 316696
rect 516134 316684 516140 316696
rect 516192 316684 516198 316736
rect 254854 316112 254860 316124
rect 254815 316084 254860 316112
rect 254854 316072 254860 316084
rect 254912 316072 254918 316124
rect 256602 316072 256608 316124
rect 256660 316112 256666 316124
rect 256694 316112 256700 316124
rect 256660 316084 256700 316112
rect 256660 316072 256666 316084
rect 256694 316072 256700 316084
rect 256752 316072 256758 316124
rect 274358 316044 274364 316056
rect 274319 316016 274364 316044
rect 274358 316004 274364 316016
rect 274416 316004 274422 316056
rect 258258 315460 258264 315512
rect 258316 315500 258322 315512
rect 285674 315500 285680 315512
rect 258316 315472 285680 315500
rect 258316 315460 258322 315472
rect 285674 315460 285680 315472
rect 285732 315460 285738 315512
rect 274082 315392 274088 315444
rect 274140 315432 274146 315444
rect 423674 315432 423680 315444
rect 274140 315404 423680 315432
rect 274140 315392 274146 315404
rect 423674 315392 423680 315404
rect 423732 315392 423738 315444
rect 143442 315324 143448 315376
rect 143500 315364 143506 315376
rect 244826 315364 244832 315376
rect 143500 315336 244832 315364
rect 143500 315324 143506 315336
rect 244826 315324 244832 315336
rect 244884 315324 244890 315376
rect 283466 315324 283472 315376
rect 283524 315364 283530 315376
rect 460934 315364 460940 315376
rect 283524 315336 460940 315364
rect 283524 315324 283530 315336
rect 460934 315324 460940 315336
rect 460992 315324 460998 315376
rect 24118 315256 24124 315308
rect 24176 315296 24182 315308
rect 232682 315296 232688 315308
rect 24176 315268 232688 315296
rect 24176 315256 24182 315268
rect 232682 315256 232688 315268
rect 232740 315256 232746 315308
rect 285214 315256 285220 315308
rect 285272 315296 285278 315308
rect 534074 315296 534080 315308
rect 285272 315268 534080 315296
rect 285272 315256 285278 315268
rect 534074 315256 534080 315268
rect 534132 315256 534138 315308
rect 260650 314684 260656 314696
rect 260611 314656 260656 314684
rect 260650 314644 260656 314656
rect 260708 314644 260714 314696
rect 262398 314644 262404 314696
rect 262456 314684 262462 314696
rect 262582 314684 262588 314696
rect 262456 314656 262588 314684
rect 262456 314644 262462 314656
rect 262582 314644 262588 314656
rect 262640 314644 262646 314696
rect 275370 314032 275376 314084
rect 275428 314072 275434 314084
rect 441614 314072 441620 314084
rect 275428 314044 441620 314072
rect 275428 314032 275434 314044
rect 441614 314032 441620 314044
rect 441672 314032 441678 314084
rect 147582 313964 147588 314016
rect 147640 314004 147646 314016
rect 245010 314004 245016 314016
rect 147640 313976 245016 314004
rect 147640 313964 147646 313976
rect 245010 313964 245016 313976
rect 245068 313964 245074 314016
rect 279418 313964 279424 314016
rect 279476 314004 279482 314016
rect 478874 314004 478880 314016
rect 279476 313976 478880 314004
rect 279476 313964 279482 313976
rect 478874 313964 478880 313976
rect 478932 313964 478938 314016
rect 31018 313896 31024 313948
rect 31076 313936 31082 313948
rect 232038 313936 232044 313948
rect 31076 313908 232044 313936
rect 31076 313896 31082 313908
rect 232038 313896 232044 313908
rect 232096 313896 232102 313948
rect 261754 313896 261760 313948
rect 261812 313936 261818 313948
rect 278774 313936 278780 313948
rect 261812 313908 278780 313936
rect 261812 313896 261818 313908
rect 278774 313896 278780 313908
rect 278832 313896 278838 313948
rect 286410 313896 286416 313948
rect 286468 313936 286474 313948
rect 545114 313936 545120 313948
rect 286468 313908 545120 313936
rect 286468 313896 286474 313908
rect 545114 313896 545120 313908
rect 545172 313896 545178 313948
rect 278406 312672 278412 312724
rect 278464 312712 278470 312724
rect 466454 312712 466460 312724
rect 278464 312684 466460 312712
rect 278464 312672 278470 312684
rect 466454 312672 466460 312684
rect 466512 312672 466518 312724
rect 158622 312604 158628 312656
rect 158680 312644 158686 312656
rect 246114 312644 246120 312656
rect 158680 312616 246120 312644
rect 158680 312604 158686 312616
rect 246114 312604 246120 312616
rect 246172 312604 246178 312656
rect 279510 312604 279516 312656
rect 279568 312644 279574 312656
rect 484394 312644 484400 312656
rect 279568 312616 484400 312644
rect 279568 312604 279574 312616
rect 484394 312604 484400 312616
rect 484452 312604 484458 312656
rect 31662 312536 31668 312588
rect 31720 312576 31726 312588
rect 233142 312576 233148 312588
rect 31720 312548 233148 312576
rect 31720 312536 31726 312548
rect 233142 312536 233148 312548
rect 233200 312536 233206 312588
rect 286778 312536 286784 312588
rect 286836 312576 286842 312588
rect 552014 312576 552020 312588
rect 286836 312548 552020 312576
rect 286836 312536 286842 312548
rect 552014 312536 552020 312548
rect 552072 312536 552078 312588
rect 245194 311828 245200 311840
rect 245155 311800 245200 311828
rect 245194 311788 245200 311800
rect 245252 311788 245258 311840
rect 500218 311788 500224 311840
rect 500276 311828 500282 311840
rect 580166 311828 580172 311840
rect 500276 311800 580172 311828
rect 500276 311788 500282 311800
rect 580166 311788 580172 311800
rect 580224 311788 580230 311840
rect 260834 311312 260840 311364
rect 260892 311352 260898 311364
rect 310514 311352 310520 311364
rect 260892 311324 310520 311352
rect 260892 311312 260898 311324
rect 310514 311312 310520 311324
rect 310572 311312 310578 311364
rect 268562 311244 268568 311296
rect 268620 311284 268626 311296
rect 378134 311284 378140 311296
rect 268620 311256 378140 311284
rect 268620 311244 268626 311256
rect 378134 311244 378140 311256
rect 378192 311244 378198 311296
rect 161382 311176 161388 311228
rect 161440 311216 161446 311228
rect 246482 311216 246488 311228
rect 161440 311188 246488 311216
rect 161440 311176 161446 311188
rect 246482 311176 246488 311188
rect 246540 311176 246546 311228
rect 273622 311176 273628 311228
rect 273680 311216 273686 311228
rect 273990 311216 273996 311228
rect 273680 311188 273996 311216
rect 273680 311176 273686 311188
rect 273990 311176 273996 311188
rect 274048 311176 274054 311228
rect 280890 311176 280896 311228
rect 280948 311216 280954 311228
rect 491294 311216 491300 311228
rect 280948 311188 491300 311216
rect 280948 311176 280954 311188
rect 491294 311176 491300 311188
rect 491352 311176 491358 311228
rect 50338 311108 50344 311160
rect 50396 311148 50402 311160
rect 235902 311148 235908 311160
rect 50396 311120 235908 311148
rect 50396 311108 50402 311120
rect 235902 311108 235908 311120
rect 235960 311108 235966 311160
rect 289446 311108 289452 311160
rect 289504 311148 289510 311160
rect 571978 311148 571984 311160
rect 289504 311120 571984 311148
rect 289504 311108 289510 311120
rect 571978 311108 571984 311120
rect 572036 311108 572042 311160
rect 229462 310808 229468 310820
rect 229423 310780 229468 310808
rect 229462 310768 229468 310780
rect 229520 310768 229526 310820
rect 277762 310088 277768 310140
rect 277820 310128 277826 310140
rect 277946 310128 277952 310140
rect 277820 310100 277952 310128
rect 277820 310088 277826 310100
rect 277946 310088 277952 310100
rect 278004 310088 278010 310140
rect 263226 309952 263232 310004
rect 263284 309992 263290 310004
rect 317414 309992 317420 310004
rect 263284 309964 317420 309992
rect 263284 309952 263290 309964
rect 317414 309952 317420 309964
rect 317472 309952 317478 310004
rect 269942 309884 269948 309936
rect 270000 309924 270006 309936
rect 389174 309924 389180 309936
rect 270000 309896 389180 309924
rect 270000 309884 270006 309896
rect 389174 309884 389180 309896
rect 389232 309884 389238 309936
rect 280982 309816 280988 309868
rect 281040 309856 281046 309868
rect 494054 309856 494060 309868
rect 281040 309828 494060 309856
rect 281040 309816 281046 309828
rect 494054 309816 494060 309828
rect 494112 309816 494118 309868
rect 107470 309748 107476 309800
rect 107528 309788 107534 309800
rect 240502 309788 240508 309800
rect 107528 309760 240508 309788
rect 107528 309748 107534 309760
rect 240502 309748 240508 309760
rect 240560 309748 240566 309800
rect 287422 309748 287428 309800
rect 287480 309788 287486 309800
rect 556798 309788 556804 309800
rect 287480 309760 556804 309788
rect 287480 309748 287486 309760
rect 556798 309748 556804 309760
rect 556856 309748 556862 309800
rect 3418 309068 3424 309120
rect 3476 309108 3482 309120
rect 211798 309108 211804 309120
rect 3476 309080 211804 309108
rect 3476 309068 3482 309080
rect 211798 309068 211804 309080
rect 211856 309068 211862 309120
rect 229462 309108 229468 309120
rect 229423 309080 229468 309108
rect 229462 309068 229468 309080
rect 229520 309068 229526 309120
rect 273622 309108 273628 309120
rect 273583 309080 273628 309108
rect 273622 309068 273628 309080
rect 273680 309068 273686 309120
rect 263962 308524 263968 308576
rect 264020 308564 264026 308576
rect 339494 308564 339500 308576
rect 264020 308536 339500 308564
rect 264020 308524 264026 308536
rect 339494 308524 339500 308536
rect 339552 308524 339558 308576
rect 281074 308456 281080 308508
rect 281132 308496 281138 308508
rect 498194 308496 498200 308508
rect 281132 308468 498200 308496
rect 281132 308456 281138 308468
rect 498194 308456 498200 308468
rect 498252 308456 498258 308508
rect 288618 308388 288624 308440
rect 288676 308428 288682 308440
rect 574830 308428 574836 308440
rect 288676 308400 574836 308428
rect 288676 308388 288682 308400
rect 574830 308388 574836 308400
rect 574888 308388 574894 308440
rect 269666 307884 269672 307896
rect 269592 307856 269672 307884
rect 233970 307708 233976 307760
rect 234028 307708 234034 307760
rect 237193 307751 237251 307757
rect 237193 307717 237205 307751
rect 237239 307748 237251 307751
rect 237282 307748 237288 307760
rect 237239 307720 237288 307748
rect 237239 307717 237251 307720
rect 237193 307711 237251 307717
rect 237282 307708 237288 307720
rect 237340 307708 237346 307760
rect 233786 307640 233792 307692
rect 233844 307680 233850 307692
rect 233988 307680 234016 307708
rect 269592 307692 269620 307856
rect 269666 307844 269672 307856
rect 269724 307844 269730 307896
rect 233844 307652 234016 307680
rect 233844 307640 233850 307652
rect 269574 307640 269580 307692
rect 269632 307640 269638 307692
rect 270954 307096 270960 307148
rect 271012 307136 271018 307148
rect 405734 307136 405740 307148
rect 271012 307108 405740 307136
rect 271012 307096 271018 307108
rect 405734 307096 405740 307108
rect 405792 307096 405798 307148
rect 43438 307028 43444 307080
rect 43496 307068 43502 307080
rect 233694 307068 233700 307080
rect 43496 307040 233700 307068
rect 43496 307028 43502 307040
rect 233694 307028 233700 307040
rect 233752 307028 233758 307080
rect 279326 307028 279332 307080
rect 279384 307068 279390 307080
rect 279786 307068 279792 307080
rect 279384 307040 279792 307068
rect 279384 307028 279390 307040
rect 279786 307028 279792 307040
rect 279844 307028 279850 307080
rect 282178 307028 282184 307080
rect 282236 307068 282242 307080
rect 511994 307068 512000 307080
rect 282236 307040 512000 307068
rect 282236 307028 282242 307040
rect 511994 307028 512000 307040
rect 512052 307028 512058 307080
rect 262582 306484 262588 306536
rect 262640 306524 262646 306536
rect 262640 306496 262720 306524
rect 262640 306484 262646 306496
rect 262692 306400 262720 306496
rect 268838 306416 268844 306468
rect 268896 306456 268902 306468
rect 269022 306456 269028 306468
rect 268896 306428 269028 306456
rect 268896 306416 268902 306428
rect 269022 306416 269028 306428
rect 269080 306416 269086 306468
rect 262674 306348 262680 306400
rect 262732 306348 262738 306400
rect 264238 306348 264244 306400
rect 264296 306388 264302 306400
rect 264330 306388 264336 306400
rect 264296 306360 264336 306388
rect 264296 306348 264302 306360
rect 264330 306348 264336 306360
rect 264388 306348 264394 306400
rect 272426 305668 272432 305720
rect 272484 305708 272490 305720
rect 412634 305708 412640 305720
rect 272484 305680 412640 305708
rect 272484 305668 272490 305680
rect 412634 305668 412640 305680
rect 412692 305668 412698 305720
rect 38470 305600 38476 305652
rect 38528 305640 38534 305652
rect 233602 305640 233608 305652
rect 38528 305612 233608 305640
rect 38528 305600 38534 305612
rect 233602 305600 233608 305612
rect 233660 305600 233666 305652
rect 284018 305600 284024 305652
rect 284076 305640 284082 305652
rect 520274 305640 520280 305652
rect 284076 305612 520280 305640
rect 284076 305600 284082 305612
rect 520274 305600 520280 305612
rect 520332 305600 520338 305652
rect 254762 304920 254768 304972
rect 254820 304960 254826 304972
rect 255038 304960 255044 304972
rect 254820 304932 255044 304960
rect 254820 304920 254826 304932
rect 255038 304920 255044 304932
rect 255096 304920 255102 304972
rect 273162 304308 273168 304360
rect 273220 304348 273226 304360
rect 419534 304348 419540 304360
rect 273220 304320 419540 304348
rect 273220 304308 273226 304320
rect 419534 304308 419540 304320
rect 419592 304308 419598 304360
rect 42702 304240 42708 304292
rect 42760 304280 42766 304292
rect 234246 304280 234252 304292
rect 42760 304252 234252 304280
rect 42760 304240 42766 304252
rect 234246 304240 234252 304252
rect 234304 304240 234310 304292
rect 283834 304240 283840 304292
rect 283892 304280 283898 304292
rect 523034 304280 523040 304292
rect 283892 304252 523040 304280
rect 283892 304240 283898 304252
rect 523034 304240 523040 304252
rect 523092 304240 523098 304292
rect 273438 302948 273444 303000
rect 273496 302988 273502 303000
rect 426434 302988 426440 303000
rect 273496 302960 426440 302988
rect 273496 302948 273502 302960
rect 426434 302948 426440 302960
rect 426492 302948 426498 303000
rect 283926 302880 283932 302932
rect 283984 302920 283990 302932
rect 527174 302920 527180 302932
rect 283984 302892 527180 302920
rect 283984 302880 283990 302892
rect 527174 302880 527180 302892
rect 527232 302880 527238 302932
rect 277762 302132 277768 302184
rect 277820 302172 277826 302184
rect 277946 302172 277952 302184
rect 277820 302144 277952 302172
rect 277820 302132 277826 302144
rect 277946 302132 277952 302144
rect 278004 302132 278010 302184
rect 235261 301971 235319 301977
rect 235261 301937 235273 301971
rect 235307 301968 235319 301971
rect 235350 301968 235356 301980
rect 235307 301940 235356 301968
rect 235307 301937 235319 301940
rect 235261 301931 235319 301937
rect 235350 301928 235356 301940
rect 235408 301928 235414 301980
rect 275554 301520 275560 301572
rect 275612 301560 275618 301572
rect 444374 301560 444380 301572
rect 275612 301532 444380 301560
rect 275612 301520 275618 301532
rect 444374 301520 444380 301532
rect 444432 301520 444438 301572
rect 285122 301452 285128 301504
rect 285180 301492 285186 301504
rect 529934 301492 529940 301504
rect 285180 301464 529940 301492
rect 285180 301452 285186 301464
rect 529934 301452 529940 301464
rect 529992 301452 529998 301504
rect 276014 300160 276020 300212
rect 276072 300200 276078 300212
rect 455414 300200 455420 300212
rect 276072 300172 455420 300200
rect 276072 300160 276078 300172
rect 455414 300160 455420 300172
rect 455472 300160 455478 300212
rect 284478 300092 284484 300144
rect 284536 300132 284542 300144
rect 536926 300132 536932 300144
rect 284536 300104 536932 300132
rect 284536 300092 284542 300104
rect 536926 300092 536932 300104
rect 536984 300092 536990 300144
rect 274450 299588 274456 299600
rect 274376 299560 274456 299588
rect 229465 299523 229523 299529
rect 229465 299489 229477 299523
rect 229511 299520 229523 299523
rect 229554 299520 229560 299532
rect 229511 299492 229560 299520
rect 229511 299489 229523 299492
rect 229465 299483 229523 299489
rect 229554 299480 229560 299492
rect 229612 299480 229618 299532
rect 266170 299480 266176 299532
rect 266228 299520 266234 299532
rect 266262 299520 266268 299532
rect 266228 299492 266268 299520
rect 266228 299480 266234 299492
rect 266262 299480 266268 299492
rect 266320 299480 266326 299532
rect 271138 299480 271144 299532
rect 271196 299520 271202 299532
rect 271506 299520 271512 299532
rect 271196 299492 271512 299520
rect 271196 299480 271202 299492
rect 271506 299480 271512 299492
rect 271564 299480 271570 299532
rect 274376 299464 274404 299560
rect 274450 299548 274456 299560
rect 274508 299548 274514 299600
rect 274358 299412 274364 299464
rect 274416 299412 274422 299464
rect 302970 299412 302976 299464
rect 303028 299452 303034 299464
rect 579798 299452 579804 299464
rect 303028 299424 579804 299452
rect 303028 299412 303034 299424
rect 579798 299412 579804 299424
rect 579856 299412 579862 299464
rect 277578 298732 277584 298784
rect 277636 298772 277642 298784
rect 473354 298772 473360 298784
rect 277636 298744 473360 298772
rect 277636 298732 277642 298744
rect 473354 298732 473360 298744
rect 473412 298732 473418 298784
rect 237190 298160 237196 298172
rect 237151 298132 237196 298160
rect 237190 298120 237196 298132
rect 237248 298120 237254 298172
rect 235350 298092 235356 298104
rect 235311 298064 235356 298092
rect 235350 298052 235356 298064
rect 235408 298052 235414 298104
rect 284573 298095 284631 298101
rect 284573 298061 284585 298095
rect 284619 298092 284631 298095
rect 284662 298092 284668 298104
rect 284619 298064 284668 298092
rect 284619 298061 284631 298064
rect 284573 298055 284631 298061
rect 284662 298052 284668 298064
rect 284720 298052 284726 298104
rect 288342 298092 288348 298104
rect 288303 298064 288348 298092
rect 288342 298052 288348 298064
rect 288400 298052 288406 298104
rect 289081 298095 289139 298101
rect 289081 298061 289093 298095
rect 289127 298092 289139 298095
rect 289262 298092 289268 298104
rect 289127 298064 289268 298092
rect 289127 298061 289139 298064
rect 289081 298055 289139 298061
rect 289262 298052 289268 298064
rect 289320 298052 289326 298104
rect 286594 297440 286600 297492
rect 286652 297480 286658 297492
rect 547874 297480 547880 297492
rect 286652 297452 547880 297480
rect 286652 297440 286658 297452
rect 547874 297440 547880 297452
rect 547932 297440 547938 297492
rect 288710 297372 288716 297424
rect 288768 297412 288774 297424
rect 570598 297412 570604 297424
rect 288768 297384 570604 297412
rect 288768 297372 288774 297384
rect 570598 297372 570604 297384
rect 570656 297372 570662 297424
rect 264238 296692 264244 296744
rect 264296 296732 264302 296744
rect 264422 296732 264428 296744
rect 264296 296704 264428 296732
rect 264296 296692 264302 296704
rect 264422 296692 264428 296704
rect 264480 296692 264486 296744
rect 273622 296732 273628 296744
rect 273583 296704 273628 296732
rect 273622 296692 273628 296704
rect 273680 296692 273686 296744
rect 252186 296624 252192 296676
rect 252244 296664 252250 296676
rect 252278 296664 252284 296676
rect 252244 296636 252284 296664
rect 252244 296624 252250 296636
rect 252278 296624 252284 296636
rect 252336 296624 252342 296676
rect 288986 296012 288992 296064
rect 289044 296052 289050 296064
rect 482278 296052 482284 296064
rect 289044 296024 482284 296052
rect 289044 296012 289050 296024
rect 482278 296012 482284 296024
rect 482336 296012 482342 296064
rect 287882 295944 287888 295996
rect 287940 295984 287946 295996
rect 563054 295984 563060 295996
rect 287940 295956 563060 295984
rect 287940 295944 287946 295956
rect 563054 295944 563060 295956
rect 563112 295944 563118 295996
rect 3050 295264 3056 295316
rect 3108 295304 3114 295316
rect 227162 295304 227168 295316
rect 3108 295276 227168 295304
rect 3108 295264 3114 295276
rect 227162 295264 227168 295276
rect 227220 295264 227226 295316
rect 254854 295304 254860 295316
rect 254815 295276 254860 295304
rect 254854 295264 254860 295276
rect 254912 295264 254918 295316
rect 255777 295307 255835 295313
rect 255777 295273 255789 295307
rect 255823 295304 255835 295307
rect 255866 295304 255872 295316
rect 255823 295276 255872 295304
rect 255823 295273 255835 295276
rect 255777 295267 255835 295273
rect 255866 295264 255872 295276
rect 255924 295264 255930 295316
rect 256418 295264 256424 295316
rect 256476 295304 256482 295316
rect 256602 295304 256608 295316
rect 256476 295276 256608 295304
rect 256476 295264 256482 295276
rect 256602 295264 256608 295276
rect 256660 295264 256666 295316
rect 287974 294584 287980 294636
rect 288032 294624 288038 294636
rect 560938 294624 560944 294636
rect 288032 294596 560944 294624
rect 288032 294584 288038 294596
rect 560938 294584 560944 294596
rect 560996 294584 561002 294636
rect 262490 293292 262496 293344
rect 262548 293332 262554 293344
rect 324314 293332 324320 293344
rect 262548 293304 324320 293332
rect 262548 293292 262554 293304
rect 324314 293292 324320 293304
rect 324372 293292 324378 293344
rect 292022 293224 292028 293276
rect 292080 293264 292086 293276
rect 572714 293264 572720 293276
rect 292080 293236 572720 293264
rect 292080 293224 292086 293236
rect 572714 293224 572720 293236
rect 572772 293224 572778 293276
rect 243538 292652 243544 292664
rect 243372 292624 243544 292652
rect 243372 292596 243400 292624
rect 243538 292612 243544 292624
rect 243596 292612 243602 292664
rect 243354 292544 243360 292596
rect 243412 292544 243418 292596
rect 272794 291864 272800 291916
rect 272852 291904 272858 291916
rect 416866 291904 416872 291916
rect 272852 291876 416872 291904
rect 272852 291864 272858 291876
rect 416866 291864 416872 291876
rect 416924 291864 416930 291916
rect 282638 291796 282644 291848
rect 282696 291836 282702 291848
rect 506474 291836 506480 291848
rect 282696 291808 506480 291836
rect 282696 291796 282702 291808
rect 506474 291796 506480 291808
rect 506532 291796 506538 291848
rect 274174 290504 274180 290556
rect 274232 290544 274238 290556
rect 430574 290544 430580 290556
rect 274232 290516 430580 290544
rect 274232 290504 274238 290516
rect 430574 290504 430580 290516
rect 430632 290504 430638 290556
rect 277118 290436 277124 290488
rect 277176 290476 277182 290488
rect 277302 290476 277308 290488
rect 277176 290448 277308 290476
rect 277176 290436 277182 290448
rect 277302 290436 277308 290448
rect 277360 290436 277366 290488
rect 285766 290436 285772 290488
rect 285824 290476 285830 290488
rect 542354 290476 542360 290488
rect 285824 290448 542360 290476
rect 285824 290436 285830 290448
rect 542354 290436 542360 290448
rect 542412 290436 542418 290488
rect 235350 289796 235356 289808
rect 235311 289768 235356 289796
rect 235350 289756 235356 289768
rect 235408 289756 235414 289808
rect 273806 289756 273812 289808
rect 273864 289796 273870 289808
rect 273898 289796 273904 289808
rect 273864 289768 273904 289796
rect 273864 289756 273870 289768
rect 273898 289756 273904 289768
rect 273956 289756 273962 289808
rect 277118 289756 277124 289808
rect 277176 289796 277182 289808
rect 277302 289796 277308 289808
rect 277176 289768 277308 289796
rect 277176 289756 277182 289768
rect 277302 289756 277308 289768
rect 277360 289756 277366 289808
rect 276842 289144 276848 289196
rect 276900 289184 276906 289196
rect 451366 289184 451372 289196
rect 276900 289156 451372 289184
rect 276900 289144 276906 289156
rect 451366 289144 451372 289156
rect 451424 289144 451430 289196
rect 255774 289116 255780 289128
rect 255735 289088 255780 289116
rect 255774 289076 255780 289088
rect 255832 289076 255838 289128
rect 288345 289119 288403 289125
rect 288345 289085 288357 289119
rect 288391 289116 288403 289119
rect 556154 289116 556160 289128
rect 288391 289088 556160 289116
rect 288391 289085 288403 289088
rect 288345 289079 288403 289085
rect 556154 289076 556160 289088
rect 556212 289076 556218 289128
rect 284570 288436 284576 288448
rect 284531 288408 284576 288436
rect 284570 288396 284576 288408
rect 284628 288396 284634 288448
rect 289078 288436 289084 288448
rect 289039 288408 289084 288436
rect 289078 288396 289084 288408
rect 289136 288396 289142 288448
rect 276934 287648 276940 287700
rect 276992 287688 276998 287700
rect 459646 287688 459652 287700
rect 276992 287660 459652 287688
rect 276992 287648 276998 287660
rect 459646 287648 459652 287660
rect 459704 287648 459710 287700
rect 257154 287036 257160 287088
rect 257212 287076 257218 287088
rect 257246 287076 257252 287088
rect 257212 287048 257252 287076
rect 257212 287036 257218 287048
rect 257246 287036 257252 287048
rect 257304 287036 257310 287088
rect 279602 286288 279608 286340
rect 279660 286328 279666 286340
rect 477494 286328 477500 286340
rect 279660 286300 477500 286328
rect 279660 286288 279666 286300
rect 477494 286288 477500 286300
rect 477552 286288 477558 286340
rect 254854 285716 254860 285728
rect 254815 285688 254860 285716
rect 254854 285676 254860 285688
rect 254912 285676 254918 285728
rect 279694 284928 279700 284980
rect 279752 284968 279758 284980
rect 480254 284968 480260 284980
rect 279752 284940 480260 284968
rect 279752 284928 279758 284940
rect 480254 284928 480260 284940
rect 480312 284928 480318 284980
rect 277026 283568 277032 283620
rect 277084 283608 277090 283620
rect 277210 283608 277216 283620
rect 277084 283580 277216 283608
rect 277084 283568 277090 283580
rect 277210 283568 277216 283580
rect 277268 283568 277274 283620
rect 279786 283568 279792 283620
rect 279844 283608 279850 283620
rect 485774 283608 485780 283620
rect 279844 283580 485780 283608
rect 279844 283568 279850 283580
rect 485774 283568 485780 283580
rect 485832 283568 485838 283620
rect 233694 282888 233700 282940
rect 233752 282928 233758 282940
rect 233878 282928 233884 282940
rect 233752 282900 233884 282928
rect 233752 282888 233758 282900
rect 233878 282888 233884 282900
rect 233936 282888 233942 282940
rect 280154 282140 280160 282192
rect 280212 282180 280218 282192
rect 488534 282180 488540 282192
rect 280212 282152 488540 282180
rect 280212 282140 280218 282152
rect 488534 282140 488540 282152
rect 488592 282140 488598 282192
rect 281258 280780 281264 280832
rect 281316 280820 281322 280832
rect 492674 280820 492680 280832
rect 281316 280792 492680 280820
rect 281316 280780 281322 280792
rect 492674 280780 492680 280792
rect 492732 280780 492738 280832
rect 250530 280168 250536 280220
rect 250588 280208 250594 280220
rect 250714 280208 250720 280220
rect 250588 280180 250720 280208
rect 250588 280168 250594 280180
rect 250714 280168 250720 280180
rect 250772 280168 250778 280220
rect 229554 280140 229560 280152
rect 229515 280112 229560 280140
rect 229554 280100 229560 280112
rect 229612 280100 229618 280152
rect 235534 280140 235540 280152
rect 235495 280112 235540 280140
rect 235534 280100 235540 280112
rect 235592 280100 235598 280152
rect 237098 280100 237104 280152
rect 237156 280140 237162 280152
rect 237190 280140 237196 280152
rect 237156 280112 237196 280140
rect 237156 280100 237162 280112
rect 237190 280100 237196 280112
rect 237248 280100 237254 280152
rect 281350 279420 281356 279472
rect 281408 279460 281414 279472
rect 495434 279460 495440 279472
rect 281408 279432 495440 279460
rect 281408 279420 281414 279432
rect 495434 279420 495440 279432
rect 495492 279420 495498 279472
rect 235166 278740 235172 278792
rect 235224 278780 235230 278792
rect 235350 278780 235356 278792
rect 235224 278752 235356 278780
rect 235224 278740 235230 278752
rect 235350 278740 235356 278752
rect 235408 278740 235414 278792
rect 284938 277992 284944 278044
rect 284996 278032 285002 278044
rect 502426 278032 502432 278044
rect 284996 278004 502432 278032
rect 284996 277992 285002 278004
rect 502426 277992 502432 278004
rect 502484 277992 502490 278044
rect 281994 276632 282000 276684
rect 282052 276672 282058 276684
rect 510614 276672 510620 276684
rect 282052 276644 510620 276672
rect 282052 276632 282058 276644
rect 510614 276632 510620 276644
rect 510672 276632 510678 276684
rect 309778 275952 309784 276004
rect 309836 275992 309842 276004
rect 580166 275992 580172 276004
rect 309836 275964 580172 275992
rect 309836 275952 309842 275964
rect 580166 275952 580172 275964
rect 580224 275952 580230 276004
rect 255774 274632 255780 274644
rect 255735 274604 255780 274632
rect 255774 274592 255780 274604
rect 255832 274592 255838 274644
rect 277210 274632 277216 274644
rect 277171 274604 277216 274632
rect 277210 274592 277216 274604
rect 277268 274592 277274 274644
rect 235169 273955 235227 273961
rect 235169 273921 235181 273955
rect 235215 273952 235227 273955
rect 235258 273952 235264 273964
rect 235215 273924 235264 273952
rect 235215 273921 235227 273924
rect 235169 273915 235227 273921
rect 235258 273912 235264 273924
rect 235316 273912 235322 273964
rect 282270 273912 282276 273964
rect 282328 273952 282334 273964
rect 513374 273952 513380 273964
rect 282328 273924 513380 273952
rect 282328 273912 282334 273924
rect 513374 273912 513380 273924
rect 513432 273912 513438 273964
rect 250254 273096 250260 273148
rect 250312 273136 250318 273148
rect 250714 273136 250720 273148
rect 250312 273108 250720 273136
rect 250312 273096 250318 273108
rect 250714 273096 250720 273108
rect 250772 273096 250778 273148
rect 283006 272484 283012 272536
rect 283064 272524 283070 272536
rect 517514 272524 517520 272536
rect 283064 272496 517520 272524
rect 283064 272484 283070 272496
rect 517514 272484 517520 272496
rect 517572 272484 517578 272536
rect 284110 271124 284116 271176
rect 284168 271164 284174 271176
rect 520366 271164 520372 271176
rect 284168 271136 520372 271164
rect 284168 271124 284174 271136
rect 520366 271124 520372 271136
rect 520424 271124 520430 271176
rect 238846 270580 238852 270632
rect 238904 270620 238910 270632
rect 259914 270620 259920 270632
rect 238904 270592 238984 270620
rect 238904 270580 238910 270592
rect 238956 270564 238984 270592
rect 259840 270592 259920 270620
rect 229557 270555 229615 270561
rect 229557 270521 229569 270555
rect 229603 270552 229615 270555
rect 229646 270552 229652 270564
rect 229603 270524 229652 270552
rect 229603 270521 229615 270524
rect 229557 270515 229615 270521
rect 229646 270512 229652 270524
rect 229704 270512 229710 270564
rect 235534 270552 235540 270564
rect 235495 270524 235540 270552
rect 235534 270512 235540 270524
rect 235592 270512 235598 270564
rect 238938 270512 238944 270564
rect 238996 270512 239002 270564
rect 259840 270496 259868 270592
rect 259914 270580 259920 270592
rect 259972 270580 259978 270632
rect 259822 270444 259828 270496
rect 259880 270444 259886 270496
rect 283190 269764 283196 269816
rect 283248 269804 283254 269816
rect 524414 269804 524420 269816
rect 283248 269776 524420 269804
rect 283248 269764 283254 269776
rect 524414 269764 524420 269776
rect 524472 269764 524478 269816
rect 285306 268336 285312 268388
rect 285364 268376 285370 268388
rect 528646 268376 528652 268388
rect 285364 268348 528652 268376
rect 285364 268336 285370 268348
rect 528646 268336 528652 268348
rect 528704 268336 528710 268388
rect 284662 266976 284668 267028
rect 284720 267016 284726 267028
rect 531314 267016 531320 267028
rect 284720 266988 531320 267016
rect 284720 266976 284726 266988
rect 531314 266976 531320 266988
rect 531372 266976 531378 267028
rect 2866 266296 2872 266348
rect 2924 266336 2930 266348
rect 209038 266336 209044 266348
rect 2924 266308 209044 266336
rect 2924 266296 2930 266308
rect 209038 266296 209044 266308
rect 209096 266296 209102 266348
rect 276934 266296 276940 266348
rect 276992 266336 276998 266348
rect 277029 266339 277087 266345
rect 277029 266336 277041 266339
rect 276992 266308 277041 266336
rect 276992 266296 276998 266308
rect 277029 266305 277041 266308
rect 277075 266305 277087 266339
rect 277029 266299 277087 266305
rect 284754 265616 284760 265668
rect 284812 265656 284818 265668
rect 535454 265656 535460 265668
rect 284812 265628 535460 265656
rect 284812 265616 284818 265628
rect 535454 265616 535460 265628
rect 535512 265616 535518 265668
rect 255774 264976 255780 264988
rect 255735 264948 255780 264976
rect 255774 264936 255780 264948
rect 255832 264936 255838 264988
rect 277210 264976 277216 264988
rect 277171 264948 277216 264976
rect 277210 264936 277216 264948
rect 277268 264936 277274 264988
rect 498838 264868 498844 264920
rect 498896 264908 498902 264920
rect 580166 264908 580172 264920
rect 498896 264880 580172 264908
rect 498896 264868 498902 264880
rect 580166 264868 580172 264880
rect 580224 264868 580230 264920
rect 288894 264188 288900 264240
rect 288952 264228 288958 264240
rect 475378 264228 475384 264240
rect 288952 264200 475384 264228
rect 288952 264188 288958 264200
rect 475378 264188 475384 264200
rect 475436 264188 475442 264240
rect 233694 263576 233700 263628
rect 233752 263616 233758 263628
rect 233878 263616 233884 263628
rect 233752 263588 233884 263616
rect 233752 263576 233758 263588
rect 233878 263576 233884 263588
rect 233936 263576 233942 263628
rect 273622 263576 273628 263628
rect 273680 263576 273686 263628
rect 273640 263548 273668 263576
rect 273714 263548 273720 263560
rect 273640 263520 273720 263548
rect 273714 263508 273720 263520
rect 273772 263508 273778 263560
rect 285950 262828 285956 262880
rect 286008 262868 286014 262880
rect 546586 262868 546592 262880
rect 286008 262840 546592 262868
rect 286008 262828 286014 262840
rect 546586 262828 546592 262840
rect 546644 262828 546650 262880
rect 286042 261468 286048 261520
rect 286100 261508 286106 261520
rect 549254 261508 549260 261520
rect 286100 261480 549260 261508
rect 286100 261468 286106 261480
rect 549254 261468 549260 261480
rect 549312 261468 549318 261520
rect 235166 260896 235172 260908
rect 235127 260868 235172 260896
rect 235166 260856 235172 260868
rect 235224 260856 235230 260908
rect 257154 260856 257160 260908
rect 257212 260896 257218 260908
rect 257246 260896 257252 260908
rect 257212 260868 257252 260896
rect 257212 260856 257218 260868
rect 257246 260856 257252 260868
rect 257304 260856 257310 260908
rect 229554 260828 229560 260840
rect 229515 260800 229560 260828
rect 229554 260788 229560 260800
rect 229612 260788 229618 260840
rect 250438 260788 250444 260840
rect 250496 260828 250502 260840
rect 250717 260831 250775 260837
rect 250717 260828 250729 260831
rect 250496 260800 250729 260828
rect 250496 260788 250502 260800
rect 250717 260797 250729 260800
rect 250763 260797 250775 260831
rect 250717 260791 250775 260797
rect 286134 260108 286140 260160
rect 286192 260148 286198 260160
rect 553394 260148 553400 260160
rect 286192 260120 553400 260148
rect 286192 260108 286198 260120
rect 553394 260108 553400 260120
rect 553452 260108 553458 260160
rect 235166 259400 235172 259412
rect 235127 259372 235172 259400
rect 235166 259360 235172 259372
rect 235224 259360 235230 259412
rect 287238 258680 287244 258732
rect 287296 258720 287302 258732
rect 560294 258720 560300 258732
rect 287296 258692 560300 258720
rect 287296 258680 287302 258692
rect 560294 258680 560300 258692
rect 560352 258680 560358 258732
rect 287330 257320 287336 257372
rect 287388 257360 287394 257372
rect 563146 257360 563152 257372
rect 287388 257332 563152 257360
rect 287388 257320 287394 257332
rect 563146 257320 563152 257332
rect 563204 257320 563210 257372
rect 277026 256748 277032 256760
rect 276987 256720 277032 256748
rect 277026 256708 277032 256720
rect 277084 256708 277090 256760
rect 276934 256680 276940 256692
rect 276895 256652 276940 256680
rect 276934 256640 276940 256652
rect 276992 256640 276998 256692
rect 291102 255960 291108 256012
rect 291160 256000 291166 256012
rect 471238 256000 471244 256012
rect 291160 255972 471244 256000
rect 291160 255960 291166 255972
rect 471238 255960 471244 255972
rect 471296 255960 471302 256012
rect 255774 255252 255780 255264
rect 255735 255224 255780 255252
rect 255774 255212 255780 255224
rect 255832 255212 255838 255264
rect 259914 255252 259920 255264
rect 259875 255224 259920 255252
rect 259914 255212 259920 255224
rect 259972 255212 259978 255264
rect 277210 255252 277216 255264
rect 277171 255224 277216 255252
rect 277210 255212 277216 255224
rect 277268 255212 277274 255264
rect 237006 253852 237012 253904
rect 237064 253892 237070 253904
rect 237190 253892 237196 253904
rect 237064 253864 237196 253892
rect 237064 253852 237070 253864
rect 237190 253852 237196 253864
rect 237248 253852 237254 253904
rect 250714 253824 250720 253836
rect 250675 253796 250720 253824
rect 250714 253784 250720 253796
rect 250772 253784 250778 253836
rect 3418 252492 3424 252544
rect 3476 252532 3482 252544
rect 225782 252532 225788 252544
rect 3476 252504 225788 252532
rect 3476 252492 3482 252504
rect 225782 252492 225788 252504
rect 225840 252492 225846 252544
rect 301590 252492 301596 252544
rect 301648 252532 301654 252544
rect 579798 252532 579804 252544
rect 301648 252504 579804 252532
rect 301648 252492 301654 252504
rect 579798 252492 579804 252504
rect 579856 252492 579862 252544
rect 252189 251311 252247 251317
rect 252189 251277 252201 251311
rect 252235 251308 252247 251311
rect 252278 251308 252284 251320
rect 252235 251280 252284 251308
rect 252235 251277 252247 251280
rect 252189 251271 252247 251277
rect 252278 251268 252284 251280
rect 252336 251268 252342 251320
rect 229557 251243 229615 251249
rect 229557 251209 229569 251243
rect 229603 251240 229615 251243
rect 229646 251240 229652 251252
rect 229603 251212 229652 251240
rect 229603 251209 229615 251212
rect 229557 251203 229615 251209
rect 229646 251200 229652 251212
rect 229704 251200 229710 251252
rect 254854 251240 254860 251252
rect 254815 251212 254860 251240
rect 254854 251200 254860 251212
rect 254912 251200 254918 251252
rect 273714 251200 273720 251252
rect 273772 251200 273778 251252
rect 237101 251175 237159 251181
rect 237101 251141 237113 251175
rect 237147 251172 237159 251175
rect 237190 251172 237196 251184
rect 237147 251144 237196 251172
rect 237147 251141 237159 251144
rect 237101 251135 237159 251141
rect 237190 251132 237196 251144
rect 237248 251132 237254 251184
rect 273732 251104 273760 251200
rect 273806 251104 273812 251116
rect 273732 251076 273812 251104
rect 273806 251064 273812 251076
rect 273864 251064 273870 251116
rect 252186 249812 252192 249824
rect 252147 249784 252192 249812
rect 252186 249772 252192 249784
rect 252244 249772 252250 249824
rect 254854 249812 254860 249824
rect 254815 249784 254860 249812
rect 254854 249772 254860 249784
rect 254912 249772 254918 249824
rect 256970 249772 256976 249824
rect 257028 249812 257034 249824
rect 257246 249812 257252 249824
rect 257028 249784 257252 249812
rect 257028 249772 257034 249784
rect 257246 249772 257252 249784
rect 257304 249772 257310 249824
rect 274174 249772 274180 249824
rect 274232 249812 274238 249824
rect 274266 249812 274272 249824
rect 274232 249784 274272 249812
rect 274232 249772 274238 249784
rect 274266 249772 274272 249784
rect 274324 249772 274330 249824
rect 276934 249744 276940 249756
rect 276895 249716 276940 249744
rect 276934 249704 276940 249716
rect 276992 249704 276998 249756
rect 260561 247027 260619 247033
rect 260561 246993 260573 247027
rect 260607 247024 260619 247027
rect 260650 247024 260656 247036
rect 260607 246996 260656 247024
rect 260607 246993 260619 246996
rect 260561 246987 260619 246993
rect 260650 246984 260656 246996
rect 260708 246984 260714 247036
rect 262490 246984 262496 247036
rect 262548 247024 262554 247036
rect 262674 247024 262680 247036
rect 262548 246996 262680 247024
rect 262548 246984 262554 246996
rect 262674 246984 262680 246996
rect 262732 246984 262738 247036
rect 274177 247027 274235 247033
rect 274177 246993 274189 247027
rect 274223 247024 274235 247027
rect 274266 247024 274272 247036
rect 274223 246996 274272 247024
rect 274223 246993 274235 246996
rect 274177 246987 274235 246993
rect 274266 246984 274272 246996
rect 274324 246984 274330 247036
rect 277210 247024 277216 247036
rect 277171 246996 277216 247024
rect 277210 246984 277216 246996
rect 277268 246984 277274 247036
rect 259914 245664 259920 245676
rect 259875 245636 259920 245664
rect 259914 245624 259920 245636
rect 259972 245624 259978 245676
rect 271506 245624 271512 245676
rect 271564 245664 271570 245676
rect 271782 245664 271788 245676
rect 271564 245636 271788 245664
rect 271564 245624 271570 245636
rect 271782 245624 271788 245636
rect 271840 245624 271846 245676
rect 233694 244264 233700 244316
rect 233752 244304 233758 244316
rect 233878 244304 233884 244316
rect 233752 244276 233884 244304
rect 233752 244264 233758 244276
rect 233878 244264 233884 244276
rect 233936 244264 233942 244316
rect 252094 244196 252100 244248
rect 252152 244236 252158 244248
rect 252278 244236 252284 244248
rect 252152 244208 252284 244236
rect 252152 244196 252158 244208
rect 252278 244196 252284 244208
rect 252336 244196 252342 244248
rect 235166 244032 235172 244044
rect 235127 244004 235172 244032
rect 235166 243992 235172 244004
rect 235224 243992 235230 244044
rect 237098 241516 237104 241528
rect 237059 241488 237104 241516
rect 237098 241476 237104 241488
rect 237156 241476 237162 241528
rect 273714 241476 273720 241528
rect 273772 241516 273778 241528
rect 273806 241516 273812 241528
rect 273772 241488 273812 241516
rect 273772 241476 273778 241488
rect 273806 241476 273812 241488
rect 273864 241476 273870 241528
rect 277210 241516 277216 241528
rect 277171 241488 277216 241516
rect 277210 241476 277216 241488
rect 277268 241476 277274 241528
rect 238938 241448 238944 241460
rect 238899 241420 238944 241448
rect 238938 241408 238944 241420
rect 238996 241408 239002 241460
rect 256510 238688 256516 238740
rect 256568 238728 256574 238740
rect 256602 238728 256608 238740
rect 256568 238700 256608 238728
rect 256568 238688 256574 238700
rect 256602 238688 256608 238700
rect 256660 238688 256666 238740
rect 255777 237439 255835 237445
rect 255777 237405 255789 237439
rect 255823 237436 255835 237439
rect 255866 237436 255872 237448
rect 255823 237408 255872 237436
rect 255823 237405 255835 237408
rect 255777 237399 255835 237405
rect 255866 237396 255872 237408
rect 255924 237396 255930 237448
rect 260558 237436 260564 237448
rect 260519 237408 260564 237436
rect 260558 237396 260564 237408
rect 260616 237396 260622 237448
rect 271598 237396 271604 237448
rect 271656 237436 271662 237448
rect 271782 237436 271788 237448
rect 271656 237408 271788 237436
rect 271656 237396 271662 237408
rect 271782 237396 271788 237408
rect 271840 237396 271846 237448
rect 274174 237436 274180 237448
rect 274135 237408 274180 237436
rect 274174 237396 274180 237408
rect 274232 237396 274238 237448
rect 277210 237436 277216 237448
rect 277171 237408 277216 237436
rect 277210 237396 277216 237408
rect 277268 237396 277274 237448
rect 264238 237368 264244 237380
rect 264199 237340 264244 237368
rect 264238 237328 264244 237340
rect 264296 237328 264302 237380
rect 262493 234719 262551 234725
rect 262493 234685 262505 234719
rect 262539 234716 262551 234719
rect 262674 234716 262680 234728
rect 262539 234688 262680 234716
rect 262539 234685 262551 234688
rect 262493 234679 262551 234685
rect 262674 234676 262680 234688
rect 262732 234676 262738 234728
rect 250714 234608 250720 234660
rect 250772 234608 250778 234660
rect 243354 234540 243360 234592
rect 243412 234580 243418 234592
rect 243538 234580 243544 234592
rect 243412 234552 243544 234580
rect 243412 234540 243418 234552
rect 243538 234540 243544 234552
rect 243596 234540 243602 234592
rect 250732 234524 250760 234608
rect 250714 234472 250720 234524
rect 250772 234472 250778 234524
rect 229646 231820 229652 231872
rect 229704 231860 229710 231872
rect 229830 231860 229836 231872
rect 229704 231832 229836 231860
rect 229704 231820 229710 231832
rect 229830 231820 229836 231832
rect 229888 231820 229894 231872
rect 234982 231820 234988 231872
rect 235040 231860 235046 231872
rect 235258 231860 235264 231872
rect 235040 231832 235264 231860
rect 235040 231820 235046 231832
rect 235258 231820 235264 231832
rect 235316 231820 235322 231872
rect 238938 231860 238944 231872
rect 238899 231832 238944 231860
rect 238938 231820 238944 231832
rect 238996 231820 239002 231872
rect 235534 230460 235540 230512
rect 235592 230500 235598 230512
rect 235718 230500 235724 230512
rect 235592 230472 235724 230500
rect 235592 230460 235598 230472
rect 235718 230460 235724 230472
rect 235776 230460 235782 230512
rect 262490 229072 262496 229084
rect 262451 229044 262496 229072
rect 262490 229032 262496 229044
rect 262548 229032 262554 229084
rect 274174 229032 274180 229084
rect 274232 229032 274238 229084
rect 276934 229032 276940 229084
rect 276992 229072 276998 229084
rect 277026 229072 277032 229084
rect 276992 229044 277032 229072
rect 276992 229032 276998 229044
rect 277026 229032 277032 229044
rect 277084 229032 277090 229084
rect 274192 229004 274220 229032
rect 274358 229004 274364 229016
rect 274192 228976 274364 229004
rect 274358 228964 274364 228976
rect 274416 228964 274422 229016
rect 328454 228080 328460 228132
rect 328512 228080 328518 228132
rect 328472 227928 328500 228080
rect 418062 227944 418068 227996
rect 418120 227984 418126 227996
rect 424962 227984 424968 227996
rect 418120 227956 424968 227984
rect 418120 227944 418126 227956
rect 424962 227944 424968 227956
rect 425020 227944 425026 227996
rect 328454 227876 328460 227928
rect 328512 227876 328518 227928
rect 495342 227876 495348 227928
rect 495400 227916 495406 227928
rect 496998 227916 497004 227928
rect 495400 227888 497004 227916
rect 495400 227876 495406 227888
rect 496998 227876 497004 227888
rect 497056 227876 497062 227928
rect 553302 227876 553308 227928
rect 553360 227916 553366 227928
rect 554590 227916 554596 227928
rect 553360 227888 554596 227916
rect 553360 227876 553366 227888
rect 554590 227876 554596 227888
rect 554648 227876 554654 227928
rect 437382 227808 437388 227860
rect 437440 227848 437446 227860
rect 444282 227848 444288 227860
rect 437440 227820 444288 227848
rect 437440 227808 437446 227820
rect 444282 227808 444288 227820
rect 444340 227808 444346 227860
rect 476022 227808 476028 227860
rect 476080 227848 476086 227860
rect 482922 227848 482928 227860
rect 476080 227820 482928 227848
rect 476080 227808 476086 227820
rect 482922 227808 482928 227820
rect 482980 227808 482986 227860
rect 514662 227808 514668 227860
rect 514720 227848 514726 227860
rect 521562 227848 521568 227860
rect 514720 227820 521568 227848
rect 514720 227808 514726 227820
rect 521562 227808 521568 227820
rect 521620 227808 521626 227860
rect 278682 227740 278688 227792
rect 278740 227780 278746 227792
rect 289722 227780 289728 227792
rect 278740 227752 289728 227780
rect 278740 227740 278746 227752
rect 289722 227740 289728 227752
rect 289780 227740 289786 227792
rect 309134 227740 309140 227792
rect 309192 227780 309198 227792
rect 312630 227780 312636 227792
rect 309192 227752 312636 227780
rect 309192 227740 309198 227752
rect 312630 227740 312636 227752
rect 312688 227740 312694 227792
rect 533982 227740 533988 227792
rect 534040 227780 534046 227792
rect 540882 227780 540888 227792
rect 534040 227752 540888 227780
rect 534040 227740 534046 227752
rect 540882 227740 540888 227752
rect 540940 227740 540946 227792
rect 233694 224952 233700 225004
rect 233752 224992 233758 225004
rect 233878 224992 233884 225004
rect 233752 224964 233884 224992
rect 233752 224952 233758 224964
rect 233878 224952 233884 224964
rect 233936 224952 233942 225004
rect 3142 223524 3148 223576
rect 3200 223564 3206 223576
rect 207658 223564 207664 223576
rect 3200 223536 207664 223564
rect 3200 223524 3206 223536
rect 207658 223524 207664 223536
rect 207716 223524 207722 223576
rect 235166 222164 235172 222216
rect 235224 222204 235230 222216
rect 235350 222204 235356 222216
rect 235224 222176 235356 222204
rect 235224 222164 235230 222176
rect 235350 222164 235356 222176
rect 235408 222164 235414 222216
rect 254762 222164 254768 222216
rect 254820 222164 254826 222216
rect 254780 222136 254808 222164
rect 254854 222136 254860 222148
rect 254780 222108 254860 222136
rect 254854 222096 254860 222108
rect 254912 222096 254918 222148
rect 256602 220912 256608 220924
rect 256436 220884 256608 220912
rect 256436 220788 256464 220884
rect 256602 220872 256608 220884
rect 256660 220872 256666 220924
rect 256418 220736 256424 220788
rect 256476 220736 256482 220788
rect 255866 219512 255872 219564
rect 255924 219552 255930 219564
rect 256050 219552 256056 219564
rect 255924 219524 256056 219552
rect 255924 219512 255930 219524
rect 256050 219512 256056 219524
rect 256108 219512 256114 219564
rect 260742 219484 260748 219496
rect 260668 219456 260748 219484
rect 260668 219428 260696 219456
rect 260742 219444 260748 219456
rect 260800 219444 260806 219496
rect 264238 219484 264244 219496
rect 264199 219456 264244 219484
rect 264238 219444 264244 219456
rect 264296 219444 264302 219496
rect 260650 219376 260656 219428
rect 260708 219376 260714 219428
rect 255866 217988 255872 218000
rect 255827 217960 255872 217988
rect 255866 217948 255872 217960
rect 255924 217948 255930 218000
rect 260650 217948 260656 218000
rect 260708 217988 260714 218000
rect 260926 217988 260932 218000
rect 260708 217960 260932 217988
rect 260708 217948 260714 217960
rect 260926 217948 260932 217960
rect 260984 217948 260990 218000
rect 262674 217988 262680 218000
rect 262635 217960 262680 217988
rect 262674 217948 262680 217960
rect 262732 217948 262738 218000
rect 264238 217988 264244 218000
rect 264199 217960 264244 217988
rect 264238 217948 264244 217960
rect 264296 217948 264302 218000
rect 413278 217948 413284 218000
rect 413336 217988 413342 218000
rect 580166 217988 580172 218000
rect 413336 217960 580172 217988
rect 413336 217948 413342 217960
rect 580166 217948 580172 217960
rect 580224 217948 580230 218000
rect 243538 215404 243544 215416
rect 243372 215376 243544 215404
rect 243372 215348 243400 215376
rect 243538 215364 243544 215376
rect 243596 215364 243602 215416
rect 243354 215296 243360 215348
rect 243412 215296 243418 215348
rect 274174 213936 274180 213988
rect 274232 213976 274238 213988
rect 274358 213976 274364 213988
rect 274232 213948 274364 213976
rect 274232 213936 274238 213948
rect 274358 213936 274364 213948
rect 274416 213936 274422 213988
rect 277578 212712 277584 212764
rect 277636 212752 277642 212764
rect 277946 212752 277952 212764
rect 277636 212724 277952 212752
rect 277636 212712 277642 212724
rect 277946 212712 277952 212724
rect 278004 212712 278010 212764
rect 229646 212508 229652 212560
rect 229704 212548 229710 212560
rect 229830 212548 229836 212560
rect 229704 212520 229836 212548
rect 229704 212508 229710 212520
rect 229830 212508 229836 212520
rect 229888 212508 229894 212560
rect 237006 212508 237012 212560
rect 237064 212508 237070 212560
rect 245010 212508 245016 212560
rect 245068 212548 245074 212560
rect 245194 212548 245200 212560
rect 245068 212520 245200 212548
rect 245068 212508 245074 212520
rect 245194 212508 245200 212520
rect 245252 212508 245258 212560
rect 237024 212424 237052 212508
rect 237006 212372 237012 212424
rect 237064 212372 237070 212424
rect 277118 209720 277124 209772
rect 277176 209760 277182 209772
rect 277210 209760 277216 209772
rect 277176 209732 277216 209760
rect 277176 209720 277182 209732
rect 277210 209720 277216 209732
rect 277268 209720 277274 209772
rect 255866 208400 255872 208412
rect 255827 208372 255872 208400
rect 255866 208360 255872 208372
rect 255924 208360 255930 208412
rect 264241 208403 264299 208409
rect 264241 208369 264253 208403
rect 264287 208400 264299 208403
rect 264422 208400 264428 208412
rect 264287 208372 264428 208400
rect 264287 208369 264299 208372
rect 264241 208363 264299 208369
rect 264422 208360 264428 208372
rect 264480 208360 264486 208412
rect 3418 208292 3424 208344
rect 3476 208332 3482 208344
rect 222930 208332 222936 208344
rect 3476 208304 222936 208332
rect 3476 208292 3482 208304
rect 222930 208292 222936 208304
rect 222988 208292 222994 208344
rect 252186 208332 252192 208344
rect 252147 208304 252192 208332
rect 252186 208292 252192 208304
rect 252244 208292 252250 208344
rect 277118 208292 277124 208344
rect 277176 208332 277182 208344
rect 277210 208332 277216 208344
rect 277176 208304 277216 208332
rect 277176 208292 277182 208304
rect 277210 208292 277216 208304
rect 277268 208292 277274 208344
rect 233694 205640 233700 205692
rect 233752 205680 233758 205692
rect 233878 205680 233884 205692
rect 233752 205652 233884 205680
rect 233752 205640 233758 205652
rect 233878 205640 233884 205652
rect 233936 205640 233942 205692
rect 259822 205640 259828 205692
rect 259880 205640 259886 205692
rect 259840 205612 259868 205640
rect 259914 205612 259920 205624
rect 259840 205584 259920 205612
rect 259914 205572 259920 205584
rect 259972 205572 259978 205624
rect 298830 205572 298836 205624
rect 298888 205612 298894 205624
rect 579798 205612 579804 205624
rect 298888 205584 579804 205612
rect 298888 205572 298894 205584
rect 579798 205572 579804 205584
rect 579856 205572 579862 205624
rect 235534 202852 235540 202904
rect 235592 202892 235598 202904
rect 235626 202892 235632 202904
rect 235592 202864 235632 202892
rect 235592 202852 235598 202864
rect 235626 202852 235632 202864
rect 235684 202852 235690 202904
rect 254854 202852 254860 202904
rect 254912 202892 254918 202904
rect 254946 202892 254952 202904
rect 254912 202864 254952 202892
rect 254912 202852 254918 202864
rect 254946 202852 254952 202864
rect 255004 202852 255010 202904
rect 273898 202852 273904 202904
rect 273956 202892 273962 202904
rect 273990 202892 273996 202904
rect 273956 202864 273996 202892
rect 273956 202852 273962 202864
rect 273990 202852 273996 202864
rect 274048 202852 274054 202904
rect 235166 202784 235172 202836
rect 235224 202824 235230 202836
rect 235258 202824 235264 202836
rect 235224 202796 235264 202824
rect 235224 202784 235230 202796
rect 235258 202784 235264 202796
rect 235316 202784 235322 202836
rect 237098 202784 237104 202836
rect 237156 202824 237162 202836
rect 237190 202824 237196 202836
rect 237156 202796 237196 202824
rect 237156 202784 237162 202796
rect 237190 202784 237196 202796
rect 237248 202784 237254 202836
rect 238938 202824 238944 202836
rect 238899 202796 238944 202824
rect 238938 202784 238944 202796
rect 238996 202784 239002 202836
rect 235258 201424 235264 201476
rect 235316 201424 235322 201476
rect 234982 201356 234988 201408
rect 235040 201396 235046 201408
rect 235276 201396 235304 201424
rect 235040 201368 235304 201396
rect 235040 201356 235046 201368
rect 268838 200064 268844 200116
rect 268896 200104 268902 200116
rect 269022 200104 269028 200116
rect 268896 200076 269028 200104
rect 268896 200064 268902 200076
rect 269022 200064 269028 200076
rect 269080 200064 269086 200116
rect 274174 200064 274180 200116
rect 274232 200064 274238 200116
rect 274192 200036 274220 200064
rect 274266 200036 274272 200048
rect 274192 200008 274272 200036
rect 274266 199996 274272 200008
rect 274324 199996 274330 200048
rect 252189 198747 252247 198753
rect 252189 198713 252201 198747
rect 252235 198744 252247 198747
rect 252278 198744 252284 198756
rect 252235 198716 252284 198744
rect 252235 198713 252247 198716
rect 252189 198707 252247 198713
rect 252278 198704 252284 198716
rect 252336 198704 252342 198756
rect 262674 198744 262680 198756
rect 262635 198716 262680 198744
rect 262674 198704 262680 198716
rect 262732 198704 262738 198756
rect 264238 198704 264244 198756
rect 264296 198744 264302 198756
rect 264422 198744 264428 198756
rect 264296 198716 264428 198744
rect 264296 198704 264302 198716
rect 264422 198704 264428 198716
rect 264480 198704 264486 198756
rect 255777 198679 255835 198685
rect 255777 198645 255789 198679
rect 255823 198676 255835 198679
rect 255866 198676 255872 198688
rect 255823 198648 255872 198676
rect 255823 198645 255835 198648
rect 255777 198639 255835 198645
rect 255866 198636 255872 198648
rect 255924 198636 255930 198688
rect 260650 198636 260656 198688
rect 260708 198676 260714 198688
rect 260742 198676 260748 198688
rect 260708 198648 260748 198676
rect 260708 198636 260714 198648
rect 260742 198636 260748 198648
rect 260800 198636 260806 198688
rect 260650 197276 260656 197328
rect 260708 197276 260714 197328
rect 277118 197316 277124 197328
rect 277079 197288 277124 197316
rect 277118 197276 277124 197288
rect 277176 197276 277182 197328
rect 260668 197189 260696 197276
rect 260653 197183 260711 197189
rect 260653 197149 260665 197183
rect 260699 197149 260711 197183
rect 260653 197143 260711 197149
rect 271598 195956 271604 195968
rect 271559 195928 271604 195956
rect 271598 195916 271604 195928
rect 271656 195916 271662 195968
rect 277762 195916 277768 195968
rect 277820 195916 277826 195968
rect 277780 195888 277808 195916
rect 277946 195888 277952 195900
rect 277780 195860 277952 195888
rect 277946 195848 277952 195860
rect 278004 195848 278010 195900
rect 229646 193196 229652 193248
rect 229704 193236 229710 193248
rect 229830 193236 229836 193248
rect 229704 193208 229836 193236
rect 229704 193196 229710 193208
rect 229830 193196 229836 193208
rect 229888 193196 229894 193248
rect 235534 193196 235540 193248
rect 235592 193236 235598 193248
rect 235626 193236 235632 193248
rect 235592 193208 235632 193236
rect 235592 193196 235598 193208
rect 235626 193196 235632 193208
rect 235684 193196 235690 193248
rect 245010 193196 245016 193248
rect 245068 193236 245074 193248
rect 245194 193236 245200 193248
rect 245068 193208 245200 193236
rect 245068 193196 245074 193208
rect 245194 193196 245200 193208
rect 245252 193196 245258 193248
rect 238938 191876 238944 191888
rect 238899 191848 238944 191876
rect 238938 191836 238944 191848
rect 238996 191836 239002 191888
rect 255774 191332 255780 191344
rect 255735 191304 255780 191332
rect 255774 191292 255780 191304
rect 255832 191292 255838 191344
rect 252094 189048 252100 189100
rect 252152 189088 252158 189100
rect 252278 189088 252284 189100
rect 252152 189060 252284 189088
rect 252152 189048 252158 189060
rect 252278 189048 252284 189060
rect 252336 189048 252342 189100
rect 254762 189020 254768 189032
rect 254723 188992 254768 189020
rect 254762 188980 254768 188992
rect 254820 188980 254826 189032
rect 255774 189020 255780 189032
rect 255735 188992 255780 189020
rect 255774 188980 255780 188992
rect 255832 188980 255838 189032
rect 262674 189020 262680 189032
rect 262635 188992 262680 189020
rect 262674 188980 262680 188992
rect 262732 188980 262738 189032
rect 264238 189020 264244 189032
rect 264199 188992 264244 189020
rect 264238 188980 264244 188992
rect 264296 188980 264302 189032
rect 260650 187728 260656 187740
rect 260611 187700 260656 187728
rect 260650 187688 260656 187700
rect 260708 187688 260714 187740
rect 277118 187728 277124 187740
rect 277079 187700 277124 187728
rect 277118 187688 277124 187700
rect 277176 187688 277182 187740
rect 233694 186328 233700 186380
rect 233752 186368 233758 186380
rect 233878 186368 233884 186380
rect 233752 186340 233884 186368
rect 233752 186328 233758 186340
rect 233878 186328 233884 186340
rect 233936 186328 233942 186380
rect 271601 186371 271659 186377
rect 271601 186337 271613 186371
rect 271647 186368 271659 186371
rect 271690 186368 271696 186380
rect 271647 186340 271696 186368
rect 271647 186337 271659 186340
rect 271601 186331 271659 186337
rect 271690 186328 271696 186340
rect 271748 186328 271754 186380
rect 252094 186300 252100 186312
rect 252055 186272 252100 186300
rect 252094 186260 252100 186272
rect 252152 186260 252158 186312
rect 273809 184263 273867 184269
rect 273809 184229 273821 184263
rect 273855 184260 273867 184263
rect 273898 184260 273904 184272
rect 273855 184232 273904 184260
rect 273855 184229 273867 184232
rect 273809 184223 273867 184229
rect 273898 184220 273904 184232
rect 273956 184220 273962 184272
rect 255777 184195 255835 184201
rect 255777 184161 255789 184195
rect 255823 184192 255835 184195
rect 255866 184192 255872 184204
rect 255823 184164 255872 184192
rect 255823 184161 255835 184164
rect 255777 184155 255835 184161
rect 255866 184152 255872 184164
rect 255924 184152 255930 184204
rect 234982 183540 234988 183592
rect 235040 183580 235046 183592
rect 235166 183580 235172 183592
rect 235040 183552 235172 183580
rect 235040 183540 235046 183552
rect 235166 183540 235172 183552
rect 235224 183540 235230 183592
rect 273714 183540 273720 183592
rect 273772 183580 273778 183592
rect 273806 183580 273812 183592
rect 273772 183552 273812 183580
rect 273772 183540 273778 183552
rect 273806 183540 273812 183552
rect 273864 183540 273870 183592
rect 276934 183540 276940 183592
rect 276992 183580 276998 183592
rect 277026 183580 277032 183592
rect 276992 183552 277032 183580
rect 276992 183540 276998 183552
rect 277026 183540 277032 183552
rect 277084 183540 277090 183592
rect 277118 183540 277124 183592
rect 277176 183540 277182 183592
rect 237098 183472 237104 183524
rect 237156 183512 237162 183524
rect 237190 183512 237196 183524
rect 237156 183484 237196 183512
rect 237156 183472 237162 183484
rect 237190 183472 237196 183484
rect 237248 183472 237254 183524
rect 277136 183444 277164 183540
rect 277210 183444 277216 183456
rect 277136 183416 277216 183444
rect 277210 183404 277216 183416
rect 277268 183404 277274 183456
rect 284846 182792 284852 182844
rect 284904 182832 284910 182844
rect 538214 182832 538220 182844
rect 284904 182804 538220 182832
rect 284904 182792 284910 182804
rect 538214 182792 538220 182804
rect 538272 182792 538278 182844
rect 308398 182112 308404 182164
rect 308456 182152 308462 182164
rect 580166 182152 580172 182164
rect 308456 182124 580172 182152
rect 308456 182112 308462 182124
rect 580166 182112 580172 182124
rect 580224 182112 580230 182164
rect 3234 180752 3240 180804
rect 3292 180792 3298 180804
rect 204898 180792 204904 180804
rect 3292 180764 204904 180792
rect 3292 180752 3298 180764
rect 204898 180752 204904 180764
rect 204956 180752 204962 180804
rect 245010 180792 245016 180804
rect 244971 180764 245016 180792
rect 245010 180752 245016 180764
rect 245068 180752 245074 180804
rect 273806 180792 273812 180804
rect 273767 180764 273812 180792
rect 273806 180752 273812 180764
rect 273864 180752 273870 180804
rect 281442 180072 281448 180124
rect 281500 180112 281506 180124
rect 499574 180112 499580 180124
rect 281500 180084 499580 180112
rect 281500 180072 281506 180084
rect 499574 180072 499580 180084
rect 499632 180072 499638 180124
rect 254765 179435 254823 179441
rect 254765 179401 254777 179435
rect 254811 179432 254823 179435
rect 254946 179432 254952 179444
rect 254811 179404 254952 179432
rect 254811 179401 254823 179404
rect 254765 179395 254823 179401
rect 254946 179392 254952 179404
rect 255004 179392 255010 179444
rect 260650 179432 260656 179444
rect 260611 179404 260656 179432
rect 260650 179392 260656 179404
rect 260708 179392 260714 179444
rect 262674 179432 262680 179444
rect 262635 179404 262680 179432
rect 262674 179392 262680 179404
rect 262732 179392 262738 179444
rect 264238 179432 264244 179444
rect 264199 179404 264244 179432
rect 264238 179392 264244 179404
rect 264296 179392 264302 179444
rect 260650 178072 260656 178084
rect 260611 178044 260656 178072
rect 260650 178032 260656 178044
rect 260708 178032 260714 178084
rect 271598 178032 271604 178084
rect 271656 178072 271662 178084
rect 271690 178072 271696 178084
rect 271656 178044 271696 178072
rect 271656 178032 271662 178044
rect 271690 178032 271696 178044
rect 271748 178032 271754 178084
rect 268838 178004 268844 178016
rect 268799 177976 268844 178004
rect 268838 177964 268844 177976
rect 268896 177964 268902 178016
rect 277210 177964 277216 178016
rect 277268 178004 277274 178016
rect 277394 178004 277400 178016
rect 277268 177976 277400 178004
rect 277268 177964 277274 177976
rect 277394 177964 277400 177976
rect 277452 177964 277458 178016
rect 252097 176715 252155 176721
rect 252097 176681 252109 176715
rect 252143 176712 252155 176715
rect 252186 176712 252192 176724
rect 252143 176684 252192 176712
rect 252143 176681 252155 176684
rect 252097 176675 252155 176681
rect 252186 176672 252192 176684
rect 252244 176672 252250 176724
rect 252186 173992 252192 174004
rect 252147 173964 252192 173992
rect 252186 173952 252192 173964
rect 252244 173952 252250 174004
rect 229646 173884 229652 173936
rect 229704 173924 229710 173936
rect 229830 173924 229836 173936
rect 229704 173896 229836 173924
rect 229704 173884 229710 173896
rect 229830 173884 229836 173896
rect 229888 173884 229894 173936
rect 234982 173884 234988 173936
rect 235040 173924 235046 173936
rect 235258 173924 235264 173936
rect 235040 173896 235264 173924
rect 235040 173884 235046 173896
rect 235258 173884 235264 173896
rect 235316 173884 235322 173936
rect 235442 173884 235448 173936
rect 235500 173924 235506 173936
rect 235534 173924 235540 173936
rect 235500 173896 235540 173924
rect 235500 173884 235506 173896
rect 235534 173884 235540 173896
rect 235592 173884 235598 173936
rect 234982 172456 234988 172508
rect 235040 172496 235046 172508
rect 235258 172496 235264 172508
rect 235040 172468 235264 172496
rect 235040 172456 235046 172468
rect 235258 172456 235264 172468
rect 235316 172456 235322 172508
rect 245013 171139 245071 171145
rect 245013 171105 245025 171139
rect 245059 171136 245071 171139
rect 245286 171136 245292 171148
rect 245059 171108 245292 171136
rect 245059 171105 245071 171108
rect 245013 171099 245071 171105
rect 245286 171096 245292 171108
rect 245344 171096 245350 171148
rect 273806 171028 273812 171080
rect 273864 171068 273870 171080
rect 273898 171068 273904 171080
rect 273864 171040 273904 171068
rect 273864 171028 273870 171040
rect 273898 171028 273904 171040
rect 273956 171028 273962 171080
rect 493318 171028 493324 171080
rect 493376 171068 493382 171080
rect 580166 171068 580172 171080
rect 493376 171040 580172 171068
rect 493376 171028 493382 171040
rect 580166 171028 580172 171040
rect 580224 171028 580230 171080
rect 259914 169776 259920 169788
rect 259748 169748 259920 169776
rect 259748 169720 259776 169748
rect 259914 169736 259920 169748
rect 259972 169736 259978 169788
rect 259730 169668 259736 169720
rect 259788 169668 259794 169720
rect 262674 169708 262680 169720
rect 262635 169680 262680 169708
rect 262674 169668 262680 169680
rect 262732 169668 262738 169720
rect 264238 169708 264244 169720
rect 264199 169680 264244 169708
rect 264238 169668 264244 169680
rect 264296 169668 264302 169720
rect 257246 169056 257252 169108
rect 257304 169096 257310 169108
rect 257430 169096 257436 169108
rect 257304 169068 257436 169096
rect 257304 169056 257310 169068
rect 257430 169056 257436 169068
rect 257488 169056 257494 169108
rect 268841 168419 268899 168425
rect 268841 168385 268853 168419
rect 268887 168416 268899 168419
rect 268930 168416 268936 168428
rect 268887 168388 268936 168416
rect 268887 168385 268899 168388
rect 268841 168379 268899 168385
rect 268930 168376 268936 168388
rect 268988 168376 268994 168428
rect 252186 168348 252192 168360
rect 252147 168320 252192 168348
rect 252186 168308 252192 168320
rect 252244 168308 252250 168360
rect 254857 168351 254915 168357
rect 254857 168317 254869 168351
rect 254903 168348 254915 168351
rect 254946 168348 254952 168360
rect 254903 168320 254952 168348
rect 254903 168317 254915 168320
rect 254857 168311 254915 168317
rect 254946 168308 254952 168320
rect 255004 168308 255010 168360
rect 233694 167016 233700 167068
rect 233752 167056 233758 167068
rect 233878 167056 233884 167068
rect 233752 167028 233884 167056
rect 233752 167016 233758 167028
rect 233878 167016 233884 167028
rect 233936 167016 233942 167068
rect 3510 165520 3516 165572
rect 3568 165560 3574 165572
rect 218698 165560 218704 165572
rect 3568 165532 218704 165560
rect 3568 165520 3574 165532
rect 218698 165520 218704 165532
rect 218756 165520 218762 165572
rect 219250 164840 219256 164892
rect 219308 164880 219314 164892
rect 252186 164880 252192 164892
rect 219308 164852 252192 164880
rect 219308 164840 219314 164852
rect 252186 164840 252192 164852
rect 252244 164840 252250 164892
rect 273622 164228 273628 164280
rect 273680 164228 273686 164280
rect 229554 164160 229560 164212
rect 229612 164200 229618 164212
rect 229830 164200 229836 164212
rect 229612 164172 229836 164200
rect 229612 164160 229618 164172
rect 229830 164160 229836 164172
rect 229888 164160 229894 164212
rect 273640 164132 273668 164228
rect 273714 164132 273720 164144
rect 273640 164104 273720 164132
rect 273714 164092 273720 164104
rect 273772 164092 273778 164144
rect 238754 162800 238760 162852
rect 238812 162840 238818 162852
rect 238938 162840 238944 162852
rect 238812 162812 238944 162840
rect 238812 162800 238818 162812
rect 238938 162800 238944 162812
rect 238996 162800 239002 162852
rect 235166 162772 235172 162784
rect 235127 162744 235172 162772
rect 235166 162732 235172 162744
rect 235224 162732 235230 162784
rect 268838 161440 268844 161492
rect 268896 161480 268902 161492
rect 268930 161480 268936 161492
rect 268896 161452 268936 161480
rect 268896 161440 268902 161452
rect 268930 161440 268936 161452
rect 268988 161440 268994 161492
rect 245013 161415 245071 161421
rect 245013 161381 245025 161415
rect 245059 161412 245071 161415
rect 245286 161412 245292 161424
rect 245059 161384 245292 161412
rect 245059 161381 245071 161384
rect 245013 161375 245071 161381
rect 245286 161372 245292 161384
rect 245344 161372 245350 161424
rect 259730 160080 259736 160132
rect 259788 160120 259794 160132
rect 259914 160120 259920 160132
rect 259788 160092 259920 160120
rect 259788 160080 259794 160092
rect 259914 160080 259920 160092
rect 259972 160080 259978 160132
rect 262674 160120 262680 160132
rect 262635 160092 262680 160120
rect 262674 160080 262680 160092
rect 262732 160080 262738 160132
rect 264238 160120 264244 160132
rect 264199 160092 264244 160120
rect 264238 160080 264244 160092
rect 264296 160080 264302 160132
rect 276842 160080 276848 160132
rect 276900 160120 276906 160132
rect 277026 160120 277032 160132
rect 276900 160092 277032 160120
rect 276900 160080 276906 160092
rect 277026 160080 277032 160092
rect 277084 160080 277090 160132
rect 277118 160080 277124 160132
rect 277176 160120 277182 160132
rect 277394 160120 277400 160132
rect 277176 160092 277400 160120
rect 277176 160080 277182 160092
rect 277394 160080 277400 160092
rect 277452 160080 277458 160132
rect 268838 160052 268844 160064
rect 268799 160024 268844 160052
rect 268838 160012 268844 160024
rect 268896 160012 268902 160064
rect 271598 160052 271604 160064
rect 271559 160024 271604 160052
rect 271598 160012 271604 160024
rect 271656 160012 271662 160064
rect 274174 160012 274180 160064
rect 274232 160012 274238 160064
rect 274192 159928 274220 160012
rect 274174 159876 274180 159928
rect 274232 159876 274238 159928
rect 254854 158760 254860 158772
rect 254815 158732 254860 158760
rect 254854 158720 254860 158732
rect 254912 158720 254918 158772
rect 260558 158692 260564 158704
rect 260519 158664 260564 158692
rect 260558 158652 260564 158664
rect 260616 158652 260622 158704
rect 277118 158652 277124 158704
rect 277176 158692 277182 158704
rect 277210 158692 277216 158704
rect 277176 158664 277216 158692
rect 277176 158652 277182 158664
rect 277210 158652 277216 158664
rect 277268 158652 277274 158704
rect 297450 158652 297456 158704
rect 297508 158692 297514 158704
rect 579798 158692 579804 158704
rect 297508 158664 579804 158692
rect 297508 158652 297514 158664
rect 579798 158652 579804 158664
rect 579856 158652 579862 158704
rect 235166 157400 235172 157412
rect 235127 157372 235172 157400
rect 235166 157360 235172 157372
rect 235224 157360 235230 157412
rect 255866 157400 255872 157412
rect 255827 157372 255872 157400
rect 255866 157360 255872 157372
rect 255924 157360 255930 157412
rect 237006 157292 237012 157344
rect 237064 157332 237070 157344
rect 237190 157332 237196 157344
rect 237064 157304 237196 157332
rect 237064 157292 237070 157304
rect 237190 157292 237196 157304
rect 237248 157292 237254 157344
rect 257246 154680 257252 154692
rect 257172 154652 257252 154680
rect 257172 154556 257200 154652
rect 257246 154640 257252 154652
rect 257304 154640 257310 154692
rect 255866 154544 255872 154556
rect 255827 154516 255872 154544
rect 255866 154504 255872 154516
rect 255924 154504 255930 154556
rect 257154 154504 257160 154556
rect 257212 154504 257218 154556
rect 245010 151824 245016 151836
rect 244971 151796 245016 151824
rect 245010 151784 245016 151796
rect 245068 151784 245074 151836
rect 3142 151716 3148 151768
rect 3200 151756 3206 151768
rect 227070 151756 227076 151768
rect 3200 151728 227076 151756
rect 3200 151716 3206 151728
rect 227070 151716 227076 151728
rect 227128 151716 227134 151768
rect 254854 150424 254860 150476
rect 254912 150464 254918 150476
rect 255038 150464 255044 150476
rect 254912 150436 255044 150464
rect 254912 150424 254918 150436
rect 255038 150424 255044 150436
rect 255096 150424 255102 150476
rect 268841 150467 268899 150473
rect 268841 150433 268853 150467
rect 268887 150464 268899 150467
rect 268930 150464 268936 150476
rect 268887 150436 268936 150464
rect 268887 150433 268899 150436
rect 268841 150427 268899 150433
rect 268930 150424 268936 150436
rect 268988 150424 268994 150476
rect 271601 149175 271659 149181
rect 271601 149141 271613 149175
rect 271647 149172 271659 149175
rect 271690 149172 271696 149184
rect 271647 149144 271696 149172
rect 271647 149141 271659 149144
rect 271601 149135 271659 149141
rect 271690 149132 271696 149144
rect 271748 149132 271754 149184
rect 260561 149107 260619 149113
rect 260561 149073 260573 149107
rect 260607 149104 260619 149107
rect 260650 149104 260656 149116
rect 260607 149076 260656 149104
rect 260607 149073 260619 149076
rect 260561 149067 260619 149073
rect 260650 149064 260656 149076
rect 260708 149064 260714 149116
rect 271598 149036 271604 149048
rect 271559 149008 271604 149036
rect 271598 148996 271604 149008
rect 271656 148996 271662 149048
rect 277118 149036 277124 149048
rect 277079 149008 277124 149036
rect 277118 148996 277124 149008
rect 277176 148996 277182 149048
rect 259822 147636 259828 147688
rect 259880 147636 259886 147688
rect 259840 147608 259868 147636
rect 259914 147608 259920 147620
rect 259840 147580 259920 147608
rect 259914 147568 259920 147580
rect 259972 147568 259978 147620
rect 237098 144916 237104 144968
rect 237156 144956 237162 144968
rect 237190 144956 237196 144968
rect 237156 144928 237196 144956
rect 237156 144916 237162 144928
rect 237190 144916 237196 144928
rect 237248 144916 237254 144968
rect 235166 144848 235172 144900
rect 235224 144848 235230 144900
rect 235534 144888 235540 144900
rect 235495 144860 235540 144888
rect 235534 144848 235540 144860
rect 235592 144848 235598 144900
rect 235184 144820 235212 144848
rect 235258 144820 235264 144832
rect 235184 144792 235264 144820
rect 235258 144780 235264 144792
rect 235316 144780 235322 144832
rect 235258 143528 235264 143540
rect 235219 143500 235264 143528
rect 235258 143488 235264 143500
rect 235316 143488 235322 143540
rect 268838 142128 268844 142180
rect 268896 142168 268902 142180
rect 268930 142168 268936 142180
rect 268896 142140 268936 142168
rect 268896 142128 268902 142140
rect 268930 142128 268936 142140
rect 268988 142128 268994 142180
rect 273622 142128 273628 142180
rect 273680 142168 273686 142180
rect 273714 142168 273720 142180
rect 273680 142140 273720 142168
rect 273680 142128 273686 142140
rect 273714 142128 273720 142140
rect 273772 142128 273778 142180
rect 273806 142128 273812 142180
rect 273864 142168 273870 142180
rect 273898 142168 273904 142180
rect 273864 142140 273904 142168
rect 273864 142128 273870 142140
rect 273898 142128 273904 142140
rect 273956 142128 273962 142180
rect 250533 140743 250591 140749
rect 250533 140709 250545 140743
rect 250579 140740 250591 140743
rect 250622 140740 250628 140752
rect 250579 140712 250628 140740
rect 250579 140709 250591 140712
rect 250533 140703 250591 140709
rect 250622 140700 250628 140712
rect 250680 140700 250686 140752
rect 254946 140700 254952 140752
rect 255004 140740 255010 140752
rect 255038 140740 255044 140752
rect 255004 140712 255044 140740
rect 255004 140700 255010 140712
rect 255038 140700 255044 140712
rect 255096 140700 255102 140752
rect 260558 140740 260564 140752
rect 260519 140712 260564 140740
rect 260558 140700 260564 140712
rect 260616 140700 260622 140752
rect 262674 140740 262680 140752
rect 262635 140712 262680 140740
rect 262674 140700 262680 140712
rect 262732 140700 262738 140752
rect 264238 140740 264244 140752
rect 264199 140712 264244 140740
rect 264238 140700 264244 140712
rect 264296 140700 264302 140752
rect 271598 139516 271604 139528
rect 271559 139488 271604 139516
rect 271598 139476 271604 139488
rect 271656 139476 271662 139528
rect 277121 139451 277179 139457
rect 277121 139417 277133 139451
rect 277167 139448 277179 139451
rect 277210 139448 277216 139460
rect 277167 139420 277216 139448
rect 277167 139417 277179 139420
rect 277121 139411 277179 139417
rect 277210 139408 277216 139420
rect 277268 139408 277274 139460
rect 271509 139383 271567 139389
rect 271509 139349 271521 139383
rect 271555 139380 271567 139383
rect 271598 139380 271604 139392
rect 271555 139352 271604 139380
rect 271555 139349 271567 139352
rect 271509 139343 271567 139349
rect 271598 139340 271604 139352
rect 271656 139340 271662 139392
rect 245194 138700 245200 138712
rect 245155 138672 245200 138700
rect 245194 138660 245200 138672
rect 245252 138660 245258 138712
rect 229554 137980 229560 138032
rect 229612 137980 229618 138032
rect 237098 137980 237104 138032
rect 237156 137980 237162 138032
rect 229462 137912 229468 137964
rect 229520 137952 229526 137964
rect 229572 137952 229600 137980
rect 229520 137924 229600 137952
rect 237116 137952 237144 137980
rect 237190 137952 237196 137964
rect 237116 137924 237196 137952
rect 229520 137912 229526 137924
rect 237190 137912 237196 137924
rect 237248 137912 237254 137964
rect 3234 136552 3240 136604
rect 3292 136592 3298 136604
rect 17218 136592 17224 136604
rect 3292 136564 17224 136592
rect 3292 136552 3298 136564
rect 17218 136552 17224 136564
rect 17276 136552 17282 136604
rect 235534 135300 235540 135312
rect 235495 135272 235540 135300
rect 235534 135260 235540 135272
rect 235592 135260 235598 135312
rect 255866 135192 255872 135244
rect 255924 135232 255930 135244
rect 256050 135232 256056 135244
rect 255924 135204 256056 135232
rect 255924 135192 255930 135204
rect 256050 135192 256056 135204
rect 256108 135192 256114 135244
rect 319438 135192 319444 135244
rect 319496 135232 319502 135244
rect 580166 135232 580172 135244
rect 319496 135204 580172 135232
rect 319496 135192 319502 135204
rect 580166 135192 580172 135204
rect 580224 135192 580230 135244
rect 245197 135167 245255 135173
rect 245197 135133 245209 135167
rect 245243 135164 245255 135167
rect 245378 135164 245384 135176
rect 245243 135136 245384 135164
rect 245243 135133 245255 135136
rect 245197 135127 245255 135133
rect 245378 135124 245384 135136
rect 245436 135124 245442 135176
rect 235258 133940 235264 133952
rect 235219 133912 235264 133940
rect 235258 133900 235264 133912
rect 235316 133900 235322 133952
rect 273806 133832 273812 133884
rect 273864 133872 273870 133884
rect 273990 133872 273996 133884
rect 273864 133844 273996 133872
rect 273864 133832 273870 133844
rect 273990 133832 273996 133844
rect 274048 133832 274054 133884
rect 276934 132472 276940 132524
rect 276992 132512 276998 132524
rect 277026 132512 277032 132524
rect 276992 132484 277032 132512
rect 276992 132472 276998 132484
rect 277026 132472 277032 132484
rect 277084 132472 277090 132524
rect 262674 131152 262680 131164
rect 262635 131124 262680 131152
rect 262674 131112 262680 131124
rect 262732 131112 262738 131164
rect 264238 131152 264244 131164
rect 264199 131124 264244 131152
rect 264238 131112 264244 131124
rect 264296 131112 264302 131164
rect 274085 131087 274143 131093
rect 274085 131053 274097 131087
rect 274131 131084 274143 131087
rect 274174 131084 274180 131096
rect 274131 131056 274180 131084
rect 274131 131053 274143 131056
rect 274085 131047 274143 131053
rect 274174 131044 274180 131056
rect 274232 131044 274238 131096
rect 257154 130364 257160 130416
rect 257212 130364 257218 130416
rect 257172 130336 257200 130364
rect 257246 130336 257252 130348
rect 257172 130308 257252 130336
rect 257246 130296 257252 130308
rect 257304 130296 257310 130348
rect 260558 129792 260564 129804
rect 260519 129764 260564 129792
rect 260558 129752 260564 129764
rect 260616 129752 260622 129804
rect 271506 129752 271512 129804
rect 271564 129792 271570 129804
rect 271564 129764 271609 129792
rect 271564 129752 271570 129764
rect 233694 128324 233700 128376
rect 233752 128364 233758 128376
rect 233878 128364 233884 128376
rect 233752 128336 233884 128364
rect 233752 128324 233758 128336
rect 233878 128324 233884 128336
rect 233936 128324 233942 128376
rect 259822 128324 259828 128376
rect 259880 128324 259886 128376
rect 250530 128296 250536 128308
rect 250491 128268 250536 128296
rect 250530 128256 250536 128268
rect 250588 128256 250594 128308
rect 259840 128296 259868 128324
rect 259914 128296 259920 128308
rect 259840 128268 259920 128296
rect 259914 128256 259920 128268
rect 259972 128256 259978 128308
rect 254946 125644 254952 125656
rect 254872 125616 254952 125644
rect 254872 125588 254900 125616
rect 254946 125604 254952 125616
rect 255004 125604 255010 125656
rect 235534 125576 235540 125588
rect 235495 125548 235540 125576
rect 235534 125536 235540 125548
rect 235592 125536 235598 125588
rect 254854 125536 254860 125588
rect 254912 125536 254918 125588
rect 245102 125468 245108 125520
rect 245160 125508 245166 125520
rect 245378 125508 245384 125520
rect 245160 125480 245384 125508
rect 245160 125468 245166 125480
rect 245378 125468 245384 125480
rect 245436 125468 245442 125520
rect 250622 125468 250628 125520
rect 250680 125508 250686 125520
rect 250714 125508 250720 125520
rect 250680 125480 250720 125508
rect 250680 125468 250686 125480
rect 250714 125468 250720 125480
rect 250772 125468 250778 125520
rect 235258 124216 235264 124228
rect 235219 124188 235264 124216
rect 235258 124176 235264 124188
rect 235316 124176 235322 124228
rect 245102 124148 245108 124160
rect 245063 124120 245108 124148
rect 245102 124108 245108 124120
rect 245160 124108 245166 124160
rect 254854 124108 254860 124160
rect 254912 124148 254918 124160
rect 255130 124148 255136 124160
rect 254912 124120 255136 124148
rect 254912 124108 254918 124120
rect 255130 124108 255136 124120
rect 255188 124108 255194 124160
rect 255866 124108 255872 124160
rect 255924 124148 255930 124160
rect 256050 124148 256056 124160
rect 255924 124120 256056 124148
rect 255924 124108 255930 124120
rect 256050 124108 256056 124120
rect 256108 124108 256114 124160
rect 257246 124148 257252 124160
rect 257207 124120 257252 124148
rect 257246 124108 257252 124120
rect 257304 124108 257310 124160
rect 312538 124108 312544 124160
rect 312596 124148 312602 124160
rect 580166 124148 580172 124160
rect 312596 124120 580172 124148
rect 312596 124108 312602 124120
rect 580166 124108 580172 124120
rect 580224 124108 580230 124160
rect 235258 122856 235264 122868
rect 235219 122828 235264 122856
rect 235258 122816 235264 122828
rect 235316 122816 235322 122868
rect 3418 122748 3424 122800
rect 3476 122788 3482 122800
rect 215938 122788 215944 122800
rect 3476 122760 215944 122788
rect 3476 122748 3482 122760
rect 215938 122748 215944 122760
rect 215996 122748 216002 122800
rect 255041 122791 255099 122797
rect 255041 122757 255053 122791
rect 255087 122788 255099 122791
rect 255130 122788 255136 122800
rect 255087 122760 255136 122788
rect 255087 122757 255099 122760
rect 255041 122751 255099 122757
rect 255130 122748 255136 122760
rect 255188 122748 255194 122800
rect 274082 121496 274088 121508
rect 274043 121468 274088 121496
rect 274082 121456 274088 121468
rect 274140 121456 274146 121508
rect 268838 121428 268844 121440
rect 268799 121400 268844 121428
rect 268838 121388 268844 121400
rect 268896 121388 268902 121440
rect 273898 120068 273904 120080
rect 273859 120040 273904 120068
rect 273898 120028 273904 120040
rect 273956 120028 273962 120080
rect 229554 118668 229560 118720
rect 229612 118668 229618 118720
rect 237098 118668 237104 118720
rect 237156 118668 237162 118720
rect 229462 118600 229468 118652
rect 229520 118640 229526 118652
rect 229572 118640 229600 118668
rect 229520 118612 229600 118640
rect 237116 118640 237144 118668
rect 237190 118640 237196 118652
rect 237116 118612 237196 118640
rect 229520 118600 229526 118612
rect 237190 118600 237196 118612
rect 237248 118600 237254 118652
rect 235534 115988 235540 116000
rect 235495 115960 235540 115988
rect 235534 115948 235540 115960
rect 235592 115948 235598 116000
rect 277210 115988 277216 116000
rect 277171 115960 277216 115988
rect 277210 115948 277216 115960
rect 277268 115948 277274 116000
rect 259822 115880 259828 115932
rect 259880 115920 259886 115932
rect 259914 115920 259920 115932
rect 259880 115892 259920 115920
rect 259880 115880 259886 115892
rect 259914 115880 259920 115892
rect 259972 115880 259978 115932
rect 245102 114560 245108 114572
rect 245063 114532 245108 114560
rect 245102 114520 245108 114532
rect 245160 114520 245166 114572
rect 257246 114560 257252 114572
rect 257207 114532 257252 114560
rect 257246 114520 257252 114532
rect 257304 114520 257310 114572
rect 235258 114452 235264 114504
rect 235316 114492 235322 114504
rect 235350 114492 235356 114504
rect 235316 114464 235356 114492
rect 235316 114452 235322 114464
rect 235350 114452 235356 114464
rect 235408 114452 235414 114504
rect 255038 113200 255044 113212
rect 254999 113172 255044 113200
rect 255038 113160 255044 113172
rect 255096 113160 255102 113212
rect 268838 111908 268844 111920
rect 268799 111880 268844 111908
rect 268838 111868 268844 111880
rect 268896 111868 268902 111920
rect 274082 111800 274088 111852
rect 274140 111840 274146 111852
rect 274266 111840 274272 111852
rect 274140 111812 274272 111840
rect 274140 111800 274146 111812
rect 274266 111800 274272 111812
rect 274324 111800 274330 111852
rect 250625 111775 250683 111781
rect 250625 111741 250637 111775
rect 250671 111772 250683 111775
rect 250714 111772 250720 111784
rect 250671 111744 250720 111772
rect 250671 111741 250683 111744
rect 250625 111735 250683 111741
rect 250714 111732 250720 111744
rect 250772 111732 250778 111784
rect 260466 111732 260472 111784
rect 260524 111772 260530 111784
rect 260558 111772 260564 111784
rect 260524 111744 260564 111772
rect 260524 111732 260530 111744
rect 260558 111732 260564 111744
rect 260616 111732 260622 111784
rect 262674 111772 262680 111784
rect 262635 111744 262680 111772
rect 262674 111732 262680 111744
rect 262732 111732 262738 111784
rect 268838 111772 268844 111784
rect 268799 111744 268844 111772
rect 268838 111732 268844 111744
rect 268896 111732 268902 111784
rect 276934 111772 276940 111784
rect 276895 111744 276940 111772
rect 276934 111732 276940 111744
rect 276992 111732 276998 111784
rect 291930 111732 291936 111784
rect 291988 111772 291994 111784
rect 579798 111772 579804 111784
rect 291988 111744 579804 111772
rect 291988 111732 291994 111744
rect 579798 111732 579804 111744
rect 579856 111732 579862 111784
rect 273901 110483 273959 110489
rect 273901 110449 273913 110483
rect 273947 110480 273959 110483
rect 273990 110480 273996 110492
rect 273947 110452 273996 110480
rect 273947 110449 273959 110452
rect 273901 110443 273959 110449
rect 273990 110440 273996 110452
rect 274048 110440 274054 110492
rect 260466 110412 260472 110424
rect 260427 110384 260472 110412
rect 260466 110372 260472 110384
rect 260524 110372 260530 110424
rect 233694 109012 233700 109064
rect 233752 109052 233758 109064
rect 233878 109052 233884 109064
rect 233752 109024 233884 109052
rect 233752 109012 233758 109024
rect 233878 109012 233884 109024
rect 233936 109012 233942 109064
rect 245102 109012 245108 109064
rect 245160 109012 245166 109064
rect 245120 108984 245148 109012
rect 245194 108984 245200 108996
rect 245120 108956 245200 108984
rect 245194 108944 245200 108956
rect 245252 108944 245258 108996
rect 233786 104836 233792 104848
rect 233747 104808 233792 104836
rect 233786 104796 233792 104808
rect 233844 104796 233850 104848
rect 254854 104836 254860 104848
rect 254815 104808 254860 104836
rect 254854 104796 254860 104808
rect 254912 104796 254918 104848
rect 256510 104836 256516 104848
rect 256471 104808 256516 104836
rect 256510 104796 256516 104808
rect 256568 104796 256574 104848
rect 262674 102252 262680 102264
rect 262635 102224 262680 102252
rect 262674 102212 262680 102224
rect 262732 102212 262738 102264
rect 277210 102252 277216 102264
rect 277171 102224 277216 102252
rect 277210 102212 277216 102224
rect 277268 102212 277274 102264
rect 250622 102184 250628 102196
rect 250583 102156 250628 102184
rect 250622 102144 250628 102156
rect 250680 102144 250686 102196
rect 276937 102187 276995 102193
rect 276937 102153 276949 102187
rect 276983 102184 276995 102187
rect 277026 102184 277032 102196
rect 276983 102156 277032 102184
rect 276983 102153 276995 102156
rect 276937 102147 276995 102153
rect 277026 102144 277032 102156
rect 277084 102144 277090 102196
rect 260469 102119 260527 102125
rect 260469 102085 260481 102119
rect 260515 102116 260527 102119
rect 260558 102116 260564 102128
rect 260515 102088 260564 102116
rect 260515 102085 260527 102088
rect 260469 102079 260527 102085
rect 260558 102076 260564 102088
rect 260616 102076 260622 102128
rect 262674 102116 262680 102128
rect 262635 102088 262680 102116
rect 262674 102076 262680 102088
rect 262732 102076 262738 102128
rect 264238 102116 264244 102128
rect 264199 102088 264244 102116
rect 264238 102076 264244 102088
rect 264296 102076 264302 102128
rect 268838 100756 268844 100768
rect 268799 100728 268844 100756
rect 268838 100716 268844 100728
rect 268896 100716 268902 100768
rect 235350 99532 235356 99544
rect 235184 99504 235356 99532
rect 235184 99408 235212 99504
rect 235350 99492 235356 99504
rect 235408 99492 235414 99544
rect 229554 99356 229560 99408
rect 229612 99356 229618 99408
rect 235166 99356 235172 99408
rect 235224 99356 235230 99408
rect 229462 99288 229468 99340
rect 229520 99328 229526 99340
rect 229572 99328 229600 99356
rect 229520 99300 229600 99328
rect 229520 99288 229526 99300
rect 243354 99288 243360 99340
rect 243412 99328 243418 99340
rect 243538 99328 243544 99340
rect 243412 99300 243544 99328
rect 243412 99288 243418 99300
rect 243538 99288 243544 99300
rect 243596 99288 243602 99340
rect 274085 99331 274143 99337
rect 274085 99297 274097 99331
rect 274131 99328 274143 99331
rect 274174 99328 274180 99340
rect 274131 99300 274180 99328
rect 274131 99297 274143 99300
rect 274085 99291 274143 99297
rect 274174 99288 274180 99300
rect 274232 99288 274238 99340
rect 255866 98676 255872 98728
rect 255924 98716 255930 98728
rect 256050 98716 256056 98728
rect 255924 98688 256056 98716
rect 255924 98676 255930 98688
rect 256050 98676 256056 98688
rect 256108 98676 256114 98728
rect 233789 95251 233847 95257
rect 233789 95217 233801 95251
rect 233835 95248 233847 95251
rect 233970 95248 233976 95260
rect 233835 95220 233976 95248
rect 233835 95217 233847 95220
rect 233789 95211 233847 95217
rect 233970 95208 233976 95220
rect 234028 95208 234034 95260
rect 254857 95251 254915 95257
rect 254857 95217 254869 95251
rect 254903 95248 254915 95251
rect 255038 95248 255044 95260
rect 254903 95220 255044 95248
rect 254903 95217 254915 95220
rect 254857 95211 254915 95217
rect 255038 95208 255044 95220
rect 255096 95208 255102 95260
rect 256513 95251 256571 95257
rect 256513 95217 256525 95251
rect 256559 95248 256571 95251
rect 256694 95248 256700 95260
rect 256559 95220 256700 95248
rect 256559 95217 256571 95220
rect 256513 95211 256571 95217
rect 256694 95208 256700 95220
rect 256752 95208 256758 95260
rect 257246 95248 257252 95260
rect 257207 95220 257252 95248
rect 257246 95208 257252 95220
rect 257304 95208 257310 95260
rect 259914 95248 259920 95260
rect 259875 95220 259920 95248
rect 259914 95208 259920 95220
rect 259972 95208 259978 95260
rect 257246 93888 257252 93900
rect 257207 93860 257252 93888
rect 257246 93848 257252 93860
rect 257304 93848 257310 93900
rect 3418 93780 3424 93832
rect 3476 93820 3482 93832
rect 203518 93820 203524 93832
rect 3476 93792 203524 93820
rect 3476 93780 3482 93792
rect 203518 93780 203524 93792
rect 203576 93780 203582 93832
rect 259914 92528 259920 92540
rect 259875 92500 259920 92528
rect 259914 92488 259920 92500
rect 259972 92488 259978 92540
rect 264238 92528 264244 92540
rect 264199 92500 264244 92528
rect 264238 92488 264244 92500
rect 264296 92488 264302 92540
rect 268838 92460 268844 92472
rect 268799 92432 268844 92460
rect 268838 92420 268844 92432
rect 268896 92420 268902 92472
rect 273806 92420 273812 92472
rect 273864 92460 273870 92472
rect 273990 92460 273996 92472
rect 273864 92432 273996 92460
rect 273864 92420 273870 92432
rect 273990 92420 273996 92432
rect 274048 92420 274054 92472
rect 262582 91060 262588 91112
rect 262640 91100 262646 91112
rect 262677 91103 262735 91109
rect 262677 91100 262689 91103
rect 262640 91072 262689 91100
rect 262640 91060 262646 91072
rect 262677 91069 262689 91072
rect 262723 91069 262735 91103
rect 262677 91063 262735 91069
rect 276934 91060 276940 91112
rect 276992 91100 276998 91112
rect 277118 91100 277124 91112
rect 276992 91072 277124 91100
rect 276992 91060 276998 91072
rect 277118 91060 277124 91072
rect 277176 91060 277182 91112
rect 305638 88272 305644 88324
rect 305696 88312 305702 88324
rect 580166 88312 580172 88324
rect 305696 88284 580172 88312
rect 305696 88272 305702 88284
rect 580166 88272 580172 88284
rect 580224 88272 580230 88324
rect 268841 87091 268899 87097
rect 268841 87057 268853 87091
rect 268887 87088 268899 87091
rect 268930 87088 268936 87100
rect 268887 87060 268936 87088
rect 268887 87057 268899 87060
rect 268841 87051 268899 87057
rect 268930 87048 268936 87060
rect 268988 87048 268994 87100
rect 235166 86912 235172 86964
rect 235224 86952 235230 86964
rect 235258 86952 235264 86964
rect 235224 86924 235264 86952
rect 235224 86912 235230 86924
rect 235258 86912 235264 86924
rect 235316 86912 235322 86964
rect 235258 85524 235264 85536
rect 235219 85496 235264 85524
rect 235258 85484 235264 85496
rect 235316 85484 235322 85536
rect 237009 85527 237067 85533
rect 237009 85493 237021 85527
rect 237055 85524 237067 85527
rect 237190 85524 237196 85536
rect 237055 85496 237196 85524
rect 237055 85493 237067 85496
rect 237009 85487 237067 85493
rect 237190 85484 237196 85496
rect 237248 85484 237254 85536
rect 245194 85524 245200 85536
rect 245155 85496 245200 85524
rect 245194 85484 245200 85496
rect 245252 85484 245258 85536
rect 277118 84164 277124 84176
rect 277079 84136 277124 84164
rect 277118 84124 277124 84136
rect 277176 84124 277182 84176
rect 274085 82875 274143 82881
rect 274085 82841 274097 82875
rect 274131 82872 274143 82875
rect 274174 82872 274180 82884
rect 274131 82844 274180 82872
rect 274131 82841 274143 82844
rect 274085 82835 274143 82841
rect 274174 82832 274180 82844
rect 274232 82832 274238 82884
rect 250622 82764 250628 82816
rect 250680 82804 250686 82816
rect 250717 82807 250775 82813
rect 250717 82804 250729 82807
rect 250680 82776 250729 82804
rect 250680 82764 250686 82776
rect 250717 82773 250729 82776
rect 250763 82773 250775 82807
rect 250717 82767 250775 82773
rect 256418 82764 256424 82816
rect 256476 82804 256482 82816
rect 256602 82804 256608 82816
rect 256476 82776 256608 82804
rect 256476 82764 256482 82776
rect 256602 82764 256608 82776
rect 256660 82764 256666 82816
rect 264238 82804 264244 82816
rect 264199 82776 264244 82804
rect 264238 82764 264244 82776
rect 264296 82764 264302 82816
rect 254762 81404 254768 81456
rect 254820 81444 254826 81456
rect 254946 81444 254952 81456
rect 254820 81416 254952 81444
rect 254820 81404 254826 81416
rect 254946 81404 254952 81416
rect 255004 81404 255010 81456
rect 255774 81404 255780 81456
rect 255832 81444 255838 81456
rect 256050 81444 256056 81456
rect 255832 81416 256056 81444
rect 255832 81404 255838 81416
rect 256050 81404 256056 81416
rect 256108 81404 256114 81456
rect 259822 81404 259828 81456
rect 259880 81444 259886 81456
rect 259914 81444 259920 81456
rect 259880 81416 259920 81444
rect 259880 81404 259886 81416
rect 259914 81404 259920 81416
rect 259972 81404 259978 81456
rect 262582 81444 262588 81456
rect 262508 81416 262588 81444
rect 262508 81388 262536 81416
rect 262582 81404 262588 81416
rect 262640 81404 262646 81456
rect 262490 81336 262496 81388
rect 262548 81336 262554 81388
rect 229554 80044 229560 80096
rect 229612 80044 229618 80096
rect 3418 79976 3424 80028
rect 3476 80016 3482 80028
rect 214558 80016 214564 80028
rect 3476 79988 214564 80016
rect 3476 79976 3482 79988
rect 214558 79976 214564 79988
rect 214616 79976 214622 80028
rect 229572 80016 229600 80044
rect 229646 80016 229652 80028
rect 229572 79988 229652 80016
rect 229646 79976 229652 79988
rect 229704 79976 229710 80028
rect 233786 77256 233792 77308
rect 233844 77296 233850 77308
rect 233878 77296 233884 77308
rect 233844 77268 233884 77296
rect 233844 77256 233850 77268
rect 233878 77256 233884 77268
rect 233936 77256 233942 77308
rect 235442 77256 235448 77308
rect 235500 77296 235506 77308
rect 235534 77296 235540 77308
rect 235500 77268 235540 77296
rect 235500 77256 235506 77268
rect 235534 77256 235540 77268
rect 235592 77256 235598 77308
rect 229557 77231 229615 77237
rect 229557 77197 229569 77231
rect 229603 77228 229615 77231
rect 229646 77228 229652 77240
rect 229603 77200 229652 77228
rect 229603 77197 229615 77200
rect 229557 77191 229615 77197
rect 229646 77188 229652 77200
rect 229704 77188 229710 77240
rect 250898 77228 250904 77240
rect 250859 77200 250904 77228
rect 250898 77188 250904 77200
rect 250956 77188 250962 77240
rect 251082 77228 251088 77240
rect 251043 77200 251088 77228
rect 251082 77188 251088 77200
rect 251140 77188 251146 77240
rect 250990 77160 250996 77172
rect 250951 77132 250996 77160
rect 250990 77120 250996 77132
rect 251048 77120 251054 77172
rect 268930 76616 268936 76628
rect 268891 76588 268936 76616
rect 268930 76576 268936 76588
rect 268988 76576 268994 76628
rect 273901 76619 273959 76625
rect 273901 76585 273913 76619
rect 273947 76616 273959 76619
rect 274082 76616 274088 76628
rect 273947 76588 274088 76616
rect 273947 76585 273959 76588
rect 273901 76579 273959 76585
rect 274082 76576 274088 76588
rect 274140 76576 274146 76628
rect 274174 76576 274180 76628
rect 274232 76616 274238 76628
rect 274450 76616 274456 76628
rect 274232 76588 274456 76616
rect 274232 76576 274238 76588
rect 274450 76576 274456 76588
rect 274508 76576 274514 76628
rect 328454 76304 328460 76356
rect 328512 76304 328518 76356
rect 328472 76152 328500 76304
rect 328454 76100 328460 76152
rect 328512 76100 328518 76152
rect 553302 76100 553308 76152
rect 553360 76140 553366 76152
rect 554590 76140 554596 76152
rect 553360 76112 554596 76140
rect 553360 76100 553366 76112
rect 554590 76100 554596 76112
rect 554648 76100 554654 76152
rect 437382 76032 437388 76084
rect 437440 76072 437446 76084
rect 444282 76072 444288 76084
rect 437440 76044 444288 76072
rect 437440 76032 437446 76044
rect 444282 76032 444288 76044
rect 444340 76032 444346 76084
rect 502242 76032 502248 76084
rect 502300 76072 502306 76084
rect 510522 76072 510528 76084
rect 502300 76044 510528 76072
rect 502300 76032 502306 76044
rect 510522 76032 510528 76044
rect 510580 76032 510586 76084
rect 533982 76032 533988 76084
rect 534040 76072 534046 76084
rect 540882 76072 540888 76084
rect 534040 76044 540888 76072
rect 534040 76032 534046 76044
rect 540882 76032 540888 76044
rect 540940 76032 540946 76084
rect 237006 76004 237012 76016
rect 236967 75976 237012 76004
rect 237006 75964 237012 75976
rect 237064 75964 237070 76016
rect 309134 75964 309140 76016
rect 309192 76004 309198 76016
rect 313918 76004 313924 76016
rect 309192 75976 313924 76004
rect 309192 75964 309198 75976
rect 313918 75964 313924 75976
rect 313976 75964 313982 76016
rect 235258 75936 235264 75948
rect 235219 75908 235264 75936
rect 235258 75896 235264 75908
rect 235316 75896 235322 75948
rect 245194 75936 245200 75948
rect 245155 75908 245200 75936
rect 245194 75896 245200 75908
rect 245252 75896 245258 75948
rect 237006 75828 237012 75880
rect 237064 75868 237070 75880
rect 237193 75871 237251 75877
rect 237193 75868 237205 75871
rect 237064 75840 237205 75868
rect 237064 75828 237070 75840
rect 237193 75837 237205 75840
rect 237239 75837 237251 75871
rect 267458 75868 267464 75880
rect 267419 75840 267464 75868
rect 237193 75831 237251 75837
rect 267458 75828 267464 75840
rect 267516 75828 267522 75880
rect 264241 75803 264299 75809
rect 264241 75769 264253 75803
rect 264287 75800 264299 75803
rect 264330 75800 264336 75812
rect 264287 75772 264336 75800
rect 264287 75769 264299 75772
rect 264241 75763 264299 75769
rect 264330 75760 264336 75772
rect 264388 75760 264394 75812
rect 273622 74536 273628 74588
rect 273680 74576 273686 74588
rect 273714 74576 273720 74588
rect 273680 74548 273720 74576
rect 273680 74536 273686 74548
rect 273714 74536 273720 74548
rect 273772 74536 273778 74588
rect 277118 74576 277124 74588
rect 277079 74548 277124 74576
rect 277118 74536 277124 74548
rect 277176 74536 277182 74588
rect 256418 73148 256424 73160
rect 256379 73120 256424 73148
rect 256418 73108 256424 73120
rect 256476 73108 256482 73160
rect 259822 73108 259828 73160
rect 259880 73148 259886 73160
rect 260098 73148 260104 73160
rect 259880 73120 260104 73148
rect 259880 73108 259886 73120
rect 260098 73108 260104 73120
rect 260156 73108 260162 73160
rect 255774 73080 255780 73092
rect 255735 73052 255780 73080
rect 255774 73040 255780 73052
rect 255832 73040 255838 73092
rect 277118 73080 277124 73092
rect 277079 73052 277124 73080
rect 277118 73040 277124 73052
rect 277176 73040 277182 73092
rect 250898 72468 250904 72480
rect 250859 72440 250904 72468
rect 250898 72428 250904 72440
rect 250956 72428 250962 72480
rect 268933 71791 268991 71797
rect 268933 71757 268945 71791
rect 268979 71788 268991 71791
rect 269022 71788 269028 71800
rect 268979 71760 269028 71788
rect 268979 71757 268991 71760
rect 268933 71751 268991 71757
rect 269022 71748 269028 71760
rect 269080 71748 269086 71800
rect 250990 71720 250996 71732
rect 250951 71692 250996 71720
rect 250990 71680 250996 71692
rect 251048 71680 251054 71732
rect 235258 70496 235264 70508
rect 235184 70468 235264 70496
rect 235184 70372 235212 70468
rect 235258 70456 235264 70468
rect 235316 70456 235322 70508
rect 245105 70499 245163 70505
rect 245105 70465 245117 70499
rect 245151 70496 245163 70499
rect 245194 70496 245200 70508
rect 245151 70468 245200 70496
rect 245151 70465 245163 70468
rect 245105 70459 245163 70465
rect 245194 70456 245200 70468
rect 245252 70456 245258 70508
rect 243354 70388 243360 70440
rect 243412 70428 243418 70440
rect 243538 70428 243544 70440
rect 243412 70400 243544 70428
rect 243412 70388 243418 70400
rect 243538 70388 243544 70400
rect 243596 70388 243602 70440
rect 251082 70428 251088 70440
rect 251043 70400 251088 70428
rect 251082 70388 251088 70400
rect 251140 70388 251146 70440
rect 235166 70320 235172 70372
rect 235224 70320 235230 70372
rect 268838 68484 268844 68536
rect 268896 68524 268902 68536
rect 269022 68524 269028 68536
rect 268896 68496 269028 68524
rect 268896 68484 268902 68496
rect 269022 68484 269028 68496
rect 269080 68484 269086 68536
rect 257157 68391 257215 68397
rect 257157 68357 257169 68391
rect 257203 68388 257215 68391
rect 257246 68388 257252 68400
rect 257203 68360 257252 68388
rect 257203 68357 257215 68360
rect 257157 68351 257215 68357
rect 257246 68348 257252 68360
rect 257304 68348 257310 68400
rect 250438 68280 250444 68332
rect 250496 68320 250502 68332
rect 250717 68323 250775 68329
rect 250717 68320 250729 68323
rect 250496 68292 250729 68320
rect 250496 68280 250502 68292
rect 250717 68289 250729 68292
rect 250763 68289 250775 68323
rect 250717 68283 250775 68289
rect 229554 67640 229560 67652
rect 229515 67612 229560 67640
rect 229554 67600 229560 67612
rect 229612 67600 229618 67652
rect 233786 67600 233792 67652
rect 233844 67640 233850 67652
rect 233878 67640 233884 67652
rect 233844 67612 233884 67640
rect 233844 67600 233850 67612
rect 233878 67600 233884 67612
rect 233936 67600 233942 67652
rect 245102 67640 245108 67652
rect 245063 67612 245108 67640
rect 245102 67600 245108 67612
rect 245160 67600 245166 67652
rect 235534 67572 235540 67584
rect 235495 67544 235540 67572
rect 235534 67532 235540 67544
rect 235592 67532 235598 67584
rect 273622 66308 273628 66360
rect 273680 66308 273686 66360
rect 264238 66240 264244 66292
rect 264296 66280 264302 66292
rect 264330 66280 264336 66292
rect 264296 66252 264336 66280
rect 264296 66240 264302 66252
rect 264330 66240 264336 66252
rect 264388 66240 264394 66292
rect 267458 66280 267464 66292
rect 267419 66252 267464 66280
rect 267458 66240 267464 66252
rect 267516 66240 267522 66292
rect 273640 66224 273668 66308
rect 271138 66172 271144 66224
rect 271196 66212 271202 66224
rect 271230 66212 271236 66224
rect 271196 66184 271236 66212
rect 271196 66172 271202 66184
rect 271230 66172 271236 66184
rect 271288 66172 271294 66224
rect 273622 66172 273628 66224
rect 273680 66172 273686 66224
rect 3326 64812 3332 64864
rect 3384 64852 3390 64864
rect 197998 64852 198004 64864
rect 3384 64824 198004 64852
rect 3384 64812 3390 64824
rect 197998 64812 198004 64824
rect 198056 64812 198062 64864
rect 294598 64812 294604 64864
rect 294656 64852 294662 64864
rect 579798 64852 579804 64864
rect 294656 64824 579804 64852
rect 294656 64812 294662 64824
rect 579798 64812 579804 64824
rect 579856 64812 579862 64864
rect 255777 63563 255835 63569
rect 255777 63529 255789 63563
rect 255823 63560 255835 63563
rect 255866 63560 255872 63572
rect 255823 63532 255872 63560
rect 255823 63529 255835 63532
rect 255777 63523 255835 63529
rect 255866 63520 255872 63532
rect 255924 63520 255930 63572
rect 256421 63563 256479 63569
rect 256421 63529 256433 63563
rect 256467 63560 256479 63563
rect 256602 63560 256608 63572
rect 256467 63532 256608 63560
rect 256467 63529 256479 63532
rect 256421 63523 256479 63529
rect 256602 63520 256608 63532
rect 256660 63520 256666 63572
rect 257154 63560 257160 63572
rect 257115 63532 257160 63560
rect 257154 63520 257160 63532
rect 257212 63520 257218 63572
rect 260006 63520 260012 63572
rect 260064 63520 260070 63572
rect 273898 63560 273904 63572
rect 273859 63532 273904 63560
rect 273898 63520 273904 63532
rect 273956 63520 273962 63572
rect 274358 63560 274364 63572
rect 274284 63532 274364 63560
rect 260024 63436 260052 63520
rect 274284 63436 274312 63532
rect 274358 63520 274364 63532
rect 274416 63520 274422 63572
rect 277121 63563 277179 63569
rect 277121 63529 277133 63563
rect 277167 63560 277179 63563
rect 277210 63560 277216 63572
rect 277167 63532 277216 63560
rect 277167 63529 277179 63532
rect 277121 63523 277179 63529
rect 277210 63520 277216 63532
rect 277268 63520 277274 63572
rect 260006 63384 260012 63436
rect 260064 63384 260070 63436
rect 274266 63384 274272 63436
rect 274324 63384 274330 63436
rect 259730 62092 259736 62144
rect 259788 62132 259794 62144
rect 259822 62132 259828 62144
rect 259788 62104 259828 62132
rect 259788 62092 259794 62104
rect 259822 62092 259828 62104
rect 259880 62092 259886 62144
rect 255774 61996 255780 62008
rect 255735 61968 255780 61996
rect 255774 61956 255780 61968
rect 255832 61956 255838 62008
rect 229462 60664 229468 60716
rect 229520 60704 229526 60716
rect 229646 60704 229652 60716
rect 229520 60676 229652 60704
rect 229520 60664 229526 60676
rect 229646 60664 229652 60676
rect 229704 60664 229710 60716
rect 254854 60596 254860 60648
rect 254912 60636 254918 60648
rect 254949 60639 255007 60645
rect 254949 60636 254961 60639
rect 254912 60608 254961 60636
rect 254912 60596 254918 60608
rect 254949 60605 254961 60608
rect 254995 60605 255007 60639
rect 254949 60599 255007 60605
rect 277578 60392 277584 60444
rect 277636 60432 277642 60444
rect 277946 60432 277952 60444
rect 277636 60404 277952 60432
rect 277636 60392 277642 60404
rect 277946 60392 277952 60404
rect 278004 60392 278010 60444
rect 273622 58624 273628 58676
rect 273680 58664 273686 58676
rect 273898 58664 273904 58676
rect 273680 58636 273904 58664
rect 273680 58624 273686 58636
rect 273898 58624 273904 58636
rect 273956 58624 273962 58676
rect 235166 57944 235172 57996
rect 235224 57984 235230 57996
rect 235258 57984 235264 57996
rect 235224 57956 235264 57984
rect 235224 57944 235230 57956
rect 235258 57944 235264 57956
rect 235316 57944 235322 57996
rect 235534 57984 235540 57996
rect 235495 57956 235540 57984
rect 235534 57944 235540 57956
rect 235592 57944 235598 57996
rect 237190 57984 237196 57996
rect 237151 57956 237196 57984
rect 237190 57944 237196 57956
rect 237248 57944 237254 57996
rect 229557 57919 229615 57925
rect 229557 57885 229569 57919
rect 229603 57916 229615 57919
rect 229646 57916 229652 57928
rect 229603 57888 229652 57916
rect 229603 57885 229615 57888
rect 229557 57879 229615 57885
rect 229646 57876 229652 57888
rect 229704 57876 229710 57928
rect 245197 57919 245255 57925
rect 245197 57885 245209 57919
rect 245243 57916 245255 57919
rect 245286 57916 245292 57928
rect 245243 57888 245292 57916
rect 245243 57885 245255 57888
rect 245197 57879 245255 57885
rect 245286 57876 245292 57888
rect 245344 57876 245350 57928
rect 269574 56556 269580 56568
rect 269535 56528 269580 56556
rect 269574 56516 269580 56528
rect 269632 56516 269638 56568
rect 276934 53796 276940 53848
rect 276992 53836 276998 53848
rect 277026 53836 277032 53848
rect 276992 53808 277032 53836
rect 276992 53796 276998 53808
rect 277026 53796 277032 53808
rect 277084 53796 277090 53848
rect 269577 53635 269635 53641
rect 269577 53601 269589 53635
rect 269623 53632 269635 53635
rect 269666 53632 269672 53644
rect 269623 53604 269672 53632
rect 269623 53601 269635 53604
rect 269577 53595 269635 53601
rect 269666 53592 269672 53604
rect 269724 53592 269730 53644
rect 255774 52476 255780 52488
rect 255735 52448 255780 52476
rect 255774 52436 255780 52448
rect 255832 52436 255838 52488
rect 256970 52436 256976 52488
rect 257028 52476 257034 52488
rect 257246 52476 257252 52488
rect 257028 52448 257252 52476
rect 257028 52436 257034 52448
rect 257246 52436 257252 52448
rect 257304 52436 257310 52488
rect 237190 51116 237196 51128
rect 237116 51088 237196 51116
rect 237116 51060 237144 51088
rect 237190 51076 237196 51088
rect 237248 51076 237254 51128
rect 254949 51119 255007 51125
rect 254949 51085 254961 51119
rect 254995 51116 255007 51119
rect 255038 51116 255044 51128
rect 254995 51088 255044 51116
rect 254995 51085 255007 51088
rect 254949 51079 255007 51085
rect 255038 51076 255044 51088
rect 255096 51076 255102 51128
rect 259822 51076 259828 51128
rect 259880 51076 259886 51128
rect 3418 51008 3424 51060
rect 3476 51048 3482 51060
rect 200758 51048 200764 51060
rect 3476 51020 200764 51048
rect 3476 51008 3482 51020
rect 200758 51008 200764 51020
rect 200816 51008 200822 51060
rect 237098 51008 237104 51060
rect 237156 51008 237162 51060
rect 259840 51048 259868 51076
rect 259914 51048 259920 51060
rect 259840 51020 259920 51048
rect 259914 51008 259920 51020
rect 259972 51008 259978 51060
rect 235166 48356 235172 48408
rect 235224 48396 235230 48408
rect 235258 48396 235264 48408
rect 235224 48368 235264 48396
rect 235224 48356 235230 48368
rect 235258 48356 235264 48368
rect 235316 48356 235322 48408
rect 229554 48328 229560 48340
rect 229515 48300 229560 48328
rect 229554 48288 229560 48300
rect 229612 48288 229618 48340
rect 245194 48328 245200 48340
rect 245155 48300 245200 48328
rect 245194 48288 245200 48300
rect 245252 48288 245258 48340
rect 257154 48288 257160 48340
rect 257212 48328 257218 48340
rect 257246 48328 257252 48340
rect 257212 48300 257252 48328
rect 257212 48288 257218 48300
rect 257246 48288 257252 48300
rect 257304 48288 257310 48340
rect 271138 48288 271144 48340
rect 271196 48328 271202 48340
rect 271230 48328 271236 48340
rect 271196 48300 271236 48328
rect 271196 48288 271202 48300
rect 271230 48288 271236 48300
rect 271288 48288 271294 48340
rect 273898 48288 273904 48340
rect 273956 48328 273962 48340
rect 273990 48328 273996 48340
rect 273956 48300 273996 48328
rect 273956 48288 273962 48300
rect 273990 48288 273996 48300
rect 274048 48288 274054 48340
rect 277118 48288 277124 48340
rect 277176 48328 277182 48340
rect 277210 48328 277216 48340
rect 277176 48300 277216 48328
rect 277176 48288 277182 48300
rect 277210 48288 277216 48300
rect 277268 48288 277274 48340
rect 235166 46900 235172 46912
rect 235127 46872 235172 46900
rect 235166 46860 235172 46872
rect 235224 46860 235230 46912
rect 260558 45500 260564 45552
rect 260616 45500 260622 45552
rect 262582 45500 262588 45552
rect 262640 45540 262646 45552
rect 262674 45540 262680 45552
rect 262640 45512 262680 45540
rect 262640 45500 262646 45512
rect 262674 45500 262680 45512
rect 262732 45500 262738 45552
rect 264238 45540 264244 45552
rect 264199 45512 264244 45540
rect 264238 45500 264244 45512
rect 264296 45500 264302 45552
rect 260576 45416 260604 45500
rect 260558 45364 260564 45416
rect 260616 45364 260622 45416
rect 276845 44999 276903 45005
rect 276845 44965 276857 44999
rect 276891 44996 276903 44999
rect 276934 44996 276940 45008
rect 276891 44968 276940 44996
rect 276891 44965 276903 44968
rect 276845 44959 276903 44965
rect 276934 44956 276940 44968
rect 276992 44956 276998 45008
rect 255774 44208 255780 44260
rect 255832 44248 255838 44260
rect 255869 44251 255927 44257
rect 255869 44248 255881 44251
rect 255832 44220 255881 44248
rect 255832 44208 255838 44220
rect 255869 44217 255881 44220
rect 255915 44217 255927 44251
rect 255869 44211 255927 44217
rect 256602 44112 256608 44124
rect 256563 44084 256608 44112
rect 256602 44072 256608 44084
rect 256660 44072 256666 44124
rect 254762 42780 254768 42832
rect 254820 42820 254826 42832
rect 255038 42820 255044 42832
rect 254820 42792 255044 42820
rect 254820 42780 254826 42792
rect 255038 42780 255044 42792
rect 255096 42780 255102 42832
rect 255866 42820 255872 42832
rect 255827 42792 255872 42820
rect 255866 42780 255872 42792
rect 255924 42780 255930 42832
rect 229462 41352 229468 41404
rect 229520 41392 229526 41404
rect 229646 41392 229652 41404
rect 229520 41364 229652 41392
rect 229520 41352 229526 41364
rect 229646 41352 229652 41364
rect 229704 41352 229710 41404
rect 237006 41352 237012 41404
rect 237064 41392 237070 41404
rect 237190 41392 237196 41404
rect 237064 41364 237196 41392
rect 237064 41352 237070 41364
rect 237190 41352 237196 41364
rect 237248 41352 237254 41404
rect 277762 41352 277768 41404
rect 277820 41352 277826 41404
rect 304258 41352 304264 41404
rect 304316 41392 304322 41404
rect 580166 41392 580172 41404
rect 304316 41364 580172 41392
rect 304316 41352 304322 41364
rect 580166 41352 580172 41364
rect 580224 41352 580230 41404
rect 277780 41324 277808 41352
rect 277946 41324 277952 41336
rect 277780 41296 277952 41324
rect 277946 41284 277952 41296
rect 278004 41284 278010 41336
rect 257154 39352 257160 39364
rect 257115 39324 257160 39352
rect 257154 39312 257160 39324
rect 257212 39312 257218 39364
rect 229557 38607 229615 38613
rect 229557 38573 229569 38607
rect 229603 38604 229615 38607
rect 229646 38604 229652 38616
rect 229603 38576 229652 38604
rect 229603 38573 229615 38576
rect 229557 38567 229615 38573
rect 229646 38564 229652 38576
rect 229704 38564 229710 38616
rect 235166 37312 235172 37324
rect 235127 37284 235172 37312
rect 235166 37272 235172 37284
rect 235224 37272 235230 37324
rect 276842 37312 276848 37324
rect 276803 37284 276848 37312
rect 276842 37272 276848 37284
rect 276900 37272 276906 37324
rect 269574 37204 269580 37256
rect 269632 37244 269638 37256
rect 269666 37244 269672 37256
rect 269632 37216 269672 37244
rect 269632 37204 269638 37216
rect 269666 37204 269672 37216
rect 269724 37204 269730 37256
rect 271598 37244 271604 37256
rect 271559 37216 271604 37244
rect 271598 37204 271604 37216
rect 271656 37204 271662 37256
rect 273622 37204 273628 37256
rect 273680 37244 273686 37256
rect 273714 37244 273720 37256
rect 273680 37216 273720 37244
rect 273680 37204 273686 37216
rect 273714 37204 273720 37216
rect 273772 37204 273778 37256
rect 264238 35952 264244 35964
rect 264199 35924 264244 35952
rect 264238 35912 264244 35924
rect 264296 35912 264302 35964
rect 3418 35844 3424 35896
rect 3476 35884 3482 35896
rect 213178 35884 213184 35896
rect 3476 35856 213184 35884
rect 3476 35844 3482 35856
rect 213178 35844 213184 35856
rect 213236 35844 213242 35896
rect 260558 34620 260564 34672
rect 260616 34620 260622 34672
rect 255774 34552 255780 34604
rect 255832 34592 255838 34604
rect 255832 34564 255912 34592
rect 255832 34552 255838 34564
rect 255884 34536 255912 34564
rect 254762 34484 254768 34536
rect 254820 34524 254826 34536
rect 254854 34524 254860 34536
rect 254820 34496 254860 34524
rect 254820 34484 254826 34496
rect 254854 34484 254860 34496
rect 254912 34484 254918 34536
rect 255866 34484 255872 34536
rect 255924 34484 255930 34536
rect 257157 34527 257215 34533
rect 257157 34493 257169 34527
rect 257203 34524 257215 34527
rect 257246 34524 257252 34536
rect 257203 34496 257252 34524
rect 257203 34493 257215 34496
rect 257157 34487 257215 34493
rect 257246 34484 257252 34496
rect 257304 34484 257310 34536
rect 260576 34524 260604 34620
rect 260650 34524 260656 34536
rect 260576 34496 260656 34524
rect 260650 34484 260656 34496
rect 260708 34484 260714 34536
rect 237190 31804 237196 31816
rect 237024 31776 237196 31804
rect 237024 31748 237052 31776
rect 237190 31764 237196 31776
rect 237248 31764 237254 31816
rect 237006 31696 237012 31748
rect 237064 31696 237070 31748
rect 398098 29248 398104 29300
rect 398156 29288 398162 29300
rect 405642 29288 405648 29300
rect 398156 29260 405648 29288
rect 398156 29248 398162 29260
rect 405642 29248 405648 29260
rect 405700 29248 405706 29300
rect 436738 29248 436744 29300
rect 436796 29288 436802 29300
rect 444282 29288 444288 29300
rect 436796 29260 444288 29288
rect 436796 29248 436802 29260
rect 444282 29248 444288 29260
rect 444340 29248 444346 29300
rect 417326 29180 417332 29232
rect 417384 29220 417390 29232
rect 424962 29220 424968 29232
rect 417384 29192 424968 29220
rect 417384 29180 417390 29192
rect 424962 29180 424968 29192
rect 425020 29180 425026 29232
rect 456702 29180 456708 29232
rect 456760 29220 456766 29232
rect 463602 29220 463608 29232
rect 456760 29192 463608 29220
rect 456760 29180 456766 29192
rect 463602 29180 463608 29192
rect 463660 29180 463666 29232
rect 475286 29180 475292 29232
rect 475344 29220 475350 29232
rect 482922 29220 482928 29232
rect 475344 29192 482928 29220
rect 475344 29180 475350 29192
rect 482922 29180 482928 29192
rect 482980 29180 482986 29232
rect 495158 29180 495164 29232
rect 495216 29220 495222 29232
rect 502242 29220 502248 29232
rect 495216 29192 502248 29220
rect 495216 29180 495222 29192
rect 502242 29180 502248 29192
rect 502300 29180 502306 29232
rect 513558 29180 513564 29232
rect 513616 29220 513622 29232
rect 521562 29220 521568 29232
rect 513616 29192 521568 29220
rect 513616 29180 513622 29192
rect 521562 29180 521568 29192
rect 521620 29180 521626 29232
rect 533798 29180 533804 29232
rect 533856 29220 533862 29232
rect 540882 29220 540888 29232
rect 533856 29192 540888 29220
rect 533856 29180 533862 29192
rect 540882 29180 540888 29192
rect 540940 29180 540946 29232
rect 552474 29180 552480 29232
rect 552532 29220 552538 29232
rect 560202 29220 560208 29232
rect 552532 29192 560208 29220
rect 552532 29180 552538 29192
rect 560202 29180 560208 29192
rect 560260 29180 560266 29232
rect 280246 29044 280252 29096
rect 280304 29084 280310 29096
rect 289722 29084 289728 29096
rect 280304 29056 289728 29084
rect 280304 29044 280310 29056
rect 289722 29044 289728 29056
rect 289780 29044 289786 29096
rect 229554 29016 229560 29028
rect 229515 28988 229560 29016
rect 229554 28976 229560 28988
rect 229612 28976 229618 29028
rect 260650 29016 260656 29028
rect 260576 28988 260656 29016
rect 260576 28960 260604 28988
rect 260650 28976 260656 28988
rect 260708 28976 260714 29028
rect 235534 28948 235540 28960
rect 235495 28920 235540 28948
rect 235534 28908 235540 28920
rect 235592 28908 235598 28960
rect 260558 28908 260564 28960
rect 260616 28908 260622 28960
rect 287606 28228 287612 28280
rect 287664 28268 287670 28280
rect 567194 28268 567200 28280
rect 287664 28240 567200 28268
rect 287664 28228 287670 28240
rect 567194 28228 567200 28240
rect 567252 28228 567258 28280
rect 257246 27588 257252 27600
rect 257207 27560 257252 27588
rect 257246 27548 257252 27560
rect 257304 27548 257310 27600
rect 259822 27548 259828 27600
rect 259880 27588 259886 27600
rect 259914 27588 259920 27600
rect 259880 27560 259920 27588
rect 259880 27548 259886 27560
rect 259914 27548 259920 27560
rect 259972 27548 259978 27600
rect 274266 27588 274272 27600
rect 274227 27560 274272 27588
rect 274266 27548 274272 27560
rect 274324 27548 274330 27600
rect 264238 26228 264244 26240
rect 264199 26200 264244 26228
rect 264238 26188 264244 26200
rect 264296 26188 264302 26240
rect 268838 26228 268844 26240
rect 268799 26200 268844 26228
rect 268838 26188 268844 26200
rect 268896 26188 268902 26240
rect 229554 22108 229560 22160
rect 229612 22108 229618 22160
rect 277762 22108 277768 22160
rect 277820 22148 277826 22160
rect 277946 22148 277952 22160
rect 277820 22120 277952 22148
rect 277820 22108 277826 22120
rect 277946 22108 277952 22120
rect 278004 22108 278010 22160
rect 3142 22040 3148 22092
rect 3200 22080 3206 22092
rect 225598 22080 225604 22092
rect 3200 22052 225604 22080
rect 3200 22040 3206 22052
rect 225598 22040 225604 22052
rect 225656 22040 225662 22092
rect 229572 22024 229600 22108
rect 229554 21972 229560 22024
rect 229612 21972 229618 22024
rect 320818 21360 320824 21412
rect 320876 21400 320882 21412
rect 561674 21400 561680 21412
rect 320876 21372 561680 21400
rect 320876 21360 320882 21372
rect 561674 21360 561680 21372
rect 561732 21360 561738 21412
rect 294690 19932 294696 19984
rect 294748 19972 294754 19984
rect 543734 19972 543740 19984
rect 294748 19944 543740 19972
rect 294748 19932 294754 19944
rect 543734 19932 543740 19944
rect 543792 19932 543798 19984
rect 235166 19320 235172 19372
rect 235224 19360 235230 19372
rect 235258 19360 235264 19372
rect 235224 19332 235264 19360
rect 235224 19320 235230 19332
rect 235258 19320 235264 19332
rect 235316 19320 235322 19372
rect 235534 19360 235540 19372
rect 235495 19332 235540 19360
rect 235534 19320 235540 19332
rect 235592 19320 235598 19372
rect 237006 19320 237012 19372
rect 237064 19360 237070 19372
rect 237098 19360 237104 19372
rect 237064 19332 237104 19360
rect 237064 19320 237070 19332
rect 237098 19320 237104 19332
rect 237156 19320 237162 19372
rect 250441 19295 250499 19301
rect 250441 19261 250453 19295
rect 250487 19292 250499 19295
rect 250530 19292 250536 19304
rect 250487 19264 250536 19292
rect 250487 19261 250499 19264
rect 250441 19255 250499 19261
rect 250530 19252 250536 19264
rect 250588 19252 250594 19304
rect 297358 18572 297364 18624
rect 297416 18612 297422 18624
rect 525794 18612 525800 18624
rect 297416 18584 525800 18612
rect 297416 18572 297422 18584
rect 525794 18572 525800 18584
rect 525852 18572 525858 18624
rect 269666 18068 269672 18080
rect 269592 18040 269672 18068
rect 269592 18012 269620 18040
rect 269666 18028 269672 18040
rect 269724 18028 269730 18080
rect 256602 18000 256608 18012
rect 256563 17972 256608 18000
rect 256602 17960 256608 17972
rect 256660 17960 256666 18012
rect 257246 18000 257252 18012
rect 257207 17972 257252 18000
rect 257246 17960 257252 17972
rect 257304 17960 257310 18012
rect 269574 17960 269580 18012
rect 269632 17960 269638 18012
rect 271598 18000 271604 18012
rect 271559 17972 271604 18000
rect 271598 17960 271604 17972
rect 271656 17960 271662 18012
rect 274266 18000 274272 18012
rect 274227 17972 274272 18000
rect 274266 17960 274272 17972
rect 274324 17960 274330 18012
rect 229094 17892 229100 17944
rect 229152 17932 229158 17944
rect 579798 17932 579804 17944
rect 229152 17904 579804 17932
rect 229152 17892 229158 17904
rect 579798 17892 579804 17904
rect 579856 17892 579862 17944
rect 117222 17212 117228 17264
rect 117280 17252 117286 17264
rect 222838 17252 222844 17264
rect 117280 17224 222844 17252
rect 117280 17212 117286 17224
rect 222838 17212 222844 17224
rect 222896 17212 222902 17264
rect 277762 17212 277768 17264
rect 277820 17252 277826 17264
rect 278130 17252 278136 17264
rect 277820 17224 278136 17252
rect 277820 17212 277826 17224
rect 278130 17212 278136 17224
rect 278188 17212 278194 17264
rect 264238 16640 264244 16652
rect 264199 16612 264244 16640
rect 264238 16600 264244 16612
rect 264296 16600 264302 16652
rect 268838 16640 268844 16652
rect 268799 16612 268844 16640
rect 268838 16600 268844 16612
rect 268896 16600 268902 16652
rect 260650 16572 260656 16584
rect 260611 16544 260656 16572
rect 260650 16532 260656 16544
rect 260708 16532 260714 16584
rect 262585 16575 262643 16581
rect 262585 16541 262597 16575
rect 262631 16572 262643 16575
rect 262674 16572 262680 16584
rect 262631 16544 262680 16572
rect 262631 16541 262643 16544
rect 262585 16535 262643 16541
rect 262674 16532 262680 16544
rect 262732 16532 262738 16584
rect 151630 15852 151636 15904
rect 151688 15892 151694 15904
rect 245286 15892 245292 15904
rect 151688 15864 245292 15892
rect 151688 15852 151694 15864
rect 245286 15852 245292 15864
rect 245344 15852 245350 15904
rect 290458 15852 290464 15904
rect 290516 15892 290522 15904
rect 514754 15892 514760 15904
rect 290516 15864 514760 15892
rect 290516 15852 290522 15864
rect 514754 15852 514760 15864
rect 514812 15852 514818 15904
rect 164142 14424 164148 14476
rect 164200 14464 164206 14476
rect 228358 14464 228364 14476
rect 164200 14436 228364 14464
rect 164200 14424 164206 14436
rect 228358 14424 228364 14436
rect 228416 14424 228422 14476
rect 298738 14424 298744 14476
rect 298796 14464 298802 14476
rect 512086 14464 512092 14476
rect 298796 14436 512092 14464
rect 298796 14424 298802 14436
rect 512086 14424 512092 14436
rect 512144 14424 512150 14476
rect 148962 13064 148968 13116
rect 149020 13104 149026 13116
rect 225690 13104 225696 13116
rect 149020 13076 225696 13104
rect 149020 13064 149026 13076
rect 225690 13064 225696 13076
rect 225748 13064 225754 13116
rect 291838 13064 291844 13116
rect 291896 13104 291902 13116
rect 507854 13104 507860 13116
rect 291896 13076 507860 13104
rect 291896 13064 291902 13076
rect 507854 13064 507860 13076
rect 507912 13064 507918 13116
rect 166902 11704 166908 11756
rect 166960 11744 166966 11756
rect 226978 11744 226984 11756
rect 166960 11716 226984 11744
rect 166960 11704 166966 11716
rect 226978 11704 226984 11716
rect 227036 11704 227042 11756
rect 228910 11704 228916 11756
rect 228968 11744 228974 11756
rect 252002 11744 252008 11756
rect 228968 11716 252008 11744
rect 228968 11704 228974 11716
rect 252002 11704 252008 11716
rect 252060 11704 252066 11756
rect 301498 11704 301504 11756
rect 301556 11744 301562 11756
rect 503714 11744 503720 11756
rect 301556 11716 503720 11744
rect 301556 11704 301562 11716
rect 503714 11704 503720 11716
rect 503772 11704 503778 11756
rect 267458 10956 267464 11008
rect 267516 10996 267522 11008
rect 356146 10996 356152 11008
rect 267516 10968 356152 10996
rect 267516 10956 267522 10968
rect 356146 10956 356152 10968
rect 356204 10956 356210 11008
rect 267274 10888 267280 10940
rect 267332 10928 267338 10940
rect 358814 10928 358820 10940
rect 267332 10900 358820 10928
rect 267332 10888 267338 10900
rect 358814 10888 358820 10900
rect 358872 10888 358878 10940
rect 267182 10820 267188 10872
rect 267240 10860 267246 10872
rect 362954 10860 362960 10872
rect 267240 10832 362960 10860
rect 267240 10820 267246 10832
rect 362954 10820 362960 10832
rect 363012 10820 363018 10872
rect 267366 10752 267372 10804
rect 267424 10792 267430 10804
rect 365714 10792 365720 10804
rect 267424 10764 365720 10792
rect 267424 10752 267430 10764
rect 365714 10752 365720 10764
rect 365772 10752 365778 10804
rect 64782 10684 64788 10736
rect 64840 10724 64846 10736
rect 236730 10724 236736 10736
rect 64840 10696 236736 10724
rect 64840 10684 64846 10696
rect 236730 10684 236736 10696
rect 236788 10684 236794 10736
rect 268838 10684 268844 10736
rect 268896 10724 268902 10736
rect 369854 10724 369860 10736
rect 268896 10696 369860 10724
rect 268896 10684 268902 10696
rect 369854 10684 369860 10696
rect 369912 10684 369918 10736
rect 60642 10616 60648 10668
rect 60700 10656 60706 10668
rect 236822 10656 236828 10668
rect 60700 10628 236828 10656
rect 60700 10616 60706 10628
rect 236822 10616 236828 10628
rect 236880 10616 236886 10668
rect 268654 10616 268660 10668
rect 268712 10656 268718 10668
rect 374086 10656 374092 10668
rect 268712 10628 374092 10656
rect 268712 10616 268718 10628
rect 374086 10616 374092 10628
rect 374144 10616 374150 10668
rect 30282 10548 30288 10600
rect 30340 10588 30346 10600
rect 233050 10588 233056 10600
rect 30340 10560 233056 10588
rect 30340 10548 30346 10560
rect 233050 10548 233056 10560
rect 233108 10548 233114 10600
rect 268746 10548 268752 10600
rect 268804 10588 268810 10600
rect 376754 10588 376760 10600
rect 268804 10560 376760 10588
rect 268804 10548 268810 10560
rect 376754 10548 376760 10560
rect 376812 10548 376818 10600
rect 27522 10480 27528 10532
rect 27580 10520 27586 10532
rect 232222 10520 232228 10532
rect 27580 10492 232228 10520
rect 27580 10480 27586 10492
rect 232222 10480 232228 10492
rect 232280 10480 232286 10532
rect 269206 10480 269212 10532
rect 269264 10520 269270 10532
rect 380894 10520 380900 10532
rect 269264 10492 380900 10520
rect 269264 10480 269270 10492
rect 380894 10480 380900 10492
rect 380952 10480 380958 10532
rect 22002 10412 22008 10464
rect 22060 10452 22066 10464
rect 232130 10452 232136 10464
rect 22060 10424 232136 10452
rect 22060 10412 22066 10424
rect 232130 10412 232136 10424
rect 232188 10412 232194 10464
rect 235994 10412 236000 10464
rect 236052 10452 236058 10464
rect 253198 10452 253204 10464
rect 236052 10424 253204 10452
rect 236052 10412 236058 10424
rect 253198 10412 253204 10424
rect 253256 10412 253262 10464
rect 270034 10412 270040 10464
rect 270092 10452 270098 10464
rect 383654 10452 383660 10464
rect 270092 10424 383660 10452
rect 270092 10412 270098 10424
rect 383654 10412 383660 10424
rect 383712 10412 383718 10464
rect 9582 10344 9588 10396
rect 9640 10384 9646 10396
rect 230842 10384 230848 10396
rect 9640 10356 230848 10384
rect 9640 10344 9646 10356
rect 230842 10344 230848 10356
rect 230900 10344 230906 10396
rect 232498 10344 232504 10396
rect 232556 10384 232562 10396
rect 252922 10384 252928 10396
rect 232556 10356 252928 10384
rect 232556 10344 232562 10356
rect 252922 10344 252928 10356
rect 252980 10344 252986 10396
rect 269114 10344 269120 10396
rect 269172 10384 269178 10396
rect 387794 10384 387800 10396
rect 269172 10356 387800 10384
rect 269172 10344 269178 10356
rect 387794 10344 387800 10356
rect 387852 10344 387858 10396
rect 3970 10276 3976 10328
rect 4028 10316 4034 10328
rect 229554 10316 229560 10328
rect 4028 10288 229560 10316
rect 4028 10276 4034 10288
rect 229554 10276 229560 10288
rect 229612 10276 229618 10328
rect 231302 10276 231308 10328
rect 231360 10316 231366 10328
rect 251174 10316 251180 10328
rect 231360 10288 251180 10316
rect 231360 10276 231366 10288
rect 251174 10276 251180 10288
rect 251232 10276 251238 10328
rect 270218 10276 270224 10328
rect 270276 10316 270282 10328
rect 390554 10316 390560 10328
rect 270276 10288 390560 10316
rect 270276 10276 270282 10288
rect 390554 10276 390560 10288
rect 390612 10276 390618 10328
rect 265986 10208 265992 10260
rect 266044 10248 266050 10260
rect 351914 10248 351920 10260
rect 266044 10220 351920 10248
rect 266044 10208 266050 10220
rect 351914 10208 351920 10220
rect 351972 10208 351978 10260
rect 265802 10140 265808 10192
rect 265860 10180 265866 10192
rect 347774 10180 347780 10192
rect 265860 10152 347780 10180
rect 265860 10140 265866 10152
rect 347774 10140 347780 10152
rect 347832 10140 347838 10192
rect 265710 10072 265716 10124
rect 265768 10112 265774 10124
rect 345014 10112 345020 10124
rect 265768 10084 345020 10112
rect 265768 10072 265774 10084
rect 345014 10072 345020 10084
rect 345072 10072 345078 10124
rect 265066 10004 265072 10056
rect 265124 10044 265130 10056
rect 340874 10044 340880 10056
rect 265124 10016 340880 10044
rect 265124 10004 265130 10016
rect 340874 10004 340880 10016
rect 340932 10004 340938 10056
rect 250438 9704 250444 9716
rect 250399 9676 250444 9704
rect 250438 9664 250444 9676
rect 250496 9664 250502 9716
rect 256510 9704 256516 9716
rect 256471 9676 256516 9704
rect 256510 9664 256516 9676
rect 256568 9664 256574 9716
rect 257154 9664 257160 9716
rect 257212 9704 257218 9716
rect 257246 9704 257252 9716
rect 257212 9676 257252 9704
rect 257212 9664 257218 9676
rect 257246 9664 257252 9676
rect 257304 9664 257310 9716
rect 90910 9596 90916 9648
rect 90968 9636 90974 9648
rect 239214 9636 239220 9648
rect 90968 9608 239220 9636
rect 90968 9596 90974 9608
rect 239214 9596 239220 9608
rect 239272 9596 239278 9648
rect 87322 9528 87328 9580
rect 87380 9568 87386 9580
rect 239030 9568 239036 9580
rect 87380 9540 239036 9568
rect 87380 9528 87386 9540
rect 239030 9528 239036 9540
rect 239088 9528 239094 9580
rect 83826 9460 83832 9512
rect 83884 9500 83890 9512
rect 238570 9500 238576 9512
rect 83884 9472 238576 9500
rect 83884 9460 83890 9472
rect 238570 9460 238576 9472
rect 238628 9460 238634 9512
rect 80238 9392 80244 9444
rect 80296 9432 80302 9444
rect 238202 9432 238208 9444
rect 80296 9404 238208 9432
rect 80296 9392 80302 9404
rect 238202 9392 238208 9404
rect 238260 9392 238266 9444
rect 76650 9324 76656 9376
rect 76708 9364 76714 9376
rect 237742 9364 237748 9376
rect 76708 9336 237748 9364
rect 76708 9324 76714 9336
rect 237742 9324 237748 9336
rect 237800 9324 237806 9376
rect 73062 9256 73068 9308
rect 73120 9296 73126 9308
rect 237650 9296 237656 9308
rect 73120 9268 237656 9296
rect 73120 9256 73126 9268
rect 237650 9256 237656 9268
rect 237708 9256 237714 9308
rect 259914 9256 259920 9308
rect 259972 9296 259978 9308
rect 291930 9296 291936 9308
rect 259972 9268 291936 9296
rect 259972 9256 259978 9268
rect 291930 9256 291936 9268
rect 291988 9256 291994 9308
rect 69474 9188 69480 9240
rect 69532 9228 69538 9240
rect 236638 9228 236644 9240
rect 69532 9200 236644 9228
rect 69532 9188 69538 9200
rect 236638 9188 236644 9200
rect 236696 9188 236702 9240
rect 260006 9188 260012 9240
rect 260064 9228 260070 9240
rect 295518 9228 295524 9240
rect 260064 9200 295524 9228
rect 260064 9188 260070 9200
rect 295518 9188 295524 9200
rect 295576 9188 295582 9240
rect 65978 9120 65984 9172
rect 66036 9160 66042 9172
rect 236454 9160 236460 9172
rect 66036 9132 236460 9160
rect 66036 9120 66042 9132
rect 236454 9120 236460 9132
rect 236512 9120 236518 9172
rect 260653 9163 260711 9169
rect 260653 9129 260665 9163
rect 260699 9160 260711 9163
rect 299106 9160 299112 9172
rect 260699 9132 299112 9160
rect 260699 9129 260711 9132
rect 260653 9123 260711 9129
rect 299106 9120 299112 9132
rect 299164 9120 299170 9172
rect 62390 9052 62396 9104
rect 62448 9092 62454 9104
rect 236546 9092 236552 9104
rect 62448 9064 236552 9092
rect 62448 9052 62454 9064
rect 236546 9052 236552 9064
rect 236604 9052 236610 9104
rect 261202 9052 261208 9104
rect 261260 9092 261266 9104
rect 306190 9092 306196 9104
rect 261260 9064 306196 9092
rect 261260 9052 261266 9064
rect 306190 9052 306196 9064
rect 306248 9052 306254 9104
rect 58802 8984 58808 9036
rect 58860 9024 58866 9036
rect 236362 9024 236368 9036
rect 58860 8996 236368 9024
rect 58860 8984 58866 8996
rect 236362 8984 236368 8996
rect 236420 8984 236426 9036
rect 261294 8984 261300 9036
rect 261352 9024 261358 9036
rect 309778 9024 309784 9036
rect 261352 8996 309784 9024
rect 261352 8984 261358 8996
rect 309778 8984 309784 8996
rect 309836 8984 309842 9036
rect 17218 8916 17224 8968
rect 17276 8956 17282 8968
rect 231670 8956 231676 8968
rect 17276 8928 231676 8956
rect 17276 8916 17282 8928
rect 231670 8916 231676 8928
rect 231728 8916 231734 8968
rect 241974 8916 241980 8968
rect 242032 8956 242038 8968
rect 251818 8956 251824 8968
rect 242032 8928 251824 8956
rect 242032 8916 242038 8928
rect 251818 8916 251824 8928
rect 251876 8916 251882 8968
rect 261386 8916 261392 8968
rect 261444 8956 261450 8968
rect 302602 8956 302608 8968
rect 261444 8928 302608 8956
rect 261444 8916 261450 8928
rect 302602 8916 302608 8928
rect 302660 8916 302666 8968
rect 302878 8916 302884 8968
rect 302936 8956 302942 8968
rect 494146 8956 494152 8968
rect 302936 8928 494152 8956
rect 302936 8916 302942 8928
rect 494146 8916 494152 8928
rect 494204 8916 494210 8968
rect 94498 8848 94504 8900
rect 94556 8888 94562 8900
rect 239674 8888 239680 8900
rect 94556 8860 239680 8888
rect 94556 8848 94562 8860
rect 239674 8848 239680 8860
rect 239732 8848 239738 8900
rect 98086 8780 98092 8832
rect 98144 8820 98150 8832
rect 239122 8820 239128 8832
rect 98144 8792 239128 8820
rect 98144 8780 98150 8792
rect 239122 8780 239128 8792
rect 239180 8780 239186 8832
rect 101582 8712 101588 8764
rect 101640 8752 101646 8764
rect 240410 8752 240416 8764
rect 101640 8724 240416 8752
rect 101640 8712 101646 8724
rect 240410 8712 240416 8724
rect 240468 8712 240474 8764
rect 105170 8644 105176 8696
rect 105228 8684 105234 8696
rect 240318 8684 240324 8696
rect 105228 8656 240324 8684
rect 105228 8644 105234 8656
rect 240318 8644 240324 8656
rect 240376 8644 240382 8696
rect 108758 8576 108764 8628
rect 108816 8616 108822 8628
rect 241146 8616 241152 8628
rect 108816 8588 241152 8616
rect 108816 8576 108822 8588
rect 241146 8576 241152 8588
rect 241204 8576 241210 8628
rect 112346 8508 112352 8560
rect 112404 8548 112410 8560
rect 241882 8548 241888 8560
rect 112404 8520 241888 8548
rect 112404 8508 112410 8520
rect 241882 8508 241888 8520
rect 241940 8508 241946 8560
rect 115934 8440 115940 8492
rect 115992 8480 115998 8492
rect 241790 8480 241796 8492
rect 115992 8452 241796 8480
rect 115992 8440 115998 8452
rect 241790 8440 241796 8452
rect 241848 8440 241854 8492
rect 119430 8372 119436 8424
rect 119488 8412 119494 8424
rect 242250 8412 242256 8424
rect 119488 8384 242256 8412
rect 119488 8372 119494 8384
rect 242250 8372 242256 8384
rect 242308 8372 242314 8424
rect 269666 8412 269672 8424
rect 269592 8384 269672 8412
rect 269592 8356 269620 8384
rect 269666 8372 269672 8384
rect 269724 8372 269730 8424
rect 123018 8304 123024 8356
rect 123076 8344 123082 8356
rect 242618 8344 242624 8356
rect 123076 8316 242624 8344
rect 123076 8304 123082 8316
rect 242618 8304 242624 8316
rect 242676 8304 242682 8356
rect 256510 8344 256516 8356
rect 256471 8316 256516 8344
rect 256510 8304 256516 8316
rect 256568 8304 256574 8356
rect 269574 8304 269580 8356
rect 269632 8304 269638 8356
rect 3418 8236 3424 8288
rect 3476 8276 3482 8288
rect 135898 8276 135904 8288
rect 3476 8248 135904 8276
rect 3476 8236 3482 8248
rect 135898 8236 135904 8248
rect 135956 8236 135962 8288
rect 200390 8236 200396 8288
rect 200448 8276 200454 8288
rect 250530 8276 250536 8288
rect 200448 8248 250536 8276
rect 200448 8236 200454 8248
rect 250530 8236 250536 8248
rect 250588 8236 250594 8288
rect 253842 8236 253848 8288
rect 253900 8276 253906 8288
rect 255866 8276 255872 8288
rect 253900 8248 255872 8276
rect 253900 8236 253906 8248
rect 255866 8236 255872 8248
rect 255924 8236 255930 8288
rect 261478 8236 261484 8288
rect 261536 8276 261542 8288
rect 266998 8276 267004 8288
rect 261536 8248 267004 8276
rect 261536 8236 261542 8248
rect 266998 8236 267004 8248
rect 267056 8236 267062 8288
rect 272518 8236 272524 8288
rect 272576 8276 272582 8288
rect 275278 8276 275284 8288
rect 272576 8248 275284 8276
rect 272576 8236 272582 8248
rect 275278 8236 275284 8248
rect 275336 8236 275342 8288
rect 196802 8168 196808 8220
rect 196860 8208 196866 8220
rect 250162 8208 250168 8220
rect 196860 8180 250168 8208
rect 196860 8168 196866 8180
rect 250162 8168 250168 8180
rect 250220 8168 250226 8220
rect 193214 8100 193220 8152
rect 193272 8140 193278 8152
rect 249886 8140 249892 8152
rect 193272 8112 249892 8140
rect 193272 8100 193278 8112
rect 249886 8100 249892 8112
rect 249944 8100 249950 8152
rect 189626 8032 189632 8084
rect 189684 8072 189690 8084
rect 249426 8072 249432 8084
rect 189684 8044 249432 8072
rect 189684 8032 189690 8044
rect 249426 8032 249432 8044
rect 249484 8032 249490 8084
rect 279970 8032 279976 8084
rect 280028 8032 280034 8084
rect 186038 7964 186044 8016
rect 186096 8004 186102 8016
rect 248690 8004 248696 8016
rect 186096 7976 248696 8004
rect 186096 7964 186102 7976
rect 248690 7964 248696 7976
rect 248748 7964 248754 8016
rect 182542 7896 182548 7948
rect 182600 7936 182606 7948
rect 248782 7936 248788 7948
rect 182600 7908 248788 7936
rect 182600 7896 182606 7908
rect 248782 7896 248788 7908
rect 248840 7896 248846 7948
rect 279988 7880 280016 8032
rect 178954 7828 178960 7880
rect 179012 7868 179018 7880
rect 247402 7868 247408 7880
rect 179012 7840 247408 7868
rect 179012 7828 179018 7840
rect 247402 7828 247408 7840
rect 247460 7828 247466 7880
rect 279970 7828 279976 7880
rect 280028 7828 280034 7880
rect 175366 7760 175372 7812
rect 175424 7800 175430 7812
rect 247310 7800 247316 7812
rect 175424 7772 247316 7800
rect 175424 7760 175430 7772
rect 247310 7760 247316 7772
rect 247368 7760 247374 7812
rect 171778 7692 171784 7744
rect 171836 7732 171842 7744
rect 247862 7732 247868 7744
rect 171836 7704 247868 7732
rect 171836 7692 171842 7704
rect 247862 7692 247868 7704
rect 247920 7692 247926 7744
rect 168190 7624 168196 7676
rect 168248 7664 168254 7676
rect 247494 7664 247500 7676
rect 168248 7636 247500 7664
rect 168248 7624 168254 7636
rect 247494 7624 247500 7636
rect 247552 7624 247558 7676
rect 132586 7556 132592 7608
rect 132644 7596 132650 7608
rect 243354 7596 243360 7608
rect 132644 7568 243360 7596
rect 132644 7556 132650 7568
rect 243354 7556 243360 7568
rect 243412 7556 243418 7608
rect 316678 7556 316684 7608
rect 316736 7596 316742 7608
rect 490558 7596 490564 7608
rect 316736 7568 490564 7596
rect 316736 7556 316742 7568
rect 490558 7556 490564 7568
rect 490616 7556 490622 7608
rect 203886 7488 203892 7540
rect 203944 7528 203950 7540
rect 250898 7528 250904 7540
rect 203944 7500 250904 7528
rect 203944 7488 203950 7500
rect 250898 7488 250904 7500
rect 250956 7488 250962 7540
rect 262582 6984 262588 6996
rect 262543 6956 262588 6984
rect 262582 6944 262588 6956
rect 262640 6944 262646 6996
rect 262950 6876 262956 6928
rect 263008 6916 263014 6928
rect 268102 6916 268108 6928
rect 263008 6888 268108 6916
rect 263008 6876 263014 6888
rect 268102 6876 268108 6888
rect 268160 6876 268166 6928
rect 279878 6876 279884 6928
rect 279936 6916 279942 6928
rect 280062 6916 280068 6928
rect 279936 6888 280068 6916
rect 279936 6876 279942 6888
rect 280062 6876 280068 6888
rect 280120 6876 280126 6928
rect 280798 6876 280804 6928
rect 280856 6916 280862 6928
rect 289538 6916 289544 6928
rect 280856 6888 289544 6916
rect 280856 6876 280862 6888
rect 289538 6876 289544 6888
rect 289596 6876 289602 6928
rect 199194 6808 199200 6860
rect 199252 6848 199258 6860
rect 250346 6848 250352 6860
rect 199252 6820 250352 6848
rect 199252 6808 199258 6820
rect 250346 6808 250352 6820
rect 250404 6808 250410 6860
rect 264238 6848 264244 6860
rect 264199 6820 264244 6848
rect 264238 6808 264244 6820
rect 264296 6808 264302 6860
rect 266814 6808 266820 6860
rect 266872 6848 266878 6860
rect 354950 6848 354956 6860
rect 266872 6820 354956 6848
rect 266872 6808 266878 6820
rect 354950 6808 354956 6820
rect 355008 6808 355014 6860
rect 195606 6740 195612 6792
rect 195664 6780 195670 6792
rect 250070 6780 250076 6792
rect 195664 6752 250076 6780
rect 195664 6740 195670 6752
rect 250070 6740 250076 6752
rect 250128 6740 250134 6792
rect 266722 6740 266728 6792
rect 266780 6780 266786 6792
rect 358538 6780 358544 6792
rect 266780 6752 358544 6780
rect 266780 6740 266786 6752
rect 358538 6740 358544 6752
rect 358596 6740 358602 6792
rect 192018 6672 192024 6724
rect 192076 6712 192082 6724
rect 249702 6712 249708 6724
rect 192076 6684 249708 6712
rect 192076 6672 192082 6684
rect 249702 6672 249708 6684
rect 249760 6672 249766 6724
rect 266538 6672 266544 6724
rect 266596 6712 266602 6724
rect 362126 6712 362132 6724
rect 266596 6684 362132 6712
rect 266596 6672 266602 6684
rect 362126 6672 362132 6684
rect 362184 6672 362190 6724
rect 188430 6604 188436 6656
rect 188488 6644 188494 6656
rect 249334 6644 249340 6656
rect 188488 6616 249340 6644
rect 188488 6604 188494 6616
rect 249334 6604 249340 6616
rect 249392 6604 249398 6656
rect 266446 6604 266452 6656
rect 266504 6644 266510 6656
rect 365806 6644 365812 6656
rect 266504 6616 365812 6644
rect 266504 6604 266510 6616
rect 365806 6604 365812 6616
rect 365864 6604 365870 6656
rect 184842 6536 184848 6588
rect 184900 6576 184906 6588
rect 248874 6576 248880 6588
rect 184900 6548 248880 6576
rect 184900 6536 184906 6548
rect 248874 6536 248880 6548
rect 248932 6536 248938 6588
rect 268286 6536 268292 6588
rect 268344 6576 268350 6588
rect 369210 6576 369216 6588
rect 268344 6548 369216 6576
rect 268344 6536 268350 6548
rect 369210 6536 369216 6548
rect 369268 6536 369274 6588
rect 181346 6468 181352 6520
rect 181404 6508 181410 6520
rect 248598 6508 248604 6520
rect 181404 6480 248604 6508
rect 181404 6468 181410 6480
rect 248598 6468 248604 6480
rect 248656 6468 248662 6520
rect 267918 6468 267924 6520
rect 267976 6508 267982 6520
rect 372798 6508 372804 6520
rect 267976 6480 372804 6508
rect 267976 6468 267982 6480
rect 372798 6468 372804 6480
rect 372856 6468 372862 6520
rect 177758 6400 177764 6452
rect 177816 6440 177822 6452
rect 248138 6440 248144 6452
rect 177816 6412 248144 6440
rect 177816 6400 177822 6412
rect 248138 6400 248144 6412
rect 248196 6400 248202 6452
rect 268010 6400 268016 6452
rect 268068 6440 268074 6452
rect 376386 6440 376392 6452
rect 268068 6412 376392 6440
rect 268068 6400 268074 6412
rect 376386 6400 376392 6412
rect 376444 6400 376450 6452
rect 174170 6332 174176 6384
rect 174228 6372 174234 6384
rect 247770 6372 247776 6384
rect 174228 6344 247776 6372
rect 174228 6332 174234 6344
rect 247770 6332 247776 6344
rect 247828 6332 247834 6384
rect 267826 6332 267832 6384
rect 267884 6372 267890 6384
rect 379974 6372 379980 6384
rect 267884 6344 379980 6372
rect 267884 6332 267890 6344
rect 379974 6332 379980 6344
rect 380032 6332 380038 6384
rect 134886 6264 134892 6316
rect 134944 6304 134950 6316
rect 243170 6304 243176 6316
rect 134944 6276 243176 6304
rect 134944 6264 134950 6276
rect 243170 6264 243176 6276
rect 243228 6264 243234 6316
rect 270126 6264 270132 6316
rect 270184 6304 270190 6316
rect 383562 6304 383568 6316
rect 270184 6276 383568 6304
rect 270184 6264 270190 6276
rect 383562 6264 383568 6276
rect 383620 6264 383626 6316
rect 131390 6196 131396 6248
rect 131448 6236 131454 6248
rect 243262 6236 243268 6248
rect 131448 6208 243268 6236
rect 131448 6196 131454 6208
rect 243262 6196 243268 6208
rect 243320 6196 243326 6248
rect 269390 6196 269396 6248
rect 269448 6236 269454 6248
rect 387058 6236 387064 6248
rect 269448 6208 387064 6236
rect 269448 6196 269454 6208
rect 387058 6196 387064 6208
rect 387116 6196 387122 6248
rect 12434 6128 12440 6180
rect 12492 6168 12498 6180
rect 230658 6168 230664 6180
rect 12492 6140 230664 6168
rect 12492 6128 12498 6140
rect 230658 6128 230664 6140
rect 230716 6128 230722 6180
rect 234798 6128 234804 6180
rect 234856 6168 234862 6180
rect 254486 6168 254492 6180
rect 234856 6140 254492 6168
rect 234856 6128 234862 6140
rect 254486 6128 254492 6140
rect 254544 6128 254550 6180
rect 269482 6128 269488 6180
rect 269540 6168 269546 6180
rect 390646 6168 390652 6180
rect 269540 6140 390652 6168
rect 269540 6128 269546 6140
rect 390646 6128 390652 6140
rect 390704 6128 390710 6180
rect 202690 6060 202696 6112
rect 202748 6100 202754 6112
rect 250806 6100 250812 6112
rect 202748 6072 250812 6100
rect 202748 6060 202754 6072
rect 250806 6060 250812 6072
rect 250864 6060 250870 6112
rect 265434 6060 265440 6112
rect 265492 6100 265498 6112
rect 351362 6100 351368 6112
rect 265492 6072 351368 6100
rect 265492 6060 265498 6072
rect 351362 6060 351368 6072
rect 351420 6060 351426 6112
rect 238386 5992 238392 6044
rect 238444 6032 238450 6044
rect 254394 6032 254400 6044
rect 238444 6004 254400 6032
rect 238444 5992 238450 6004
rect 254394 5992 254400 6004
rect 254452 5992 254458 6044
rect 266078 5992 266084 6044
rect 266136 6032 266142 6044
rect 347866 6032 347872 6044
rect 266136 6004 347872 6032
rect 266136 5992 266142 6004
rect 347866 5992 347872 6004
rect 347924 5992 347930 6044
rect 266170 5924 266176 5976
rect 266228 5964 266234 5976
rect 344278 5964 344284 5976
rect 266228 5936 344284 5964
rect 266228 5924 266234 5936
rect 344278 5924 344284 5936
rect 344336 5924 344342 5976
rect 264974 5856 264980 5908
rect 265032 5896 265038 5908
rect 340690 5896 340696 5908
rect 265032 5868 340696 5896
rect 265032 5856 265038 5868
rect 340690 5856 340696 5868
rect 340748 5856 340754 5908
rect 264146 5788 264152 5840
rect 264204 5828 264210 5840
rect 337102 5828 337108 5840
rect 264204 5800 337108 5828
rect 264204 5788 264210 5800
rect 337102 5788 337108 5800
rect 337160 5788 337166 5840
rect 264054 5720 264060 5772
rect 264112 5760 264118 5772
rect 333606 5760 333612 5772
rect 264112 5732 333612 5760
rect 264112 5720 264118 5732
rect 333606 5720 333612 5732
rect 333664 5720 333670 5772
rect 264241 5695 264299 5701
rect 264241 5661 264253 5695
rect 264287 5692 264299 5695
rect 330018 5692 330024 5704
rect 264287 5664 330024 5692
rect 264287 5661 264299 5664
rect 264241 5655 264299 5661
rect 330018 5652 330024 5664
rect 330076 5652 330082 5704
rect 262674 5584 262680 5636
rect 262732 5624 262738 5636
rect 326430 5624 326436 5636
rect 262732 5596 326436 5624
rect 262732 5584 262738 5596
rect 326430 5584 326436 5596
rect 326488 5584 326494 5636
rect 262766 5516 262772 5568
rect 262824 5556 262830 5568
rect 322842 5556 322848 5568
rect 262824 5528 322848 5556
rect 262824 5516 262830 5528
rect 322842 5516 322848 5528
rect 322900 5516 322906 5568
rect 197998 5448 198004 5500
rect 198056 5488 198062 5500
rect 198056 5460 244412 5488
rect 198056 5448 198062 5460
rect 194410 5380 194416 5432
rect 194468 5420 194474 5432
rect 244277 5423 244335 5429
rect 244277 5420 244289 5423
rect 194468 5392 244289 5420
rect 194468 5380 194474 5392
rect 244277 5389 244289 5392
rect 244323 5389 244335 5423
rect 244384 5420 244412 5460
rect 257798 5448 257804 5500
rect 257856 5488 257862 5500
rect 270586 5488 270592 5500
rect 257856 5460 270592 5488
rect 257856 5448 257862 5460
rect 270586 5448 270592 5460
rect 270644 5448 270650 5500
rect 249794 5420 249800 5432
rect 244384 5392 249800 5420
rect 244277 5383 244335 5389
rect 249794 5380 249800 5392
rect 249852 5380 249858 5432
rect 258626 5380 258632 5432
rect 258684 5420 258690 5432
rect 274082 5420 274088 5432
rect 258684 5392 274088 5420
rect 258684 5380 258690 5392
rect 274082 5380 274088 5392
rect 274140 5380 274146 5432
rect 190822 5312 190828 5364
rect 190880 5352 190886 5364
rect 249518 5352 249524 5364
rect 190880 5324 249524 5352
rect 190880 5312 190886 5324
rect 249518 5312 249524 5324
rect 249576 5312 249582 5364
rect 257982 5312 257988 5364
rect 258040 5352 258046 5364
rect 272886 5352 272892 5364
rect 258040 5324 272892 5352
rect 258040 5312 258046 5324
rect 272886 5312 272892 5324
rect 272944 5312 272950 5364
rect 137278 5244 137284 5296
rect 137336 5284 137342 5296
rect 137336 5256 143948 5284
rect 137336 5244 137342 5256
rect 140866 5176 140872 5228
rect 140924 5216 140930 5228
rect 142062 5216 142068 5228
rect 140924 5188 142068 5216
rect 140924 5176 140930 5188
rect 142062 5176 142068 5188
rect 142120 5176 142126 5228
rect 143920 5216 143948 5256
rect 187234 5244 187240 5296
rect 187292 5284 187298 5296
rect 249610 5284 249616 5296
rect 187292 5256 249616 5284
rect 187292 5244 187298 5256
rect 249610 5244 249616 5256
rect 249668 5244 249674 5296
rect 258902 5244 258908 5296
rect 258960 5284 258966 5296
rect 276474 5284 276480 5296
rect 258960 5256 276480 5284
rect 258960 5244 258966 5256
rect 276474 5244 276480 5256
rect 276532 5244 276538 5296
rect 243998 5216 244004 5228
rect 143920 5188 244004 5216
rect 243998 5176 244004 5188
rect 244056 5176 244062 5228
rect 244277 5219 244335 5225
rect 244277 5185 244289 5219
rect 244323 5216 244335 5219
rect 249978 5216 249984 5228
rect 244323 5188 249984 5216
rect 244323 5185 244335 5188
rect 244277 5179 244335 5185
rect 249978 5176 249984 5188
rect 250036 5176 250042 5228
rect 258442 5176 258448 5228
rect 258500 5216 258506 5228
rect 277670 5216 277676 5228
rect 258500 5188 277676 5216
rect 258500 5176 258506 5188
rect 277670 5176 277676 5188
rect 277728 5176 277734 5228
rect 133782 5108 133788 5160
rect 133840 5148 133846 5160
rect 243722 5148 243728 5160
rect 133840 5120 243728 5148
rect 133840 5108 133846 5120
rect 243722 5108 243728 5120
rect 243780 5108 243786 5160
rect 244366 5108 244372 5160
rect 244424 5148 244430 5160
rect 247678 5148 247684 5160
rect 244424 5120 247684 5148
rect 244424 5108 244430 5120
rect 247678 5108 247684 5120
rect 247736 5108 247742 5160
rect 259086 5108 259092 5160
rect 259144 5148 259150 5160
rect 280062 5148 280068 5160
rect 259144 5120 280068 5148
rect 259144 5108 259150 5120
rect 280062 5108 280068 5120
rect 280120 5108 280126 5160
rect 130194 5040 130200 5092
rect 130252 5080 130258 5092
rect 243446 5080 243452 5092
rect 130252 5052 243452 5080
rect 130252 5040 130258 5052
rect 243446 5040 243452 5052
rect 243504 5040 243510 5092
rect 259270 5040 259276 5092
rect 259328 5080 259334 5092
rect 281258 5080 281264 5092
rect 259328 5052 281264 5080
rect 259328 5040 259334 5052
rect 281258 5040 281264 5052
rect 281316 5040 281322 5092
rect 7650 4972 7656 5024
rect 7708 5012 7714 5024
rect 224129 5015 224187 5021
rect 224129 5012 224141 5015
rect 7708 4984 224141 5012
rect 7708 4972 7714 4984
rect 224129 4981 224141 4984
rect 224175 4981 224187 5015
rect 224129 4975 224187 4981
rect 224221 5015 224279 5021
rect 224221 4981 224233 5015
rect 224267 5012 224279 5015
rect 229278 5012 229284 5024
rect 224267 4984 229284 5012
rect 224267 4981 224279 4984
rect 224221 4975 224279 4981
rect 229278 4972 229284 4984
rect 229336 4972 229342 5024
rect 259178 4972 259184 5024
rect 259236 5012 259242 5024
rect 284754 5012 284760 5024
rect 259236 4984 284760 5012
rect 259236 4972 259242 4984
rect 284754 4972 284760 4984
rect 284812 4972 284818 5024
rect 2866 4904 2872 4956
rect 2924 4944 2930 4956
rect 229186 4944 229192 4956
rect 2924 4916 229192 4944
rect 2924 4904 2930 4916
rect 229186 4904 229192 4916
rect 229244 4904 229250 4956
rect 240778 4904 240784 4956
rect 240836 4944 240842 4956
rect 254302 4944 254308 4956
rect 240836 4916 254308 4944
rect 240836 4904 240842 4916
rect 254302 4904 254308 4916
rect 254360 4904 254366 4956
rect 260282 4904 260288 4956
rect 260340 4944 260346 4956
rect 278041 4947 278099 4953
rect 278041 4944 278053 4947
rect 260340 4916 278053 4944
rect 260340 4904 260346 4916
rect 278041 4913 278053 4916
rect 278087 4913 278099 4947
rect 278041 4907 278099 4913
rect 283558 4904 283564 4956
rect 283616 4944 283622 4956
rect 283616 4916 291884 4944
rect 283616 4904 283622 4916
rect 1670 4836 1676 4888
rect 1728 4876 1734 4888
rect 1728 4848 224356 4876
rect 1728 4836 1734 4848
rect 566 4768 572 4820
rect 624 4808 630 4820
rect 224221 4811 224279 4817
rect 224221 4808 224233 4811
rect 624 4780 224233 4808
rect 624 4768 630 4780
rect 224221 4777 224233 4780
rect 224267 4777 224279 4811
rect 224328 4808 224356 4848
rect 237282 4836 237288 4888
rect 237340 4876 237346 4888
rect 254118 4876 254124 4888
rect 237340 4848 254124 4876
rect 237340 4836 237346 4848
rect 254118 4836 254124 4848
rect 254176 4836 254182 4888
rect 258350 4836 258356 4888
rect 258408 4876 258414 4888
rect 283650 4876 283656 4888
rect 258408 4848 283656 4876
rect 258408 4836 258414 4848
rect 283650 4836 283656 4848
rect 283708 4836 283714 4888
rect 291856 4876 291884 4916
rect 332410 4876 332416 4888
rect 291856 4848 332416 4876
rect 332410 4836 332416 4848
rect 332468 4836 332474 4888
rect 229370 4808 229376 4820
rect 224328 4780 229376 4808
rect 224221 4771 224279 4777
rect 229370 4768 229376 4780
rect 229428 4768 229434 4820
rect 233694 4768 233700 4820
rect 233752 4808 233758 4820
rect 254210 4808 254216 4820
rect 233752 4780 254216 4808
rect 233752 4768 233758 4780
rect 254210 4768 254216 4780
rect 254268 4768 254274 4820
rect 260190 4768 260196 4820
rect 260248 4808 260254 4820
rect 290734 4808 290740 4820
rect 260248 4780 290740 4808
rect 260248 4768 260254 4780
rect 290734 4768 290740 4780
rect 290792 4768 290798 4820
rect 315298 4768 315304 4820
rect 315356 4808 315362 4820
rect 486970 4808 486976 4820
rect 315356 4780 486976 4808
rect 315356 4768 315362 4780
rect 486970 4768 486976 4780
rect 487028 4768 487034 4820
rect 489178 4768 489184 4820
rect 489236 4808 489242 4820
rect 497734 4808 497740 4820
rect 489236 4780 497740 4808
rect 489236 4768 489242 4780
rect 497734 4768 497740 4780
rect 497792 4768 497798 4820
rect 201494 4700 201500 4752
rect 201552 4740 201558 4752
rect 251082 4740 251088 4752
rect 201552 4712 251088 4740
rect 201552 4700 201558 4712
rect 251082 4700 251088 4712
rect 251140 4700 251146 4752
rect 257614 4700 257620 4752
rect 257672 4740 257678 4752
rect 269298 4740 269304 4752
rect 257672 4712 269304 4740
rect 257672 4700 257678 4712
rect 269298 4700 269304 4712
rect 269356 4700 269362 4752
rect 278041 4743 278099 4749
rect 278041 4709 278053 4743
rect 278087 4740 278099 4743
rect 287146 4740 287152 4752
rect 278087 4712 287152 4740
rect 278087 4709 278099 4712
rect 278041 4703 278099 4709
rect 287146 4700 287152 4712
rect 287204 4700 287210 4752
rect 205082 4632 205088 4684
rect 205140 4672 205146 4684
rect 250990 4672 250996 4684
rect 205140 4644 250996 4672
rect 205140 4632 205146 4644
rect 250990 4632 250996 4644
rect 251048 4632 251054 4684
rect 224129 4607 224187 4613
rect 224129 4573 224141 4607
rect 224175 4604 224187 4607
rect 230750 4604 230756 4616
rect 224175 4576 230756 4604
rect 224175 4573 224187 4576
rect 224129 4567 224187 4573
rect 230750 4564 230756 4576
rect 230808 4564 230814 4616
rect 124214 4156 124220 4208
rect 124272 4196 124278 4208
rect 125410 4196 125416 4208
rect 124272 4168 125416 4196
rect 124272 4156 124278 4168
rect 125410 4156 125416 4168
rect 125468 4156 125474 4208
rect 150434 4156 150440 4208
rect 150492 4196 150498 4208
rect 151630 4196 151636 4208
rect 150492 4168 151636 4196
rect 150492 4156 150498 4168
rect 151630 4156 151636 4168
rect 151688 4156 151694 4208
rect 158714 4156 158720 4208
rect 158772 4196 158778 4208
rect 160002 4196 160008 4208
rect 158772 4168 160008 4196
rect 158772 4156 158778 4168
rect 160002 4156 160008 4168
rect 160060 4156 160066 4208
rect 167086 4156 167092 4208
rect 167144 4196 167150 4208
rect 168282 4196 168288 4208
rect 167144 4168 168288 4196
rect 167144 4156 167150 4168
rect 168282 4156 168288 4168
rect 168340 4156 168346 4208
rect 209866 4156 209872 4208
rect 209924 4196 209930 4208
rect 211062 4196 211068 4208
rect 209924 4168 211068 4196
rect 209924 4156 209930 4168
rect 211062 4156 211068 4168
rect 211120 4156 211126 4208
rect 265342 4156 265348 4208
rect 265400 4196 265406 4208
rect 265802 4196 265808 4208
rect 265400 4168 265808 4196
rect 265400 4156 265406 4168
rect 265802 4156 265808 4168
rect 265860 4156 265866 4208
rect 287054 4156 287060 4208
rect 287112 4196 287118 4208
rect 288342 4196 288348 4208
rect 287112 4168 288348 4196
rect 287112 4156 287118 4168
rect 288342 4156 288348 4168
rect 288400 4156 288406 4208
rect 296714 4156 296720 4208
rect 296772 4196 296778 4208
rect 297910 4196 297916 4208
rect 296772 4168 297916 4196
rect 296772 4156 296778 4168
rect 297910 4156 297916 4168
rect 297968 4156 297974 4208
rect 313366 4156 313372 4208
rect 313424 4196 313430 4208
rect 314562 4196 314568 4208
rect 313424 4168 314568 4196
rect 313424 4156 313430 4168
rect 314562 4156 314568 4168
rect 314620 4156 314626 4208
rect 347774 4156 347780 4208
rect 347832 4196 347838 4208
rect 349062 4196 349068 4208
rect 347832 4168 349068 4196
rect 347832 4156 347838 4168
rect 349062 4156 349068 4168
rect 349120 4156 349126 4208
rect 356054 4156 356060 4208
rect 356112 4196 356118 4208
rect 357342 4196 357348 4208
rect 356112 4168 357348 4196
rect 356112 4156 356118 4168
rect 357342 4156 357348 4168
rect 357400 4156 357406 4208
rect 365714 4156 365720 4208
rect 365772 4196 365778 4208
rect 366910 4196 366916 4208
rect 365772 4168 366916 4196
rect 365772 4156 365778 4168
rect 366910 4156 366916 4168
rect 366968 4156 366974 4208
rect 373994 4156 374000 4208
rect 374052 4196 374058 4208
rect 375190 4196 375196 4208
rect 374052 4168 375196 4196
rect 374052 4156 374058 4168
rect 375190 4156 375196 4168
rect 375248 4156 375254 4208
rect 20714 4088 20720 4140
rect 20772 4128 20778 4140
rect 28258 4128 28264 4140
rect 20772 4100 28264 4128
rect 20772 4088 20778 4100
rect 28258 4088 28264 4100
rect 28316 4088 28322 4140
rect 79042 4088 79048 4140
rect 79100 4128 79106 4140
rect 238018 4128 238024 4140
rect 79100 4100 238024 4128
rect 79100 4088 79106 4100
rect 238018 4088 238024 4100
rect 238076 4088 238082 4140
rect 239582 4088 239588 4140
rect 239640 4128 239646 4140
rect 240042 4128 240048 4140
rect 239640 4100 240048 4128
rect 239640 4088 239646 4100
rect 240042 4088 240048 4100
rect 240100 4088 240106 4140
rect 255038 4088 255044 4140
rect 255096 4128 255102 4140
rect 256142 4128 256148 4140
rect 255096 4100 256148 4128
rect 255096 4088 255102 4100
rect 256142 4088 256148 4100
rect 256200 4088 256206 4140
rect 258534 4088 258540 4140
rect 258592 4128 258598 4140
rect 259822 4128 259828 4140
rect 258592 4100 259828 4128
rect 258592 4088 258598 4100
rect 259822 4088 259828 4100
rect 259880 4088 259886 4140
rect 262858 4088 262864 4140
rect 262916 4128 262922 4140
rect 264606 4128 264612 4140
rect 262916 4100 264612 4128
rect 262916 4088 262922 4100
rect 264606 4088 264612 4100
rect 264664 4088 264670 4140
rect 273806 4088 273812 4140
rect 273864 4128 273870 4140
rect 425054 4128 425060 4140
rect 273864 4100 425060 4128
rect 273864 4088 273870 4100
rect 425054 4088 425060 4100
rect 425112 4088 425118 4140
rect 556798 4088 556804 4140
rect 556856 4128 556862 4140
rect 559558 4128 559564 4140
rect 556856 4100 559564 4128
rect 556856 4088 556862 4100
rect 559558 4088 559564 4100
rect 559616 4088 559622 4140
rect 84102 4020 84108 4072
rect 84160 4060 84166 4072
rect 238478 4060 238484 4072
rect 84160 4032 238484 4060
rect 84160 4020 84166 4032
rect 238478 4020 238484 4032
rect 238536 4020 238542 4072
rect 243170 4020 243176 4072
rect 243228 4060 243234 4072
rect 254854 4060 254860 4072
rect 243228 4032 254860 4060
rect 243228 4020 243234 4032
rect 254854 4020 254860 4032
rect 254912 4020 254918 4072
rect 257338 4020 257344 4072
rect 257396 4060 257402 4072
rect 258626 4060 258632 4072
rect 257396 4032 258632 4060
rect 257396 4020 257402 4032
rect 258626 4020 258632 4032
rect 258684 4020 258690 4072
rect 273622 4020 273628 4072
rect 273680 4060 273686 4072
rect 428734 4060 428740 4072
rect 273680 4032 428740 4060
rect 273680 4020 273686 4032
rect 428734 4020 428740 4032
rect 428792 4020 428798 4072
rect 71866 3952 71872 4004
rect 71924 3992 71930 4004
rect 236270 3992 236276 4004
rect 71924 3964 236276 3992
rect 71924 3952 71930 3964
rect 236270 3952 236276 3964
rect 236328 3952 236334 4004
rect 257706 3952 257712 4004
rect 257764 3992 257770 4004
rect 261018 3992 261024 4004
rect 257764 3964 261024 3992
rect 257764 3952 257770 3964
rect 261018 3952 261024 3964
rect 261076 3952 261082 4004
rect 273530 3952 273536 4004
rect 273588 3992 273594 4004
rect 432322 3992 432328 4004
rect 273588 3964 432328 3992
rect 273588 3952 273594 3964
rect 432322 3952 432328 3964
rect 432380 3952 432386 4004
rect 68278 3884 68284 3936
rect 68336 3924 68342 3936
rect 236178 3924 236184 3936
rect 68336 3896 236184 3924
rect 68336 3884 68342 3896
rect 236178 3884 236184 3896
rect 236236 3884 236242 3936
rect 257154 3884 257160 3936
rect 257212 3924 257218 3936
rect 262214 3924 262220 3936
rect 257212 3896 262220 3924
rect 257212 3884 257218 3896
rect 262214 3884 262220 3896
rect 262272 3884 262278 3936
rect 275738 3884 275744 3936
rect 275796 3924 275802 3936
rect 435818 3924 435824 3936
rect 275796 3896 435824 3924
rect 275796 3884 275802 3896
rect 435818 3884 435824 3896
rect 435876 3884 435882 3936
rect 64690 3816 64696 3868
rect 64748 3856 64754 3868
rect 225233 3859 225291 3865
rect 225233 3856 225245 3859
rect 64748 3828 225245 3856
rect 64748 3816 64754 3828
rect 225233 3825 225245 3828
rect 225279 3825 225291 3859
rect 225233 3819 225291 3825
rect 225322 3816 225328 3868
rect 225380 3856 225386 3868
rect 226242 3856 226248 3868
rect 225380 3828 226248 3856
rect 225380 3816 225386 3828
rect 226242 3816 226248 3828
rect 226300 3816 226306 3868
rect 226518 3816 226524 3868
rect 226576 3856 226582 3868
rect 227622 3856 227628 3868
rect 226576 3828 227628 3856
rect 226576 3816 226582 3828
rect 227622 3816 227628 3828
rect 227680 3816 227686 3868
rect 227714 3816 227720 3868
rect 227772 3856 227778 3868
rect 229002 3856 229008 3868
rect 227772 3828 229008 3856
rect 227772 3816 227778 3828
rect 229002 3816 229008 3828
rect 229060 3816 229066 3868
rect 229741 3859 229799 3865
rect 229741 3825 229753 3859
rect 229787 3856 229799 3859
rect 235534 3856 235540 3868
rect 229787 3828 235540 3856
rect 229787 3825 229799 3828
rect 229741 3819 229799 3825
rect 235534 3816 235540 3828
rect 235592 3816 235598 3868
rect 250346 3816 250352 3868
rect 250404 3856 250410 3868
rect 255958 3856 255964 3868
rect 250404 3828 255964 3856
rect 250404 3816 250410 3828
rect 255958 3816 255964 3828
rect 256016 3816 256022 3868
rect 257062 3816 257068 3868
rect 257120 3856 257126 3868
rect 263410 3856 263416 3868
rect 257120 3828 263416 3856
rect 257120 3816 257126 3828
rect 263410 3816 263416 3828
rect 263468 3816 263474 3868
rect 275094 3816 275100 3868
rect 275152 3856 275158 3868
rect 439406 3856 439412 3868
rect 275152 3828 439412 3856
rect 275152 3816 275158 3828
rect 439406 3816 439412 3828
rect 439464 3816 439470 3868
rect 61194 3748 61200 3800
rect 61252 3788 61258 3800
rect 236086 3788 236092 3800
rect 61252 3760 236092 3788
rect 61252 3748 61258 3760
rect 236086 3748 236092 3760
rect 236144 3748 236150 3800
rect 275370 3748 275376 3800
rect 275428 3788 275434 3800
rect 442994 3788 443000 3800
rect 275428 3760 443000 3788
rect 275428 3748 275434 3760
rect 442994 3748 443000 3760
rect 443052 3748 443058 3800
rect 44542 3680 44548 3732
rect 44600 3720 44606 3732
rect 46198 3720 46204 3732
rect 44600 3692 46204 3720
rect 44600 3680 44606 3692
rect 46198 3680 46204 3692
rect 46256 3680 46262 3732
rect 57606 3680 57612 3732
rect 57664 3720 57670 3732
rect 229741 3723 229799 3729
rect 229741 3720 229753 3723
rect 57664 3692 229753 3720
rect 57664 3680 57670 3692
rect 229741 3689 229753 3692
rect 229787 3689 229799 3723
rect 229741 3683 229799 3689
rect 229833 3723 229891 3729
rect 229833 3689 229845 3723
rect 229879 3720 229891 3723
rect 241330 3720 241336 3732
rect 229879 3692 241336 3720
rect 229879 3689 229891 3692
rect 229833 3683 229891 3689
rect 241330 3680 241336 3692
rect 241388 3680 241394 3732
rect 275002 3680 275008 3732
rect 275060 3720 275066 3732
rect 446582 3720 446588 3732
rect 275060 3692 446588 3720
rect 275060 3680 275066 3692
rect 446582 3680 446588 3692
rect 446640 3680 446646 3732
rect 571426 3680 571432 3732
rect 571484 3720 571490 3732
rect 572622 3720 572628 3732
rect 571484 3692 572628 3720
rect 571484 3680 571490 3692
rect 572622 3680 572628 3692
rect 572680 3680 572686 3732
rect 573358 3680 573364 3732
rect 573416 3720 573422 3732
rect 579798 3720 579804 3732
rect 573416 3692 579804 3720
rect 573416 3680 573422 3692
rect 579798 3680 579804 3692
rect 579856 3680 579862 3732
rect 46934 3612 46940 3664
rect 46992 3652 46998 3664
rect 46992 3624 53880 3652
rect 46992 3612 46998 3624
rect 34974 3544 34980 3596
rect 35032 3584 35038 3596
rect 35032 3556 37320 3584
rect 35032 3544 35038 3556
rect 8846 3476 8852 3528
rect 8904 3516 8910 3528
rect 9582 3516 9588 3528
rect 8904 3488 9588 3516
rect 8904 3476 8910 3488
rect 9582 3476 9588 3488
rect 9640 3476 9646 3528
rect 10042 3476 10048 3528
rect 10100 3516 10106 3528
rect 14458 3516 14464 3528
rect 10100 3488 14464 3516
rect 10100 3476 10106 3488
rect 14458 3476 14464 3488
rect 14516 3476 14522 3528
rect 18322 3476 18328 3528
rect 18380 3516 18386 3528
rect 19978 3516 19984 3528
rect 18380 3488 19984 3516
rect 18380 3476 18386 3488
rect 19978 3476 19984 3488
rect 20036 3476 20042 3528
rect 23106 3476 23112 3528
rect 23164 3516 23170 3528
rect 24118 3516 24124 3528
rect 23164 3488 24124 3516
rect 23164 3476 23170 3488
rect 24118 3476 24124 3488
rect 24176 3476 24182 3528
rect 26694 3476 26700 3528
rect 26752 3516 26758 3528
rect 27522 3516 27528 3528
rect 26752 3488 27528 3516
rect 26752 3476 26758 3488
rect 27522 3476 27528 3488
rect 27580 3476 27586 3528
rect 32398 3516 32404 3528
rect 28736 3488 32404 3516
rect 5258 3408 5264 3460
rect 5316 3448 5322 3460
rect 10318 3448 10324 3460
rect 5316 3420 10324 3448
rect 5316 3408 5322 3420
rect 10318 3408 10324 3420
rect 10376 3408 10382 3460
rect 19518 3408 19524 3460
rect 19576 3448 19582 3460
rect 28736 3448 28764 3488
rect 32398 3476 32404 3488
rect 32456 3476 32462 3528
rect 33870 3476 33876 3528
rect 33928 3516 33934 3528
rect 34422 3516 34428 3528
rect 33928 3488 34428 3516
rect 33928 3476 33934 3488
rect 34422 3476 34428 3488
rect 34480 3476 34486 3528
rect 37292 3516 37320 3556
rect 37366 3544 37372 3596
rect 37424 3584 37430 3596
rect 38562 3584 38568 3596
rect 37424 3556 38568 3584
rect 37424 3544 37430 3556
rect 38562 3544 38568 3556
rect 38620 3544 38626 3596
rect 43438 3584 43444 3596
rect 38672 3556 43444 3584
rect 38672 3516 38700 3556
rect 43438 3544 43444 3556
rect 43496 3544 43502 3596
rect 50522 3544 50528 3596
rect 50580 3584 50586 3596
rect 50982 3584 50988 3596
rect 50580 3556 50988 3584
rect 50580 3544 50586 3556
rect 50982 3544 50988 3556
rect 51040 3544 51046 3596
rect 51626 3544 51632 3596
rect 51684 3584 51690 3596
rect 52362 3584 52368 3596
rect 51684 3556 52368 3584
rect 51684 3544 51690 3556
rect 52362 3544 52368 3556
rect 52420 3544 52426 3596
rect 52822 3544 52828 3596
rect 52880 3584 52886 3596
rect 53742 3584 53748 3596
rect 52880 3556 53748 3584
rect 52880 3544 52886 3556
rect 53742 3544 53748 3556
rect 53800 3544 53806 3596
rect 53852 3584 53880 3624
rect 54018 3612 54024 3664
rect 54076 3652 54082 3664
rect 235166 3652 235172 3664
rect 54076 3624 235172 3652
rect 54076 3612 54082 3624
rect 235166 3612 235172 3624
rect 235224 3612 235230 3664
rect 247954 3612 247960 3664
rect 248012 3652 248018 3664
rect 254578 3652 254584 3664
rect 248012 3624 254584 3652
rect 248012 3612 248018 3624
rect 254578 3612 254584 3624
rect 254636 3612 254642 3664
rect 276566 3612 276572 3664
rect 276624 3652 276630 3664
rect 450170 3652 450176 3664
rect 276624 3624 450176 3652
rect 276624 3612 276630 3624
rect 450170 3612 450176 3624
rect 450228 3612 450234 3664
rect 502426 3612 502432 3664
rect 502484 3652 502490 3664
rect 503622 3652 503628 3664
rect 502484 3624 503628 3652
rect 502484 3612 502490 3624
rect 503622 3612 503628 3624
rect 503680 3612 503686 3664
rect 536926 3612 536932 3664
rect 536984 3652 536990 3664
rect 538122 3652 538128 3664
rect 536984 3624 538128 3652
rect 536984 3612 536990 3624
rect 538122 3612 538128 3624
rect 538180 3612 538186 3664
rect 546494 3612 546500 3664
rect 546552 3652 546558 3664
rect 547690 3652 547696 3664
rect 546552 3624 547696 3652
rect 546552 3612 546558 3624
rect 547690 3612 547696 3624
rect 547748 3612 547754 3664
rect 563146 3612 563152 3664
rect 563204 3652 563210 3664
rect 564342 3652 564348 3664
rect 563204 3624 564348 3652
rect 563204 3612 563210 3624
rect 564342 3612 564348 3624
rect 564400 3612 564406 3664
rect 571978 3612 571984 3664
rect 572036 3652 572042 3664
rect 580994 3652 581000 3664
rect 572036 3624 581000 3652
rect 572036 3612 572042 3624
rect 580994 3612 581000 3624
rect 581052 3612 581058 3664
rect 225049 3587 225107 3593
rect 225049 3584 225061 3587
rect 53852 3556 225061 3584
rect 225049 3553 225061 3556
rect 225095 3553 225107 3587
rect 226153 3587 226211 3593
rect 226153 3584 226165 3587
rect 225049 3547 225107 3553
rect 225156 3556 226165 3584
rect 37292 3488 38700 3516
rect 40954 3476 40960 3528
rect 41012 3516 41018 3528
rect 42058 3516 42064 3528
rect 41012 3488 42064 3516
rect 41012 3476 41018 3488
rect 42058 3476 42064 3488
rect 42116 3476 42122 3528
rect 42150 3476 42156 3528
rect 42208 3516 42214 3528
rect 42702 3516 42708 3528
rect 42208 3488 42708 3516
rect 42208 3476 42214 3488
rect 42702 3476 42708 3488
rect 42760 3476 42766 3528
rect 43346 3476 43352 3528
rect 43404 3516 43410 3528
rect 225156 3516 225184 3556
rect 226153 3553 226165 3556
rect 226199 3553 226211 3587
rect 226153 3547 226211 3553
rect 226245 3587 226303 3593
rect 226245 3553 226257 3587
rect 226291 3584 226303 3587
rect 229833 3587 229891 3593
rect 229833 3584 229845 3587
rect 226291 3556 229845 3584
rect 226291 3553 226303 3556
rect 226245 3547 226303 3553
rect 229833 3553 229845 3556
rect 229879 3553 229891 3587
rect 229833 3547 229891 3553
rect 234157 3587 234215 3593
rect 234157 3553 234169 3587
rect 234203 3584 234215 3587
rect 238938 3584 238944 3596
rect 234203 3556 238944 3584
rect 234203 3553 234215 3556
rect 234157 3547 234215 3553
rect 238938 3544 238944 3556
rect 238996 3544 239002 3596
rect 245562 3544 245568 3596
rect 245620 3584 245626 3596
rect 255222 3584 255228 3596
rect 245620 3556 255228 3584
rect 245620 3544 245626 3556
rect 255222 3544 255228 3556
rect 255280 3544 255286 3596
rect 276382 3544 276388 3596
rect 276440 3584 276446 3596
rect 453666 3584 453672 3596
rect 276440 3556 453672 3584
rect 276440 3544 276446 3556
rect 453666 3544 453672 3556
rect 453724 3544 453730 3596
rect 482278 3544 482284 3596
rect 482336 3584 482342 3596
rect 567749 3587 567807 3593
rect 567749 3584 567761 3587
rect 482336 3556 567761 3584
rect 482336 3544 482342 3556
rect 567749 3553 567761 3556
rect 567795 3553 567807 3587
rect 567749 3547 567807 3553
rect 567838 3544 567844 3596
rect 567896 3584 567902 3596
rect 570230 3584 570236 3596
rect 567896 3556 570236 3584
rect 567896 3544 567902 3556
rect 570230 3544 570236 3556
rect 570288 3544 570294 3596
rect 570598 3544 570604 3596
rect 570656 3584 570662 3596
rect 571426 3584 571432 3596
rect 570656 3556 571432 3584
rect 570656 3544 570662 3556
rect 571426 3544 571432 3556
rect 571484 3544 571490 3596
rect 574738 3544 574744 3596
rect 574796 3584 574802 3596
rect 576210 3584 576216 3596
rect 574796 3556 576216 3584
rect 574796 3544 574802 3556
rect 576210 3544 576216 3556
rect 576268 3544 576274 3596
rect 43404 3488 225184 3516
rect 225233 3519 225291 3525
rect 43404 3476 43410 3488
rect 225233 3485 225245 3519
rect 225279 3516 225291 3519
rect 229649 3519 229707 3525
rect 229649 3516 229661 3519
rect 225279 3488 229661 3516
rect 225279 3485 225291 3488
rect 225233 3479 225291 3485
rect 229649 3485 229661 3488
rect 229695 3485 229707 3519
rect 229649 3479 229707 3485
rect 229738 3476 229744 3528
rect 229796 3516 229802 3528
rect 234062 3516 234068 3528
rect 229796 3488 234068 3516
rect 229796 3476 229802 3488
rect 234062 3476 234068 3488
rect 234120 3476 234126 3528
rect 277118 3476 277124 3528
rect 277176 3516 277182 3528
rect 457254 3516 457260 3528
rect 277176 3488 457260 3516
rect 277176 3476 277182 3488
rect 457254 3476 457260 3488
rect 457312 3476 457318 3528
rect 467834 3476 467840 3528
rect 467892 3516 467898 3528
rect 469122 3516 469128 3528
rect 467892 3488 469128 3516
rect 467892 3476 467898 3488
rect 469122 3476 469128 3488
rect 469180 3476 469186 3528
rect 475378 3476 475384 3528
rect 475436 3516 475442 3528
rect 578602 3516 578608 3528
rect 475436 3488 578608 3516
rect 475436 3476 475442 3488
rect 578602 3476 578608 3488
rect 578660 3476 578666 3528
rect 19576 3420 28764 3448
rect 19576 3408 19582 3420
rect 29086 3408 29092 3460
rect 29144 3448 29150 3460
rect 35158 3448 35164 3460
rect 29144 3420 35164 3448
rect 29144 3408 29150 3420
rect 35158 3408 35164 3420
rect 35216 3408 35222 3460
rect 39758 3408 39764 3460
rect 39816 3448 39822 3460
rect 224954 3448 224960 3460
rect 39816 3420 224960 3448
rect 39816 3408 39822 3420
rect 224954 3408 224960 3420
rect 225012 3408 225018 3460
rect 225049 3451 225107 3457
rect 225049 3417 225061 3451
rect 225095 3448 225107 3451
rect 235074 3448 235080 3460
rect 225095 3420 235080 3448
rect 225095 3417 225107 3420
rect 225049 3411 225107 3417
rect 235074 3408 235080 3420
rect 235132 3408 235138 3460
rect 252646 3408 252652 3460
rect 252704 3448 252710 3460
rect 255498 3448 255504 3460
rect 252704 3420 255504 3448
rect 252704 3408 252710 3420
rect 255498 3408 255504 3420
rect 255556 3408 255562 3460
rect 276842 3408 276848 3460
rect 276900 3448 276906 3460
rect 460842 3448 460848 3460
rect 276900 3420 460848 3448
rect 276900 3408 276906 3420
rect 460842 3408 460848 3420
rect 460900 3408 460906 3460
rect 471238 3408 471244 3460
rect 471296 3448 471302 3460
rect 582190 3448 582196 3460
rect 471296 3420 582196 3448
rect 471296 3408 471302 3420
rect 582190 3408 582196 3420
rect 582248 3408 582254 3460
rect 55214 3340 55220 3392
rect 55272 3380 55278 3392
rect 56502 3380 56508 3392
rect 55272 3352 56508 3380
rect 55272 3340 55278 3352
rect 56502 3340 56508 3352
rect 56560 3340 56566 3392
rect 59998 3340 60004 3392
rect 60056 3380 60062 3392
rect 60642 3380 60648 3392
rect 60056 3352 60648 3380
rect 60056 3340 60062 3352
rect 60642 3340 60648 3352
rect 60700 3340 60706 3392
rect 63586 3340 63592 3392
rect 63644 3380 63650 3392
rect 64782 3380 64788 3392
rect 63644 3352 64788 3380
rect 63644 3340 63650 3352
rect 64782 3340 64788 3352
rect 64840 3340 64846 3392
rect 70670 3340 70676 3392
rect 70728 3380 70734 3392
rect 71682 3380 71688 3392
rect 70728 3352 71688 3380
rect 70728 3340 70734 3352
rect 71682 3340 71688 3352
rect 71740 3340 71746 3392
rect 77846 3340 77852 3392
rect 77904 3380 77910 3392
rect 78582 3380 78588 3392
rect 77904 3352 78588 3380
rect 77904 3340 77910 3352
rect 78582 3340 78588 3352
rect 78640 3340 78646 3392
rect 81434 3340 81440 3392
rect 81492 3380 81498 3392
rect 82722 3380 82728 3392
rect 81492 3352 82728 3380
rect 81492 3340 81498 3352
rect 82722 3340 82728 3352
rect 82780 3340 82786 3392
rect 225141 3383 225199 3389
rect 82832 3352 225092 3380
rect 27890 3204 27896 3256
rect 27948 3244 27954 3256
rect 31018 3244 31024 3256
rect 27948 3216 31024 3244
rect 27948 3204 27954 3216
rect 31018 3204 31024 3216
rect 31076 3204 31082 3256
rect 36170 3204 36176 3256
rect 36228 3244 36234 3256
rect 39298 3244 39304 3256
rect 36228 3216 39304 3244
rect 36228 3204 36234 3216
rect 39298 3204 39304 3216
rect 39356 3204 39362 3256
rect 82630 3204 82636 3256
rect 82688 3244 82694 3256
rect 82832 3244 82860 3352
rect 84930 3272 84936 3324
rect 84988 3312 84994 3324
rect 85482 3312 85488 3324
rect 84988 3284 85488 3312
rect 84988 3272 84994 3284
rect 85482 3272 85488 3284
rect 85540 3272 85546 3324
rect 225064 3321 225092 3352
rect 225141 3349 225153 3383
rect 225187 3380 225199 3383
rect 229097 3383 229155 3389
rect 229097 3380 229109 3383
rect 225187 3352 229109 3380
rect 225187 3349 225199 3352
rect 225141 3343 225199 3349
rect 229097 3349 229109 3352
rect 229143 3349 229155 3383
rect 229097 3343 229155 3349
rect 229649 3383 229707 3389
rect 229649 3349 229661 3383
rect 229695 3380 229707 3383
rect 237006 3380 237012 3392
rect 229695 3352 237012 3380
rect 229695 3349 229707 3352
rect 229649 3343 229707 3349
rect 237006 3340 237012 3352
rect 237064 3340 237070 3392
rect 246758 3340 246764 3392
rect 246816 3380 246822 3392
rect 255590 3380 255596 3392
rect 246816 3352 255596 3380
rect 246816 3340 246822 3352
rect 255590 3340 255596 3352
rect 255648 3340 255654 3392
rect 274266 3340 274272 3392
rect 274324 3380 274330 3392
rect 421558 3380 421564 3392
rect 274324 3352 421564 3380
rect 274324 3340 274330 3352
rect 421558 3340 421564 3352
rect 421616 3340 421622 3392
rect 433334 3340 433340 3392
rect 433392 3380 433398 3392
rect 434622 3380 434628 3392
rect 433392 3352 434628 3380
rect 433392 3340 433398 3352
rect 434622 3340 434628 3352
rect 434680 3340 434686 3392
rect 494054 3340 494060 3392
rect 494112 3380 494118 3392
rect 495342 3380 495348 3392
rect 494112 3352 495348 3380
rect 494112 3340 494118 3352
rect 495342 3340 495348 3352
rect 495400 3340 495406 3392
rect 511994 3340 512000 3392
rect 512052 3380 512058 3392
rect 513190 3380 513196 3392
rect 512052 3352 513196 3380
rect 512052 3340 512058 3352
rect 513190 3340 513196 3352
rect 513248 3340 513254 3392
rect 528554 3340 528560 3392
rect 528612 3380 528618 3392
rect 529842 3380 529848 3392
rect 528612 3352 529848 3380
rect 528612 3340 528618 3352
rect 529842 3340 529848 3352
rect 529900 3340 529906 3392
rect 567749 3383 567807 3389
rect 567749 3349 567761 3383
rect 567795 3380 567807 3383
rect 575014 3380 575020 3392
rect 567795 3352 575020 3380
rect 567795 3349 567807 3352
rect 567749 3343 567807 3349
rect 575014 3340 575020 3352
rect 575072 3340 575078 3392
rect 224957 3315 225015 3321
rect 224957 3312 224969 3315
rect 89640 3284 224969 3312
rect 82688 3216 82860 3244
rect 82688 3204 82694 3216
rect 86126 3204 86132 3256
rect 86184 3244 86190 3256
rect 89640 3244 89668 3284
rect 224957 3281 224969 3284
rect 225003 3281 225015 3315
rect 224957 3275 225015 3281
rect 225049 3315 225107 3321
rect 225049 3281 225061 3315
rect 225095 3281 225107 3315
rect 229741 3315 229799 3321
rect 229741 3312 229753 3315
rect 225049 3275 225107 3281
rect 225156 3284 229753 3312
rect 86184 3216 89668 3244
rect 86184 3204 86190 3216
rect 89714 3204 89720 3256
rect 89772 3244 89778 3256
rect 225156 3244 225184 3284
rect 229741 3281 229753 3284
rect 229787 3281 229799 3315
rect 229741 3275 229799 3281
rect 229830 3272 229836 3324
rect 229888 3312 229894 3324
rect 234430 3312 234436 3324
rect 229888 3284 234436 3312
rect 229888 3272 229894 3284
rect 234430 3272 234436 3284
rect 234488 3272 234494 3324
rect 272150 3272 272156 3324
rect 272208 3312 272214 3324
rect 417970 3312 417976 3324
rect 272208 3284 417976 3312
rect 272208 3272 272214 3284
rect 417970 3272 417976 3284
rect 418028 3272 418034 3324
rect 574830 3272 574836 3324
rect 574888 3312 574894 3324
rect 577406 3312 577412 3324
rect 574888 3284 577412 3312
rect 574888 3272 574894 3284
rect 577406 3272 577412 3284
rect 577464 3272 577470 3324
rect 89772 3216 225184 3244
rect 225233 3247 225291 3253
rect 89772 3204 89778 3216
rect 225233 3213 225245 3247
rect 225279 3244 225291 3247
rect 238110 3244 238116 3256
rect 225279 3216 238116 3244
rect 225279 3213 225291 3216
rect 225233 3207 225291 3213
rect 238110 3204 238116 3216
rect 238168 3204 238174 3256
rect 272334 3204 272340 3256
rect 272392 3244 272398 3256
rect 414474 3244 414480 3256
rect 272392 3216 414480 3244
rect 272392 3204 272398 3216
rect 414474 3204 414480 3216
rect 414532 3204 414538 3256
rect 75454 3136 75460 3188
rect 75512 3176 75518 3188
rect 84102 3176 84108 3188
rect 75512 3148 84108 3176
rect 75512 3136 75518 3148
rect 84102 3136 84108 3148
rect 84160 3136 84166 3188
rect 88518 3136 88524 3188
rect 88576 3176 88582 3188
rect 89622 3176 89628 3188
rect 88576 3148 89628 3176
rect 88576 3136 88582 3148
rect 89622 3136 89628 3148
rect 89680 3136 89686 3188
rect 93302 3136 93308 3188
rect 93360 3176 93366 3188
rect 239490 3176 239496 3188
rect 93360 3148 239496 3176
rect 93360 3136 93366 3148
rect 239490 3136 239496 3148
rect 239548 3136 239554 3188
rect 271966 3136 271972 3188
rect 272024 3176 272030 3188
rect 410886 3176 410892 3188
rect 272024 3148 410892 3176
rect 272024 3136 272030 3148
rect 410886 3136 410892 3148
rect 410944 3136 410950 3188
rect 95694 3068 95700 3120
rect 95752 3108 95758 3120
rect 96522 3108 96528 3120
rect 95752 3080 96528 3108
rect 95752 3068 95758 3080
rect 96522 3068 96528 3080
rect 96580 3068 96586 3120
rect 102778 3068 102784 3120
rect 102836 3108 102842 3120
rect 103422 3108 103428 3120
rect 102836 3080 103428 3108
rect 102836 3068 102842 3080
rect 103422 3068 103428 3080
rect 103480 3068 103486 3120
rect 106366 3068 106372 3120
rect 106424 3108 106430 3120
rect 107470 3108 107476 3120
rect 106424 3080 107476 3108
rect 106424 3068 106430 3080
rect 107470 3068 107476 3080
rect 107528 3068 107534 3120
rect 239674 3108 239680 3120
rect 108316 3080 239680 3108
rect 11238 3000 11244 3052
rect 11296 3040 11302 3052
rect 15838 3040 15844 3052
rect 11296 3012 15844 3040
rect 11296 3000 11302 3012
rect 15838 3000 15844 3012
rect 15896 3000 15902 3052
rect 96890 3000 96896 3052
rect 96948 3040 96954 3052
rect 108316 3040 108344 3080
rect 239674 3068 239680 3080
rect 239732 3068 239738 3120
rect 272242 3068 272248 3120
rect 272300 3108 272306 3120
rect 407298 3108 407304 3120
rect 272300 3080 407304 3108
rect 272300 3068 272306 3080
rect 407298 3068 407304 3080
rect 407356 3068 407362 3120
rect 226429 3043 226487 3049
rect 96948 3012 108344 3040
rect 108408 3012 226380 3040
rect 96948 3000 96954 3012
rect 45738 2864 45744 2916
rect 45796 2904 45802 2916
rect 50338 2904 50344 2916
rect 45796 2876 50344 2904
rect 45796 2864 45802 2876
rect 50338 2864 50344 2876
rect 50396 2864 50402 2916
rect 103974 2864 103980 2916
rect 104032 2904 104038 2916
rect 108408 2904 108436 3012
rect 113542 2932 113548 2984
rect 113600 2972 113606 2984
rect 114462 2972 114468 2984
rect 113600 2944 114468 2972
rect 113600 2932 113606 2944
rect 114462 2932 114468 2944
rect 114520 2932 114526 2984
rect 226245 2975 226303 2981
rect 226245 2972 226257 2975
rect 114572 2944 226257 2972
rect 104032 2876 108436 2904
rect 104032 2864 104038 2876
rect 111150 2864 111156 2916
rect 111208 2904 111214 2916
rect 114572 2904 114600 2944
rect 226245 2941 226257 2944
rect 226291 2941 226303 2975
rect 226352 2972 226380 3012
rect 226429 3009 226441 3043
rect 226475 3040 226487 3043
rect 229646 3040 229652 3052
rect 226475 3012 229652 3040
rect 226475 3009 226487 3012
rect 226429 3003 226487 3009
rect 229646 3000 229652 3012
rect 229704 3000 229710 3052
rect 229741 3043 229799 3049
rect 229741 3009 229753 3043
rect 229787 3040 229799 3043
rect 239950 3040 239956 3052
rect 229787 3012 239956 3040
rect 229787 3009 229799 3012
rect 229741 3003 229799 3009
rect 239950 3000 239956 3012
rect 240008 3000 240014 3052
rect 271138 3000 271144 3052
rect 271196 3040 271202 3052
rect 403710 3040 403716 3052
rect 271196 3012 403716 3040
rect 271196 3000 271202 3012
rect 403710 3000 403716 3012
rect 403768 3000 403774 3052
rect 560938 3000 560944 3052
rect 560996 3040 561002 3052
rect 566734 3040 566740 3052
rect 560996 3012 566740 3040
rect 560996 3000 561002 3012
rect 566734 3000 566740 3012
rect 566792 3000 566798 3052
rect 241054 2972 241060 2984
rect 226352 2944 241060 2972
rect 226245 2935 226303 2941
rect 241054 2932 241060 2944
rect 241112 2932 241118 2984
rect 249150 2932 249156 2984
rect 249208 2972 249214 2984
rect 255682 2972 255688 2984
rect 249208 2944 255688 2972
rect 249208 2932 249214 2944
rect 255682 2932 255688 2944
rect 255740 2932 255746 2984
rect 271046 2932 271052 2984
rect 271104 2972 271110 2984
rect 400214 2972 400220 2984
rect 271104 2944 400220 2972
rect 271104 2932 271110 2944
rect 400214 2932 400220 2944
rect 400272 2932 400278 2984
rect 111208 2876 114600 2904
rect 111208 2864 111214 2876
rect 114738 2864 114744 2916
rect 114796 2904 114802 2916
rect 115842 2904 115848 2916
rect 114796 2876 115848 2904
rect 114796 2864 114802 2876
rect 115842 2864 115848 2876
rect 115900 2864 115906 2916
rect 120626 2864 120632 2916
rect 120684 2904 120690 2916
rect 121362 2904 121368 2916
rect 120684 2876 121368 2904
rect 120684 2864 120690 2876
rect 121362 2864 121368 2876
rect 121420 2864 121426 2916
rect 242066 2904 242072 2916
rect 121472 2876 242072 2904
rect 118234 2796 118240 2848
rect 118292 2836 118298 2848
rect 121472 2836 121500 2876
rect 242066 2864 242072 2876
rect 242124 2864 242130 2916
rect 271598 2864 271604 2916
rect 271656 2904 271662 2916
rect 396626 2904 396632 2916
rect 271656 2876 396632 2904
rect 271656 2864 271662 2876
rect 396626 2864 396632 2876
rect 396684 2864 396690 2916
rect 425146 2864 425152 2916
rect 425204 2904 425210 2916
rect 426342 2904 426348 2916
rect 425204 2876 426348 2904
rect 425204 2864 425210 2876
rect 426342 2864 426348 2876
rect 426400 2864 426406 2916
rect 118292 2808 121500 2836
rect 118292 2796 118298 2808
rect 121822 2796 121828 2848
rect 121880 2836 121886 2848
rect 242158 2836 242164 2848
rect 121880 2808 242164 2836
rect 121880 2796 121886 2808
rect 242158 2796 242164 2808
rect 242216 2796 242222 2848
rect 269574 2796 269580 2848
rect 269632 2836 269638 2848
rect 269632 2808 390508 2836
rect 269632 2796 269638 2808
rect 229097 2771 229155 2777
rect 229097 2737 229109 2771
rect 229143 2768 229155 2771
rect 234157 2771 234215 2777
rect 234157 2768 234169 2771
rect 229143 2740 234169 2768
rect 229143 2737 229155 2740
rect 229097 2731 229155 2737
rect 234157 2737 234169 2740
rect 234203 2737 234215 2771
rect 390480 2768 390508 2808
rect 390554 2796 390560 2848
rect 390612 2836 390618 2848
rect 391842 2836 391848 2848
rect 390612 2808 391848 2836
rect 390612 2796 390618 2808
rect 391842 2796 391848 2808
rect 391900 2796 391906 2848
rect 393038 2836 393044 2848
rect 391952 2808 393044 2836
rect 391952 2768 391980 2808
rect 393038 2796 393044 2808
rect 393096 2796 393102 2848
rect 390480 2740 391980 2768
rect 234157 2731 234215 2737
rect 256510 1844 256516 1896
rect 256568 1884 256574 1896
rect 257430 1884 257436 1896
rect 256568 1856 257436 1884
rect 256568 1844 256574 1856
rect 257430 1844 257436 1856
rect 257488 1844 257494 1896
rect 270494 1368 270500 1420
rect 270552 1408 270558 1420
rect 271690 1408 271696 1420
rect 270552 1380 271696 1408
rect 270552 1368 270558 1380
rect 271690 1368 271696 1380
rect 271748 1368 271754 1420
rect 74258 552 74264 604
rect 74316 592 74322 604
rect 74442 592 74448 604
rect 74316 564 74448 592
rect 74316 552 74322 564
rect 74442 552 74448 564
rect 74500 552 74506 604
rect 92106 552 92112 604
rect 92164 592 92170 604
rect 92382 592 92388 604
rect 92164 564 92388 592
rect 92164 552 92170 564
rect 92382 552 92388 564
rect 92440 552 92446 604
rect 109954 552 109960 604
rect 110012 592 110018 604
rect 110322 592 110328 604
rect 110012 564 110328 592
rect 110012 552 110018 564
rect 110322 552 110328 564
rect 110380 552 110386 604
rect 183738 552 183744 604
rect 183796 592 183802 604
rect 184750 592 184756 604
rect 183796 564 184756 592
rect 183796 552 183802 564
rect 184750 552 184756 564
rect 184808 552 184814 604
rect 206278 552 206284 604
rect 206336 592 206342 604
rect 206922 592 206928 604
rect 206336 564 206928 592
rect 206336 552 206342 564
rect 206922 552 206928 564
rect 206980 552 206986 604
rect 207474 552 207480 604
rect 207532 592 207538 604
rect 208302 592 208308 604
rect 207532 564 208308 592
rect 207532 552 207538 564
rect 208302 552 208308 564
rect 208360 552 208366 604
rect 208670 552 208676 604
rect 208728 592 208734 604
rect 209682 592 209688 604
rect 208728 564 209688 592
rect 208728 552 208734 564
rect 209682 552 209688 564
rect 209740 552 209746 604
rect 230106 552 230112 604
rect 230164 592 230170 604
rect 230382 592 230388 604
rect 230164 564 230388 592
rect 230164 552 230170 564
rect 230382 552 230388 564
rect 230440 552 230446 604
rect 251450 552 251456 604
rect 251508 592 251514 604
rect 254670 592 254676 604
rect 251508 564 254676 592
rect 251508 552 251514 564
rect 254670 552 254676 564
rect 254728 552 254734 604
rect 281534 552 281540 604
rect 281592 592 281598 604
rect 282454 592 282460 604
rect 281592 564 282460 592
rect 281592 552 281598 564
rect 282454 552 282460 564
rect 282512 552 282518 604
rect 285674 552 285680 604
rect 285732 592 285738 604
rect 285950 592 285956 604
rect 285732 564 285956 592
rect 285732 552 285738 564
rect 285950 552 285956 564
rect 286008 552 286014 604
rect 299474 552 299480 604
rect 299532 592 299538 604
rect 300302 592 300308 604
rect 299532 564 300308 592
rect 299532 552 299538 564
rect 300302 552 300308 564
rect 300360 552 300366 604
rect 300854 552 300860 604
rect 300912 592 300918 604
rect 301406 592 301412 604
rect 300912 564 301412 592
rect 300912 552 300918 564
rect 301406 552 301412 564
rect 301464 552 301470 604
rect 303614 552 303620 604
rect 303672 592 303678 604
rect 303798 592 303804 604
rect 303672 564 303804 592
rect 303672 552 303678 564
rect 303798 552 303804 564
rect 303856 552 303862 604
rect 492674 552 492680 604
rect 492732 592 492738 604
rect 492950 592 492956 604
rect 492732 564 492956 592
rect 492732 552 492738 564
rect 492950 552 492956 564
rect 493008 552 493014 604
rect 495434 552 495440 604
rect 495492 592 495498 604
rect 496538 592 496544 604
rect 495492 564 496544 592
rect 495492 552 495498 564
rect 496538 552 496544 564
rect 496596 552 496602 604
rect 498194 552 498200 604
rect 498252 592 498258 604
rect 498930 592 498936 604
rect 498252 564 498936 592
rect 498252 552 498258 564
rect 498930 552 498936 564
rect 498988 552 498994 604
<< via1 >>
rect 257896 700952 257948 701004
rect 397460 700952 397512 701004
rect 259276 700884 259328 700936
rect 413652 700884 413704 700936
rect 257988 700816 258040 700868
rect 429844 700816 429896 700868
rect 72976 700748 73028 700800
rect 265072 700748 265124 700800
rect 256424 700680 256476 700732
rect 462320 700680 462372 700732
rect 256516 700612 256568 700664
rect 478512 700612 478564 700664
rect 256608 700544 256660 700596
rect 494796 700544 494848 700596
rect 8116 700476 8168 700528
rect 266544 700476 266596 700528
rect 255228 700408 255280 700460
rect 527180 700408 527232 700460
rect 40500 700340 40552 700392
rect 41328 700340 41380 700392
rect 255136 700340 255188 700392
rect 543464 700340 543516 700392
rect 253848 700272 253900 700324
rect 559656 700272 559708 700324
rect 137836 700204 137888 700256
rect 263784 700204 263836 700256
rect 259368 700136 259420 700188
rect 364984 700136 365036 700188
rect 260656 700068 260708 700120
rect 348792 700068 348844 700120
rect 259184 700000 259236 700052
rect 332508 700000 332560 700052
rect 202788 699932 202840 699984
rect 262220 699932 262272 699984
rect 262128 699864 262180 699916
rect 283840 699864 283892 699916
rect 24308 699660 24360 699712
rect 24768 699660 24820 699712
rect 89168 699660 89220 699712
rect 89628 699660 89680 699712
rect 105452 699660 105504 699712
rect 106188 699660 106240 699712
rect 170312 699660 170364 699712
rect 171048 699660 171100 699712
rect 235172 699660 235224 699712
rect 235908 699660 235960 699712
rect 260748 699660 260800 699712
rect 267648 699660 267700 699712
rect 253756 696940 253808 696992
rect 580172 696940 580224 696992
rect 154120 695512 154172 695564
rect 154212 695512 154264 695564
rect 219164 695444 219216 695496
rect 154212 688576 154264 688628
rect 154396 688576 154448 688628
rect 299664 688576 299716 688628
rect 300124 688576 300176 688628
rect 219072 685899 219124 685908
rect 219072 685865 219081 685899
rect 219081 685865 219115 685899
rect 219115 685865 219124 685899
rect 219072 685856 219124 685865
rect 253664 685856 253716 685908
rect 580172 685856 580224 685908
rect 154396 685788 154448 685840
rect 299572 684428 299624 684480
rect 154304 676243 154356 676252
rect 154304 676209 154313 676243
rect 154313 676209 154347 676243
rect 154347 676209 154356 676243
rect 154304 676200 154356 676209
rect 218980 676175 219032 676184
rect 218980 676141 218989 676175
rect 218989 676141 219023 676175
rect 219023 676141 219032 676175
rect 218980 676132 219032 676141
rect 154304 673480 154356 673532
rect 154488 673480 154540 673532
rect 252468 673480 252520 673532
rect 580172 673480 580224 673532
rect 3516 667904 3568 667956
rect 262864 667904 262916 667956
rect 219072 666544 219124 666596
rect 299940 666544 299992 666596
rect 219164 659608 219216 659660
rect 219348 659608 219400 659660
rect 219348 656820 219400 656872
rect 154304 654100 154356 654152
rect 154488 654100 154540 654152
rect 3056 652740 3108 652792
rect 267832 652740 267884 652792
rect 252376 650020 252428 650072
rect 580172 650020 580224 650072
rect 219256 647275 219308 647284
rect 219256 647241 219265 647275
rect 219265 647241 219299 647275
rect 219299 647241 219308 647275
rect 219256 647232 219308 647241
rect 299664 647232 299716 647284
rect 299756 647232 299808 647284
rect 219256 640364 219308 640416
rect 299664 640364 299716 640416
rect 299756 640364 299808 640416
rect 219072 640228 219124 640280
rect 252284 638936 252336 638988
rect 580172 638936 580224 638988
rect 219072 637508 219124 637560
rect 219164 637508 219216 637560
rect 154304 634788 154356 634840
rect 154488 634788 154540 634840
rect 299572 630640 299624 630692
rect 299756 630640 299808 630692
rect 251088 626560 251140 626612
rect 580172 626560 580224 626612
rect 219348 626535 219400 626544
rect 219348 626501 219357 626535
rect 219357 626501 219391 626535
rect 219391 626501 219400 626535
rect 219348 626492 219400 626501
rect 219348 616879 219400 616888
rect 219348 616845 219357 616879
rect 219357 616845 219391 616879
rect 219391 616845 219400 616879
rect 219348 616836 219400 616845
rect 154304 615476 154356 615528
rect 154488 615476 154540 615528
rect 219348 611396 219400 611448
rect 299572 611328 299624 611380
rect 299756 611328 299808 611380
rect 3608 609968 3660 610020
rect 264244 609968 264296 610020
rect 219072 608719 219124 608728
rect 219072 608685 219081 608719
rect 219081 608685 219115 608719
rect 219115 608685 219124 608719
rect 219072 608676 219124 608685
rect 219072 608540 219124 608592
rect 299664 608583 299716 608592
rect 299664 608549 299673 608583
rect 299673 608549 299707 608583
rect 299707 608549 299716 608583
rect 299664 608540 299716 608549
rect 249708 603100 249760 603152
rect 580172 603100 580224 603152
rect 299848 601672 299900 601724
rect 219256 601579 219308 601588
rect 219256 601545 219265 601579
rect 219265 601545 219299 601579
rect 219299 601545 219308 601579
rect 219256 601536 219308 601545
rect 219256 598884 219308 598936
rect 299848 598927 299900 598936
rect 299848 598893 299857 598927
rect 299857 598893 299891 598927
rect 299891 598893 299900 598927
rect 299848 598884 299900 598893
rect 154304 596164 154356 596216
rect 154488 596164 154540 596216
rect 3332 594804 3384 594856
rect 269304 594804 269356 594856
rect 250996 592016 251048 592068
rect 580172 592016 580224 592068
rect 219164 589339 219216 589348
rect 219164 589305 219173 589339
rect 219173 589305 219207 589339
rect 219207 589305 219216 589339
rect 219164 589296 219216 589305
rect 299940 589296 299992 589348
rect 154304 589271 154356 589280
rect 154304 589237 154313 589271
rect 154313 589237 154347 589271
rect 154347 589237 154356 589271
rect 154304 589228 154356 589237
rect 218980 582360 219032 582412
rect 219164 582360 219216 582412
rect 299940 582428 299992 582480
rect 299848 582292 299900 582344
rect 154304 579751 154356 579760
rect 154304 579717 154313 579751
rect 154313 579717 154347 579751
rect 154347 579717 154356 579751
rect 154304 579708 154356 579717
rect 249616 579640 249668 579692
rect 580172 579640 580224 579692
rect 154212 579572 154264 579624
rect 154396 579572 154448 579624
rect 218980 579572 219032 579624
rect 218888 569959 218940 569968
rect 218888 569925 218897 569959
rect 218897 569925 218931 569959
rect 218931 569925 218940 569959
rect 218888 569916 218940 569925
rect 299572 563116 299624 563168
rect 218888 563048 218940 563100
rect 154212 562912 154264 562964
rect 154396 562912 154448 562964
rect 299572 562980 299624 563032
rect 218980 562912 219032 562964
rect 248328 556180 248380 556232
rect 580172 556180 580224 556232
rect 218888 553435 218940 553444
rect 218888 553401 218897 553435
rect 218897 553401 218931 553435
rect 218931 553401 218940 553435
rect 218888 553392 218940 553401
rect 299572 553460 299624 553512
rect 299480 553324 299532 553376
rect 3332 552032 3384 552084
rect 265624 552032 265676 552084
rect 218888 550647 218940 550656
rect 218888 550613 218897 550647
rect 218897 550613 218931 550647
rect 218931 550613 218940 550647
rect 218888 550604 218940 550613
rect 249524 545096 249576 545148
rect 580172 545096 580224 545148
rect 218888 543736 218940 543788
rect 299296 543668 299348 543720
rect 299480 543668 299532 543720
rect 218980 543600 219032 543652
rect 3240 538228 3292 538280
rect 270776 538228 270828 538280
rect 248236 532720 248288 532772
rect 580172 532720 580224 532772
rect 299572 531292 299624 531344
rect 299756 531292 299808 531344
rect 154396 531267 154448 531276
rect 154396 531233 154405 531267
rect 154405 531233 154439 531267
rect 154439 531233 154448 531267
rect 154396 531224 154448 531233
rect 299756 524424 299808 524476
rect 299848 524356 299900 524408
rect 218980 524288 219032 524340
rect 219164 524288 219216 524340
rect 154488 521636 154540 521688
rect 218796 514632 218848 514684
rect 219072 514632 219124 514684
rect 299664 511980 299716 512032
rect 299940 511980 299992 512032
rect 154396 511955 154448 511964
rect 154396 511921 154405 511955
rect 154405 511921 154439 511955
rect 154439 511921 154448 511955
rect 154396 511912 154448 511921
rect 219072 510595 219124 510604
rect 219072 510561 219081 510595
rect 219081 510561 219115 510595
rect 219115 510561 219124 510595
rect 219072 510552 219124 510561
rect 246948 509260 247000 509312
rect 580172 509260 580224 509312
rect 219072 505087 219124 505096
rect 219072 505053 219081 505087
rect 219081 505053 219115 505087
rect 219115 505053 219124 505087
rect 219072 505044 219124 505053
rect 154488 502324 154540 502376
rect 299756 502324 299808 502376
rect 299940 502324 299992 502376
rect 248144 498176 248196 498228
rect 580172 498176 580224 498228
rect 3332 495456 3384 495508
rect 267004 495456 267056 495508
rect 219072 492668 219124 492720
rect 219164 492668 219216 492720
rect 154212 492600 154264 492652
rect 154396 492600 154448 492652
rect 299664 492643 299716 492652
rect 299664 492609 299673 492643
rect 299673 492609 299707 492643
rect 299707 492609 299716 492643
rect 299664 492600 299716 492609
rect 219164 485800 219216 485852
rect 246856 485800 246908 485852
rect 580172 485800 580224 485852
rect 299664 485775 299716 485784
rect 299664 485741 299673 485775
rect 299673 485741 299707 485775
rect 299707 485741 299716 485775
rect 299664 485732 299716 485741
rect 219256 485664 219308 485716
rect 2964 480224 3016 480276
rect 272524 480224 272576 480276
rect 299572 476076 299624 476128
rect 299756 476076 299808 476128
rect 299664 473331 299716 473340
rect 299664 473297 299673 473331
rect 299673 473297 299707 473331
rect 299707 473297 299716 473331
rect 299664 473288 299716 473297
rect 154304 466420 154356 466472
rect 154488 466420 154540 466472
rect 218980 466420 219032 466472
rect 299664 466395 299716 466404
rect 299664 466361 299673 466395
rect 299673 466361 299707 466395
rect 299707 466361 299716 466395
rect 299664 466352 299716 466361
rect 219348 466284 219400 466336
rect 245568 462340 245620 462392
rect 580172 462340 580224 462392
rect 299388 460844 299440 460896
rect 299756 460844 299808 460896
rect 154304 453976 154356 454028
rect 219072 453976 219124 454028
rect 245476 451256 245528 451308
rect 580172 451256 580224 451308
rect 299480 449871 299532 449880
rect 299480 449837 299489 449871
rect 299489 449837 299523 449871
rect 299523 449837 299532 449871
rect 299480 449828 299532 449837
rect 154212 444431 154264 444440
rect 154212 444397 154221 444431
rect 154221 444397 154255 444431
rect 154255 444397 154264 444431
rect 154212 444388 154264 444397
rect 218980 444431 219032 444440
rect 218980 444397 218989 444431
rect 218989 444397 219023 444431
rect 219023 444397 219032 444431
rect 218980 444388 219032 444397
rect 299572 440240 299624 440292
rect 245384 438880 245436 438932
rect 580172 438880 580224 438932
rect 3332 437452 3384 437504
rect 269764 437452 269816 437504
rect 299572 436815 299624 436824
rect 299572 436781 299581 436815
rect 299581 436781 299615 436815
rect 299615 436781 299624 436815
rect 299572 436772 299624 436781
rect 154396 434707 154448 434716
rect 154396 434673 154405 434707
rect 154405 434673 154439 434707
rect 154439 434673 154448 434707
rect 154396 434664 154448 434673
rect 218980 434664 219032 434716
rect 219072 434664 219124 434716
rect 154396 427771 154448 427780
rect 154396 427737 154405 427771
rect 154405 427737 154439 427771
rect 154439 427737 154448 427771
rect 154396 427728 154448 427737
rect 299572 427771 299624 427780
rect 299572 427737 299581 427771
rect 299581 427737 299615 427771
rect 299615 427737 299624 427771
rect 299572 427728 299624 427737
rect 3332 423648 3384 423700
rect 273904 423648 273956 423700
rect 244188 415420 244240 415472
rect 580172 415420 580224 415472
rect 154304 415395 154356 415404
rect 154304 415361 154313 415395
rect 154313 415361 154347 415395
rect 154347 415361 154356 415395
rect 154304 415352 154356 415361
rect 299756 415352 299808 415404
rect 258448 407736 258500 407788
rect 259276 407736 259328 407788
rect 154396 405696 154448 405748
rect 299664 405739 299716 405748
rect 299664 405705 299673 405739
rect 299673 405705 299707 405739
rect 299707 405705 299716 405739
rect 299664 405696 299716 405705
rect 243820 404336 243872 404388
rect 580172 404336 580224 404388
rect 171048 402908 171100 402960
rect 263324 402908 263376 402960
rect 269212 402908 269264 402960
rect 154396 402840 154448 402892
rect 264336 402840 264388 402892
rect 106188 402772 106240 402824
rect 89628 402704 89680 402756
rect 264244 402772 264296 402824
rect 270684 402772 270736 402824
rect 41328 402636 41380 402688
rect 264888 402704 264940 402756
rect 265624 402704 265676 402756
rect 272248 402704 272300 402756
rect 24768 402568 24820 402620
rect 258080 402568 258132 402620
rect 265900 402636 265952 402688
rect 260196 402568 260248 402620
rect 266452 402568 266504 402620
rect 267004 402568 267056 402620
rect 273812 402568 273864 402620
rect 3424 402500 3476 402552
rect 3516 402432 3568 402484
rect 261208 402432 261260 402484
rect 267556 402500 267608 402552
rect 262956 402432 263008 402484
rect 269120 402432 269172 402484
rect 3700 402364 3752 402416
rect 271236 402364 271288 402416
rect 3884 402296 3936 402348
rect 272800 402296 272852 402348
rect 4068 402228 4120 402280
rect 274364 402228 274416 402280
rect 219348 402160 219400 402212
rect 262772 402160 262824 402212
rect 269764 402160 269816 402212
rect 275376 402160 275428 402212
rect 240692 402092 240744 402144
rect 248604 402092 248656 402144
rect 249524 402092 249576 402144
rect 250168 402092 250220 402144
rect 250996 402092 251048 402144
rect 251180 402092 251232 402144
rect 252376 402092 252428 402144
rect 252744 402092 252796 402144
rect 253756 402092 253808 402144
rect 254400 402092 254452 402144
rect 255228 402092 255280 402144
rect 255412 402092 255464 402144
rect 256608 402092 256660 402144
rect 256976 402092 257028 402144
rect 257988 402092 258040 402144
rect 235908 402024 235960 402076
rect 261760 402092 261812 402144
rect 299664 402092 299716 402144
rect 258540 402024 258592 402076
rect 259368 402024 259420 402076
rect 259644 402024 259696 402076
rect 260656 402024 260708 402076
rect 261208 402024 261260 402076
rect 262128 402024 262180 402076
rect 268016 402024 268068 402076
rect 272524 402024 272576 402076
rect 273260 402024 273312 402076
rect 273904 402024 273956 402076
rect 274916 402024 274968 402076
rect 493324 401956 493376 402008
rect 235908 401888 235960 401940
rect 239128 401888 239180 401940
rect 244924 401888 244976 401940
rect 245568 401888 245620 401940
rect 243268 401820 243320 401872
rect 244188 401820 244240 401872
rect 244372 401820 244424 401872
rect 245384 401820 245436 401872
rect 245936 401820 245988 401872
rect 246856 401820 246908 401872
rect 247040 401888 247092 401940
rect 248144 401888 248196 401940
rect 500224 401888 500276 401940
rect 498844 401820 498896 401872
rect 3976 401752 4028 401804
rect 278596 401752 278648 401804
rect 3792 401684 3844 401736
rect 280160 401684 280212 401736
rect 3608 401616 3660 401668
rect 281724 401616 281776 401668
rect 13084 401276 13136 401328
rect 277492 401276 277544 401328
rect 226984 401208 227036 401260
rect 276480 401208 276532 401260
rect 241244 401140 241296 401192
rect 290464 401140 290516 401192
rect 225788 401072 225840 401124
rect 280712 401072 280764 401124
rect 227076 401004 227128 401056
rect 284852 401004 284904 401056
rect 234896 400936 234948 400988
rect 297456 400936 297508 400988
rect 231768 400868 231820 400920
rect 294604 400868 294656 400920
rect 238024 400800 238076 400852
rect 301596 400800 301648 400852
rect 218704 400732 218756 400784
rect 283840 400732 283892 400784
rect 211804 400664 211856 400716
rect 278044 400664 278096 400716
rect 214564 400596 214616 400648
rect 286968 400596 287020 400648
rect 207664 400528 207716 400580
rect 281172 400528 281224 400580
rect 230664 400460 230716 400512
rect 304264 400460 304316 400512
rect 235448 400392 235500 400444
rect 308404 400392 308456 400444
rect 203524 400324 203576 400376
rect 285956 400324 286008 400376
rect 237564 400256 237616 400308
rect 413284 400256 413336 400308
rect 240140 400188 240192 400240
rect 290556 400188 290608 400240
rect 10968 399916 11020 399968
rect 275652 399916 275704 399968
rect 242072 399891 242124 399900
rect 242072 399857 242081 399891
rect 242081 399857 242115 399891
rect 242115 399857 242124 399891
rect 242072 399848 242124 399857
rect 242900 399848 242952 399900
rect 290648 399848 290700 399900
rect 227168 399780 227220 399832
rect 278780 399780 278832 399832
rect 222936 399712 222988 399764
rect 281908 399712 281960 399764
rect 233608 399644 233660 399696
rect 291936 399644 291988 399696
rect 236736 399576 236788 399628
rect 298836 399576 298888 399628
rect 225604 399508 225656 399560
rect 289268 399508 289320 399560
rect 232504 399440 232556 399492
rect 239864 399440 239916 399492
rect 302976 399440 303028 399492
rect 215944 399372 215996 399424
rect 285036 399372 285088 399424
rect 209044 399304 209096 399356
rect 279332 399304 279384 399356
rect 282460 399347 282512 399356
rect 282460 399313 282469 399347
rect 282469 399313 282503 399347
rect 282503 399313 282512 399347
rect 282460 399304 282512 399313
rect 288348 399347 288400 399356
rect 288348 399313 288357 399347
rect 288357 399313 288391 399347
rect 288391 399313 288400 399347
rect 288348 399304 288400 399313
rect 288716 399347 288768 399356
rect 288716 399313 288725 399347
rect 288725 399313 288759 399347
rect 288759 399313 288768 399347
rect 288716 399304 288768 399313
rect 234160 399279 234212 399288
rect 234160 399245 234169 399279
rect 234169 399245 234203 399279
rect 234203 399245 234212 399279
rect 234160 399236 234212 399245
rect 234528 399279 234580 399288
rect 234528 399245 234537 399279
rect 234537 399245 234571 399279
rect 234571 399245 234580 399279
rect 234528 399236 234580 399245
rect 305644 399236 305696 399288
rect 213184 399168 213236 399220
rect 204904 399100 204956 399152
rect 312544 399032 312596 399084
rect 319444 398964 319496 399016
rect 135904 398896 135956 398948
rect 291844 398828 291896 398880
rect 3148 395972 3200 396024
rect 10968 395972 11020 396024
rect 290648 393252 290700 393304
rect 579804 393252 579856 393304
rect 3424 380808 3476 380860
rect 225696 380808 225748 380860
rect 291844 369792 291896 369844
rect 580172 369792 580224 369844
rect 2964 367004 3016 367056
rect 226984 367004 227036 367056
rect 326344 358708 326396 358760
rect 580080 358708 580132 358760
rect 290464 346332 290516 346384
rect 579804 346332 579856 346384
rect 277032 338555 277084 338564
rect 277032 338521 277041 338555
rect 277041 338521 277075 338555
rect 277075 338521 277084 338555
rect 277032 338512 277084 338521
rect 263600 338376 263652 338428
rect 265900 338376 265952 338428
rect 247408 338172 247460 338224
rect 247684 338172 247736 338224
rect 253020 338104 253072 338156
rect 253204 338104 253256 338156
rect 270868 338104 270920 338156
rect 3424 338036 3476 338088
rect 13084 338036 13136 338088
rect 125508 338036 125560 338088
rect 107568 337968 107620 338020
rect 240968 338036 241020 338088
rect 247684 338036 247736 338088
rect 255044 338036 255096 338088
rect 261300 338036 261352 338088
rect 271972 338036 272024 338088
rect 240232 337968 240284 338020
rect 262772 337968 262824 338020
rect 279700 338036 279752 338088
rect 282276 338036 282328 338088
rect 291200 338036 291252 338088
rect 115848 337900 115900 337952
rect 100668 337832 100720 337884
rect 253204 337900 253256 337952
rect 254216 337900 254268 337952
rect 263968 337900 264020 337952
rect 268108 337900 268160 337952
rect 240232 337832 240284 337884
rect 246580 337832 246632 337884
rect 280712 337968 280764 338020
rect 281172 337968 281224 338020
rect 287060 337968 287112 338020
rect 283012 337900 283064 337952
rect 297364 337968 297416 338020
rect 290832 337900 290884 337952
rect 35164 337764 35216 337816
rect 232872 337764 232924 337816
rect 241704 337764 241756 337816
rect 264152 337764 264204 337816
rect 39304 337696 39356 337748
rect 233608 337696 233660 337748
rect 242808 337696 242860 337748
rect 265256 337696 265308 337748
rect 32404 337628 32456 337680
rect 231952 337628 232004 337680
rect 258264 337628 258316 337680
rect 277492 337832 277544 337884
rect 284116 337832 284168 337884
rect 288072 337832 288124 337884
rect 298744 337832 298796 337884
rect 302884 337832 302936 337884
rect 276020 337764 276072 337816
rect 280068 337764 280120 337816
rect 28264 337560 28316 337612
rect 232044 337560 232096 337612
rect 233608 337560 233660 337612
rect 234896 337560 234948 337612
rect 246948 337560 247000 337612
rect 257160 337560 257212 337612
rect 14464 337492 14516 337544
rect 230940 337492 230992 337544
rect 240324 337492 240376 337544
rect 242992 337492 243044 337544
rect 257528 337492 257580 337544
rect 15844 337424 15896 337476
rect 231032 337424 231084 337476
rect 231860 337424 231912 337476
rect 235264 337424 235316 337476
rect 242900 337424 242952 337476
rect 251364 337424 251416 337476
rect 257252 337424 257304 337476
rect 10324 337356 10376 337408
rect 230480 337356 230532 337408
rect 231952 337356 232004 337408
rect 253020 337356 253072 337408
rect 260564 337356 260616 337408
rect 266360 337492 266412 337544
rect 266636 337492 266688 337544
rect 266728 337492 266780 337544
rect 280344 337560 280396 337612
rect 280804 337603 280856 337612
rect 280804 337569 280813 337603
rect 280813 337569 280847 337603
rect 280847 337569 280856 337603
rect 280804 337560 280856 337569
rect 287704 337764 287756 337816
rect 301504 337764 301556 337816
rect 289544 337739 289596 337748
rect 289544 337705 289553 337739
rect 289553 337705 289587 337739
rect 289587 337705 289596 337739
rect 289544 337696 289596 337705
rect 284484 337628 284536 337680
rect 287796 337628 287848 337680
rect 320824 337628 320876 337680
rect 283012 337492 283064 337544
rect 283748 337492 283800 337544
rect 284116 337492 284168 337544
rect 284852 337560 284904 337612
rect 285496 337560 285548 337612
rect 316684 337560 316736 337612
rect 315304 337492 315356 337544
rect 265624 337424 265676 337476
rect 346400 337424 346452 337476
rect 273260 337356 273312 337408
rect 273444 337356 273496 337408
rect 276940 337356 276992 337408
rect 277216 337356 277268 337408
rect 280436 337356 280488 337408
rect 285956 337356 286008 337408
rect 226984 337288 227036 337340
rect 258632 337288 258684 337340
rect 264336 337288 264388 337340
rect 264796 337288 264848 337340
rect 268016 337288 268068 337340
rect 269028 337288 269080 337340
rect 281080 337288 281132 337340
rect 222844 337220 222896 337272
rect 241980 337220 242032 337272
rect 242992 337220 243044 337272
rect 246212 337220 246264 337272
rect 259644 337220 259696 337272
rect 262220 337220 262272 337272
rect 266728 337220 266780 337272
rect 267556 337220 267608 337272
rect 277032 337220 277084 337272
rect 277400 337220 277452 337272
rect 290464 337220 290516 337272
rect 225696 337152 225748 337204
rect 245108 337152 245160 337204
rect 260104 337152 260156 337204
rect 260748 337152 260800 337204
rect 262496 337152 262548 337204
rect 262956 337152 263008 337204
rect 268016 337152 268068 337204
rect 268660 337152 268712 337204
rect 277860 337152 277912 337204
rect 279240 337152 279292 337204
rect 280712 337152 280764 337204
rect 281172 337152 281224 337204
rect 281540 337152 281592 337204
rect 228364 337084 228416 337136
rect 254584 337084 254636 337136
rect 257436 337084 257488 337136
rect 246764 337016 246816 337068
rect 246948 337016 247000 337068
rect 252928 337016 252980 337068
rect 256700 337016 256752 337068
rect 258540 337016 258592 337068
rect 248512 336948 248564 337000
rect 251272 336948 251324 337000
rect 252192 336948 252244 337000
rect 252560 336948 252612 337000
rect 256792 336880 256844 336932
rect 257712 336880 257764 336932
rect 258264 336880 258316 336932
rect 259092 336880 259144 336932
rect 251272 336812 251324 336864
rect 253756 336812 253808 336864
rect 256516 336812 256568 336864
rect 257344 336812 257396 336864
rect 258908 336812 258960 336864
rect 259276 336812 259328 336864
rect 259736 337084 259788 337136
rect 263692 337084 263744 337136
rect 263968 337084 264020 337136
rect 264888 337084 264940 337136
rect 267740 337084 267792 337136
rect 277400 337084 277452 337136
rect 278596 337084 278648 337136
rect 282920 337152 282972 337204
rect 283288 337152 283340 337204
rect 283380 337152 283432 337204
rect 284024 337152 284076 337204
rect 284392 337152 284444 337204
rect 285404 337152 285456 337204
rect 287428 337152 287480 337204
rect 287796 337152 287848 337204
rect 291844 337152 291896 337204
rect 289268 337084 289320 337136
rect 289544 337084 289596 337136
rect 260196 337016 260248 337068
rect 269120 337016 269172 337068
rect 269856 337016 269908 337068
rect 273352 337016 273404 337068
rect 274364 337016 274416 337068
rect 274916 337016 274968 337068
rect 263784 336948 263836 337000
rect 264428 336948 264480 337000
rect 266360 336948 266412 337000
rect 267188 336948 267240 337000
rect 269396 336948 269448 337000
rect 261208 336880 261260 336932
rect 261852 336880 261904 336932
rect 269488 336880 269540 336932
rect 270040 336880 270092 336932
rect 230388 336744 230440 336796
rect 231308 336744 231360 336796
rect 237104 336744 237156 336796
rect 239036 336744 239088 336796
rect 240968 336744 241020 336796
rect 241612 336744 241664 336796
rect 244280 336744 244332 336796
rect 245844 336744 245896 336796
rect 254584 336744 254636 336796
rect 255412 336744 255464 336796
rect 257436 336744 257488 336796
rect 257896 336744 257948 336796
rect 258172 336744 258224 336796
rect 258632 336744 258684 336796
rect 258724 336744 258776 336796
rect 259092 336744 259144 336796
rect 259460 336744 259512 336796
rect 260380 336744 260432 336796
rect 233792 336608 233844 336660
rect 236828 336608 236880 336660
rect 262864 336812 262916 336864
rect 263232 336812 263284 336864
rect 264152 336812 264204 336864
rect 264612 336812 264664 336864
rect 265348 336812 265400 336864
rect 266268 336812 266320 336864
rect 267096 336812 267148 336864
rect 267464 336812 267516 336864
rect 267832 336812 267884 336864
rect 268384 336812 268436 336864
rect 269580 336812 269632 336864
rect 270132 336812 270184 336864
rect 261024 336744 261076 336796
rect 261484 336744 261536 336796
rect 262772 336744 262824 336796
rect 263140 336744 263192 336796
rect 265624 336787 265676 336796
rect 265624 336753 265633 336787
rect 265633 336753 265667 336787
rect 265667 336753 265676 336787
rect 265624 336744 265676 336753
rect 266636 336744 266688 336796
rect 262864 336719 262916 336728
rect 262864 336685 262873 336719
rect 262873 336685 262907 336719
rect 262907 336685 262916 336719
rect 262864 336676 262916 336685
rect 266268 336719 266320 336728
rect 266268 336685 266277 336719
rect 266277 336685 266311 336719
rect 266311 336685 266320 336719
rect 266268 336676 266320 336685
rect 266912 336744 266964 336796
rect 267372 336744 267424 336796
rect 267740 336744 267792 336796
rect 268292 336744 268344 336796
rect 267832 336676 267884 336728
rect 268936 336744 268988 336796
rect 269396 336744 269448 336796
rect 269764 336744 269816 336796
rect 273536 336948 273588 337000
rect 274088 336948 274140 337000
rect 275284 336948 275336 337000
rect 275560 336948 275612 337000
rect 276020 336948 276072 337000
rect 276848 336948 276900 337000
rect 273352 336880 273404 336932
rect 273812 336880 273864 336932
rect 273628 336812 273680 336864
rect 274180 336812 274232 336864
rect 276204 336812 276256 336864
rect 277124 336812 277176 336864
rect 271972 336744 272024 336796
rect 272248 336744 272300 336796
rect 272340 336744 272392 336796
rect 272616 336744 272668 336796
rect 272708 336744 272760 336796
rect 269028 336719 269080 336728
rect 269028 336685 269037 336719
rect 269037 336685 269071 336719
rect 269071 336685 269080 336719
rect 269028 336676 269080 336685
rect 270132 336676 270184 336728
rect 261024 336608 261076 336660
rect 272892 336744 272944 336796
rect 273076 336744 273128 336796
rect 273444 336744 273496 336796
rect 273904 336744 273956 336796
rect 273168 336719 273220 336728
rect 273168 336685 273177 336719
rect 273177 336685 273211 336719
rect 273211 336685 273220 336719
rect 273168 336676 273220 336685
rect 273536 336676 273588 336728
rect 274456 336744 274508 336796
rect 275008 336744 275060 336796
rect 275192 336744 275244 336796
rect 275284 336744 275336 336796
rect 275468 336744 275520 336796
rect 276480 336744 276532 336796
rect 276848 336744 276900 336796
rect 277860 337016 277912 337068
rect 278688 337016 278740 337068
rect 281816 337016 281868 337068
rect 282368 337016 282420 337068
rect 284484 337016 284536 337068
rect 285312 337016 285364 337068
rect 285588 337059 285640 337068
rect 285588 337025 285597 337059
rect 285597 337025 285631 337059
rect 285631 337025 285640 337059
rect 285588 337016 285640 337025
rect 286324 337016 286376 337068
rect 286968 337016 287020 337068
rect 277584 336948 277636 337000
rect 278596 336948 278648 337000
rect 280712 336948 280764 337000
rect 281356 336948 281408 337000
rect 282092 336948 282144 337000
rect 282644 336948 282696 337000
rect 288532 336948 288584 337000
rect 290740 336948 290792 337000
rect 282276 336880 282328 336932
rect 282828 336880 282880 336932
rect 277492 336812 277544 336864
rect 278320 336812 278372 336864
rect 279148 336812 279200 336864
rect 280068 336812 280120 336864
rect 280620 336812 280672 336864
rect 281356 336812 281408 336864
rect 281908 336812 281960 336864
rect 282460 336812 282512 336864
rect 282920 336812 282972 336864
rect 274364 336719 274416 336728
rect 274364 336685 274373 336719
rect 274373 336685 274407 336719
rect 274407 336685 274416 336719
rect 274364 336676 274416 336685
rect 277584 336744 277636 336796
rect 277860 336744 277912 336796
rect 277952 336744 278004 336796
rect 278412 336744 278464 336796
rect 279516 336744 279568 336796
rect 279976 336744 280028 336796
rect 280160 336744 280212 336796
rect 280436 336744 280488 336796
rect 280988 336744 281040 336796
rect 281448 336744 281500 336796
rect 282184 336744 282236 336796
rect 282736 336744 282788 336796
rect 288992 336880 289044 336932
rect 292028 336880 292080 336932
rect 283288 336812 283340 336864
rect 283932 336812 283984 336864
rect 284576 336812 284628 336864
rect 285128 336812 285180 336864
rect 285404 336855 285456 336864
rect 285404 336821 285413 336855
rect 285413 336821 285447 336855
rect 285447 336821 285456 336855
rect 285404 336812 285456 336821
rect 286232 336812 286284 336864
rect 286508 336812 286560 336864
rect 287336 336812 287388 336864
rect 287980 336812 288032 336864
rect 288900 336812 288952 336864
rect 290648 336812 290700 336864
rect 283104 336744 283156 336796
rect 283656 336744 283708 336796
rect 284300 336744 284352 336796
rect 278688 336676 278740 336728
rect 284944 336744 284996 336796
rect 285220 336744 285272 336796
rect 287244 336744 287296 336796
rect 287612 336744 287664 336796
rect 285312 336676 285364 336728
rect 294696 336676 294748 336728
rect 489184 336676 489236 336728
rect 273076 336608 273128 336660
rect 280344 336608 280396 336660
rect 293960 336608 294012 336660
rect 240324 336540 240376 336592
rect 296720 336540 296772 336592
rect 230480 336472 230532 336524
rect 253572 336472 253624 336524
rect 260932 336472 260984 336524
rect 219348 336404 219400 336456
rect 252468 336404 252520 336456
rect 262496 336404 262548 336456
rect 314660 336404 314712 336456
rect 209688 336336 209740 336388
rect 242900 336336 242952 336388
rect 268108 336336 268160 336388
rect 331220 336336 331272 336388
rect 180708 336268 180760 336320
rect 248420 336268 248472 336320
rect 262496 336311 262548 336320
rect 262496 336277 262505 336311
rect 262505 336277 262539 336311
rect 262539 336277 262548 336311
rect 262496 336268 262548 336277
rect 265992 336268 266044 336320
rect 349160 336268 349212 336320
rect 169668 336200 169720 336252
rect 247316 336200 247368 336252
rect 275652 336200 275704 336252
rect 443092 336200 443144 336252
rect 126888 336132 126940 336184
rect 71688 336064 71740 336116
rect 237196 336132 237248 336184
rect 291200 336132 291252 336184
rect 483020 336132 483072 336184
rect 236552 336064 236604 336116
rect 236920 336064 236972 336116
rect 284116 336064 284168 336116
rect 521660 336064 521712 336116
rect 48228 335996 48280 336048
rect 233608 335996 233660 336048
rect 287796 335996 287848 336048
rect 557540 335996 557592 336048
rect 233240 335928 233292 335980
rect 234160 335928 234212 335980
rect 251732 335971 251784 335980
rect 251732 335937 251741 335971
rect 251741 335937 251775 335971
rect 251775 335937 251784 335971
rect 251732 335928 251784 335937
rect 300860 335928 300912 335980
rect 232228 335860 232280 335912
rect 232688 335860 232740 335912
rect 232044 335792 232096 335844
rect 232780 335792 232832 335844
rect 233424 335792 233476 335844
rect 234160 335792 234212 335844
rect 236460 335792 236512 335844
rect 236644 335792 236696 335844
rect 242900 335792 242952 335844
rect 243176 335792 243228 335844
rect 254124 335792 254176 335844
rect 254492 335792 254544 335844
rect 232504 335724 232556 335776
rect 232964 335724 233016 335776
rect 248880 335724 248932 335776
rect 255780 335724 255832 335776
rect 258356 335724 258408 335776
rect 258908 335724 258960 335776
rect 262588 335724 262640 335776
rect 263416 335724 263468 335776
rect 232228 335656 232280 335708
rect 232596 335656 232648 335708
rect 233424 335656 233476 335708
rect 233700 335656 233752 335708
rect 234068 335656 234120 335708
rect 234436 335656 234488 335708
rect 236092 335656 236144 335708
rect 236368 335656 236420 335708
rect 229192 335588 229244 335640
rect 230204 335588 230256 335640
rect 230664 335588 230716 335640
rect 231124 335588 231176 335640
rect 232320 335588 232372 335640
rect 232780 335588 232832 335640
rect 234620 335588 234672 335640
rect 235908 335588 235960 335640
rect 230572 335452 230624 335504
rect 231124 335452 231176 335504
rect 230296 335384 230348 335436
rect 227628 335316 227680 335368
rect 231952 335316 232004 335368
rect 237656 335656 237708 335708
rect 238484 335656 238536 335708
rect 239128 335656 239180 335708
rect 239956 335656 240008 335708
rect 240324 335656 240376 335708
rect 240784 335656 240836 335708
rect 243176 335656 243228 335708
rect 243820 335656 243872 335708
rect 244832 335656 244884 335708
rect 245108 335656 245160 335708
rect 248788 335699 248840 335708
rect 248788 335665 248797 335699
rect 248797 335665 248831 335699
rect 248831 335665 248840 335699
rect 248788 335656 248840 335665
rect 256056 335656 256108 335708
rect 266084 335656 266136 335708
rect 266544 335656 266596 335708
rect 267464 335656 267516 335708
rect 268016 335656 268068 335708
rect 268568 335656 268620 335708
rect 268936 335656 268988 335708
rect 276388 335656 276440 335708
rect 277216 335656 277268 335708
rect 280344 335656 280396 335708
rect 280712 335656 280764 335708
rect 280804 335656 280856 335708
rect 284024 335656 284076 335708
rect 286048 335656 286100 335708
rect 286324 335656 286376 335708
rect 289360 335656 289412 335708
rect 236552 335588 236604 335640
rect 236644 335588 236696 335640
rect 237012 335588 237064 335640
rect 238116 335588 238168 335640
rect 238392 335588 238444 335640
rect 239588 335588 239640 335640
rect 239864 335588 239916 335640
rect 240692 335588 240744 335640
rect 241060 335588 241112 335640
rect 242164 335588 242216 335640
rect 242440 335588 242492 335640
rect 242532 335588 242584 335640
rect 242716 335588 242768 335640
rect 243268 335588 243320 335640
rect 243452 335588 243504 335640
rect 244924 335588 244976 335640
rect 245568 335588 245620 335640
rect 245936 335588 245988 335640
rect 246856 335588 246908 335640
rect 247592 335588 247644 335640
rect 247868 335588 247920 335640
rect 248880 335588 248932 335640
rect 249248 335588 249300 335640
rect 249616 335588 249668 335640
rect 250720 335588 250772 335640
rect 251088 335588 251140 335640
rect 251180 335588 251232 335640
rect 251548 335588 251600 335640
rect 252928 335588 252980 335640
rect 253848 335588 253900 335640
rect 254308 335588 254360 335640
rect 254676 335588 254728 335640
rect 239128 335520 239180 335572
rect 240048 335520 240100 335572
rect 255872 335520 255924 335572
rect 236276 335452 236328 335504
rect 237288 335452 237340 335504
rect 248696 335452 248748 335504
rect 249064 335452 249116 335504
rect 249800 335452 249852 335504
rect 250260 335452 250312 335504
rect 251456 335452 251508 335504
rect 251732 335452 251784 335504
rect 240048 335427 240100 335436
rect 240048 335393 240057 335427
rect 240057 335393 240091 335427
rect 240091 335393 240100 335427
rect 240048 335384 240100 335393
rect 236184 335316 236236 335368
rect 236828 335316 236880 335368
rect 251640 335248 251692 335300
rect 236828 335180 236880 335232
rect 236000 335112 236052 335164
rect 236368 335112 236420 335164
rect 224868 335044 224920 335096
rect 246948 335044 247000 335096
rect 251732 335044 251784 335096
rect 255504 335044 255556 335096
rect 269488 335588 269540 335640
rect 270316 335588 270368 335640
rect 272340 335588 272392 335640
rect 272524 335588 272576 335640
rect 265716 335452 265768 335504
rect 266084 335452 266136 335504
rect 268016 335452 268068 335504
rect 268568 335452 268620 335504
rect 268844 335452 268896 335504
rect 272524 335495 272576 335504
rect 272524 335461 272533 335495
rect 272533 335461 272567 335495
rect 272567 335461 272576 335495
rect 272524 335452 272576 335461
rect 279056 335452 279108 335504
rect 279608 335452 279660 335504
rect 280712 335452 280764 335504
rect 283472 335452 283524 335504
rect 284024 335452 284076 335504
rect 284208 335452 284260 335504
rect 288624 335452 288676 335504
rect 289268 335452 289320 335504
rect 277032 335427 277084 335436
rect 277032 335393 277041 335427
rect 277041 335393 277075 335427
rect 277075 335393 277084 335427
rect 277032 335384 277084 335393
rect 278964 335384 279016 335436
rect 279516 335384 279568 335436
rect 283564 335384 283616 335436
rect 284116 335384 284168 335436
rect 265164 335359 265216 335368
rect 265164 335325 265173 335359
rect 265173 335325 265207 335359
rect 265207 335325 265216 335359
rect 265164 335316 265216 335325
rect 265440 335316 265492 335368
rect 265532 335316 265584 335368
rect 266360 335316 266412 335368
rect 267004 335316 267056 335368
rect 280344 335316 280396 335368
rect 280528 335359 280580 335368
rect 280528 335325 280537 335359
rect 280537 335325 280571 335359
rect 280571 335325 280580 335359
rect 280528 335316 280580 335325
rect 282920 335316 282972 335368
rect 283288 335316 283340 335368
rect 286140 335316 286192 335368
rect 286876 335316 286928 335368
rect 278780 335180 278832 335232
rect 279148 335180 279200 335232
rect 283472 335180 283524 335232
rect 281080 335112 281132 335164
rect 305000 335112 305052 335164
rect 260748 335044 260800 335096
rect 292580 335044 292632 335096
rect 223488 334976 223540 335028
rect 252836 334976 252888 335028
rect 262036 334976 262088 335028
rect 311900 334976 311952 335028
rect 212448 334908 212500 334960
rect 265900 334908 265952 334960
rect 327080 334908 327132 334960
rect 176568 334840 176620 334892
rect 248052 334840 248104 334892
rect 353300 334840 353352 334892
rect 162768 334772 162820 334824
rect 240232 334772 240284 334824
rect 273260 334772 273312 334824
rect 422300 334772 422352 334824
rect 160008 334704 160060 334756
rect 242992 334704 243044 334756
rect 500960 334704 501012 334756
rect 74448 334636 74500 334688
rect 237564 334636 237616 334688
rect 256884 334636 256936 334688
rect 257160 334636 257212 334688
rect 285496 334636 285548 334688
rect 532700 334636 532752 334688
rect 52368 334568 52420 334620
rect 231860 334568 231912 334620
rect 240232 334568 240284 334620
rect 240508 334568 240560 334620
rect 262220 334568 262272 334620
rect 287060 334568 287112 334620
rect 289636 334568 289688 334620
rect 573364 334568 573416 334620
rect 240692 334364 240744 334416
rect 241244 334364 241296 334416
rect 233332 334296 233384 334348
rect 245752 334092 245804 334144
rect 246212 334092 246264 334144
rect 270776 334092 270828 334144
rect 271788 334092 271840 334144
rect 276296 334092 276348 334144
rect 276480 334092 276532 334144
rect 251916 333956 251968 334008
rect 252376 333956 252428 334008
rect 254952 333888 255004 333940
rect 233608 333820 233660 333872
rect 234068 333820 234120 333872
rect 241520 333752 241572 333804
rect 241888 333752 241940 333804
rect 220728 333616 220780 333668
rect 252652 333752 252704 333804
rect 261668 333752 261720 333804
rect 216588 333548 216640 333600
rect 252468 333684 252520 333736
rect 307760 333752 307812 333804
rect 247408 333616 247460 333668
rect 262956 333616 263008 333668
rect 316040 333616 316092 333668
rect 173808 333480 173860 333532
rect 261024 333548 261076 333600
rect 261576 333548 261628 333600
rect 264704 333548 264756 333600
rect 338120 333548 338172 333600
rect 254032 333480 254084 333532
rect 254216 333480 254268 333532
rect 268936 333480 268988 333532
rect 374000 333480 374052 333532
rect 142068 333412 142120 333464
rect 244464 333412 244516 333464
rect 247316 333412 247368 333464
rect 247960 333412 248012 333464
rect 262496 333412 262548 333464
rect 262864 333412 262916 333464
rect 271236 333412 271288 333464
rect 400312 333412 400364 333464
rect 129648 333344 129700 333396
rect 242900 333344 242952 333396
rect 247408 333344 247460 333396
rect 248328 333344 248380 333396
rect 259828 333344 259880 333396
rect 260196 333344 260248 333396
rect 275560 333344 275612 333396
rect 440240 333344 440292 333396
rect 92388 333276 92440 333328
rect 239404 333276 239456 333328
rect 250536 333319 250588 333328
rect 250536 333285 250545 333319
rect 250545 333285 250579 333319
rect 250579 333285 250588 333319
rect 250536 333276 250588 333285
rect 261300 333276 261352 333328
rect 261760 333276 261812 333328
rect 271880 333276 271932 333328
rect 272248 333276 272300 333328
rect 276112 333276 276164 333328
rect 276572 333276 276624 333328
rect 277860 333276 277912 333328
rect 278504 333276 278556 333328
rect 284208 333276 284260 333328
rect 518900 333276 518952 333328
rect 56508 333208 56560 333260
rect 235632 333208 235684 333260
rect 286968 333208 287020 333260
rect 546500 333208 546552 333260
rect 274824 333004 274876 333056
rect 275744 333004 275796 333056
rect 261208 332936 261260 332988
rect 261392 332936 261444 332988
rect 231492 332596 231544 332648
rect 231768 332596 231820 332648
rect 244372 332596 244424 332648
rect 245476 332596 245528 332648
rect 264796 332392 264848 332444
rect 260472 332324 260524 332376
rect 296812 332324 296864 332376
rect 211068 332188 211120 332240
rect 251364 332188 251416 332240
rect 270868 332188 270920 332240
rect 271328 332188 271380 332240
rect 184848 332120 184900 332172
rect 270960 332120 271012 332172
rect 271696 332120 271748 332172
rect 281172 332256 281224 332308
rect 318800 332256 318852 332308
rect 333980 332188 334032 332240
rect 356060 332120 356112 332172
rect 153108 332052 153160 332104
rect 245660 332052 245712 332104
rect 271604 332052 271656 332104
rect 404360 332052 404412 332104
rect 144828 331984 144880 332036
rect 245108 331984 245160 332036
rect 266452 331984 266504 332036
rect 266728 331984 266780 332036
rect 278228 331984 278280 332036
rect 467840 331984 467892 332036
rect 89628 331916 89680 331968
rect 237104 331916 237156 331968
rect 285404 331916 285456 331968
rect 528560 331916 528612 331968
rect 49608 331848 49660 331900
rect 234988 331848 235040 331900
rect 289544 331848 289596 331900
rect 574744 331848 574796 331900
rect 234068 331780 234120 331832
rect 234344 331780 234396 331832
rect 234804 331644 234856 331696
rect 235080 331644 235132 331696
rect 235540 331576 235592 331628
rect 235816 331576 235868 331628
rect 262680 331304 262732 331356
rect 235724 331236 235776 331288
rect 233516 331168 233568 331220
rect 233700 331168 233752 331220
rect 261944 331236 261996 331288
rect 263232 331236 263284 331288
rect 275836 331304 275888 331356
rect 281724 331304 281776 331356
rect 277308 331279 277360 331288
rect 277308 331245 277317 331279
rect 277317 331245 277351 331279
rect 277351 331245 277360 331279
rect 277308 331236 277360 331245
rect 258264 331168 258316 331220
rect 259368 331168 259420 331220
rect 260840 331168 260892 331220
rect 275008 331168 275060 331220
rect 235724 331100 235776 331152
rect 287428 331236 287480 331288
rect 287980 331168 288032 331220
rect 284944 331100 284996 331152
rect 287152 331100 287204 331152
rect 287704 331100 287756 331152
rect 229008 330828 229060 330880
rect 253296 330828 253348 330880
rect 262128 330828 262180 330880
rect 313280 330828 313332 330880
rect 208308 330760 208360 330812
rect 248420 330760 248472 330812
rect 270500 330760 270552 330812
rect 393320 330760 393372 330812
rect 151728 330692 151780 330744
rect 244372 330692 244424 330744
rect 272616 330692 272668 330744
rect 411260 330692 411312 330744
rect 128268 330624 128320 330676
rect 243084 330624 243136 330676
rect 277216 330624 277268 330676
rect 451280 330624 451332 330676
rect 78588 330556 78640 330608
rect 237932 330556 237984 330608
rect 278596 330556 278648 330608
rect 462320 330556 462372 330608
rect 34428 330488 34480 330540
rect 234160 330488 234212 330540
rect 285588 330488 285640 330540
rect 536840 330488 536892 330540
rect 288624 329579 288676 329588
rect 288624 329545 288633 329579
rect 288633 329545 288667 329579
rect 288667 329545 288676 329579
rect 288624 329536 288676 329545
rect 263508 329400 263560 329452
rect 322940 329400 322992 329452
rect 206928 329332 206980 329384
rect 251548 329332 251600 329384
rect 265624 329332 265676 329384
rect 342260 329332 342312 329384
rect 157248 329264 157300 329316
rect 246028 329264 246080 329316
rect 280344 329264 280396 329316
rect 397460 329264 397512 329316
rect 155868 329196 155920 329248
rect 244280 329196 244332 329248
rect 273352 329196 273404 329248
rect 425152 329196 425204 329248
rect 85488 329128 85540 329180
rect 238668 329128 238720 329180
rect 277400 329128 277452 329180
rect 471980 329128 472032 329180
rect 38568 329060 38620 329112
rect 233424 329060 233476 329112
rect 539600 329060 539652 329112
rect 251824 328992 251876 329044
rect 254860 328992 254912 329044
rect 229560 328491 229612 328500
rect 229560 328457 229569 328491
rect 229569 328457 229603 328491
rect 229603 328457 229612 328491
rect 229560 328448 229612 328457
rect 250628 328448 250680 328500
rect 252008 328448 252060 328500
rect 253480 328448 253532 328500
rect 254676 328491 254728 328500
rect 254676 328457 254685 328491
rect 254685 328457 254719 328491
rect 254719 328457 254728 328491
rect 254676 328448 254728 328457
rect 255872 328491 255924 328500
rect 255872 328457 255881 328491
rect 255881 328457 255915 328491
rect 255915 328457 255924 328491
rect 255872 328448 255924 328457
rect 261760 328491 261812 328500
rect 261760 328457 261769 328491
rect 261769 328457 261803 328491
rect 261803 328457 261812 328491
rect 261760 328448 261812 328457
rect 237012 328423 237064 328432
rect 237012 328389 237021 328423
rect 237021 328389 237055 328423
rect 237055 328389 237064 328423
rect 237012 328380 237064 328389
rect 245384 328380 245436 328432
rect 257160 328380 257212 328432
rect 257252 328380 257304 328432
rect 256424 328108 256476 328160
rect 256700 328108 256752 328160
rect 260932 328108 260984 328160
rect 299480 328108 299532 328160
rect 264428 328040 264480 328092
rect 328460 328040 328512 328092
rect 215208 327972 215260 328024
rect 251640 327972 251692 328024
rect 269304 327972 269356 328024
rect 382280 327972 382332 328024
rect 168288 327904 168340 327956
rect 247132 327904 247184 327956
rect 283288 327904 283340 327956
rect 408500 327904 408552 327956
rect 139308 327836 139360 327888
rect 244188 327836 244240 327888
rect 273628 327836 273680 327888
rect 429200 327836 429252 327888
rect 96528 327768 96580 327820
rect 239772 327768 239824 327820
rect 281908 327768 281960 327820
rect 509240 327768 509292 327820
rect 53748 327700 53800 327752
rect 235356 327700 235408 327752
rect 259000 327700 259052 327752
rect 281540 327700 281592 327752
rect 286692 327700 286744 327752
rect 550640 327700 550692 327752
rect 265440 327403 265492 327412
rect 265440 327369 265449 327403
rect 265449 327369 265483 327403
rect 265483 327369 265492 327403
rect 265440 327360 265492 327369
rect 233976 327131 234028 327140
rect 233976 327097 233985 327131
rect 233985 327097 234019 327131
rect 234019 327097 234028 327131
rect 233976 327088 234028 327097
rect 266268 327131 266320 327140
rect 266268 327097 266277 327131
rect 266277 327097 266311 327131
rect 266311 327097 266320 327131
rect 266268 327088 266320 327097
rect 269028 327131 269080 327140
rect 269028 327097 269037 327131
rect 269037 327097 269071 327131
rect 269071 327097 269080 327131
rect 269028 327088 269080 327097
rect 273168 327131 273220 327140
rect 273168 327097 273177 327131
rect 273177 327097 273211 327131
rect 273211 327097 273220 327131
rect 273168 327088 273220 327097
rect 274364 327131 274416 327140
rect 274364 327097 274373 327131
rect 274373 327097 274407 327131
rect 274407 327097 274416 327131
rect 274364 327088 274416 327097
rect 265164 327020 265216 327072
rect 265256 327020 265308 327072
rect 265532 327020 265584 327072
rect 265624 327020 265676 327072
rect 277032 327020 277084 327072
rect 277124 327020 277176 327072
rect 263876 326952 263928 327004
rect 264336 326952 264388 327004
rect 269580 326952 269632 327004
rect 269488 326748 269540 326800
rect 274732 326748 274784 326800
rect 347780 326748 347832 326800
rect 263324 326680 263376 326732
rect 320180 326680 320232 326732
rect 222108 326612 222160 326664
rect 252744 326612 252796 326664
rect 266360 326612 266412 326664
rect 360200 326612 360252 326664
rect 171048 326544 171100 326596
rect 247592 326544 247644 326596
rect 273076 326544 273128 326596
rect 415400 326544 415452 326596
rect 159916 326476 159968 326528
rect 246396 326476 246448 326528
rect 279792 326476 279844 326528
rect 433340 326476 433392 326528
rect 56416 326408 56468 326460
rect 235724 326408 235776 326460
rect 19984 326340 20036 326392
rect 231492 326340 231544 326392
rect 251916 326340 251968 326392
rect 252100 326340 252152 326392
rect 264060 326340 264112 326392
rect 264244 326340 264296 326392
rect 266636 326340 266688 326392
rect 266820 326340 266872 326392
rect 267372 326340 267424 326392
rect 267648 326340 267700 326392
rect 267740 326340 267792 326392
rect 267924 326340 267976 326392
rect 272156 326340 272208 326392
rect 272984 326340 273036 326392
rect 279332 326340 279384 326392
rect 279516 326340 279568 326392
rect 261668 326272 261720 326324
rect 279516 326204 279568 326256
rect 282092 326340 282144 326392
rect 282368 326340 282420 326392
rect 284760 326340 284812 326392
rect 285036 326340 285088 326392
rect 287428 326340 287480 326392
rect 287796 326340 287848 326392
rect 284392 326272 284444 326324
rect 284852 326272 284904 326324
rect 287612 326272 287664 326324
rect 288348 326272 288400 326324
rect 347780 326408 347832 326460
rect 465080 326408 465132 326460
rect 290832 326340 290884 326392
rect 554780 326340 554832 326392
rect 279240 326136 279292 326188
rect 261668 326068 261720 326120
rect 278964 326068 279016 326120
rect 279976 326068 280028 326120
rect 280252 326068 280304 326120
rect 281448 326068 281500 326120
rect 274364 325635 274416 325644
rect 274364 325601 274373 325635
rect 274373 325601 274407 325635
rect 274407 325601 274416 325635
rect 274364 325592 274416 325601
rect 261852 325252 261904 325304
rect 303620 325252 303672 325304
rect 268384 325184 268436 325236
rect 367100 325184 367152 325236
rect 213828 325116 213880 325168
rect 251456 325116 251508 325168
rect 270776 325116 270828 325168
rect 398840 325116 398892 325168
rect 141976 325048 142028 325100
rect 244740 325048 244792 325100
rect 272892 325048 272944 325100
rect 418160 325048 418212 325100
rect 103428 324980 103480 325032
rect 240232 324980 240284 325032
rect 281816 324980 281868 325032
rect 502340 324980 502392 325032
rect 42064 324912 42116 324964
rect 233332 324912 233384 324964
rect 288164 324912 288216 324964
rect 564440 324912 564492 324964
rect 260380 324300 260432 324352
rect 260656 324300 260708 324352
rect 262680 324300 262732 324352
rect 263600 324300 263652 324352
rect 277400 324300 277452 324352
rect 262312 323892 262364 323944
rect 313372 323892 313424 323944
rect 269764 323824 269816 323876
rect 385040 323824 385092 323876
rect 217968 323756 218020 323808
rect 252376 323756 252428 323808
rect 279148 323756 279200 323808
rect 436100 323756 436152 323808
rect 165528 323688 165580 323740
rect 245936 323688 245988 323740
rect 275192 323688 275244 323740
rect 437480 323688 437532 323740
rect 114468 323620 114520 323672
rect 240784 323620 240836 323672
rect 285680 323620 285732 323672
rect 540980 323620 541032 323672
rect 46204 323552 46256 323604
rect 234528 323552 234580 323604
rect 289176 323595 289228 323604
rect 289176 323561 289185 323595
rect 289185 323561 289219 323595
rect 289219 323561 289228 323595
rect 289176 323552 289228 323561
rect 290740 323552 290792 323604
rect 568580 323552 568632 323604
rect 287980 322872 288032 322924
rect 288256 322872 288308 322924
rect 290556 322872 290608 322924
rect 580172 322872 580224 322924
rect 226248 322396 226300 322448
rect 253112 322396 253164 322448
rect 263048 322396 263100 322448
rect 321560 322396 321612 322448
rect 146208 322328 146260 322380
rect 245568 322328 245620 322380
rect 276756 322328 276808 322380
rect 454040 322328 454092 322380
rect 121368 322260 121420 322312
rect 242348 322260 242400 322312
rect 277492 322260 277544 322312
rect 469220 322260 469272 322312
rect 67548 322192 67600 322244
rect 233884 322192 233936 322244
rect 289268 322192 289320 322244
rect 567844 322192 567896 322244
rect 260656 321895 260708 321904
rect 260656 321861 260665 321895
rect 260665 321861 260699 321895
rect 260699 321861 260708 321895
rect 260656 321852 260708 321861
rect 233516 321580 233568 321632
rect 233700 321580 233752 321632
rect 289084 321648 289136 321700
rect 288992 321512 289044 321564
rect 270592 321036 270644 321088
rect 394700 321036 394752 321088
rect 150348 320968 150400 321020
rect 245200 320968 245252 321020
rect 276572 320968 276624 321020
rect 448520 320968 448572 321020
rect 125416 320900 125468 320952
rect 242532 320900 242584 320952
rect 279332 320900 279384 320952
rect 476120 320900 476172 320952
rect 82728 320832 82780 320884
rect 238300 320832 238352 320884
rect 290648 320832 290700 320884
rect 571432 320832 571484 320884
rect 245200 320331 245252 320340
rect 245200 320297 245209 320331
rect 245209 320297 245243 320331
rect 245243 320297 245252 320331
rect 245200 320288 245252 320297
rect 261668 319676 261720 319728
rect 306380 319676 306432 319728
rect 267096 319608 267148 319660
rect 364340 319608 364392 319660
rect 210976 319540 211028 319592
rect 251732 319540 251784 319592
rect 274548 319540 274600 319592
rect 433432 319540 433484 319592
rect 154488 319472 154540 319524
rect 246212 319472 246264 319524
rect 280712 319472 280764 319524
rect 487160 319472 487212 319524
rect 13728 319404 13780 319456
rect 229744 319404 229796 319456
rect 287704 319404 287756 319456
rect 554872 319404 554924 319456
rect 233976 318860 234028 318912
rect 237104 318792 237156 318844
rect 267464 318835 267516 318844
rect 267464 318801 267473 318835
rect 267473 318801 267507 318835
rect 267507 318801 267516 318835
rect 267464 318792 267516 318801
rect 289268 318792 289320 318844
rect 229560 318724 229612 318776
rect 233976 318724 234028 318776
rect 245200 318767 245252 318776
rect 245200 318733 245209 318767
rect 245209 318733 245243 318767
rect 245243 318733 245252 318767
rect 245200 318724 245252 318733
rect 264520 318248 264572 318300
rect 335360 318248 335412 318300
rect 136548 318180 136600 318232
rect 243912 318180 243964 318232
rect 270868 318180 270920 318232
rect 401600 318180 401652 318232
rect 99288 318112 99340 318164
rect 240140 318112 240192 318164
rect 280528 318112 280580 318164
rect 447140 318112 447192 318164
rect 50988 318044 51040 318096
rect 234896 318044 234948 318096
rect 257436 318044 257488 318096
rect 270500 318044 270552 318096
rect 282368 318044 282420 318096
rect 505100 318044 505152 318096
rect 267464 317475 267516 317484
rect 267464 317441 267473 317475
rect 267473 317441 267507 317475
rect 267507 317441 267516 317475
rect 267464 317432 267516 317441
rect 235172 317364 235224 317416
rect 268292 316888 268344 316940
rect 371240 316888 371292 316940
rect 272064 316820 272116 316872
rect 408592 316820 408644 316872
rect 140688 316752 140740 316804
rect 244556 316752 244608 316804
rect 276296 316752 276348 316804
rect 458180 316752 458232 316804
rect 110328 316684 110380 316736
rect 240692 316684 240744 316736
rect 279332 316684 279384 316736
rect 279792 316684 279844 316736
rect 283656 316684 283708 316736
rect 516140 316684 516192 316736
rect 254860 316115 254912 316124
rect 254860 316081 254869 316115
rect 254869 316081 254903 316115
rect 254903 316081 254912 316115
rect 254860 316072 254912 316081
rect 256608 316072 256660 316124
rect 256700 316072 256752 316124
rect 274364 316047 274416 316056
rect 274364 316013 274373 316047
rect 274373 316013 274407 316047
rect 274407 316013 274416 316047
rect 274364 316004 274416 316013
rect 258264 315460 258316 315512
rect 285680 315460 285732 315512
rect 274088 315392 274140 315444
rect 423680 315392 423732 315444
rect 143448 315324 143500 315376
rect 244832 315324 244884 315376
rect 283472 315324 283524 315376
rect 460940 315324 460992 315376
rect 24124 315256 24176 315308
rect 232688 315256 232740 315308
rect 285220 315256 285272 315308
rect 534080 315256 534132 315308
rect 260656 314687 260708 314696
rect 260656 314653 260665 314687
rect 260665 314653 260699 314687
rect 260699 314653 260708 314687
rect 260656 314644 260708 314653
rect 262404 314644 262456 314696
rect 262588 314644 262640 314696
rect 275376 314032 275428 314084
rect 441620 314032 441672 314084
rect 147588 313964 147640 314016
rect 245016 313964 245068 314016
rect 279424 313964 279476 314016
rect 478880 313964 478932 314016
rect 31024 313896 31076 313948
rect 232044 313896 232096 313948
rect 261760 313896 261812 313948
rect 278780 313896 278832 313948
rect 286416 313896 286468 313948
rect 545120 313896 545172 313948
rect 278412 312672 278464 312724
rect 466460 312672 466512 312724
rect 158628 312604 158680 312656
rect 246120 312604 246172 312656
rect 279516 312604 279568 312656
rect 484400 312604 484452 312656
rect 31668 312536 31720 312588
rect 233148 312536 233200 312588
rect 286784 312536 286836 312588
rect 552020 312536 552072 312588
rect 245200 311831 245252 311840
rect 245200 311797 245209 311831
rect 245209 311797 245243 311831
rect 245243 311797 245252 311831
rect 245200 311788 245252 311797
rect 500224 311788 500276 311840
rect 580172 311788 580224 311840
rect 260840 311312 260892 311364
rect 310520 311312 310572 311364
rect 268568 311244 268620 311296
rect 378140 311244 378192 311296
rect 161388 311176 161440 311228
rect 246488 311176 246540 311228
rect 273628 311176 273680 311228
rect 273996 311176 274048 311228
rect 280896 311176 280948 311228
rect 491300 311176 491352 311228
rect 50344 311108 50396 311160
rect 235908 311108 235960 311160
rect 289452 311108 289504 311160
rect 571984 311108 572036 311160
rect 229468 310811 229520 310820
rect 229468 310777 229477 310811
rect 229477 310777 229511 310811
rect 229511 310777 229520 310811
rect 229468 310768 229520 310777
rect 277768 310088 277820 310140
rect 277952 310088 278004 310140
rect 263232 309952 263284 310004
rect 317420 309952 317472 310004
rect 269948 309884 270000 309936
rect 389180 309884 389232 309936
rect 280988 309816 281040 309868
rect 494060 309816 494112 309868
rect 107476 309748 107528 309800
rect 240508 309748 240560 309800
rect 287428 309748 287480 309800
rect 556804 309748 556856 309800
rect 3424 309068 3476 309120
rect 211804 309068 211856 309120
rect 229468 309111 229520 309120
rect 229468 309077 229477 309111
rect 229477 309077 229511 309111
rect 229511 309077 229520 309111
rect 229468 309068 229520 309077
rect 273628 309111 273680 309120
rect 273628 309077 273637 309111
rect 273637 309077 273671 309111
rect 273671 309077 273680 309111
rect 273628 309068 273680 309077
rect 263968 308524 264020 308576
rect 339500 308524 339552 308576
rect 281080 308456 281132 308508
rect 498200 308456 498252 308508
rect 288624 308388 288676 308440
rect 574836 308388 574888 308440
rect 233976 307708 234028 307760
rect 237288 307708 237340 307760
rect 233792 307640 233844 307692
rect 269672 307844 269724 307896
rect 269580 307640 269632 307692
rect 270960 307096 271012 307148
rect 405740 307096 405792 307148
rect 43444 307028 43496 307080
rect 233700 307028 233752 307080
rect 279332 307028 279384 307080
rect 279792 307028 279844 307080
rect 282184 307028 282236 307080
rect 512000 307028 512052 307080
rect 262588 306484 262640 306536
rect 268844 306416 268896 306468
rect 269028 306416 269080 306468
rect 262680 306348 262732 306400
rect 264244 306348 264296 306400
rect 264336 306348 264388 306400
rect 272432 305668 272484 305720
rect 412640 305668 412692 305720
rect 38476 305600 38528 305652
rect 233608 305600 233660 305652
rect 284024 305600 284076 305652
rect 520280 305600 520332 305652
rect 254768 304920 254820 304972
rect 255044 304920 255096 304972
rect 273168 304308 273220 304360
rect 419540 304308 419592 304360
rect 42708 304240 42760 304292
rect 234252 304240 234304 304292
rect 283840 304240 283892 304292
rect 523040 304240 523092 304292
rect 273444 302948 273496 303000
rect 426440 302948 426492 303000
rect 283932 302880 283984 302932
rect 527180 302880 527232 302932
rect 277768 302132 277820 302184
rect 277952 302132 278004 302184
rect 235356 301928 235408 301980
rect 275560 301520 275612 301572
rect 444380 301520 444432 301572
rect 285128 301452 285180 301504
rect 529940 301452 529992 301504
rect 276020 300160 276072 300212
rect 455420 300160 455472 300212
rect 284484 300092 284536 300144
rect 536932 300092 536984 300144
rect 229560 299480 229612 299532
rect 266176 299480 266228 299532
rect 266268 299480 266320 299532
rect 271144 299480 271196 299532
rect 271512 299480 271564 299532
rect 274456 299548 274508 299600
rect 274364 299412 274416 299464
rect 302976 299412 303028 299464
rect 579804 299412 579856 299464
rect 277584 298732 277636 298784
rect 473360 298732 473412 298784
rect 237196 298163 237248 298172
rect 237196 298129 237205 298163
rect 237205 298129 237239 298163
rect 237239 298129 237248 298163
rect 237196 298120 237248 298129
rect 235356 298095 235408 298104
rect 235356 298061 235365 298095
rect 235365 298061 235399 298095
rect 235399 298061 235408 298095
rect 235356 298052 235408 298061
rect 284668 298052 284720 298104
rect 288348 298095 288400 298104
rect 288348 298061 288357 298095
rect 288357 298061 288391 298095
rect 288391 298061 288400 298095
rect 288348 298052 288400 298061
rect 289268 298052 289320 298104
rect 286600 297440 286652 297492
rect 547880 297440 547932 297492
rect 288716 297372 288768 297424
rect 570604 297372 570656 297424
rect 264244 296692 264296 296744
rect 264428 296692 264480 296744
rect 273628 296735 273680 296744
rect 273628 296701 273637 296735
rect 273637 296701 273671 296735
rect 273671 296701 273680 296735
rect 273628 296692 273680 296701
rect 252192 296624 252244 296676
rect 252284 296624 252336 296676
rect 288992 296012 289044 296064
rect 482284 296012 482336 296064
rect 287888 295944 287940 295996
rect 563060 295944 563112 295996
rect 3056 295264 3108 295316
rect 227168 295264 227220 295316
rect 254860 295307 254912 295316
rect 254860 295273 254869 295307
rect 254869 295273 254903 295307
rect 254903 295273 254912 295307
rect 254860 295264 254912 295273
rect 255872 295264 255924 295316
rect 256424 295264 256476 295316
rect 256608 295264 256660 295316
rect 287980 294584 288032 294636
rect 560944 294584 560996 294636
rect 262496 293292 262548 293344
rect 324320 293292 324372 293344
rect 292028 293224 292080 293276
rect 572720 293224 572772 293276
rect 243544 292612 243596 292664
rect 243360 292544 243412 292596
rect 272800 291864 272852 291916
rect 416872 291864 416924 291916
rect 282644 291796 282696 291848
rect 506480 291796 506532 291848
rect 274180 290504 274232 290556
rect 430580 290504 430632 290556
rect 277124 290436 277176 290488
rect 277308 290436 277360 290488
rect 285772 290436 285824 290488
rect 542360 290436 542412 290488
rect 235356 289799 235408 289808
rect 235356 289765 235365 289799
rect 235365 289765 235399 289799
rect 235399 289765 235408 289799
rect 235356 289756 235408 289765
rect 273812 289756 273864 289808
rect 273904 289756 273956 289808
rect 277124 289756 277176 289808
rect 277308 289756 277360 289808
rect 276848 289144 276900 289196
rect 451372 289144 451424 289196
rect 255780 289119 255832 289128
rect 255780 289085 255789 289119
rect 255789 289085 255823 289119
rect 255823 289085 255832 289119
rect 255780 289076 255832 289085
rect 556160 289076 556212 289128
rect 284576 288439 284628 288448
rect 284576 288405 284585 288439
rect 284585 288405 284619 288439
rect 284619 288405 284628 288439
rect 284576 288396 284628 288405
rect 289084 288439 289136 288448
rect 289084 288405 289093 288439
rect 289093 288405 289127 288439
rect 289127 288405 289136 288439
rect 289084 288396 289136 288405
rect 276940 287648 276992 287700
rect 459652 287648 459704 287700
rect 257160 287036 257212 287088
rect 257252 287036 257304 287088
rect 279608 286288 279660 286340
rect 477500 286288 477552 286340
rect 254860 285719 254912 285728
rect 254860 285685 254869 285719
rect 254869 285685 254903 285719
rect 254903 285685 254912 285719
rect 254860 285676 254912 285685
rect 279700 284928 279752 284980
rect 480260 284928 480312 284980
rect 277032 283568 277084 283620
rect 277216 283568 277268 283620
rect 279792 283568 279844 283620
rect 485780 283568 485832 283620
rect 233700 282888 233752 282940
rect 233884 282888 233936 282940
rect 280160 282140 280212 282192
rect 488540 282140 488592 282192
rect 281264 280780 281316 280832
rect 492680 280780 492732 280832
rect 250536 280168 250588 280220
rect 250720 280168 250772 280220
rect 229560 280143 229612 280152
rect 229560 280109 229569 280143
rect 229569 280109 229603 280143
rect 229603 280109 229612 280143
rect 229560 280100 229612 280109
rect 235540 280143 235592 280152
rect 235540 280109 235549 280143
rect 235549 280109 235583 280143
rect 235583 280109 235592 280143
rect 235540 280100 235592 280109
rect 237104 280100 237156 280152
rect 237196 280100 237248 280152
rect 281356 279420 281408 279472
rect 495440 279420 495492 279472
rect 235172 278740 235224 278792
rect 235356 278740 235408 278792
rect 284944 277992 284996 278044
rect 502432 277992 502484 278044
rect 282000 276632 282052 276684
rect 510620 276632 510672 276684
rect 309784 275952 309836 276004
rect 580172 275952 580224 276004
rect 255780 274635 255832 274644
rect 255780 274601 255789 274635
rect 255789 274601 255823 274635
rect 255823 274601 255832 274635
rect 255780 274592 255832 274601
rect 277216 274635 277268 274644
rect 277216 274601 277225 274635
rect 277225 274601 277259 274635
rect 277259 274601 277268 274635
rect 277216 274592 277268 274601
rect 235264 273912 235316 273964
rect 282276 273912 282328 273964
rect 513380 273912 513432 273964
rect 250260 273096 250312 273148
rect 250720 273096 250772 273148
rect 283012 272484 283064 272536
rect 517520 272484 517572 272536
rect 284116 271124 284168 271176
rect 520372 271124 520424 271176
rect 238852 270580 238904 270632
rect 229652 270512 229704 270564
rect 235540 270555 235592 270564
rect 235540 270521 235549 270555
rect 235549 270521 235583 270555
rect 235583 270521 235592 270555
rect 235540 270512 235592 270521
rect 238944 270512 238996 270564
rect 259920 270580 259972 270632
rect 259828 270444 259880 270496
rect 283196 269764 283248 269816
rect 524420 269764 524472 269816
rect 285312 268336 285364 268388
rect 528652 268336 528704 268388
rect 284668 266976 284720 267028
rect 531320 266976 531372 267028
rect 2872 266296 2924 266348
rect 209044 266296 209096 266348
rect 276940 266296 276992 266348
rect 284760 265616 284812 265668
rect 535460 265616 535512 265668
rect 255780 264979 255832 264988
rect 255780 264945 255789 264979
rect 255789 264945 255823 264979
rect 255823 264945 255832 264979
rect 255780 264936 255832 264945
rect 277216 264979 277268 264988
rect 277216 264945 277225 264979
rect 277225 264945 277259 264979
rect 277259 264945 277268 264979
rect 277216 264936 277268 264945
rect 498844 264868 498896 264920
rect 580172 264868 580224 264920
rect 288900 264188 288952 264240
rect 475384 264188 475436 264240
rect 233700 263576 233752 263628
rect 233884 263576 233936 263628
rect 273628 263576 273680 263628
rect 273720 263508 273772 263560
rect 285956 262828 286008 262880
rect 546592 262828 546644 262880
rect 286048 261468 286100 261520
rect 549260 261468 549312 261520
rect 235172 260899 235224 260908
rect 235172 260865 235181 260899
rect 235181 260865 235215 260899
rect 235215 260865 235224 260899
rect 235172 260856 235224 260865
rect 257160 260856 257212 260908
rect 257252 260856 257304 260908
rect 229560 260831 229612 260840
rect 229560 260797 229569 260831
rect 229569 260797 229603 260831
rect 229603 260797 229612 260831
rect 229560 260788 229612 260797
rect 250444 260788 250496 260840
rect 286140 260108 286192 260160
rect 553400 260108 553452 260160
rect 235172 259403 235224 259412
rect 235172 259369 235181 259403
rect 235181 259369 235215 259403
rect 235215 259369 235224 259403
rect 235172 259360 235224 259369
rect 287244 258680 287296 258732
rect 560300 258680 560352 258732
rect 287336 257320 287388 257372
rect 563152 257320 563204 257372
rect 277032 256751 277084 256760
rect 277032 256717 277041 256751
rect 277041 256717 277075 256751
rect 277075 256717 277084 256751
rect 277032 256708 277084 256717
rect 276940 256683 276992 256692
rect 276940 256649 276949 256683
rect 276949 256649 276983 256683
rect 276983 256649 276992 256683
rect 276940 256640 276992 256649
rect 291108 255960 291160 256012
rect 471244 255960 471296 256012
rect 255780 255255 255832 255264
rect 255780 255221 255789 255255
rect 255789 255221 255823 255255
rect 255823 255221 255832 255255
rect 255780 255212 255832 255221
rect 259920 255255 259972 255264
rect 259920 255221 259929 255255
rect 259929 255221 259963 255255
rect 259963 255221 259972 255255
rect 259920 255212 259972 255221
rect 277216 255255 277268 255264
rect 277216 255221 277225 255255
rect 277225 255221 277259 255255
rect 277259 255221 277268 255255
rect 277216 255212 277268 255221
rect 237012 253852 237064 253904
rect 237196 253852 237248 253904
rect 250720 253827 250772 253836
rect 250720 253793 250729 253827
rect 250729 253793 250763 253827
rect 250763 253793 250772 253827
rect 250720 253784 250772 253793
rect 3424 252492 3476 252544
rect 225788 252492 225840 252544
rect 301596 252492 301648 252544
rect 579804 252492 579856 252544
rect 252284 251268 252336 251320
rect 229652 251200 229704 251252
rect 254860 251243 254912 251252
rect 254860 251209 254869 251243
rect 254869 251209 254903 251243
rect 254903 251209 254912 251243
rect 254860 251200 254912 251209
rect 273720 251200 273772 251252
rect 237196 251132 237248 251184
rect 273812 251064 273864 251116
rect 252192 249815 252244 249824
rect 252192 249781 252201 249815
rect 252201 249781 252235 249815
rect 252235 249781 252244 249815
rect 252192 249772 252244 249781
rect 254860 249815 254912 249824
rect 254860 249781 254869 249815
rect 254869 249781 254903 249815
rect 254903 249781 254912 249815
rect 254860 249772 254912 249781
rect 256976 249772 257028 249824
rect 257252 249772 257304 249824
rect 274180 249772 274232 249824
rect 274272 249772 274324 249824
rect 276940 249747 276992 249756
rect 276940 249713 276949 249747
rect 276949 249713 276983 249747
rect 276983 249713 276992 249747
rect 276940 249704 276992 249713
rect 260656 246984 260708 247036
rect 262496 246984 262548 247036
rect 262680 246984 262732 247036
rect 274272 246984 274324 247036
rect 277216 247027 277268 247036
rect 277216 246993 277225 247027
rect 277225 246993 277259 247027
rect 277259 246993 277268 247027
rect 277216 246984 277268 246993
rect 259920 245667 259972 245676
rect 259920 245633 259929 245667
rect 259929 245633 259963 245667
rect 259963 245633 259972 245667
rect 259920 245624 259972 245633
rect 271512 245624 271564 245676
rect 271788 245624 271840 245676
rect 233700 244264 233752 244316
rect 233884 244264 233936 244316
rect 252100 244196 252152 244248
rect 252284 244196 252336 244248
rect 235172 244035 235224 244044
rect 235172 244001 235181 244035
rect 235181 244001 235215 244035
rect 235215 244001 235224 244035
rect 235172 243992 235224 244001
rect 237104 241519 237156 241528
rect 237104 241485 237113 241519
rect 237113 241485 237147 241519
rect 237147 241485 237156 241519
rect 237104 241476 237156 241485
rect 273720 241476 273772 241528
rect 273812 241476 273864 241528
rect 277216 241519 277268 241528
rect 277216 241485 277225 241519
rect 277225 241485 277259 241519
rect 277259 241485 277268 241519
rect 277216 241476 277268 241485
rect 238944 241451 238996 241460
rect 238944 241417 238953 241451
rect 238953 241417 238987 241451
rect 238987 241417 238996 241451
rect 238944 241408 238996 241417
rect 256516 238688 256568 238740
rect 256608 238688 256660 238740
rect 255872 237396 255924 237448
rect 260564 237439 260616 237448
rect 260564 237405 260573 237439
rect 260573 237405 260607 237439
rect 260607 237405 260616 237439
rect 260564 237396 260616 237405
rect 271604 237396 271656 237448
rect 271788 237396 271840 237448
rect 274180 237439 274232 237448
rect 274180 237405 274189 237439
rect 274189 237405 274223 237439
rect 274223 237405 274232 237439
rect 274180 237396 274232 237405
rect 277216 237439 277268 237448
rect 277216 237405 277225 237439
rect 277225 237405 277259 237439
rect 277259 237405 277268 237439
rect 277216 237396 277268 237405
rect 264244 237371 264296 237380
rect 264244 237337 264253 237371
rect 264253 237337 264287 237371
rect 264287 237337 264296 237371
rect 264244 237328 264296 237337
rect 262680 234676 262732 234728
rect 250720 234608 250772 234660
rect 243360 234540 243412 234592
rect 243544 234540 243596 234592
rect 250720 234472 250772 234524
rect 229652 231820 229704 231872
rect 229836 231820 229888 231872
rect 234988 231820 235040 231872
rect 235264 231820 235316 231872
rect 238944 231863 238996 231872
rect 238944 231829 238953 231863
rect 238953 231829 238987 231863
rect 238987 231829 238996 231863
rect 238944 231820 238996 231829
rect 235540 230460 235592 230512
rect 235724 230460 235776 230512
rect 262496 229075 262548 229084
rect 262496 229041 262505 229075
rect 262505 229041 262539 229075
rect 262539 229041 262548 229075
rect 262496 229032 262548 229041
rect 274180 229032 274232 229084
rect 276940 229032 276992 229084
rect 277032 229032 277084 229084
rect 274364 228964 274416 229016
rect 328460 228080 328512 228132
rect 418068 227944 418120 227996
rect 424968 227944 425020 227996
rect 328460 227876 328512 227928
rect 495348 227876 495400 227928
rect 497004 227876 497056 227928
rect 553308 227876 553360 227928
rect 554596 227876 554648 227928
rect 437388 227808 437440 227860
rect 444288 227808 444340 227860
rect 476028 227808 476080 227860
rect 482928 227808 482980 227860
rect 514668 227808 514720 227860
rect 521568 227808 521620 227860
rect 278688 227740 278740 227792
rect 289728 227740 289780 227792
rect 309140 227740 309192 227792
rect 312636 227740 312688 227792
rect 533988 227740 534040 227792
rect 540888 227740 540940 227792
rect 233700 224952 233752 225004
rect 233884 224952 233936 225004
rect 3148 223524 3200 223576
rect 207664 223524 207716 223576
rect 235172 222164 235224 222216
rect 235356 222164 235408 222216
rect 254768 222164 254820 222216
rect 254860 222096 254912 222148
rect 256608 220872 256660 220924
rect 256424 220736 256476 220788
rect 255872 219512 255924 219564
rect 256056 219512 256108 219564
rect 260748 219444 260800 219496
rect 264244 219487 264296 219496
rect 264244 219453 264253 219487
rect 264253 219453 264287 219487
rect 264287 219453 264296 219487
rect 264244 219444 264296 219453
rect 260656 219376 260708 219428
rect 255872 217991 255924 218000
rect 255872 217957 255881 217991
rect 255881 217957 255915 217991
rect 255915 217957 255924 217991
rect 255872 217948 255924 217957
rect 260656 217948 260708 218000
rect 260932 217948 260984 218000
rect 262680 217991 262732 218000
rect 262680 217957 262689 217991
rect 262689 217957 262723 217991
rect 262723 217957 262732 217991
rect 262680 217948 262732 217957
rect 264244 217991 264296 218000
rect 264244 217957 264253 217991
rect 264253 217957 264287 217991
rect 264287 217957 264296 217991
rect 264244 217948 264296 217957
rect 413284 217948 413336 218000
rect 580172 217948 580224 218000
rect 243544 215364 243596 215416
rect 243360 215296 243412 215348
rect 274180 213936 274232 213988
rect 274364 213936 274416 213988
rect 277584 212712 277636 212764
rect 277952 212712 278004 212764
rect 229652 212508 229704 212560
rect 229836 212508 229888 212560
rect 237012 212508 237064 212560
rect 245016 212508 245068 212560
rect 245200 212508 245252 212560
rect 237012 212372 237064 212424
rect 277124 209720 277176 209772
rect 277216 209720 277268 209772
rect 255872 208403 255924 208412
rect 255872 208369 255881 208403
rect 255881 208369 255915 208403
rect 255915 208369 255924 208403
rect 255872 208360 255924 208369
rect 264428 208360 264480 208412
rect 3424 208292 3476 208344
rect 222936 208292 222988 208344
rect 252192 208335 252244 208344
rect 252192 208301 252201 208335
rect 252201 208301 252235 208335
rect 252235 208301 252244 208335
rect 252192 208292 252244 208301
rect 277124 208292 277176 208344
rect 277216 208292 277268 208344
rect 233700 205640 233752 205692
rect 233884 205640 233936 205692
rect 259828 205640 259880 205692
rect 259920 205572 259972 205624
rect 298836 205572 298888 205624
rect 579804 205572 579856 205624
rect 235540 202852 235592 202904
rect 235632 202852 235684 202904
rect 254860 202852 254912 202904
rect 254952 202852 255004 202904
rect 273904 202852 273956 202904
rect 273996 202852 274048 202904
rect 235172 202784 235224 202836
rect 235264 202784 235316 202836
rect 237104 202784 237156 202836
rect 237196 202784 237248 202836
rect 238944 202827 238996 202836
rect 238944 202793 238953 202827
rect 238953 202793 238987 202827
rect 238987 202793 238996 202827
rect 238944 202784 238996 202793
rect 235264 201424 235316 201476
rect 234988 201356 235040 201408
rect 268844 200064 268896 200116
rect 269028 200064 269080 200116
rect 274180 200064 274232 200116
rect 274272 199996 274324 200048
rect 252284 198704 252336 198756
rect 262680 198747 262732 198756
rect 262680 198713 262689 198747
rect 262689 198713 262723 198747
rect 262723 198713 262732 198747
rect 262680 198704 262732 198713
rect 264244 198704 264296 198756
rect 264428 198704 264480 198756
rect 255872 198636 255924 198688
rect 260656 198636 260708 198688
rect 260748 198636 260800 198688
rect 260656 197276 260708 197328
rect 277124 197319 277176 197328
rect 277124 197285 277133 197319
rect 277133 197285 277167 197319
rect 277167 197285 277176 197319
rect 277124 197276 277176 197285
rect 271604 195959 271656 195968
rect 271604 195925 271613 195959
rect 271613 195925 271647 195959
rect 271647 195925 271656 195959
rect 271604 195916 271656 195925
rect 277768 195916 277820 195968
rect 277952 195848 278004 195900
rect 229652 193196 229704 193248
rect 229836 193196 229888 193248
rect 235540 193196 235592 193248
rect 235632 193196 235684 193248
rect 245016 193196 245068 193248
rect 245200 193196 245252 193248
rect 238944 191879 238996 191888
rect 238944 191845 238953 191879
rect 238953 191845 238987 191879
rect 238987 191845 238996 191879
rect 238944 191836 238996 191845
rect 255780 191335 255832 191344
rect 255780 191301 255789 191335
rect 255789 191301 255823 191335
rect 255823 191301 255832 191335
rect 255780 191292 255832 191301
rect 252100 189048 252152 189100
rect 252284 189048 252336 189100
rect 254768 189023 254820 189032
rect 254768 188989 254777 189023
rect 254777 188989 254811 189023
rect 254811 188989 254820 189023
rect 254768 188980 254820 188989
rect 255780 189023 255832 189032
rect 255780 188989 255789 189023
rect 255789 188989 255823 189023
rect 255823 188989 255832 189023
rect 255780 188980 255832 188989
rect 262680 189023 262732 189032
rect 262680 188989 262689 189023
rect 262689 188989 262723 189023
rect 262723 188989 262732 189023
rect 262680 188980 262732 188989
rect 264244 189023 264296 189032
rect 264244 188989 264253 189023
rect 264253 188989 264287 189023
rect 264287 188989 264296 189023
rect 264244 188980 264296 188989
rect 260656 187731 260708 187740
rect 260656 187697 260665 187731
rect 260665 187697 260699 187731
rect 260699 187697 260708 187731
rect 260656 187688 260708 187697
rect 277124 187731 277176 187740
rect 277124 187697 277133 187731
rect 277133 187697 277167 187731
rect 277167 187697 277176 187731
rect 277124 187688 277176 187697
rect 233700 186328 233752 186380
rect 233884 186328 233936 186380
rect 271696 186328 271748 186380
rect 252100 186303 252152 186312
rect 252100 186269 252109 186303
rect 252109 186269 252143 186303
rect 252143 186269 252152 186303
rect 252100 186260 252152 186269
rect 273904 184220 273956 184272
rect 255872 184152 255924 184204
rect 234988 183540 235040 183592
rect 235172 183540 235224 183592
rect 273720 183540 273772 183592
rect 273812 183540 273864 183592
rect 276940 183540 276992 183592
rect 277032 183540 277084 183592
rect 277124 183540 277176 183592
rect 237104 183472 237156 183524
rect 237196 183472 237248 183524
rect 277216 183404 277268 183456
rect 284852 182792 284904 182844
rect 538220 182792 538272 182844
rect 308404 182112 308456 182164
rect 580172 182112 580224 182164
rect 3240 180752 3292 180804
rect 204904 180752 204956 180804
rect 245016 180795 245068 180804
rect 245016 180761 245025 180795
rect 245025 180761 245059 180795
rect 245059 180761 245068 180795
rect 245016 180752 245068 180761
rect 273812 180795 273864 180804
rect 273812 180761 273821 180795
rect 273821 180761 273855 180795
rect 273855 180761 273864 180795
rect 273812 180752 273864 180761
rect 281448 180072 281500 180124
rect 499580 180072 499632 180124
rect 254952 179392 255004 179444
rect 260656 179435 260708 179444
rect 260656 179401 260665 179435
rect 260665 179401 260699 179435
rect 260699 179401 260708 179435
rect 260656 179392 260708 179401
rect 262680 179435 262732 179444
rect 262680 179401 262689 179435
rect 262689 179401 262723 179435
rect 262723 179401 262732 179435
rect 262680 179392 262732 179401
rect 264244 179435 264296 179444
rect 264244 179401 264253 179435
rect 264253 179401 264287 179435
rect 264287 179401 264296 179435
rect 264244 179392 264296 179401
rect 260656 178075 260708 178084
rect 260656 178041 260665 178075
rect 260665 178041 260699 178075
rect 260699 178041 260708 178075
rect 260656 178032 260708 178041
rect 271604 178032 271656 178084
rect 271696 178032 271748 178084
rect 268844 178007 268896 178016
rect 268844 177973 268853 178007
rect 268853 177973 268887 178007
rect 268887 177973 268896 178007
rect 268844 177964 268896 177973
rect 277216 177964 277268 178016
rect 277400 177964 277452 178016
rect 252192 176672 252244 176724
rect 252192 173995 252244 174004
rect 252192 173961 252201 173995
rect 252201 173961 252235 173995
rect 252235 173961 252244 173995
rect 252192 173952 252244 173961
rect 229652 173884 229704 173936
rect 229836 173884 229888 173936
rect 234988 173884 235040 173936
rect 235264 173884 235316 173936
rect 235448 173884 235500 173936
rect 235540 173884 235592 173936
rect 234988 172456 235040 172508
rect 235264 172456 235316 172508
rect 245292 171096 245344 171148
rect 273812 171028 273864 171080
rect 273904 171028 273956 171080
rect 493324 171028 493376 171080
rect 580172 171028 580224 171080
rect 259920 169736 259972 169788
rect 259736 169668 259788 169720
rect 262680 169711 262732 169720
rect 262680 169677 262689 169711
rect 262689 169677 262723 169711
rect 262723 169677 262732 169711
rect 262680 169668 262732 169677
rect 264244 169711 264296 169720
rect 264244 169677 264253 169711
rect 264253 169677 264287 169711
rect 264287 169677 264296 169711
rect 264244 169668 264296 169677
rect 257252 169056 257304 169108
rect 257436 169056 257488 169108
rect 268936 168376 268988 168428
rect 252192 168351 252244 168360
rect 252192 168317 252201 168351
rect 252201 168317 252235 168351
rect 252235 168317 252244 168351
rect 252192 168308 252244 168317
rect 254952 168308 255004 168360
rect 233700 167016 233752 167068
rect 233884 167016 233936 167068
rect 3516 165520 3568 165572
rect 218704 165520 218756 165572
rect 219256 164840 219308 164892
rect 252192 164840 252244 164892
rect 273628 164228 273680 164280
rect 229560 164160 229612 164212
rect 229836 164160 229888 164212
rect 273720 164092 273772 164144
rect 238760 162800 238812 162852
rect 238944 162800 238996 162852
rect 235172 162775 235224 162784
rect 235172 162741 235181 162775
rect 235181 162741 235215 162775
rect 235215 162741 235224 162775
rect 235172 162732 235224 162741
rect 268844 161440 268896 161492
rect 268936 161440 268988 161492
rect 245292 161372 245344 161424
rect 259736 160080 259788 160132
rect 259920 160080 259972 160132
rect 262680 160123 262732 160132
rect 262680 160089 262689 160123
rect 262689 160089 262723 160123
rect 262723 160089 262732 160123
rect 262680 160080 262732 160089
rect 264244 160123 264296 160132
rect 264244 160089 264253 160123
rect 264253 160089 264287 160123
rect 264287 160089 264296 160123
rect 264244 160080 264296 160089
rect 276848 160080 276900 160132
rect 277032 160080 277084 160132
rect 277124 160080 277176 160132
rect 277400 160080 277452 160132
rect 268844 160055 268896 160064
rect 268844 160021 268853 160055
rect 268853 160021 268887 160055
rect 268887 160021 268896 160055
rect 268844 160012 268896 160021
rect 271604 160055 271656 160064
rect 271604 160021 271613 160055
rect 271613 160021 271647 160055
rect 271647 160021 271656 160055
rect 271604 160012 271656 160021
rect 274180 160012 274232 160064
rect 274180 159876 274232 159928
rect 254860 158763 254912 158772
rect 254860 158729 254869 158763
rect 254869 158729 254903 158763
rect 254903 158729 254912 158763
rect 254860 158720 254912 158729
rect 260564 158695 260616 158704
rect 260564 158661 260573 158695
rect 260573 158661 260607 158695
rect 260607 158661 260616 158695
rect 260564 158652 260616 158661
rect 277124 158652 277176 158704
rect 277216 158652 277268 158704
rect 297456 158652 297508 158704
rect 579804 158652 579856 158704
rect 235172 157403 235224 157412
rect 235172 157369 235181 157403
rect 235181 157369 235215 157403
rect 235215 157369 235224 157403
rect 235172 157360 235224 157369
rect 255872 157403 255924 157412
rect 255872 157369 255881 157403
rect 255881 157369 255915 157403
rect 255915 157369 255924 157403
rect 255872 157360 255924 157369
rect 237012 157292 237064 157344
rect 237196 157292 237248 157344
rect 257252 154640 257304 154692
rect 255872 154547 255924 154556
rect 255872 154513 255881 154547
rect 255881 154513 255915 154547
rect 255915 154513 255924 154547
rect 255872 154504 255924 154513
rect 257160 154504 257212 154556
rect 245016 151827 245068 151836
rect 245016 151793 245025 151827
rect 245025 151793 245059 151827
rect 245059 151793 245068 151827
rect 245016 151784 245068 151793
rect 3148 151716 3200 151768
rect 227076 151716 227128 151768
rect 254860 150424 254912 150476
rect 255044 150424 255096 150476
rect 268936 150424 268988 150476
rect 271696 149132 271748 149184
rect 260656 149064 260708 149116
rect 271604 149039 271656 149048
rect 271604 149005 271613 149039
rect 271613 149005 271647 149039
rect 271647 149005 271656 149039
rect 271604 148996 271656 149005
rect 277124 149039 277176 149048
rect 277124 149005 277133 149039
rect 277133 149005 277167 149039
rect 277167 149005 277176 149039
rect 277124 148996 277176 149005
rect 259828 147636 259880 147688
rect 259920 147568 259972 147620
rect 237104 144916 237156 144968
rect 237196 144916 237248 144968
rect 235172 144848 235224 144900
rect 235540 144891 235592 144900
rect 235540 144857 235549 144891
rect 235549 144857 235583 144891
rect 235583 144857 235592 144891
rect 235540 144848 235592 144857
rect 235264 144780 235316 144832
rect 235264 143531 235316 143540
rect 235264 143497 235273 143531
rect 235273 143497 235307 143531
rect 235307 143497 235316 143531
rect 235264 143488 235316 143497
rect 268844 142128 268896 142180
rect 268936 142128 268988 142180
rect 273628 142128 273680 142180
rect 273720 142128 273772 142180
rect 273812 142128 273864 142180
rect 273904 142128 273956 142180
rect 250628 140700 250680 140752
rect 254952 140700 255004 140752
rect 255044 140700 255096 140752
rect 260564 140743 260616 140752
rect 260564 140709 260573 140743
rect 260573 140709 260607 140743
rect 260607 140709 260616 140743
rect 260564 140700 260616 140709
rect 262680 140743 262732 140752
rect 262680 140709 262689 140743
rect 262689 140709 262723 140743
rect 262723 140709 262732 140743
rect 262680 140700 262732 140709
rect 264244 140743 264296 140752
rect 264244 140709 264253 140743
rect 264253 140709 264287 140743
rect 264287 140709 264296 140743
rect 264244 140700 264296 140709
rect 271604 139519 271656 139528
rect 271604 139485 271613 139519
rect 271613 139485 271647 139519
rect 271647 139485 271656 139519
rect 271604 139476 271656 139485
rect 277216 139408 277268 139460
rect 271604 139340 271656 139392
rect 245200 138703 245252 138712
rect 245200 138669 245209 138703
rect 245209 138669 245243 138703
rect 245243 138669 245252 138703
rect 245200 138660 245252 138669
rect 229560 137980 229612 138032
rect 237104 137980 237156 138032
rect 229468 137912 229520 137964
rect 237196 137912 237248 137964
rect 3240 136552 3292 136604
rect 17224 136552 17276 136604
rect 235540 135303 235592 135312
rect 235540 135269 235549 135303
rect 235549 135269 235583 135303
rect 235583 135269 235592 135303
rect 235540 135260 235592 135269
rect 255872 135192 255924 135244
rect 256056 135192 256108 135244
rect 319444 135192 319496 135244
rect 580172 135192 580224 135244
rect 245384 135124 245436 135176
rect 235264 133943 235316 133952
rect 235264 133909 235273 133943
rect 235273 133909 235307 133943
rect 235307 133909 235316 133943
rect 235264 133900 235316 133909
rect 273812 133832 273864 133884
rect 273996 133832 274048 133884
rect 276940 132472 276992 132524
rect 277032 132472 277084 132524
rect 262680 131155 262732 131164
rect 262680 131121 262689 131155
rect 262689 131121 262723 131155
rect 262723 131121 262732 131155
rect 262680 131112 262732 131121
rect 264244 131155 264296 131164
rect 264244 131121 264253 131155
rect 264253 131121 264287 131155
rect 264287 131121 264296 131155
rect 264244 131112 264296 131121
rect 274180 131044 274232 131096
rect 257160 130364 257212 130416
rect 257252 130296 257304 130348
rect 260564 129795 260616 129804
rect 260564 129761 260573 129795
rect 260573 129761 260607 129795
rect 260607 129761 260616 129795
rect 260564 129752 260616 129761
rect 271512 129795 271564 129804
rect 271512 129761 271521 129795
rect 271521 129761 271555 129795
rect 271555 129761 271564 129795
rect 271512 129752 271564 129761
rect 233700 128324 233752 128376
rect 233884 128324 233936 128376
rect 259828 128324 259880 128376
rect 250536 128299 250588 128308
rect 250536 128265 250545 128299
rect 250545 128265 250579 128299
rect 250579 128265 250588 128299
rect 250536 128256 250588 128265
rect 259920 128256 259972 128308
rect 254952 125604 255004 125656
rect 235540 125579 235592 125588
rect 235540 125545 235549 125579
rect 235549 125545 235583 125579
rect 235583 125545 235592 125579
rect 235540 125536 235592 125545
rect 254860 125536 254912 125588
rect 245108 125468 245160 125520
rect 245384 125468 245436 125520
rect 250628 125468 250680 125520
rect 250720 125468 250772 125520
rect 235264 124219 235316 124228
rect 235264 124185 235273 124219
rect 235273 124185 235307 124219
rect 235307 124185 235316 124219
rect 235264 124176 235316 124185
rect 245108 124151 245160 124160
rect 245108 124117 245117 124151
rect 245117 124117 245151 124151
rect 245151 124117 245160 124151
rect 245108 124108 245160 124117
rect 254860 124108 254912 124160
rect 255136 124108 255188 124160
rect 255872 124108 255924 124160
rect 256056 124108 256108 124160
rect 257252 124151 257304 124160
rect 257252 124117 257261 124151
rect 257261 124117 257295 124151
rect 257295 124117 257304 124151
rect 257252 124108 257304 124117
rect 312544 124108 312596 124160
rect 580172 124108 580224 124160
rect 235264 122859 235316 122868
rect 235264 122825 235273 122859
rect 235273 122825 235307 122859
rect 235307 122825 235316 122859
rect 235264 122816 235316 122825
rect 3424 122748 3476 122800
rect 215944 122748 215996 122800
rect 255136 122748 255188 122800
rect 274088 121499 274140 121508
rect 274088 121465 274097 121499
rect 274097 121465 274131 121499
rect 274131 121465 274140 121499
rect 274088 121456 274140 121465
rect 268844 121431 268896 121440
rect 268844 121397 268853 121431
rect 268853 121397 268887 121431
rect 268887 121397 268896 121431
rect 268844 121388 268896 121397
rect 273904 120071 273956 120080
rect 273904 120037 273913 120071
rect 273913 120037 273947 120071
rect 273947 120037 273956 120071
rect 273904 120028 273956 120037
rect 229560 118668 229612 118720
rect 237104 118668 237156 118720
rect 229468 118600 229520 118652
rect 237196 118600 237248 118652
rect 235540 115991 235592 116000
rect 235540 115957 235549 115991
rect 235549 115957 235583 115991
rect 235583 115957 235592 115991
rect 235540 115948 235592 115957
rect 277216 115991 277268 116000
rect 277216 115957 277225 115991
rect 277225 115957 277259 115991
rect 277259 115957 277268 115991
rect 277216 115948 277268 115957
rect 259828 115880 259880 115932
rect 259920 115880 259972 115932
rect 245108 114563 245160 114572
rect 245108 114529 245117 114563
rect 245117 114529 245151 114563
rect 245151 114529 245160 114563
rect 245108 114520 245160 114529
rect 257252 114563 257304 114572
rect 257252 114529 257261 114563
rect 257261 114529 257295 114563
rect 257295 114529 257304 114563
rect 257252 114520 257304 114529
rect 235264 114452 235316 114504
rect 235356 114452 235408 114504
rect 255044 113203 255096 113212
rect 255044 113169 255053 113203
rect 255053 113169 255087 113203
rect 255087 113169 255096 113203
rect 255044 113160 255096 113169
rect 268844 111911 268896 111920
rect 268844 111877 268853 111911
rect 268853 111877 268887 111911
rect 268887 111877 268896 111911
rect 268844 111868 268896 111877
rect 274088 111800 274140 111852
rect 274272 111800 274324 111852
rect 250720 111732 250772 111784
rect 260472 111732 260524 111784
rect 260564 111732 260616 111784
rect 262680 111775 262732 111784
rect 262680 111741 262689 111775
rect 262689 111741 262723 111775
rect 262723 111741 262732 111775
rect 262680 111732 262732 111741
rect 268844 111775 268896 111784
rect 268844 111741 268853 111775
rect 268853 111741 268887 111775
rect 268887 111741 268896 111775
rect 268844 111732 268896 111741
rect 276940 111775 276992 111784
rect 276940 111741 276949 111775
rect 276949 111741 276983 111775
rect 276983 111741 276992 111775
rect 276940 111732 276992 111741
rect 291936 111732 291988 111784
rect 579804 111732 579856 111784
rect 273996 110440 274048 110492
rect 260472 110415 260524 110424
rect 260472 110381 260481 110415
rect 260481 110381 260515 110415
rect 260515 110381 260524 110415
rect 260472 110372 260524 110381
rect 233700 109012 233752 109064
rect 233884 109012 233936 109064
rect 245108 109012 245160 109064
rect 245200 108944 245252 108996
rect 233792 104839 233844 104848
rect 233792 104805 233801 104839
rect 233801 104805 233835 104839
rect 233835 104805 233844 104839
rect 233792 104796 233844 104805
rect 254860 104839 254912 104848
rect 254860 104805 254869 104839
rect 254869 104805 254903 104839
rect 254903 104805 254912 104839
rect 254860 104796 254912 104805
rect 256516 104839 256568 104848
rect 256516 104805 256525 104839
rect 256525 104805 256559 104839
rect 256559 104805 256568 104839
rect 256516 104796 256568 104805
rect 262680 102255 262732 102264
rect 262680 102221 262689 102255
rect 262689 102221 262723 102255
rect 262723 102221 262732 102255
rect 262680 102212 262732 102221
rect 277216 102255 277268 102264
rect 277216 102221 277225 102255
rect 277225 102221 277259 102255
rect 277259 102221 277268 102255
rect 277216 102212 277268 102221
rect 250628 102187 250680 102196
rect 250628 102153 250637 102187
rect 250637 102153 250671 102187
rect 250671 102153 250680 102187
rect 250628 102144 250680 102153
rect 277032 102144 277084 102196
rect 260564 102076 260616 102128
rect 262680 102119 262732 102128
rect 262680 102085 262689 102119
rect 262689 102085 262723 102119
rect 262723 102085 262732 102119
rect 262680 102076 262732 102085
rect 264244 102119 264296 102128
rect 264244 102085 264253 102119
rect 264253 102085 264287 102119
rect 264287 102085 264296 102119
rect 264244 102076 264296 102085
rect 268844 100759 268896 100768
rect 268844 100725 268853 100759
rect 268853 100725 268887 100759
rect 268887 100725 268896 100759
rect 268844 100716 268896 100725
rect 235356 99492 235408 99544
rect 229560 99356 229612 99408
rect 235172 99356 235224 99408
rect 229468 99288 229520 99340
rect 243360 99288 243412 99340
rect 243544 99288 243596 99340
rect 274180 99288 274232 99340
rect 255872 98676 255924 98728
rect 256056 98676 256108 98728
rect 233976 95208 234028 95260
rect 255044 95208 255096 95260
rect 256700 95208 256752 95260
rect 257252 95251 257304 95260
rect 257252 95217 257261 95251
rect 257261 95217 257295 95251
rect 257295 95217 257304 95251
rect 257252 95208 257304 95217
rect 259920 95251 259972 95260
rect 259920 95217 259929 95251
rect 259929 95217 259963 95251
rect 259963 95217 259972 95251
rect 259920 95208 259972 95217
rect 257252 93891 257304 93900
rect 257252 93857 257261 93891
rect 257261 93857 257295 93891
rect 257295 93857 257304 93891
rect 257252 93848 257304 93857
rect 3424 93780 3476 93832
rect 203524 93780 203576 93832
rect 259920 92531 259972 92540
rect 259920 92497 259929 92531
rect 259929 92497 259963 92531
rect 259963 92497 259972 92531
rect 259920 92488 259972 92497
rect 264244 92531 264296 92540
rect 264244 92497 264253 92531
rect 264253 92497 264287 92531
rect 264287 92497 264296 92531
rect 264244 92488 264296 92497
rect 268844 92463 268896 92472
rect 268844 92429 268853 92463
rect 268853 92429 268887 92463
rect 268887 92429 268896 92463
rect 268844 92420 268896 92429
rect 273812 92420 273864 92472
rect 273996 92420 274048 92472
rect 262588 91060 262640 91112
rect 276940 91060 276992 91112
rect 277124 91060 277176 91112
rect 305644 88272 305696 88324
rect 580172 88272 580224 88324
rect 268936 87048 268988 87100
rect 235172 86912 235224 86964
rect 235264 86912 235316 86964
rect 235264 85527 235316 85536
rect 235264 85493 235273 85527
rect 235273 85493 235307 85527
rect 235307 85493 235316 85527
rect 235264 85484 235316 85493
rect 237196 85484 237248 85536
rect 245200 85527 245252 85536
rect 245200 85493 245209 85527
rect 245209 85493 245243 85527
rect 245243 85493 245252 85527
rect 245200 85484 245252 85493
rect 277124 84167 277176 84176
rect 277124 84133 277133 84167
rect 277133 84133 277167 84167
rect 277167 84133 277176 84167
rect 277124 84124 277176 84133
rect 274180 82832 274232 82884
rect 250628 82764 250680 82816
rect 256424 82764 256476 82816
rect 256608 82764 256660 82816
rect 264244 82807 264296 82816
rect 264244 82773 264253 82807
rect 264253 82773 264287 82807
rect 264287 82773 264296 82807
rect 264244 82764 264296 82773
rect 254768 81404 254820 81456
rect 254952 81404 255004 81456
rect 255780 81404 255832 81456
rect 256056 81404 256108 81456
rect 259828 81404 259880 81456
rect 259920 81404 259972 81456
rect 262588 81404 262640 81456
rect 262496 81336 262548 81388
rect 229560 80044 229612 80096
rect 3424 79976 3476 80028
rect 214564 79976 214616 80028
rect 229652 79976 229704 80028
rect 233792 77256 233844 77308
rect 233884 77256 233936 77308
rect 235448 77256 235500 77308
rect 235540 77256 235592 77308
rect 229652 77188 229704 77240
rect 250904 77231 250956 77240
rect 250904 77197 250913 77231
rect 250913 77197 250947 77231
rect 250947 77197 250956 77231
rect 250904 77188 250956 77197
rect 251088 77231 251140 77240
rect 251088 77197 251097 77231
rect 251097 77197 251131 77231
rect 251131 77197 251140 77231
rect 251088 77188 251140 77197
rect 250996 77163 251048 77172
rect 250996 77129 251005 77163
rect 251005 77129 251039 77163
rect 251039 77129 251048 77163
rect 250996 77120 251048 77129
rect 268936 76619 268988 76628
rect 268936 76585 268945 76619
rect 268945 76585 268979 76619
rect 268979 76585 268988 76619
rect 268936 76576 268988 76585
rect 274088 76576 274140 76628
rect 274180 76576 274232 76628
rect 274456 76576 274508 76628
rect 328460 76304 328512 76356
rect 328460 76100 328512 76152
rect 553308 76100 553360 76152
rect 554596 76100 554648 76152
rect 437388 76032 437440 76084
rect 444288 76032 444340 76084
rect 502248 76032 502300 76084
rect 510528 76032 510580 76084
rect 533988 76032 534040 76084
rect 540888 76032 540940 76084
rect 237012 76007 237064 76016
rect 237012 75973 237021 76007
rect 237021 75973 237055 76007
rect 237055 75973 237064 76007
rect 237012 75964 237064 75973
rect 309140 75964 309192 76016
rect 313924 75964 313976 76016
rect 235264 75939 235316 75948
rect 235264 75905 235273 75939
rect 235273 75905 235307 75939
rect 235307 75905 235316 75939
rect 235264 75896 235316 75905
rect 245200 75939 245252 75948
rect 245200 75905 245209 75939
rect 245209 75905 245243 75939
rect 245243 75905 245252 75939
rect 245200 75896 245252 75905
rect 237012 75828 237064 75880
rect 267464 75871 267516 75880
rect 267464 75837 267473 75871
rect 267473 75837 267507 75871
rect 267507 75837 267516 75871
rect 267464 75828 267516 75837
rect 264336 75760 264388 75812
rect 273628 74536 273680 74588
rect 273720 74536 273772 74588
rect 277124 74579 277176 74588
rect 277124 74545 277133 74579
rect 277133 74545 277167 74579
rect 277167 74545 277176 74579
rect 277124 74536 277176 74545
rect 256424 73151 256476 73160
rect 256424 73117 256433 73151
rect 256433 73117 256467 73151
rect 256467 73117 256476 73151
rect 256424 73108 256476 73117
rect 259828 73108 259880 73160
rect 260104 73108 260156 73160
rect 255780 73083 255832 73092
rect 255780 73049 255789 73083
rect 255789 73049 255823 73083
rect 255823 73049 255832 73083
rect 255780 73040 255832 73049
rect 277124 73083 277176 73092
rect 277124 73049 277133 73083
rect 277133 73049 277167 73083
rect 277167 73049 277176 73083
rect 277124 73040 277176 73049
rect 250904 72471 250956 72480
rect 250904 72437 250913 72471
rect 250913 72437 250947 72471
rect 250947 72437 250956 72471
rect 250904 72428 250956 72437
rect 269028 71748 269080 71800
rect 250996 71723 251048 71732
rect 250996 71689 251005 71723
rect 251005 71689 251039 71723
rect 251039 71689 251048 71723
rect 250996 71680 251048 71689
rect 235264 70456 235316 70508
rect 245200 70456 245252 70508
rect 243360 70388 243412 70440
rect 243544 70388 243596 70440
rect 251088 70431 251140 70440
rect 251088 70397 251097 70431
rect 251097 70397 251131 70431
rect 251131 70397 251140 70431
rect 251088 70388 251140 70397
rect 235172 70320 235224 70372
rect 268844 68484 268896 68536
rect 269028 68484 269080 68536
rect 257252 68348 257304 68400
rect 250444 68280 250496 68332
rect 229560 67643 229612 67652
rect 229560 67609 229569 67643
rect 229569 67609 229603 67643
rect 229603 67609 229612 67643
rect 229560 67600 229612 67609
rect 233792 67600 233844 67652
rect 233884 67600 233936 67652
rect 245108 67643 245160 67652
rect 245108 67609 245117 67643
rect 245117 67609 245151 67643
rect 245151 67609 245160 67643
rect 245108 67600 245160 67609
rect 235540 67575 235592 67584
rect 235540 67541 235549 67575
rect 235549 67541 235583 67575
rect 235583 67541 235592 67575
rect 235540 67532 235592 67541
rect 273628 66308 273680 66360
rect 264244 66240 264296 66292
rect 264336 66240 264388 66292
rect 267464 66283 267516 66292
rect 267464 66249 267473 66283
rect 267473 66249 267507 66283
rect 267507 66249 267516 66283
rect 267464 66240 267516 66249
rect 271144 66172 271196 66224
rect 271236 66172 271288 66224
rect 273628 66172 273680 66224
rect 3332 64812 3384 64864
rect 198004 64812 198056 64864
rect 294604 64812 294656 64864
rect 579804 64812 579856 64864
rect 255872 63520 255924 63572
rect 256608 63520 256660 63572
rect 257160 63563 257212 63572
rect 257160 63529 257169 63563
rect 257169 63529 257203 63563
rect 257203 63529 257212 63563
rect 257160 63520 257212 63529
rect 260012 63520 260064 63572
rect 273904 63563 273956 63572
rect 273904 63529 273913 63563
rect 273913 63529 273947 63563
rect 273947 63529 273956 63563
rect 273904 63520 273956 63529
rect 274364 63520 274416 63572
rect 277216 63520 277268 63572
rect 260012 63384 260064 63436
rect 274272 63384 274324 63436
rect 259736 62092 259788 62144
rect 259828 62092 259880 62144
rect 255780 61999 255832 62008
rect 255780 61965 255789 61999
rect 255789 61965 255823 61999
rect 255823 61965 255832 61999
rect 255780 61956 255832 61965
rect 229468 60664 229520 60716
rect 229652 60664 229704 60716
rect 254860 60596 254912 60648
rect 277584 60392 277636 60444
rect 277952 60392 278004 60444
rect 273628 58624 273680 58676
rect 273904 58624 273956 58676
rect 235172 57944 235224 57996
rect 235264 57944 235316 57996
rect 235540 57987 235592 57996
rect 235540 57953 235549 57987
rect 235549 57953 235583 57987
rect 235583 57953 235592 57987
rect 235540 57944 235592 57953
rect 237196 57987 237248 57996
rect 237196 57953 237205 57987
rect 237205 57953 237239 57987
rect 237239 57953 237248 57987
rect 237196 57944 237248 57953
rect 229652 57876 229704 57928
rect 245292 57876 245344 57928
rect 269580 56559 269632 56568
rect 269580 56525 269589 56559
rect 269589 56525 269623 56559
rect 269623 56525 269632 56559
rect 269580 56516 269632 56525
rect 276940 53796 276992 53848
rect 277032 53796 277084 53848
rect 269672 53592 269724 53644
rect 255780 52479 255832 52488
rect 255780 52445 255789 52479
rect 255789 52445 255823 52479
rect 255823 52445 255832 52479
rect 255780 52436 255832 52445
rect 256976 52436 257028 52488
rect 257252 52436 257304 52488
rect 237196 51076 237248 51128
rect 255044 51076 255096 51128
rect 259828 51076 259880 51128
rect 3424 51008 3476 51060
rect 200764 51008 200816 51060
rect 237104 51008 237156 51060
rect 259920 51008 259972 51060
rect 235172 48356 235224 48408
rect 235264 48356 235316 48408
rect 229560 48331 229612 48340
rect 229560 48297 229569 48331
rect 229569 48297 229603 48331
rect 229603 48297 229612 48331
rect 229560 48288 229612 48297
rect 245200 48331 245252 48340
rect 245200 48297 245209 48331
rect 245209 48297 245243 48331
rect 245243 48297 245252 48331
rect 245200 48288 245252 48297
rect 257160 48288 257212 48340
rect 257252 48288 257304 48340
rect 271144 48288 271196 48340
rect 271236 48288 271288 48340
rect 273904 48288 273956 48340
rect 273996 48288 274048 48340
rect 277124 48288 277176 48340
rect 277216 48288 277268 48340
rect 235172 46903 235224 46912
rect 235172 46869 235181 46903
rect 235181 46869 235215 46903
rect 235215 46869 235224 46903
rect 235172 46860 235224 46869
rect 260564 45500 260616 45552
rect 262588 45500 262640 45552
rect 262680 45500 262732 45552
rect 264244 45543 264296 45552
rect 264244 45509 264253 45543
rect 264253 45509 264287 45543
rect 264287 45509 264296 45543
rect 264244 45500 264296 45509
rect 260564 45364 260616 45416
rect 276940 44956 276992 45008
rect 255780 44208 255832 44260
rect 256608 44115 256660 44124
rect 256608 44081 256617 44115
rect 256617 44081 256651 44115
rect 256651 44081 256660 44115
rect 256608 44072 256660 44081
rect 254768 42780 254820 42832
rect 255044 42780 255096 42832
rect 255872 42823 255924 42832
rect 255872 42789 255881 42823
rect 255881 42789 255915 42823
rect 255915 42789 255924 42823
rect 255872 42780 255924 42789
rect 229468 41352 229520 41404
rect 229652 41352 229704 41404
rect 237012 41352 237064 41404
rect 237196 41352 237248 41404
rect 277768 41352 277820 41404
rect 304264 41352 304316 41404
rect 580172 41352 580224 41404
rect 277952 41284 278004 41336
rect 257160 39355 257212 39364
rect 257160 39321 257169 39355
rect 257169 39321 257203 39355
rect 257203 39321 257212 39355
rect 257160 39312 257212 39321
rect 229652 38564 229704 38616
rect 235172 37315 235224 37324
rect 235172 37281 235181 37315
rect 235181 37281 235215 37315
rect 235215 37281 235224 37315
rect 235172 37272 235224 37281
rect 276848 37315 276900 37324
rect 276848 37281 276857 37315
rect 276857 37281 276891 37315
rect 276891 37281 276900 37315
rect 276848 37272 276900 37281
rect 269580 37204 269632 37256
rect 269672 37204 269724 37256
rect 271604 37247 271656 37256
rect 271604 37213 271613 37247
rect 271613 37213 271647 37247
rect 271647 37213 271656 37247
rect 271604 37204 271656 37213
rect 273628 37204 273680 37256
rect 273720 37204 273772 37256
rect 264244 35955 264296 35964
rect 264244 35921 264253 35955
rect 264253 35921 264287 35955
rect 264287 35921 264296 35955
rect 264244 35912 264296 35921
rect 3424 35844 3476 35896
rect 213184 35844 213236 35896
rect 260564 34620 260616 34672
rect 255780 34552 255832 34604
rect 254768 34484 254820 34536
rect 254860 34484 254912 34536
rect 255872 34484 255924 34536
rect 257252 34484 257304 34536
rect 260656 34484 260708 34536
rect 237196 31764 237248 31816
rect 237012 31696 237064 31748
rect 398104 29248 398156 29300
rect 405648 29248 405700 29300
rect 436744 29248 436796 29300
rect 444288 29248 444340 29300
rect 417332 29180 417384 29232
rect 424968 29180 425020 29232
rect 456708 29180 456760 29232
rect 463608 29180 463660 29232
rect 475292 29180 475344 29232
rect 482928 29180 482980 29232
rect 495164 29180 495216 29232
rect 502248 29180 502300 29232
rect 513564 29180 513616 29232
rect 521568 29180 521620 29232
rect 533804 29180 533856 29232
rect 540888 29180 540940 29232
rect 552480 29180 552532 29232
rect 560208 29180 560260 29232
rect 280252 29044 280304 29096
rect 289728 29044 289780 29096
rect 229560 29019 229612 29028
rect 229560 28985 229569 29019
rect 229569 28985 229603 29019
rect 229603 28985 229612 29019
rect 229560 28976 229612 28985
rect 260656 28976 260708 29028
rect 235540 28951 235592 28960
rect 235540 28917 235549 28951
rect 235549 28917 235583 28951
rect 235583 28917 235592 28951
rect 235540 28908 235592 28917
rect 260564 28908 260616 28960
rect 287612 28228 287664 28280
rect 567200 28228 567252 28280
rect 257252 27591 257304 27600
rect 257252 27557 257261 27591
rect 257261 27557 257295 27591
rect 257295 27557 257304 27591
rect 257252 27548 257304 27557
rect 259828 27548 259880 27600
rect 259920 27548 259972 27600
rect 274272 27591 274324 27600
rect 274272 27557 274281 27591
rect 274281 27557 274315 27591
rect 274315 27557 274324 27591
rect 274272 27548 274324 27557
rect 264244 26231 264296 26240
rect 264244 26197 264253 26231
rect 264253 26197 264287 26231
rect 264287 26197 264296 26231
rect 264244 26188 264296 26197
rect 268844 26231 268896 26240
rect 268844 26197 268853 26231
rect 268853 26197 268887 26231
rect 268887 26197 268896 26231
rect 268844 26188 268896 26197
rect 229560 22108 229612 22160
rect 277768 22108 277820 22160
rect 277952 22108 278004 22160
rect 3148 22040 3200 22092
rect 225604 22040 225656 22092
rect 229560 21972 229612 22024
rect 320824 21360 320876 21412
rect 561680 21360 561732 21412
rect 294696 19932 294748 19984
rect 543740 19932 543792 19984
rect 235172 19320 235224 19372
rect 235264 19320 235316 19372
rect 235540 19363 235592 19372
rect 235540 19329 235549 19363
rect 235549 19329 235583 19363
rect 235583 19329 235592 19363
rect 235540 19320 235592 19329
rect 237012 19320 237064 19372
rect 237104 19320 237156 19372
rect 250536 19252 250588 19304
rect 297364 18572 297416 18624
rect 525800 18572 525852 18624
rect 269672 18028 269724 18080
rect 256608 18003 256660 18012
rect 256608 17969 256617 18003
rect 256617 17969 256651 18003
rect 256651 17969 256660 18003
rect 256608 17960 256660 17969
rect 257252 18003 257304 18012
rect 257252 17969 257261 18003
rect 257261 17969 257295 18003
rect 257295 17969 257304 18003
rect 257252 17960 257304 17969
rect 269580 17960 269632 18012
rect 271604 18003 271656 18012
rect 271604 17969 271613 18003
rect 271613 17969 271647 18003
rect 271647 17969 271656 18003
rect 271604 17960 271656 17969
rect 274272 18003 274324 18012
rect 274272 17969 274281 18003
rect 274281 17969 274315 18003
rect 274315 17969 274324 18003
rect 274272 17960 274324 17969
rect 229100 17892 229152 17944
rect 579804 17892 579856 17944
rect 117228 17212 117280 17264
rect 222844 17212 222896 17264
rect 277768 17212 277820 17264
rect 278136 17212 278188 17264
rect 264244 16643 264296 16652
rect 264244 16609 264253 16643
rect 264253 16609 264287 16643
rect 264287 16609 264296 16643
rect 264244 16600 264296 16609
rect 268844 16643 268896 16652
rect 268844 16609 268853 16643
rect 268853 16609 268887 16643
rect 268887 16609 268896 16643
rect 268844 16600 268896 16609
rect 260656 16575 260708 16584
rect 260656 16541 260665 16575
rect 260665 16541 260699 16575
rect 260699 16541 260708 16575
rect 260656 16532 260708 16541
rect 262680 16532 262732 16584
rect 151636 15852 151688 15904
rect 245292 15852 245344 15904
rect 290464 15852 290516 15904
rect 514760 15852 514812 15904
rect 164148 14424 164200 14476
rect 228364 14424 228416 14476
rect 298744 14424 298796 14476
rect 512092 14424 512144 14476
rect 148968 13064 149020 13116
rect 225696 13064 225748 13116
rect 291844 13064 291896 13116
rect 507860 13064 507912 13116
rect 166908 11704 166960 11756
rect 226984 11704 227036 11756
rect 228916 11704 228968 11756
rect 252008 11704 252060 11756
rect 301504 11704 301556 11756
rect 503720 11704 503772 11756
rect 267464 10956 267516 11008
rect 356152 10956 356204 11008
rect 267280 10888 267332 10940
rect 358820 10888 358872 10940
rect 267188 10820 267240 10872
rect 362960 10820 363012 10872
rect 267372 10752 267424 10804
rect 365720 10752 365772 10804
rect 64788 10684 64840 10736
rect 236736 10684 236788 10736
rect 268844 10684 268896 10736
rect 369860 10684 369912 10736
rect 60648 10616 60700 10668
rect 236828 10616 236880 10668
rect 268660 10616 268712 10668
rect 374092 10616 374144 10668
rect 30288 10548 30340 10600
rect 233056 10548 233108 10600
rect 268752 10548 268804 10600
rect 376760 10548 376812 10600
rect 27528 10480 27580 10532
rect 232228 10480 232280 10532
rect 269212 10480 269264 10532
rect 380900 10480 380952 10532
rect 22008 10412 22060 10464
rect 232136 10412 232188 10464
rect 236000 10412 236052 10464
rect 253204 10412 253256 10464
rect 270040 10412 270092 10464
rect 383660 10412 383712 10464
rect 9588 10344 9640 10396
rect 230848 10344 230900 10396
rect 232504 10344 232556 10396
rect 252928 10344 252980 10396
rect 269120 10344 269172 10396
rect 387800 10344 387852 10396
rect 3976 10276 4028 10328
rect 229560 10276 229612 10328
rect 231308 10276 231360 10328
rect 251180 10276 251232 10328
rect 270224 10276 270276 10328
rect 390560 10276 390612 10328
rect 265992 10208 266044 10260
rect 351920 10208 351972 10260
rect 265808 10140 265860 10192
rect 347780 10140 347832 10192
rect 265716 10072 265768 10124
rect 345020 10072 345072 10124
rect 265072 10004 265124 10056
rect 340880 10004 340932 10056
rect 250444 9707 250496 9716
rect 250444 9673 250453 9707
rect 250453 9673 250487 9707
rect 250487 9673 250496 9707
rect 250444 9664 250496 9673
rect 256516 9707 256568 9716
rect 256516 9673 256525 9707
rect 256525 9673 256559 9707
rect 256559 9673 256568 9707
rect 256516 9664 256568 9673
rect 257160 9664 257212 9716
rect 257252 9664 257304 9716
rect 90916 9596 90968 9648
rect 239220 9596 239272 9648
rect 87328 9528 87380 9580
rect 239036 9528 239088 9580
rect 83832 9460 83884 9512
rect 238576 9460 238628 9512
rect 80244 9392 80296 9444
rect 238208 9392 238260 9444
rect 76656 9324 76708 9376
rect 237748 9324 237800 9376
rect 73068 9256 73120 9308
rect 237656 9256 237708 9308
rect 259920 9256 259972 9308
rect 291936 9256 291988 9308
rect 69480 9188 69532 9240
rect 236644 9188 236696 9240
rect 260012 9188 260064 9240
rect 295524 9188 295576 9240
rect 65984 9120 66036 9172
rect 236460 9120 236512 9172
rect 299112 9120 299164 9172
rect 62396 9052 62448 9104
rect 236552 9052 236604 9104
rect 261208 9052 261260 9104
rect 306196 9052 306248 9104
rect 58808 8984 58860 9036
rect 236368 8984 236420 9036
rect 261300 8984 261352 9036
rect 309784 8984 309836 9036
rect 17224 8916 17276 8968
rect 231676 8916 231728 8968
rect 241980 8916 242032 8968
rect 251824 8916 251876 8968
rect 261392 8916 261444 8968
rect 302608 8916 302660 8968
rect 302884 8916 302936 8968
rect 494152 8916 494204 8968
rect 94504 8848 94556 8900
rect 239680 8848 239732 8900
rect 98092 8780 98144 8832
rect 239128 8780 239180 8832
rect 101588 8712 101640 8764
rect 240416 8712 240468 8764
rect 105176 8644 105228 8696
rect 240324 8644 240376 8696
rect 108764 8576 108816 8628
rect 241152 8576 241204 8628
rect 112352 8508 112404 8560
rect 241888 8508 241940 8560
rect 115940 8440 115992 8492
rect 241796 8440 241848 8492
rect 119436 8372 119488 8424
rect 242256 8372 242308 8424
rect 269672 8372 269724 8424
rect 123024 8304 123076 8356
rect 242624 8304 242676 8356
rect 256516 8347 256568 8356
rect 256516 8313 256525 8347
rect 256525 8313 256559 8347
rect 256559 8313 256568 8347
rect 256516 8304 256568 8313
rect 269580 8304 269632 8356
rect 3424 8236 3476 8288
rect 135904 8236 135956 8288
rect 200396 8236 200448 8288
rect 250536 8236 250588 8288
rect 253848 8236 253900 8288
rect 255872 8236 255924 8288
rect 261484 8236 261536 8288
rect 267004 8236 267056 8288
rect 272524 8236 272576 8288
rect 275284 8236 275336 8288
rect 196808 8168 196860 8220
rect 250168 8168 250220 8220
rect 193220 8100 193272 8152
rect 249892 8100 249944 8152
rect 189632 8032 189684 8084
rect 249432 8032 249484 8084
rect 279976 8032 280028 8084
rect 186044 7964 186096 8016
rect 248696 7964 248748 8016
rect 182548 7896 182600 7948
rect 248788 7896 248840 7948
rect 178960 7828 179012 7880
rect 247408 7828 247460 7880
rect 279976 7828 280028 7880
rect 175372 7760 175424 7812
rect 247316 7760 247368 7812
rect 171784 7692 171836 7744
rect 247868 7692 247920 7744
rect 168196 7624 168248 7676
rect 247500 7624 247552 7676
rect 132592 7556 132644 7608
rect 243360 7556 243412 7608
rect 316684 7556 316736 7608
rect 490564 7556 490616 7608
rect 203892 7488 203944 7540
rect 250904 7488 250956 7540
rect 262588 6987 262640 6996
rect 262588 6953 262597 6987
rect 262597 6953 262631 6987
rect 262631 6953 262640 6987
rect 262588 6944 262640 6953
rect 262956 6876 263008 6928
rect 268108 6876 268160 6928
rect 279884 6876 279936 6928
rect 280068 6876 280120 6928
rect 280804 6876 280856 6928
rect 289544 6876 289596 6928
rect 199200 6808 199252 6860
rect 250352 6808 250404 6860
rect 264244 6851 264296 6860
rect 264244 6817 264253 6851
rect 264253 6817 264287 6851
rect 264287 6817 264296 6851
rect 264244 6808 264296 6817
rect 266820 6808 266872 6860
rect 354956 6808 355008 6860
rect 195612 6740 195664 6792
rect 250076 6740 250128 6792
rect 266728 6740 266780 6792
rect 358544 6740 358596 6792
rect 192024 6672 192076 6724
rect 249708 6672 249760 6724
rect 266544 6672 266596 6724
rect 362132 6672 362184 6724
rect 188436 6604 188488 6656
rect 249340 6604 249392 6656
rect 266452 6604 266504 6656
rect 365812 6604 365864 6656
rect 184848 6536 184900 6588
rect 248880 6536 248932 6588
rect 268292 6536 268344 6588
rect 369216 6536 369268 6588
rect 181352 6468 181404 6520
rect 248604 6468 248656 6520
rect 267924 6468 267976 6520
rect 372804 6468 372856 6520
rect 177764 6400 177816 6452
rect 248144 6400 248196 6452
rect 268016 6400 268068 6452
rect 376392 6400 376444 6452
rect 174176 6332 174228 6384
rect 247776 6332 247828 6384
rect 267832 6332 267884 6384
rect 379980 6332 380032 6384
rect 134892 6264 134944 6316
rect 243176 6264 243228 6316
rect 270132 6264 270184 6316
rect 383568 6264 383620 6316
rect 131396 6196 131448 6248
rect 243268 6196 243320 6248
rect 269396 6196 269448 6248
rect 387064 6196 387116 6248
rect 12440 6128 12492 6180
rect 230664 6128 230716 6180
rect 234804 6128 234856 6180
rect 254492 6128 254544 6180
rect 269488 6128 269540 6180
rect 390652 6128 390704 6180
rect 202696 6060 202748 6112
rect 250812 6060 250864 6112
rect 265440 6060 265492 6112
rect 351368 6060 351420 6112
rect 238392 5992 238444 6044
rect 254400 5992 254452 6044
rect 266084 5992 266136 6044
rect 347872 5992 347924 6044
rect 266176 5924 266228 5976
rect 344284 5924 344336 5976
rect 264980 5856 265032 5908
rect 340696 5856 340748 5908
rect 264152 5788 264204 5840
rect 337108 5788 337160 5840
rect 264060 5720 264112 5772
rect 333612 5720 333664 5772
rect 330024 5652 330076 5704
rect 262680 5584 262732 5636
rect 326436 5584 326488 5636
rect 262772 5516 262824 5568
rect 322848 5516 322900 5568
rect 198004 5448 198056 5500
rect 194416 5380 194468 5432
rect 257804 5448 257856 5500
rect 270592 5448 270644 5500
rect 249800 5380 249852 5432
rect 258632 5380 258684 5432
rect 274088 5380 274140 5432
rect 190828 5312 190880 5364
rect 249524 5312 249576 5364
rect 257988 5312 258040 5364
rect 272892 5312 272944 5364
rect 137284 5244 137336 5296
rect 140872 5176 140924 5228
rect 142068 5176 142120 5228
rect 187240 5244 187292 5296
rect 249616 5244 249668 5296
rect 258908 5244 258960 5296
rect 276480 5244 276532 5296
rect 244004 5176 244056 5228
rect 249984 5176 250036 5228
rect 258448 5176 258500 5228
rect 277676 5176 277728 5228
rect 133788 5108 133840 5160
rect 243728 5108 243780 5160
rect 244372 5108 244424 5160
rect 247684 5108 247736 5160
rect 259092 5108 259144 5160
rect 280068 5108 280120 5160
rect 130200 5040 130252 5092
rect 243452 5040 243504 5092
rect 259276 5040 259328 5092
rect 281264 5040 281316 5092
rect 7656 4972 7708 5024
rect 229284 4972 229336 5024
rect 259184 4972 259236 5024
rect 284760 4972 284812 5024
rect 2872 4904 2924 4956
rect 229192 4904 229244 4956
rect 240784 4904 240836 4956
rect 254308 4904 254360 4956
rect 260288 4904 260340 4956
rect 283564 4904 283616 4956
rect 1676 4836 1728 4888
rect 572 4768 624 4820
rect 237288 4836 237340 4888
rect 254124 4836 254176 4888
rect 258356 4836 258408 4888
rect 283656 4836 283708 4888
rect 332416 4836 332468 4888
rect 229376 4768 229428 4820
rect 233700 4768 233752 4820
rect 254216 4768 254268 4820
rect 260196 4768 260248 4820
rect 290740 4768 290792 4820
rect 315304 4768 315356 4820
rect 486976 4768 487028 4820
rect 489184 4768 489236 4820
rect 497740 4768 497792 4820
rect 201500 4700 201552 4752
rect 251088 4700 251140 4752
rect 257620 4700 257672 4752
rect 269304 4700 269356 4752
rect 287152 4700 287204 4752
rect 205088 4632 205140 4684
rect 250996 4632 251048 4684
rect 230756 4564 230808 4616
rect 124220 4156 124272 4208
rect 125416 4156 125468 4208
rect 150440 4156 150492 4208
rect 151636 4156 151688 4208
rect 158720 4156 158772 4208
rect 160008 4156 160060 4208
rect 167092 4156 167144 4208
rect 168288 4156 168340 4208
rect 209872 4156 209924 4208
rect 211068 4156 211120 4208
rect 265348 4156 265400 4208
rect 265808 4156 265860 4208
rect 287060 4156 287112 4208
rect 288348 4156 288400 4208
rect 296720 4156 296772 4208
rect 297916 4156 297968 4208
rect 313372 4156 313424 4208
rect 314568 4156 314620 4208
rect 347780 4156 347832 4208
rect 349068 4156 349120 4208
rect 356060 4156 356112 4208
rect 357348 4156 357400 4208
rect 365720 4156 365772 4208
rect 366916 4156 366968 4208
rect 374000 4156 374052 4208
rect 375196 4156 375248 4208
rect 20720 4088 20772 4140
rect 28264 4088 28316 4140
rect 79048 4088 79100 4140
rect 238024 4088 238076 4140
rect 239588 4088 239640 4140
rect 240048 4088 240100 4140
rect 255044 4088 255096 4140
rect 256148 4088 256200 4140
rect 258540 4088 258592 4140
rect 259828 4088 259880 4140
rect 262864 4088 262916 4140
rect 264612 4088 264664 4140
rect 273812 4088 273864 4140
rect 425060 4088 425112 4140
rect 556804 4088 556856 4140
rect 559564 4088 559616 4140
rect 84108 4020 84160 4072
rect 238484 4020 238536 4072
rect 243176 4020 243228 4072
rect 254860 4020 254912 4072
rect 257344 4020 257396 4072
rect 258632 4020 258684 4072
rect 273628 4020 273680 4072
rect 428740 4020 428792 4072
rect 71872 3952 71924 4004
rect 236276 3952 236328 4004
rect 257712 3952 257764 4004
rect 261024 3952 261076 4004
rect 273536 3952 273588 4004
rect 432328 3952 432380 4004
rect 68284 3884 68336 3936
rect 236184 3884 236236 3936
rect 257160 3884 257212 3936
rect 262220 3884 262272 3936
rect 275744 3884 275796 3936
rect 435824 3884 435876 3936
rect 64696 3816 64748 3868
rect 225328 3816 225380 3868
rect 226248 3816 226300 3868
rect 226524 3816 226576 3868
rect 227628 3816 227680 3868
rect 227720 3816 227772 3868
rect 229008 3816 229060 3868
rect 235540 3816 235592 3868
rect 250352 3816 250404 3868
rect 255964 3816 256016 3868
rect 257068 3816 257120 3868
rect 263416 3816 263468 3868
rect 275100 3816 275152 3868
rect 439412 3816 439464 3868
rect 61200 3748 61252 3800
rect 236092 3748 236144 3800
rect 275376 3748 275428 3800
rect 443000 3748 443052 3800
rect 44548 3680 44600 3732
rect 46204 3680 46256 3732
rect 57612 3680 57664 3732
rect 241336 3680 241388 3732
rect 275008 3680 275060 3732
rect 446588 3680 446640 3732
rect 571432 3680 571484 3732
rect 572628 3680 572680 3732
rect 573364 3680 573416 3732
rect 579804 3680 579856 3732
rect 46940 3612 46992 3664
rect 34980 3544 35032 3596
rect 8852 3476 8904 3528
rect 9588 3476 9640 3528
rect 10048 3476 10100 3528
rect 14464 3476 14516 3528
rect 18328 3476 18380 3528
rect 19984 3476 20036 3528
rect 23112 3476 23164 3528
rect 24124 3476 24176 3528
rect 26700 3476 26752 3528
rect 27528 3476 27580 3528
rect 5264 3408 5316 3460
rect 10324 3408 10376 3460
rect 19524 3408 19576 3460
rect 32404 3476 32456 3528
rect 33876 3476 33928 3528
rect 34428 3476 34480 3528
rect 37372 3544 37424 3596
rect 38568 3544 38620 3596
rect 43444 3544 43496 3596
rect 50528 3544 50580 3596
rect 50988 3544 51040 3596
rect 51632 3544 51684 3596
rect 52368 3544 52420 3596
rect 52828 3544 52880 3596
rect 53748 3544 53800 3596
rect 54024 3612 54076 3664
rect 235172 3612 235224 3664
rect 247960 3612 248012 3664
rect 254584 3612 254636 3664
rect 276572 3612 276624 3664
rect 450176 3612 450228 3664
rect 502432 3612 502484 3664
rect 503628 3612 503680 3664
rect 536932 3612 536984 3664
rect 538128 3612 538180 3664
rect 546500 3612 546552 3664
rect 547696 3612 547748 3664
rect 563152 3612 563204 3664
rect 564348 3612 564400 3664
rect 571984 3612 572036 3664
rect 581000 3612 581052 3664
rect 40960 3476 41012 3528
rect 42064 3476 42116 3528
rect 42156 3476 42208 3528
rect 42708 3476 42760 3528
rect 43352 3476 43404 3528
rect 238944 3544 238996 3596
rect 245568 3544 245620 3596
rect 255228 3544 255280 3596
rect 276388 3544 276440 3596
rect 453672 3544 453724 3596
rect 482284 3544 482336 3596
rect 567844 3544 567896 3596
rect 570236 3544 570288 3596
rect 570604 3544 570656 3596
rect 571432 3544 571484 3596
rect 574744 3544 574796 3596
rect 576216 3544 576268 3596
rect 229744 3476 229796 3528
rect 234068 3476 234120 3528
rect 277124 3476 277176 3528
rect 457260 3476 457312 3528
rect 467840 3476 467892 3528
rect 469128 3476 469180 3528
rect 475384 3476 475436 3528
rect 578608 3476 578660 3528
rect 29092 3408 29144 3460
rect 35164 3408 35216 3460
rect 39764 3408 39816 3460
rect 224960 3408 225012 3460
rect 235080 3408 235132 3460
rect 252652 3408 252704 3460
rect 255504 3408 255556 3460
rect 276848 3408 276900 3460
rect 460848 3408 460900 3460
rect 471244 3408 471296 3460
rect 582196 3408 582248 3460
rect 55220 3340 55272 3392
rect 56508 3340 56560 3392
rect 60004 3340 60056 3392
rect 60648 3340 60700 3392
rect 63592 3340 63644 3392
rect 64788 3340 64840 3392
rect 70676 3340 70728 3392
rect 71688 3340 71740 3392
rect 77852 3340 77904 3392
rect 78588 3340 78640 3392
rect 81440 3340 81492 3392
rect 82728 3340 82780 3392
rect 27896 3204 27948 3256
rect 31024 3204 31076 3256
rect 36176 3204 36228 3256
rect 39304 3204 39356 3256
rect 82636 3204 82688 3256
rect 84936 3272 84988 3324
rect 85488 3272 85540 3324
rect 237012 3340 237064 3392
rect 246764 3340 246816 3392
rect 255596 3340 255648 3392
rect 274272 3340 274324 3392
rect 421564 3340 421616 3392
rect 433340 3340 433392 3392
rect 434628 3340 434680 3392
rect 494060 3340 494112 3392
rect 495348 3340 495400 3392
rect 512000 3340 512052 3392
rect 513196 3340 513248 3392
rect 528560 3340 528612 3392
rect 529848 3340 529900 3392
rect 575020 3340 575072 3392
rect 86132 3204 86184 3256
rect 89720 3204 89772 3256
rect 229836 3272 229888 3324
rect 234436 3272 234488 3324
rect 272156 3272 272208 3324
rect 417976 3272 418028 3324
rect 574836 3272 574888 3324
rect 577412 3272 577464 3324
rect 238116 3204 238168 3256
rect 272340 3204 272392 3256
rect 414480 3204 414532 3256
rect 75460 3136 75512 3188
rect 84108 3136 84160 3188
rect 88524 3136 88576 3188
rect 89628 3136 89680 3188
rect 93308 3136 93360 3188
rect 239496 3136 239548 3188
rect 271972 3136 272024 3188
rect 410892 3136 410944 3188
rect 95700 3068 95752 3120
rect 96528 3068 96580 3120
rect 102784 3068 102836 3120
rect 103428 3068 103480 3120
rect 106372 3068 106424 3120
rect 107476 3068 107528 3120
rect 11244 3000 11296 3052
rect 15844 3000 15896 3052
rect 96896 3000 96948 3052
rect 239680 3068 239732 3120
rect 272248 3068 272300 3120
rect 407304 3068 407356 3120
rect 45744 2864 45796 2916
rect 50344 2864 50396 2916
rect 103980 2864 104032 2916
rect 113548 2932 113600 2984
rect 114468 2932 114520 2984
rect 111156 2864 111208 2916
rect 229652 3000 229704 3052
rect 239956 3000 240008 3052
rect 271144 3000 271196 3052
rect 403716 3000 403768 3052
rect 560944 3000 560996 3052
rect 566740 3000 566792 3052
rect 241060 2932 241112 2984
rect 249156 2932 249208 2984
rect 255688 2932 255740 2984
rect 271052 2932 271104 2984
rect 400220 2932 400272 2984
rect 114744 2864 114796 2916
rect 115848 2864 115900 2916
rect 120632 2864 120684 2916
rect 121368 2864 121420 2916
rect 118240 2796 118292 2848
rect 242072 2864 242124 2916
rect 271604 2864 271656 2916
rect 396632 2864 396684 2916
rect 425152 2864 425204 2916
rect 426348 2864 426400 2916
rect 121828 2796 121880 2848
rect 242164 2796 242216 2848
rect 269580 2796 269632 2848
rect 390560 2796 390612 2848
rect 391848 2796 391900 2848
rect 393044 2796 393096 2848
rect 256516 1844 256568 1896
rect 257436 1844 257488 1896
rect 270500 1368 270552 1420
rect 271696 1368 271748 1420
rect 74264 552 74316 604
rect 74448 552 74500 604
rect 92112 552 92164 604
rect 92388 552 92440 604
rect 109960 552 110012 604
rect 110328 552 110380 604
rect 183744 552 183796 604
rect 184756 552 184808 604
rect 206284 552 206336 604
rect 206928 552 206980 604
rect 207480 552 207532 604
rect 208308 552 208360 604
rect 208676 552 208728 604
rect 209688 552 209740 604
rect 230112 552 230164 604
rect 230388 552 230440 604
rect 251456 552 251508 604
rect 254676 552 254728 604
rect 281540 552 281592 604
rect 282460 552 282512 604
rect 285680 552 285732 604
rect 285956 552 286008 604
rect 299480 552 299532 604
rect 300308 552 300360 604
rect 300860 552 300912 604
rect 301412 552 301464 604
rect 303620 552 303672 604
rect 303804 552 303856 604
rect 492680 552 492732 604
rect 492956 552 493008 604
rect 495440 552 495492 604
rect 496544 552 496596 604
rect 498200 552 498252 604
rect 498936 552 498988 604
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 8128 700534 8156 703520
rect 8116 700528 8168 700534
rect 8116 700470 8168 700476
rect 24320 699718 24348 703520
rect 40512 700398 40540 703520
rect 72988 700806 73016 703520
rect 72976 700800 73028 700806
rect 72976 700742 73028 700748
rect 40500 700392 40552 700398
rect 40500 700334 40552 700340
rect 41328 700392 41380 700398
rect 41328 700334 41380 700340
rect 24308 699712 24360 699718
rect 24308 699654 24360 699660
rect 24768 699712 24820 699718
rect 24768 699654 24820 699660
rect 3422 682272 3478 682281
rect 3422 682207 3478 682216
rect 3054 653576 3110 653585
rect 3054 653511 3110 653520
rect 3068 652798 3096 653511
rect 3056 652792 3108 652798
rect 3056 652734 3108 652740
rect 3330 596048 3386 596057
rect 3330 595983 3386 595992
rect 3344 594862 3372 595983
rect 3332 594856 3384 594862
rect 3332 594798 3384 594804
rect 3330 553072 3386 553081
rect 3330 553007 3386 553016
rect 3344 552090 3372 553007
rect 3332 552084 3384 552090
rect 3332 552026 3384 552032
rect 3238 538656 3294 538665
rect 3238 538591 3294 538600
rect 3252 538286 3280 538591
rect 3240 538280 3292 538286
rect 3240 538222 3292 538228
rect 3330 495544 3386 495553
rect 3330 495479 3332 495488
rect 3384 495479 3386 495488
rect 3332 495450 3384 495456
rect 2962 481128 3018 481137
rect 2962 481063 3018 481072
rect 2976 480282 3004 481063
rect 2964 480276 3016 480282
rect 2964 480218 3016 480224
rect 3330 438016 3386 438025
rect 3330 437951 3386 437960
rect 3344 437510 3372 437951
rect 3332 437504 3384 437510
rect 3332 437446 3384 437452
rect 3330 423736 3386 423745
rect 3330 423671 3332 423680
rect 3384 423671 3386 423680
rect 3332 423642 3384 423648
rect 3436 402558 3464 682207
rect 3514 667992 3570 668001
rect 3514 667927 3516 667936
rect 3568 667927 3570 667936
rect 3516 667898 3568 667904
rect 3514 624880 3570 624889
rect 3514 624815 3570 624824
rect 3424 402552 3476 402558
rect 3424 402494 3476 402500
rect 3528 402490 3556 624815
rect 3606 610464 3662 610473
rect 3606 610399 3662 610408
rect 3620 610026 3648 610399
rect 3608 610020 3660 610026
rect 3608 609962 3660 609968
rect 3698 567352 3754 567361
rect 3698 567287 3754 567296
rect 3516 402484 3568 402490
rect 3516 402426 3568 402432
rect 3712 402422 3740 567287
rect 3882 509960 3938 509969
rect 3882 509895 3938 509904
rect 3700 402416 3752 402422
rect 3700 402358 3752 402364
rect 3896 402354 3924 509895
rect 4066 452432 4122 452441
rect 4066 452367 4122 452376
rect 3884 402348 3936 402354
rect 3884 402290 3936 402296
rect 4080 402286 4108 452367
rect 24780 402626 24808 699654
rect 41340 402694 41368 700334
rect 89180 699718 89208 703520
rect 105464 699718 105492 703520
rect 137848 700262 137876 703520
rect 137836 700256 137888 700262
rect 137836 700198 137888 700204
rect 89168 699712 89220 699718
rect 89168 699654 89220 699660
rect 89628 699712 89680 699718
rect 89628 699654 89680 699660
rect 105452 699712 105504 699718
rect 105452 699654 105504 699660
rect 106188 699712 106240 699718
rect 106188 699654 106240 699660
rect 89640 402762 89668 699654
rect 106200 402830 106228 699654
rect 154132 695570 154160 703520
rect 170324 699718 170352 703520
rect 202800 699990 202828 703520
rect 218992 703474 219020 703520
rect 218900 703446 219020 703474
rect 202788 699984 202840 699990
rect 202788 699926 202840 699932
rect 170312 699712 170364 699718
rect 170312 699654 170364 699660
rect 171048 699712 171100 699718
rect 171048 699654 171100 699660
rect 154120 695564 154172 695570
rect 154120 695506 154172 695512
rect 154212 695564 154264 695570
rect 154212 695506 154264 695512
rect 154224 688634 154252 695506
rect 154212 688628 154264 688634
rect 154212 688570 154264 688576
rect 154396 688628 154448 688634
rect 154396 688570 154448 688576
rect 154408 685846 154436 688570
rect 154396 685840 154448 685846
rect 154396 685782 154448 685788
rect 154304 676252 154356 676258
rect 154304 676194 154356 676200
rect 154316 673538 154344 676194
rect 154304 673532 154356 673538
rect 154304 673474 154356 673480
rect 154488 673532 154540 673538
rect 154488 673474 154540 673480
rect 154500 663762 154528 673474
rect 154316 663734 154528 663762
rect 154316 654158 154344 663734
rect 154304 654152 154356 654158
rect 154304 654094 154356 654100
rect 154488 654152 154540 654158
rect 154488 654094 154540 654100
rect 154500 644450 154528 654094
rect 154316 644422 154528 644450
rect 154316 634846 154344 644422
rect 154304 634840 154356 634846
rect 154304 634782 154356 634788
rect 154488 634840 154540 634846
rect 154488 634782 154540 634788
rect 154500 625138 154528 634782
rect 154316 625110 154528 625138
rect 154316 615534 154344 625110
rect 154304 615528 154356 615534
rect 154304 615470 154356 615476
rect 154488 615528 154540 615534
rect 154488 615470 154540 615476
rect 154500 605826 154528 615470
rect 154316 605798 154528 605826
rect 154316 596222 154344 605798
rect 154304 596216 154356 596222
rect 154488 596216 154540 596222
rect 154304 596158 154356 596164
rect 154408 596164 154488 596170
rect 154408 596158 154540 596164
rect 154408 596142 154528 596158
rect 154408 591954 154436 596142
rect 154316 591926 154436 591954
rect 154316 589286 154344 591926
rect 154304 589280 154356 589286
rect 154304 589222 154356 589228
rect 154304 579760 154356 579766
rect 154224 579708 154304 579714
rect 154224 579702 154356 579708
rect 154224 579686 154344 579702
rect 154224 579630 154252 579686
rect 154212 579624 154264 579630
rect 154212 579566 154264 579572
rect 154396 579624 154448 579630
rect 154396 579566 154448 579572
rect 154408 562970 154436 579566
rect 154212 562964 154264 562970
rect 154212 562906 154264 562912
rect 154396 562964 154448 562970
rect 154396 562906 154448 562912
rect 154224 553330 154252 562906
rect 154224 553302 154344 553330
rect 154316 543810 154344 553302
rect 154316 543782 154528 543810
rect 154500 534018 154528 543782
rect 154408 533990 154528 534018
rect 154408 531282 154436 533990
rect 154396 531276 154448 531282
rect 154396 531218 154448 531224
rect 154488 521688 154540 521694
rect 154488 521630 154540 521636
rect 154500 514706 154528 521630
rect 154408 514678 154528 514706
rect 154408 511970 154436 514678
rect 154396 511964 154448 511970
rect 154396 511906 154448 511912
rect 154488 502376 154540 502382
rect 154488 502318 154540 502324
rect 154500 495394 154528 502318
rect 154408 495366 154528 495394
rect 154408 492658 154436 495366
rect 154212 492652 154264 492658
rect 154212 492594 154264 492600
rect 154396 492652 154448 492658
rect 154396 492594 154448 492600
rect 154224 483041 154252 492594
rect 154210 483032 154266 483041
rect 154210 482967 154266 482976
rect 154486 483032 154542 483041
rect 154486 482967 154542 482976
rect 154500 476082 154528 482967
rect 154316 476054 154528 476082
rect 154316 466478 154344 476054
rect 154304 466472 154356 466478
rect 154304 466414 154356 466420
rect 154488 466472 154540 466478
rect 154488 466414 154540 466420
rect 154500 456770 154528 466414
rect 154316 456742 154528 456770
rect 154316 454034 154344 456742
rect 154304 454028 154356 454034
rect 154304 453970 154356 453976
rect 154212 444440 154264 444446
rect 154212 444382 154264 444388
rect 154224 437458 154252 444382
rect 154224 437430 154436 437458
rect 154408 434722 154436 437430
rect 154396 434716 154448 434722
rect 154396 434658 154448 434664
rect 154396 427780 154448 427786
rect 154396 427722 154448 427728
rect 154408 425082 154436 427722
rect 154408 425054 154528 425082
rect 154500 418146 154528 425054
rect 154316 418118 154528 418146
rect 154316 415410 154344 418118
rect 154304 415404 154356 415410
rect 154304 415346 154356 415352
rect 154396 405748 154448 405754
rect 154396 405690 154448 405696
rect 154408 402898 154436 405690
rect 171060 402966 171088 699654
rect 218900 695745 218928 703446
rect 235184 699718 235212 703520
rect 257896 701004 257948 701010
rect 257896 700946 257948 700952
rect 256424 700732 256476 700738
rect 256424 700674 256476 700680
rect 255228 700460 255280 700466
rect 255228 700402 255280 700408
rect 255136 700392 255188 700398
rect 255136 700334 255188 700340
rect 253848 700324 253900 700330
rect 253848 700266 253900 700272
rect 235172 699712 235224 699718
rect 235172 699654 235224 699660
rect 235908 699712 235960 699718
rect 235908 699654 235960 699660
rect 218886 695736 218942 695745
rect 218886 695671 218942 695680
rect 219254 695600 219310 695609
rect 219176 695558 219254 695586
rect 219176 695502 219204 695558
rect 219254 695535 219310 695544
rect 219164 695496 219216 695502
rect 219164 695438 219216 695444
rect 219072 685908 219124 685914
rect 219072 685850 219124 685856
rect 219084 678994 219112 685850
rect 218992 678966 219112 678994
rect 218992 676190 219020 678966
rect 218980 676184 219032 676190
rect 218980 676126 219032 676132
rect 219072 666596 219124 666602
rect 219072 666538 219124 666544
rect 219084 659682 219112 666538
rect 219084 659666 219204 659682
rect 219084 659660 219216 659666
rect 219084 659654 219164 659660
rect 219164 659602 219216 659608
rect 219348 659660 219400 659666
rect 219348 659602 219400 659608
rect 219360 656878 219388 659602
rect 219348 656872 219400 656878
rect 219348 656814 219400 656820
rect 219256 647284 219308 647290
rect 219256 647226 219308 647232
rect 219268 640422 219296 647226
rect 219256 640416 219308 640422
rect 219256 640358 219308 640364
rect 219072 640280 219124 640286
rect 219072 640222 219124 640228
rect 219084 637566 219112 640222
rect 219072 637560 219124 637566
rect 219072 637502 219124 637508
rect 219164 637560 219216 637566
rect 219164 637502 219216 637508
rect 219176 630578 219204 637502
rect 219176 630550 219388 630578
rect 219360 626550 219388 630550
rect 219348 626544 219400 626550
rect 219348 626486 219400 626492
rect 219348 616888 219400 616894
rect 219348 616830 219400 616836
rect 219360 611454 219388 616830
rect 219348 611448 219400 611454
rect 219348 611390 219400 611396
rect 219072 608728 219124 608734
rect 219072 608670 219124 608676
rect 219084 608598 219112 608670
rect 219072 608592 219124 608598
rect 219072 608534 219124 608540
rect 219256 601588 219308 601594
rect 219256 601530 219308 601536
rect 219268 598942 219296 601530
rect 219256 598936 219308 598942
rect 219256 598878 219308 598884
rect 219164 589348 219216 589354
rect 219164 589290 219216 589296
rect 219176 582418 219204 589290
rect 218980 582412 219032 582418
rect 218980 582354 219032 582360
rect 219164 582412 219216 582418
rect 219164 582354 219216 582360
rect 218992 579630 219020 582354
rect 218980 579624 219032 579630
rect 218980 579566 219032 579572
rect 218888 569968 218940 569974
rect 218888 569910 218940 569916
rect 218900 563106 218928 569910
rect 218888 563100 218940 563106
rect 218888 563042 218940 563048
rect 218980 562964 219032 562970
rect 218980 562906 219032 562912
rect 218992 560266 219020 562906
rect 218900 560238 219020 560266
rect 218900 553450 218928 560238
rect 218888 553444 218940 553450
rect 218888 553386 218940 553392
rect 218888 550656 218940 550662
rect 218888 550598 218940 550604
rect 218900 543794 218928 550598
rect 218888 543788 218940 543794
rect 218888 543730 218940 543736
rect 218980 543652 219032 543658
rect 218980 543594 219032 543600
rect 218992 540977 219020 543594
rect 218978 540968 219034 540977
rect 218978 540903 219034 540912
rect 219162 540968 219218 540977
rect 219162 540903 219218 540912
rect 219176 533882 219204 540903
rect 218992 533854 219204 533882
rect 218992 531321 219020 533854
rect 218978 531312 219034 531321
rect 218978 531247 219034 531256
rect 219162 531312 219218 531321
rect 219162 531247 219218 531256
rect 219176 524346 219204 531247
rect 218980 524340 219032 524346
rect 218980 524282 219032 524288
rect 219164 524340 219216 524346
rect 219164 524282 219216 524288
rect 218992 521665 219020 524282
rect 218794 521656 218850 521665
rect 218794 521591 218850 521600
rect 218978 521656 219034 521665
rect 218978 521591 219034 521600
rect 218808 514690 218836 521591
rect 218796 514684 218848 514690
rect 218796 514626 218848 514632
rect 219072 514684 219124 514690
rect 219072 514626 219124 514632
rect 219084 510610 219112 514626
rect 219072 510604 219124 510610
rect 219072 510546 219124 510552
rect 219072 505096 219124 505102
rect 219072 505038 219124 505044
rect 219084 492726 219112 505038
rect 219072 492720 219124 492726
rect 219072 492662 219124 492668
rect 219164 492720 219216 492726
rect 219164 492662 219216 492668
rect 219176 485858 219204 492662
rect 219164 485852 219216 485858
rect 219164 485794 219216 485800
rect 219256 485716 219308 485722
rect 219256 485658 219308 485664
rect 219268 473385 219296 485658
rect 218978 473376 219034 473385
rect 218978 473311 219034 473320
rect 219254 473376 219310 473385
rect 219254 473311 219310 473320
rect 218992 466478 219020 473311
rect 218980 466472 219032 466478
rect 218980 466414 219032 466420
rect 219348 466336 219400 466342
rect 219348 466278 219400 466284
rect 219360 456770 219388 466278
rect 219084 456742 219388 456770
rect 219084 454034 219112 456742
rect 219072 454028 219124 454034
rect 219072 453970 219124 453976
rect 218980 444440 219032 444446
rect 218980 444382 219032 444388
rect 218992 437458 219020 444382
rect 218992 437430 219112 437458
rect 219084 434722 219112 437430
rect 218980 434716 219032 434722
rect 218980 434658 219032 434664
rect 219072 434716 219124 434722
rect 219072 434658 219124 434664
rect 218992 425105 219020 434658
rect 218978 425096 219034 425105
rect 218978 425031 219034 425040
rect 219346 425096 219402 425105
rect 219346 425031 219402 425040
rect 171048 402960 171100 402966
rect 171048 402902 171100 402908
rect 154396 402892 154448 402898
rect 154396 402834 154448 402840
rect 106188 402824 106240 402830
rect 106188 402766 106240 402772
rect 89628 402756 89680 402762
rect 89628 402698 89680 402704
rect 41328 402688 41380 402694
rect 41328 402630 41380 402636
rect 24768 402620 24820 402626
rect 24768 402562 24820 402568
rect 4068 402280 4120 402286
rect 4068 402222 4120 402228
rect 219360 402218 219388 425031
rect 219348 402212 219400 402218
rect 219348 402154 219400 402160
rect 235920 402082 235948 699654
rect 253756 696992 253808 696998
rect 253756 696934 253808 696940
rect 253664 685908 253716 685914
rect 253664 685850 253716 685856
rect 252468 673532 252520 673538
rect 252468 673474 252520 673480
rect 252376 650072 252428 650078
rect 252376 650014 252428 650020
rect 252284 638988 252336 638994
rect 252284 638930 252336 638936
rect 251088 626612 251140 626618
rect 251088 626554 251140 626560
rect 249708 603152 249760 603158
rect 249708 603094 249760 603100
rect 249616 579692 249668 579698
rect 249616 579634 249668 579640
rect 248328 556232 248380 556238
rect 248328 556174 248380 556180
rect 248236 532772 248288 532778
rect 248236 532714 248288 532720
rect 246948 509312 247000 509318
rect 246948 509254 247000 509260
rect 246856 485852 246908 485858
rect 246856 485794 246908 485800
rect 245568 462392 245620 462398
rect 245568 462334 245620 462340
rect 245476 451308 245528 451314
rect 245476 451250 245528 451256
rect 245384 438932 245436 438938
rect 245384 438874 245436 438880
rect 244188 415472 244240 415478
rect 244188 415414 244240 415420
rect 243820 404388 243872 404394
rect 243820 404330 243872 404336
rect 240692 402144 240744 402150
rect 240692 402086 240744 402092
rect 235908 402076 235960 402082
rect 235908 402018 235960 402024
rect 235908 401940 235960 401946
rect 235908 401882 235960 401888
rect 239128 401940 239180 401946
rect 239128 401882 239180 401888
rect 3976 401804 4028 401810
rect 3976 401746 4028 401752
rect 3792 401736 3844 401742
rect 3792 401678 3844 401684
rect 3608 401668 3660 401674
rect 3608 401610 3660 401616
rect 3148 396024 3200 396030
rect 3148 395966 3200 395972
rect 3160 395049 3188 395966
rect 3146 395040 3202 395049
rect 3146 394975 3202 394984
rect 3424 380860 3476 380866
rect 3424 380802 3476 380808
rect 3436 380633 3464 380802
rect 3422 380624 3478 380633
rect 3422 380559 3478 380568
rect 2964 367056 3016 367062
rect 2964 366998 3016 367004
rect 2976 366217 3004 366998
rect 2962 366208 3018 366217
rect 2962 366143 3018 366152
rect 3424 338088 3476 338094
rect 3424 338030 3476 338036
rect 3436 337521 3464 338030
rect 3422 337512 3478 337521
rect 3422 337447 3478 337456
rect 3424 309120 3476 309126
rect 3424 309062 3476 309068
rect 3436 308825 3464 309062
rect 3422 308816 3478 308825
rect 3422 308751 3478 308760
rect 3056 295316 3108 295322
rect 3056 295258 3108 295264
rect 3068 294409 3096 295258
rect 3054 294400 3110 294409
rect 3054 294335 3110 294344
rect 2872 266348 2924 266354
rect 2872 266290 2924 266296
rect 2884 265713 2912 266290
rect 2870 265704 2926 265713
rect 2870 265639 2926 265648
rect 3424 252544 3476 252550
rect 3424 252486 3476 252492
rect 3436 251297 3464 252486
rect 3422 251288 3478 251297
rect 3422 251223 3478 251232
rect 3620 237017 3648 401610
rect 3804 280129 3832 401678
rect 3988 323105 4016 401746
rect 13084 401328 13136 401334
rect 13084 401270 13136 401276
rect 10968 399968 11020 399974
rect 10968 399910 11020 399916
rect 10980 396030 11008 399910
rect 10968 396024 11020 396030
rect 10968 395966 11020 395972
rect 13096 338094 13124 401270
rect 226984 401260 227036 401266
rect 226984 401202 227036 401208
rect 225788 401124 225840 401130
rect 225788 401066 225840 401072
rect 218704 400784 218756 400790
rect 218704 400726 218756 400732
rect 211804 400716 211856 400722
rect 211804 400658 211856 400664
rect 207664 400580 207716 400586
rect 207664 400522 207716 400528
rect 203524 400376 203576 400382
rect 203524 400318 203576 400324
rect 135904 398948 135956 398954
rect 135904 398890 135956 398896
rect 17222 398032 17278 398041
rect 17222 397967 17278 397976
rect 13084 338088 13136 338094
rect 13084 338030 13136 338036
rect 14464 337544 14516 337550
rect 14464 337486 14516 337492
rect 10324 337408 10376 337414
rect 10324 337350 10376 337356
rect 3974 323096 4030 323105
rect 3974 323031 4030 323040
rect 3790 280120 3846 280129
rect 3790 280055 3846 280064
rect 3606 237008 3662 237017
rect 3606 236943 3662 236952
rect 3148 223576 3200 223582
rect 3148 223518 3200 223524
rect 3160 222601 3188 223518
rect 3146 222592 3202 222601
rect 3146 222527 3202 222536
rect 3424 208344 3476 208350
rect 3424 208286 3476 208292
rect 3436 208185 3464 208286
rect 3422 208176 3478 208185
rect 3422 208111 3478 208120
rect 3330 194576 3386 194585
rect 3330 194511 3386 194520
rect 3344 193905 3372 194511
rect 3330 193896 3386 193905
rect 3330 193831 3386 193840
rect 3240 180804 3292 180810
rect 3240 180746 3292 180752
rect 3252 179489 3280 180746
rect 3238 179480 3294 179489
rect 3238 179415 3294 179424
rect 3516 165572 3568 165578
rect 3516 165514 3568 165520
rect 3528 165073 3556 165514
rect 3514 165064 3570 165073
rect 3514 164999 3570 165008
rect 3148 151768 3200 151774
rect 3148 151710 3200 151716
rect 3160 150793 3188 151710
rect 3146 150784 3202 150793
rect 3146 150719 3202 150728
rect 3240 136604 3292 136610
rect 3240 136546 3292 136552
rect 3252 136377 3280 136546
rect 3238 136368 3294 136377
rect 3238 136303 3294 136312
rect 3424 122800 3476 122806
rect 3424 122742 3476 122748
rect 3436 122097 3464 122742
rect 3422 122088 3478 122097
rect 3422 122023 3478 122032
rect 3422 109032 3478 109041
rect 3422 108967 3478 108976
rect 3436 107681 3464 108967
rect 3422 107672 3478 107681
rect 3422 107607 3478 107616
rect 3424 93832 3476 93838
rect 3424 93774 3476 93780
rect 3436 93265 3464 93774
rect 3422 93256 3478 93265
rect 3422 93191 3478 93200
rect 3424 80028 3476 80034
rect 3424 79970 3476 79976
rect 3436 78985 3464 79970
rect 3422 78976 3478 78985
rect 3422 78911 3478 78920
rect 3332 64864 3384 64870
rect 3332 64806 3384 64812
rect 3344 64569 3372 64806
rect 3330 64560 3386 64569
rect 3330 64495 3386 64504
rect 3424 51060 3476 51066
rect 3424 51002 3476 51008
rect 3436 50153 3464 51002
rect 3422 50144 3478 50153
rect 3422 50079 3478 50088
rect 3424 35896 3476 35902
rect 3422 35864 3424 35873
rect 3476 35864 3478 35873
rect 3422 35799 3478 35808
rect 3148 22092 3200 22098
rect 3148 22034 3200 22040
rect 3160 21457 3188 22034
rect 3146 21448 3202 21457
rect 3146 21383 3202 21392
rect 9588 10396 9640 10402
rect 9588 10338 9640 10344
rect 3976 10328 4028 10334
rect 3976 10270 4028 10276
rect 3424 8288 3476 8294
rect 3424 8230 3476 8236
rect 3436 7177 3464 8230
rect 3422 7168 3478 7177
rect 3422 7103 3478 7112
rect 2872 4956 2924 4962
rect 2872 4898 2924 4904
rect 1676 4888 1728 4894
rect 1676 4830 1728 4836
rect 572 4820 624 4826
rect 572 4762 624 4768
rect 584 480 612 4762
rect 1688 480 1716 4830
rect 2884 480 2912 4898
rect 3988 626 4016 10270
rect 7656 5024 7708 5030
rect 7656 4966 7708 4972
rect 5264 3460 5316 3466
rect 5264 3402 5316 3408
rect 3988 598 4108 626
rect 4080 480 4108 598
rect 5276 480 5304 3402
rect 6458 3360 6514 3369
rect 6458 3295 6514 3304
rect 6472 480 6500 3295
rect 7668 480 7696 4966
rect 9600 3534 9628 10338
rect 8852 3528 8904 3534
rect 8852 3470 8904 3476
rect 9588 3528 9640 3534
rect 9588 3470 9640 3476
rect 10048 3528 10100 3534
rect 10048 3470 10100 3476
rect 8864 480 8892 3470
rect 10060 480 10088 3470
rect 10336 3466 10364 337350
rect 13728 319456 13780 319462
rect 13728 319398 13780 319404
rect 12440 6180 12492 6186
rect 12440 6122 12492 6128
rect 10324 3460 10376 3466
rect 10324 3402 10376 3408
rect 11244 3052 11296 3058
rect 11244 2994 11296 3000
rect 11256 480 11284 2994
rect 12452 480 12480 6122
rect 13740 3482 13768 319398
rect 14476 3534 14504 337486
rect 15844 337476 15896 337482
rect 15844 337418 15896 337424
rect 13648 3454 13768 3482
rect 14464 3528 14516 3534
rect 14464 3470 14516 3476
rect 14830 3496 14886 3505
rect 13648 480 13676 3454
rect 14830 3431 14886 3440
rect 14844 480 14872 3431
rect 15856 3058 15884 337418
rect 17236 136610 17264 397967
rect 125508 338088 125560 338094
rect 125508 338030 125560 338036
rect 107568 338020 107620 338026
rect 107568 337962 107620 337968
rect 100668 337884 100720 337890
rect 100668 337826 100720 337832
rect 35164 337816 35216 337822
rect 35164 337758 35216 337764
rect 32404 337680 32456 337686
rect 32404 337622 32456 337628
rect 28264 337612 28316 337618
rect 28264 337554 28316 337560
rect 19984 326392 20036 326398
rect 19984 326334 20036 326340
rect 17224 136604 17276 136610
rect 17224 136546 17276 136552
rect 17224 8968 17276 8974
rect 17224 8910 17276 8916
rect 16026 3632 16082 3641
rect 16026 3567 16082 3576
rect 15844 3052 15896 3058
rect 15844 2994 15896 3000
rect 16040 480 16068 3567
rect 17236 480 17264 8910
rect 19996 3534 20024 326334
rect 24124 315308 24176 315314
rect 24124 315250 24176 315256
rect 22008 10464 22060 10470
rect 22008 10406 22060 10412
rect 20720 4140 20772 4146
rect 20720 4082 20772 4088
rect 18328 3528 18380 3534
rect 18328 3470 18380 3476
rect 19984 3528 20036 3534
rect 19984 3470 20036 3476
rect 18340 480 18368 3470
rect 19524 3460 19576 3466
rect 19524 3402 19576 3408
rect 19536 480 19564 3402
rect 20732 480 20760 4082
rect 22020 626 22048 10406
rect 24136 3534 24164 315250
rect 27528 10532 27580 10538
rect 27528 10474 27580 10480
rect 25502 3904 25558 3913
rect 25502 3839 25558 3848
rect 24306 3768 24362 3777
rect 24306 3703 24362 3712
rect 23112 3528 23164 3534
rect 23112 3470 23164 3476
rect 24124 3528 24176 3534
rect 24124 3470 24176 3476
rect 21928 598 22048 626
rect 21928 480 21956 598
rect 23124 480 23152 3470
rect 24320 480 24348 3703
rect 25516 480 25544 3839
rect 27540 3534 27568 10474
rect 28276 4146 28304 337554
rect 31024 313948 31076 313954
rect 31024 313890 31076 313896
rect 30288 10600 30340 10606
rect 30288 10542 30340 10548
rect 28264 4140 28316 4146
rect 28264 4082 28316 4088
rect 26700 3528 26752 3534
rect 26700 3470 26752 3476
rect 27528 3528 27580 3534
rect 27528 3470 27580 3476
rect 26712 480 26740 3470
rect 29092 3460 29144 3466
rect 29092 3402 29144 3408
rect 27896 3256 27948 3262
rect 27896 3198 27948 3204
rect 27908 480 27936 3198
rect 29104 480 29132 3402
rect 30300 480 30328 10542
rect 31036 3262 31064 313890
rect 31668 312588 31720 312594
rect 31668 312530 31720 312536
rect 31680 3482 31708 312530
rect 32416 3534 32444 337622
rect 34428 330540 34480 330546
rect 34428 330482 34480 330488
rect 32678 4040 32734 4049
rect 32678 3975 32734 3984
rect 31496 3454 31708 3482
rect 32404 3528 32456 3534
rect 32404 3470 32456 3476
rect 31024 3256 31076 3262
rect 31024 3198 31076 3204
rect 31496 480 31524 3454
rect 32692 480 32720 3975
rect 34440 3534 34468 330482
rect 34980 3596 35032 3602
rect 34980 3538 35032 3544
rect 33876 3528 33928 3534
rect 33876 3470 33928 3476
rect 34428 3528 34480 3534
rect 34428 3470 34480 3476
rect 33888 480 33916 3470
rect 34992 480 35020 3538
rect 35176 3466 35204 337758
rect 39304 337748 39356 337754
rect 39304 337690 39356 337696
rect 38568 329112 38620 329118
rect 38568 329054 38620 329060
rect 38476 305652 38528 305658
rect 38476 305594 38528 305600
rect 37372 3596 37424 3602
rect 37372 3538 37424 3544
rect 35164 3460 35216 3466
rect 35164 3402 35216 3408
rect 36176 3256 36228 3262
rect 36176 3198 36228 3204
rect 36188 480 36216 3198
rect 37384 480 37412 3538
rect 38488 3482 38516 305594
rect 38580 3602 38608 329054
rect 38568 3596 38620 3602
rect 38568 3538 38620 3544
rect 38488 3454 38608 3482
rect 38580 480 38608 3454
rect 39316 3262 39344 337690
rect 71688 336116 71740 336122
rect 71688 336058 71740 336064
rect 48228 336048 48280 336054
rect 48228 335990 48280 335996
rect 42064 324964 42116 324970
rect 42064 324906 42116 324912
rect 42076 3534 42104 324906
rect 46204 323604 46256 323610
rect 46204 323546 46256 323552
rect 43444 307080 43496 307086
rect 43444 307022 43496 307028
rect 42708 304292 42760 304298
rect 42708 304234 42760 304240
rect 42720 3534 42748 304234
rect 43456 3602 43484 307022
rect 46216 3738 46244 323546
rect 44548 3732 44600 3738
rect 44548 3674 44600 3680
rect 46204 3732 46256 3738
rect 46204 3674 46256 3680
rect 43444 3596 43496 3602
rect 43444 3538 43496 3544
rect 40960 3528 41012 3534
rect 40960 3470 41012 3476
rect 42064 3528 42116 3534
rect 42064 3470 42116 3476
rect 42156 3528 42208 3534
rect 42156 3470 42208 3476
rect 42708 3528 42760 3534
rect 42708 3470 42760 3476
rect 43352 3528 43404 3534
rect 43352 3470 43404 3476
rect 39764 3460 39816 3466
rect 39764 3402 39816 3408
rect 39304 3256 39356 3262
rect 39304 3198 39356 3204
rect 39776 480 39804 3402
rect 40972 480 41000 3470
rect 42168 480 42196 3470
rect 43364 480 43392 3470
rect 44560 480 44588 3674
rect 46940 3664 46992 3670
rect 46940 3606 46992 3612
rect 45744 2916 45796 2922
rect 45744 2858 45796 2864
rect 45756 480 45784 2858
rect 46952 480 46980 3606
rect 48240 3482 48268 335990
rect 52368 334620 52420 334626
rect 52368 334562 52420 334568
rect 49608 331900 49660 331906
rect 49608 331842 49660 331848
rect 49620 3482 49648 331842
rect 50988 318096 51040 318102
rect 50988 318038 51040 318044
rect 50344 311160 50396 311166
rect 50344 311102 50396 311108
rect 48148 3454 48268 3482
rect 49344 3454 49648 3482
rect 48148 480 48176 3454
rect 49344 480 49372 3454
rect 50356 2922 50384 311102
rect 51000 3602 51028 318038
rect 52380 3602 52408 334562
rect 56508 333260 56560 333266
rect 56508 333202 56560 333208
rect 53748 327752 53800 327758
rect 53748 327694 53800 327700
rect 53760 3602 53788 327694
rect 56416 326460 56468 326466
rect 56416 326402 56468 326408
rect 54024 3664 54076 3670
rect 54024 3606 54076 3612
rect 50528 3596 50580 3602
rect 50528 3538 50580 3544
rect 50988 3596 51040 3602
rect 50988 3538 51040 3544
rect 51632 3596 51684 3602
rect 51632 3538 51684 3544
rect 52368 3596 52420 3602
rect 52368 3538 52420 3544
rect 52828 3596 52880 3602
rect 52828 3538 52880 3544
rect 53748 3596 53800 3602
rect 53748 3538 53800 3544
rect 50344 2916 50396 2922
rect 50344 2858 50396 2864
rect 50540 480 50568 3538
rect 51644 480 51672 3538
rect 52840 480 52868 3538
rect 54036 480 54064 3606
rect 55220 3392 55272 3398
rect 55220 3334 55272 3340
rect 55232 480 55260 3334
rect 56428 480 56456 326402
rect 56520 3398 56548 333202
rect 67548 322244 67600 322250
rect 67548 322186 67600 322192
rect 64788 10736 64840 10742
rect 64788 10678 64840 10684
rect 60648 10668 60700 10674
rect 60648 10610 60700 10616
rect 58808 9036 58860 9042
rect 58808 8978 58860 8984
rect 57612 3732 57664 3738
rect 57612 3674 57664 3680
rect 56508 3392 56560 3398
rect 56508 3334 56560 3340
rect 57624 480 57652 3674
rect 58820 480 58848 8978
rect 60660 3398 60688 10610
rect 62396 9104 62448 9110
rect 62396 9046 62448 9052
rect 61200 3800 61252 3806
rect 61200 3742 61252 3748
rect 60004 3392 60056 3398
rect 60004 3334 60056 3340
rect 60648 3392 60700 3398
rect 60648 3334 60700 3340
rect 60016 480 60044 3334
rect 61212 480 61240 3742
rect 62408 480 62436 9046
rect 64696 3868 64748 3874
rect 64696 3810 64748 3816
rect 63592 3392 63644 3398
rect 63592 3334 63644 3340
rect 63604 480 63632 3334
rect 64708 1986 64736 3810
rect 64800 3398 64828 10678
rect 65984 9172 66036 9178
rect 65984 9114 66036 9120
rect 64788 3392 64840 3398
rect 64788 3334 64840 3340
rect 64708 1958 64828 1986
rect 64800 480 64828 1958
rect 65996 480 66024 9114
rect 67560 626 67588 322186
rect 69480 9240 69532 9246
rect 69480 9182 69532 9188
rect 68284 3936 68336 3942
rect 68284 3878 68336 3884
rect 67192 598 67588 626
rect 67192 480 67220 598
rect 68296 480 68324 3878
rect 69492 480 69520 9182
rect 71700 3398 71728 336058
rect 74448 334688 74500 334694
rect 74448 334630 74500 334636
rect 73068 9308 73120 9314
rect 73068 9250 73120 9256
rect 71872 4004 71924 4010
rect 71872 3946 71924 3952
rect 70676 3392 70728 3398
rect 70676 3334 70728 3340
rect 71688 3392 71740 3398
rect 71688 3334 71740 3340
rect 70688 480 70716 3334
rect 71884 480 71912 3946
rect 73080 480 73108 9250
rect 74460 610 74488 334630
rect 92388 333328 92440 333334
rect 92388 333270 92440 333276
rect 89628 331968 89680 331974
rect 89628 331910 89680 331916
rect 78588 330608 78640 330614
rect 78588 330550 78640 330556
rect 76656 9376 76708 9382
rect 76656 9318 76708 9324
rect 75460 3188 75512 3194
rect 75460 3130 75512 3136
rect 74264 604 74316 610
rect 74264 546 74316 552
rect 74448 604 74500 610
rect 74448 546 74500 552
rect 74276 480 74304 546
rect 75472 480 75500 3130
rect 76668 480 76696 9318
rect 78600 3398 78628 330550
rect 85488 329180 85540 329186
rect 85488 329122 85540 329128
rect 82728 320884 82780 320890
rect 82728 320826 82780 320832
rect 80244 9444 80296 9450
rect 80244 9386 80296 9392
rect 79048 4140 79100 4146
rect 79048 4082 79100 4088
rect 77852 3392 77904 3398
rect 77852 3334 77904 3340
rect 78588 3392 78640 3398
rect 78588 3334 78640 3340
rect 77864 480 77892 3334
rect 79060 480 79088 4082
rect 80256 480 80284 9386
rect 82740 3398 82768 320826
rect 83832 9512 83884 9518
rect 83832 9454 83884 9460
rect 81440 3392 81492 3398
rect 81440 3334 81492 3340
rect 82728 3392 82780 3398
rect 82728 3334 82780 3340
rect 81452 480 81480 3334
rect 82636 3256 82688 3262
rect 82636 3198 82688 3204
rect 82648 480 82676 3198
rect 83844 480 83872 9454
rect 84108 4072 84160 4078
rect 84108 4014 84160 4020
rect 84120 3194 84148 4014
rect 85500 3330 85528 329122
rect 87328 9580 87380 9586
rect 87328 9522 87380 9528
rect 84936 3324 84988 3330
rect 84936 3266 84988 3272
rect 85488 3324 85540 3330
rect 85488 3266 85540 3272
rect 84108 3188 84160 3194
rect 84108 3130 84160 3136
rect 84948 480 84976 3266
rect 86132 3256 86184 3262
rect 86132 3198 86184 3204
rect 86144 480 86172 3198
rect 87340 480 87368 9522
rect 89640 3194 89668 331910
rect 90916 9648 90968 9654
rect 90916 9590 90968 9596
rect 89720 3256 89772 3262
rect 89720 3198 89772 3204
rect 88524 3188 88576 3194
rect 88524 3130 88576 3136
rect 89628 3188 89680 3194
rect 89628 3130 89680 3136
rect 88536 480 88564 3130
rect 89732 480 89760 3198
rect 90928 480 90956 9590
rect 92400 610 92428 333270
rect 96528 327820 96580 327826
rect 96528 327762 96580 327768
rect 94504 8900 94556 8906
rect 94504 8842 94556 8848
rect 93308 3188 93360 3194
rect 93308 3130 93360 3136
rect 92112 604 92164 610
rect 92112 546 92164 552
rect 92388 604 92440 610
rect 92388 546 92440 552
rect 92124 480 92152 546
rect 93320 480 93348 3130
rect 94516 480 94544 8842
rect 96540 3126 96568 327762
rect 99288 318164 99340 318170
rect 99288 318106 99340 318112
rect 98092 8832 98144 8838
rect 98092 8774 98144 8780
rect 95700 3120 95752 3126
rect 95700 3062 95752 3068
rect 96528 3120 96580 3126
rect 96528 3062 96580 3068
rect 95712 480 95740 3062
rect 96896 3052 96948 3058
rect 96896 2994 96948 3000
rect 96908 480 96936 2994
rect 98104 480 98132 8774
rect 99300 480 99328 318106
rect 100680 4842 100708 337826
rect 103428 325032 103480 325038
rect 103428 324974 103480 324980
rect 101588 8764 101640 8770
rect 101588 8706 101640 8712
rect 100496 4814 100708 4842
rect 100496 480 100524 4814
rect 101600 480 101628 8706
rect 103440 3126 103468 324974
rect 107476 309800 107528 309806
rect 107476 309742 107528 309748
rect 105176 8696 105228 8702
rect 105176 8638 105228 8644
rect 102784 3120 102836 3126
rect 102784 3062 102836 3068
rect 103428 3120 103480 3126
rect 103428 3062 103480 3068
rect 102796 480 102824 3062
rect 103980 2916 104032 2922
rect 103980 2858 104032 2864
rect 103992 480 104020 2858
rect 105188 480 105216 8638
rect 107488 3126 107516 309742
rect 106372 3120 106424 3126
rect 106372 3062 106424 3068
rect 107476 3120 107528 3126
rect 107476 3062 107528 3068
rect 106384 480 106412 3062
rect 107580 480 107608 337962
rect 115848 337952 115900 337958
rect 115848 337894 115900 337900
rect 114468 323672 114520 323678
rect 114468 323614 114520 323620
rect 110328 316736 110380 316742
rect 110328 316678 110380 316684
rect 108764 8628 108816 8634
rect 108764 8570 108816 8576
rect 108776 480 108804 8570
rect 110340 610 110368 316678
rect 112352 8560 112404 8566
rect 112352 8502 112404 8508
rect 111156 2916 111208 2922
rect 111156 2858 111208 2864
rect 109960 604 110012 610
rect 109960 546 110012 552
rect 110328 604 110380 610
rect 110328 546 110380 552
rect 109972 480 110000 546
rect 111168 480 111196 2858
rect 112364 480 112392 8502
rect 114480 2990 114508 323614
rect 113548 2984 113600 2990
rect 113548 2926 113600 2932
rect 114468 2984 114520 2990
rect 114468 2926 114520 2932
rect 113560 480 113588 2926
rect 115860 2922 115888 337894
rect 121368 322312 121420 322318
rect 121368 322254 121420 322260
rect 117228 17264 117280 17270
rect 117228 17206 117280 17212
rect 115940 8492 115992 8498
rect 115940 8434 115992 8440
rect 114744 2916 114796 2922
rect 114744 2858 114796 2864
rect 115848 2916 115900 2922
rect 115848 2858 115900 2864
rect 114756 480 114784 2858
rect 115952 480 115980 8434
rect 117240 4842 117268 17206
rect 119436 8424 119488 8430
rect 119436 8366 119488 8372
rect 117148 4814 117268 4842
rect 117148 480 117176 4814
rect 118240 2848 118292 2854
rect 118240 2790 118292 2796
rect 118252 480 118280 2790
rect 119448 480 119476 8366
rect 121380 2922 121408 322254
rect 125416 320952 125468 320958
rect 125416 320894 125468 320900
rect 123024 8356 123076 8362
rect 123024 8298 123076 8304
rect 120632 2916 120684 2922
rect 120632 2858 120684 2864
rect 121368 2916 121420 2922
rect 121368 2858 121420 2864
rect 120644 480 120672 2858
rect 121828 2848 121880 2854
rect 121828 2790 121880 2796
rect 121840 480 121868 2790
rect 123036 480 123064 8298
rect 125428 4214 125456 320894
rect 124220 4208 124272 4214
rect 124220 4150 124272 4156
rect 125416 4208 125468 4214
rect 125416 4150 125468 4156
rect 124232 480 124260 4150
rect 125520 3482 125548 338030
rect 126888 336184 126940 336190
rect 126888 336126 126940 336132
rect 126900 3482 126928 336126
rect 129648 333396 129700 333402
rect 129648 333338 129700 333344
rect 128268 330676 128320 330682
rect 128268 330618 128320 330624
rect 128280 3482 128308 330618
rect 129660 3482 129688 333338
rect 135916 8294 135944 398890
rect 200762 398304 200818 398313
rect 200762 398239 200818 398248
rect 198002 398168 198058 398177
rect 198002 398103 198058 398112
rect 180708 336320 180760 336326
rect 180708 336262 180760 336268
rect 169668 336252 169720 336258
rect 169668 336194 169720 336200
rect 162768 334824 162820 334830
rect 162768 334766 162820 334772
rect 160008 334756 160060 334762
rect 160008 334698 160060 334704
rect 142068 333464 142120 333470
rect 142068 333406 142120 333412
rect 139308 327888 139360 327894
rect 139308 327830 139360 327836
rect 136548 318232 136600 318238
rect 136548 318174 136600 318180
rect 135904 8288 135956 8294
rect 135904 8230 135956 8236
rect 132592 7608 132644 7614
rect 132592 7550 132644 7556
rect 131396 6248 131448 6254
rect 131396 6190 131448 6196
rect 130200 5092 130252 5098
rect 130200 5034 130252 5040
rect 125428 3454 125548 3482
rect 126624 3454 126928 3482
rect 127820 3454 128308 3482
rect 129016 3454 129688 3482
rect 125428 480 125456 3454
rect 126624 480 126652 3454
rect 127820 480 127848 3454
rect 129016 480 129044 3454
rect 130212 480 130240 5034
rect 131408 480 131436 6190
rect 132604 480 132632 7550
rect 134892 6316 134944 6322
rect 134892 6258 134944 6264
rect 133788 5160 133840 5166
rect 133788 5102 133840 5108
rect 133800 480 133828 5102
rect 134904 480 134932 6258
rect 136560 4842 136588 318174
rect 137284 5296 137336 5302
rect 137284 5238 137336 5244
rect 136100 4814 136588 4842
rect 136100 480 136128 4814
rect 137296 480 137324 5238
rect 139320 4842 139348 327830
rect 141976 325100 142028 325106
rect 141976 325042 142028 325048
rect 140688 316804 140740 316810
rect 140688 316746 140740 316752
rect 140700 4842 140728 316746
rect 140872 5228 140924 5234
rect 140872 5170 140924 5176
rect 138492 4814 139348 4842
rect 139688 4814 140728 4842
rect 138492 480 138520 4814
rect 139688 480 139716 4814
rect 140884 480 140912 5170
rect 141988 4842 142016 325042
rect 142080 5234 142108 333406
rect 153108 332104 153160 332110
rect 153108 332046 153160 332052
rect 144828 332036 144880 332042
rect 144828 331978 144880 331984
rect 143448 315376 143500 315382
rect 143448 315318 143500 315324
rect 142068 5228 142120 5234
rect 142068 5170 142120 5176
rect 141988 4814 142108 4842
rect 142080 480 142108 4814
rect 143460 3346 143488 315318
rect 144840 3346 144868 331978
rect 151728 330744 151780 330750
rect 151728 330686 151780 330692
rect 146208 322380 146260 322386
rect 146208 322322 146260 322328
rect 146220 3346 146248 322322
rect 150348 321020 150400 321026
rect 150348 320962 150400 320968
rect 147588 314016 147640 314022
rect 147588 313958 147640 313964
rect 147600 3346 147628 313958
rect 148968 13116 149020 13122
rect 148968 13058 149020 13064
rect 148980 3346 149008 13058
rect 150360 3346 150388 320962
rect 151636 15904 151688 15910
rect 151636 15846 151688 15852
rect 151648 4214 151676 15846
rect 150440 4208 150492 4214
rect 150440 4150 150492 4156
rect 151636 4208 151688 4214
rect 151636 4150 151688 4156
rect 143276 3318 143488 3346
rect 144472 3318 144868 3346
rect 145668 3318 146248 3346
rect 146864 3318 147628 3346
rect 148060 3318 149008 3346
rect 149256 3318 150388 3346
rect 143276 480 143304 3318
rect 144472 480 144500 3318
rect 145668 480 145696 3318
rect 146864 480 146892 3318
rect 148060 480 148088 3318
rect 149256 480 149284 3318
rect 150452 480 150480 4150
rect 151740 3482 151768 330686
rect 153120 3618 153148 332046
rect 157248 329316 157300 329322
rect 157248 329258 157300 329264
rect 155868 329248 155920 329254
rect 155868 329190 155920 329196
rect 154488 319524 154540 319530
rect 154488 319466 154540 319472
rect 154500 3618 154528 319466
rect 155880 3618 155908 329190
rect 157260 3618 157288 329258
rect 159916 326528 159968 326534
rect 159916 326470 159968 326476
rect 158628 312656 158680 312662
rect 158628 312598 158680 312604
rect 158640 3618 158668 312598
rect 158720 4208 158772 4214
rect 158720 4150 158772 4156
rect 151556 3454 151768 3482
rect 152752 3590 153148 3618
rect 153948 3590 154528 3618
rect 155144 3590 155908 3618
rect 156340 3590 157288 3618
rect 157536 3590 158668 3618
rect 151556 480 151584 3454
rect 152752 480 152780 3590
rect 153948 480 153976 3590
rect 155144 480 155172 3590
rect 156340 480 156368 3590
rect 157536 480 157564 3590
rect 158732 480 158760 4150
rect 159928 480 159956 326470
rect 160020 4214 160048 334698
rect 161388 311228 161440 311234
rect 161388 311170 161440 311176
rect 160008 4208 160060 4214
rect 160008 4150 160060 4156
rect 161400 3618 161428 311170
rect 161124 3590 161428 3618
rect 161124 480 161152 3590
rect 162780 3482 162808 334766
rect 168288 327956 168340 327962
rect 168288 327898 168340 327904
rect 165528 323740 165580 323746
rect 165528 323682 165580 323688
rect 164148 14476 164200 14482
rect 164148 14418 164200 14424
rect 164160 3482 164188 14418
rect 165540 3482 165568 323682
rect 166908 11756 166960 11762
rect 166908 11698 166960 11704
rect 166920 3482 166948 11698
rect 168196 7676 168248 7682
rect 168196 7618 168248 7624
rect 167092 4208 167144 4214
rect 167092 4150 167144 4156
rect 162320 3454 162808 3482
rect 163516 3454 164188 3482
rect 164712 3454 165568 3482
rect 165908 3454 166948 3482
rect 162320 480 162348 3454
rect 163516 480 163544 3454
rect 164712 480 164740 3454
rect 165908 480 165936 3454
rect 167104 480 167132 4150
rect 168208 480 168236 7618
rect 168300 4214 168328 327898
rect 168288 4208 168340 4214
rect 168288 4150 168340 4156
rect 169680 3482 169708 336194
rect 176568 334892 176620 334898
rect 176568 334834 176620 334840
rect 173808 333532 173860 333538
rect 173808 333474 173860 333480
rect 171048 326596 171100 326602
rect 171048 326538 171100 326544
rect 171060 3482 171088 326538
rect 171784 7744 171836 7750
rect 171784 7686 171836 7692
rect 169404 3454 169708 3482
rect 170600 3454 171088 3482
rect 169404 480 169432 3454
rect 170600 480 170628 3454
rect 171796 480 171824 7686
rect 173820 4842 173848 333474
rect 175372 7812 175424 7818
rect 175372 7754 175424 7760
rect 174176 6384 174228 6390
rect 174176 6326 174228 6332
rect 172992 4814 173848 4842
rect 172992 480 173020 4814
rect 174188 480 174216 6326
rect 175384 480 175412 7754
rect 176580 480 176608 334834
rect 178960 7880 179012 7886
rect 178960 7822 179012 7828
rect 177764 6452 177816 6458
rect 177764 6394 177816 6400
rect 177776 480 177804 6394
rect 178972 480 179000 7822
rect 180720 4842 180748 336262
rect 184848 332172 184900 332178
rect 184848 332114 184900 332120
rect 182548 7948 182600 7954
rect 182548 7890 182600 7896
rect 181352 6520 181404 6526
rect 181352 6462 181404 6468
rect 180168 4814 180748 4842
rect 180168 480 180196 4814
rect 181364 480 181392 6462
rect 182560 480 182588 7890
rect 184860 6746 184888 332114
rect 198016 64870 198044 398103
rect 198004 64864 198056 64870
rect 198004 64806 198056 64812
rect 200776 51066 200804 398239
rect 203536 93838 203564 400318
rect 204904 399152 204956 399158
rect 204904 399094 204956 399100
rect 204916 180810 204944 399094
rect 206928 329384 206980 329390
rect 206928 329326 206980 329332
rect 204904 180804 204956 180810
rect 204904 180746 204956 180752
rect 203524 93832 203576 93838
rect 203524 93774 203576 93780
rect 200764 51060 200816 51066
rect 200764 51002 200816 51008
rect 200396 8288 200448 8294
rect 200396 8230 200448 8236
rect 196808 8220 196860 8226
rect 196808 8162 196860 8168
rect 193220 8152 193272 8158
rect 193220 8094 193272 8100
rect 189632 8084 189684 8090
rect 189632 8026 189684 8032
rect 186044 8016 186096 8022
rect 186044 7958 186096 7964
rect 184768 6718 184888 6746
rect 184768 610 184796 6718
rect 184848 6588 184900 6594
rect 184848 6530 184900 6536
rect 183744 604 183796 610
rect 183744 546 183796 552
rect 184756 604 184808 610
rect 184756 546 184808 552
rect 183756 480 183784 546
rect 184860 480 184888 6530
rect 186056 480 186084 7958
rect 188436 6656 188488 6662
rect 188436 6598 188488 6604
rect 187240 5296 187292 5302
rect 187240 5238 187292 5244
rect 187252 480 187280 5238
rect 188448 480 188476 6598
rect 189644 480 189672 8026
rect 192024 6724 192076 6730
rect 192024 6666 192076 6672
rect 190828 5364 190880 5370
rect 190828 5306 190880 5312
rect 190840 480 190868 5306
rect 192036 480 192064 6666
rect 193232 480 193260 8094
rect 195612 6792 195664 6798
rect 195612 6734 195664 6740
rect 194416 5432 194468 5438
rect 194416 5374 194468 5380
rect 194428 480 194456 5374
rect 195624 480 195652 6734
rect 196820 480 196848 8162
rect 199200 6860 199252 6866
rect 199200 6802 199252 6808
rect 198004 5500 198056 5506
rect 198004 5442 198056 5448
rect 198016 480 198044 5442
rect 199212 480 199240 6802
rect 200408 480 200436 8230
rect 203892 7540 203944 7546
rect 203892 7482 203944 7488
rect 202696 6112 202748 6118
rect 202696 6054 202748 6060
rect 201500 4752 201552 4758
rect 201500 4694 201552 4700
rect 201512 480 201540 4694
rect 202708 480 202736 6054
rect 203904 480 203932 7482
rect 205088 4684 205140 4690
rect 205088 4626 205140 4632
rect 205100 480 205128 4626
rect 206940 610 206968 329326
rect 207676 223582 207704 400522
rect 209044 399356 209096 399362
rect 209044 399298 209096 399304
rect 208308 330812 208360 330818
rect 208308 330754 208360 330760
rect 207664 223576 207716 223582
rect 207664 223518 207716 223524
rect 208320 610 208348 330754
rect 209056 266354 209084 399298
rect 209688 336388 209740 336394
rect 209688 336330 209740 336336
rect 209044 266348 209096 266354
rect 209044 266290 209096 266296
rect 209700 610 209728 336330
rect 211068 332240 211120 332246
rect 211068 332182 211120 332188
rect 210976 319592 211028 319598
rect 210976 319534 211028 319540
rect 209872 4208 209924 4214
rect 209872 4150 209924 4156
rect 206284 604 206336 610
rect 206284 546 206336 552
rect 206928 604 206980 610
rect 206928 546 206980 552
rect 207480 604 207532 610
rect 207480 546 207532 552
rect 208308 604 208360 610
rect 208308 546 208360 552
rect 208676 604 208728 610
rect 208676 546 208728 552
rect 209688 604 209740 610
rect 209688 546 209740 552
rect 206296 480 206324 546
rect 207492 480 207520 546
rect 208688 480 208716 546
rect 209884 480 209912 4150
rect 210988 3482 211016 319534
rect 211080 4214 211108 332182
rect 211816 309126 211844 400658
rect 214564 400648 214616 400654
rect 214564 400590 214616 400596
rect 213184 399220 213236 399226
rect 213184 399162 213236 399168
rect 212448 334960 212500 334966
rect 212448 334902 212500 334908
rect 211804 309120 211856 309126
rect 211804 309062 211856 309068
rect 211068 4208 211120 4214
rect 211068 4150 211120 4156
rect 212460 3618 212488 334902
rect 213196 35902 213224 399162
rect 213828 325168 213880 325174
rect 213828 325110 213880 325116
rect 213184 35896 213236 35902
rect 213184 35838 213236 35844
rect 213840 3618 213868 325110
rect 214576 80034 214604 400590
rect 215944 399424 215996 399430
rect 215944 399366 215996 399372
rect 215208 328024 215260 328030
rect 215208 327966 215260 327972
rect 214564 80028 214616 80034
rect 214564 79970 214616 79976
rect 215220 3618 215248 327966
rect 215956 122806 215984 399366
rect 216588 333600 216640 333606
rect 216588 333542 216640 333548
rect 215944 122800 215996 122806
rect 215944 122742 215996 122748
rect 216600 3618 216628 333542
rect 217968 323808 218020 323814
rect 217968 323750 218020 323756
rect 217980 3618 218008 323750
rect 218716 165578 218744 400726
rect 222936 399764 222988 399770
rect 222936 399706 222988 399712
rect 222844 337272 222896 337278
rect 222844 337214 222896 337220
rect 219348 336456 219400 336462
rect 219348 336398 219400 336404
rect 218704 165572 218756 165578
rect 218704 165514 218756 165520
rect 219256 164892 219308 164898
rect 219256 164834 219308 164840
rect 219268 3618 219296 164834
rect 212276 3590 212488 3618
rect 213472 3590 213868 3618
rect 214668 3590 215248 3618
rect 215864 3590 216628 3618
rect 217060 3590 218008 3618
rect 218164 3590 219296 3618
rect 210988 3454 211108 3482
rect 211080 480 211108 3454
rect 212276 480 212304 3590
rect 213472 480 213500 3590
rect 214668 480 214696 3590
rect 215864 480 215892 3590
rect 217060 480 217088 3590
rect 218164 480 218192 3590
rect 219360 480 219388 336398
rect 220728 333668 220780 333674
rect 220728 333610 220780 333616
rect 220740 3346 220768 333610
rect 222108 326664 222160 326670
rect 222108 326606 222160 326612
rect 222120 3346 222148 326606
rect 222856 17270 222884 337214
rect 222948 208350 222976 399706
rect 225604 399560 225656 399566
rect 225604 399502 225656 399508
rect 224868 335096 224920 335102
rect 224868 335038 224920 335044
rect 223488 335028 223540 335034
rect 223488 334970 223540 334976
rect 222936 208344 222988 208350
rect 222936 208286 222988 208292
rect 222844 17264 222896 17270
rect 222844 17206 222896 17212
rect 223500 3346 223528 334970
rect 224880 3346 224908 335038
rect 225616 22098 225644 399502
rect 225694 398712 225750 398721
rect 225694 398647 225750 398656
rect 225708 380866 225736 398647
rect 225696 380860 225748 380866
rect 225696 380802 225748 380808
rect 225696 337204 225748 337210
rect 225696 337146 225748 337152
rect 225604 22092 225656 22098
rect 225604 22034 225656 22040
rect 225708 13122 225736 337146
rect 225800 252550 225828 401066
rect 226996 367062 227024 401202
rect 227076 401056 227128 401062
rect 227076 400998 227128 401004
rect 226984 367056 227036 367062
rect 226984 366998 227036 367004
rect 226984 337340 227036 337346
rect 226984 337282 227036 337288
rect 226248 322448 226300 322454
rect 226248 322390 226300 322396
rect 225788 252544 225840 252550
rect 225788 252486 225840 252492
rect 225696 13116 225748 13122
rect 225696 13058 225748 13064
rect 226260 3874 226288 322390
rect 226996 11762 227024 337282
rect 227088 151774 227116 400998
rect 234896 400988 234948 400994
rect 234896 400930 234948 400936
rect 231768 400920 231820 400926
rect 231768 400862 231820 400868
rect 230664 400512 230716 400518
rect 230664 400454 230716 400460
rect 230676 399908 230704 400454
rect 231780 399908 231808 400862
rect 234908 399908 234936 400930
rect 235448 400444 235500 400450
rect 235448 400386 235500 400392
rect 235460 399908 235488 400386
rect 235920 399908 235948 401882
rect 238024 400852 238076 400858
rect 238024 400794 238076 400800
rect 237564 400308 237616 400314
rect 237564 400250 237616 400256
rect 237576 399908 237604 400250
rect 238036 399908 238064 400794
rect 239140 399908 239168 401882
rect 240140 400240 240192 400246
rect 240140 400182 240192 400188
rect 240152 399908 240180 400182
rect 240704 399908 240732 402086
rect 243268 401872 243320 401878
rect 243268 401814 243320 401820
rect 241244 401192 241296 401198
rect 241244 401134 241296 401140
rect 241256 399908 241284 401134
rect 241730 399906 242112 399922
rect 242834 399906 242940 399922
rect 243280 399908 243308 401814
rect 243832 399908 243860 404330
rect 244200 401878 244228 415414
rect 244924 401940 244976 401946
rect 244924 401882 244976 401888
rect 244188 401872 244240 401878
rect 244188 401814 244240 401820
rect 244372 401872 244424 401878
rect 244372 401814 244424 401820
rect 244384 399908 244412 401814
rect 244936 399908 244964 401882
rect 245396 401878 245424 438874
rect 245384 401872 245436 401878
rect 245384 401814 245436 401820
rect 245488 399922 245516 451250
rect 245580 401946 245608 462334
rect 245568 401940 245620 401946
rect 245568 401882 245620 401888
rect 246868 401878 246896 485794
rect 245936 401872 245988 401878
rect 245936 401814 245988 401820
rect 246856 401872 246908 401878
rect 246856 401814 246908 401820
rect 241730 399900 242124 399906
rect 241730 399894 242072 399900
rect 242834 399900 242952 399906
rect 242834 399894 242900 399900
rect 242072 399842 242124 399848
rect 245410 399894 245516 399922
rect 245948 399908 245976 401814
rect 246960 399922 246988 509254
rect 248144 498228 248196 498234
rect 248144 498170 248196 498176
rect 248156 401946 248184 498170
rect 247040 401940 247092 401946
rect 247040 401882 247092 401888
rect 248144 401940 248196 401946
rect 248144 401882 248196 401888
rect 246514 399894 246988 399922
rect 247052 399908 247080 401882
rect 248248 400058 248276 532714
rect 247880 400030 248276 400058
rect 247880 399922 247908 400030
rect 248340 399922 248368 556174
rect 249524 545148 249576 545154
rect 249524 545090 249576 545096
rect 249536 402150 249564 545090
rect 248604 402144 248656 402150
rect 248604 402086 248656 402092
rect 249524 402144 249576 402150
rect 249524 402086 249576 402092
rect 247526 399894 247908 399922
rect 248078 399894 248368 399922
rect 248616 399908 248644 402086
rect 249628 400330 249656 579634
rect 249536 400302 249656 400330
rect 249536 399922 249564 400302
rect 249720 399922 249748 603094
rect 250996 592068 251048 592074
rect 250996 592010 251048 592016
rect 251008 402150 251036 592010
rect 250168 402144 250220 402150
rect 250168 402086 250220 402092
rect 250996 402144 251048 402150
rect 250996 402086 251048 402092
rect 249090 399894 249564 399922
rect 249642 399894 249748 399922
rect 250180 399908 250208 402086
rect 251100 399922 251128 626554
rect 251180 402144 251232 402150
rect 251180 402086 251232 402092
rect 250746 399894 251128 399922
rect 251192 399908 251220 402086
rect 252296 400330 252324 638930
rect 252388 402150 252416 650014
rect 252376 402144 252428 402150
rect 252376 402086 252428 402092
rect 252204 400302 252324 400330
rect 242900 399842 242952 399848
rect 227168 399832 227220 399838
rect 252204 399786 252232 400302
rect 252480 399922 252508 673474
rect 252744 402144 252796 402150
rect 252744 402086 252796 402092
rect 252310 399894 252508 399922
rect 252756 399908 252784 402086
rect 253676 399922 253704 685850
rect 253768 402150 253796 696934
rect 253756 402144 253808 402150
rect 253756 402086 253808 402092
rect 253322 399894 253704 399922
rect 253860 399908 253888 700266
rect 254400 402144 254452 402150
rect 254400 402086 254452 402092
rect 254412 399908 254440 402086
rect 255148 399922 255176 700334
rect 255240 402150 255268 700402
rect 255228 402144 255280 402150
rect 255228 402086 255280 402092
rect 255412 402144 255464 402150
rect 255412 402086 255464 402092
rect 254886 399894 255176 399922
rect 255424 399908 255452 402086
rect 256436 400330 256464 700674
rect 256516 700664 256568 700670
rect 256516 700606 256568 700612
rect 256160 400302 256464 400330
rect 256160 399922 256188 400302
rect 256528 399922 256556 700606
rect 256608 700596 256660 700602
rect 256608 700538 256660 700544
rect 256620 402150 256648 700538
rect 256608 402144 256660 402150
rect 256608 402086 256660 402092
rect 256976 402144 257028 402150
rect 256976 402086 257028 402092
rect 255990 399894 256188 399922
rect 256450 399894 256556 399922
rect 256988 399908 257016 402086
rect 257908 399922 257936 700946
rect 259276 700936 259328 700942
rect 259276 700878 259328 700884
rect 257988 700868 258040 700874
rect 257988 700810 258040 700816
rect 258000 402150 258028 700810
rect 259184 700052 259236 700058
rect 259184 699994 259236 700000
rect 258448 407788 258500 407794
rect 258448 407730 258500 407736
rect 258080 402620 258132 402626
rect 258080 402562 258132 402568
rect 258092 402529 258120 402562
rect 258078 402520 258134 402529
rect 258078 402455 258134 402464
rect 257988 402144 258040 402150
rect 257988 402086 258040 402092
rect 258460 399922 258488 407730
rect 258540 402076 258592 402082
rect 258540 402018 258592 402024
rect 257554 399894 257936 399922
rect 258106 399894 258488 399922
rect 258552 399908 258580 402018
rect 259196 399922 259224 699994
rect 259288 407794 259316 700878
rect 265072 700800 265124 700806
rect 265072 700742 265124 700748
rect 263784 700256 263836 700262
rect 263784 700198 263836 700204
rect 259368 700188 259420 700194
rect 259368 700130 259420 700136
rect 259276 407788 259328 407794
rect 259276 407730 259328 407736
rect 259380 402082 259408 700130
rect 260656 700120 260708 700126
rect 260656 700062 260708 700068
rect 260196 402620 260248 402626
rect 260196 402562 260248 402568
rect 259368 402076 259420 402082
rect 259368 402018 259420 402024
rect 259644 402076 259696 402082
rect 259644 402018 259696 402024
rect 259118 399894 259224 399922
rect 259656 399908 259684 402018
rect 260208 399908 260236 402562
rect 260668 402082 260696 700062
rect 262220 699984 262272 699990
rect 262220 699926 262272 699932
rect 262128 699916 262180 699922
rect 262128 699858 262180 699864
rect 260748 699712 260800 699718
rect 260748 699654 260800 699660
rect 260656 402076 260708 402082
rect 260656 402018 260708 402024
rect 260760 399922 260788 699654
rect 261206 402520 261262 402529
rect 261206 402455 261208 402464
rect 261260 402455 261262 402464
rect 261208 402426 261260 402432
rect 261760 402144 261812 402150
rect 261760 402086 261812 402092
rect 261208 402076 261260 402082
rect 261208 402018 261260 402024
rect 260682 399894 260788 399922
rect 261220 399908 261248 402018
rect 261772 399908 261800 402086
rect 262140 402082 262168 699858
rect 262128 402076 262180 402082
rect 262128 402018 262180 402024
rect 262232 399908 262260 699926
rect 262864 667956 262916 667962
rect 262864 667898 262916 667904
rect 262876 402778 262904 667898
rect 263324 402960 263376 402966
rect 263324 402902 263376 402908
rect 262876 402750 262996 402778
rect 262968 402490 262996 402750
rect 262956 402484 263008 402490
rect 262956 402426 263008 402432
rect 262772 402212 262824 402218
rect 262772 402154 262824 402160
rect 262784 399908 262812 402154
rect 263336 399908 263364 402902
rect 263796 399922 263824 700198
rect 264244 610020 264296 610026
rect 264244 609962 264296 609968
rect 264256 402830 264284 609962
rect 264336 402892 264388 402898
rect 264336 402834 264388 402840
rect 264244 402824 264296 402830
rect 264244 402766 264296 402772
rect 263796 399894 263902 399922
rect 264348 399908 264376 402834
rect 264888 402756 264940 402762
rect 264888 402698 264940 402704
rect 264900 399908 264928 402698
rect 265084 399922 265112 700742
rect 266544 700528 266596 700534
rect 266544 700470 266596 700476
rect 265624 552084 265676 552090
rect 265624 552026 265676 552032
rect 265636 402762 265664 552026
rect 265624 402756 265676 402762
rect 265624 402698 265676 402704
rect 265900 402688 265952 402694
rect 265900 402630 265952 402636
rect 265084 399894 265466 399922
rect 265912 399908 265940 402630
rect 266452 402620 266504 402626
rect 266452 402562 266504 402568
rect 266464 399908 266492 402562
rect 266556 399922 266584 700470
rect 267660 699718 267688 703520
rect 283852 699922 283880 703520
rect 283840 699916 283892 699922
rect 283840 699858 283892 699864
rect 267648 699712 267700 699718
rect 267648 699654 267700 699660
rect 300136 688634 300164 703520
rect 332520 700058 332548 703520
rect 348804 700126 348832 703520
rect 364996 700194 365024 703520
rect 397472 701010 397500 703520
rect 397460 701004 397512 701010
rect 397460 700946 397512 700952
rect 413664 700942 413692 703520
rect 413652 700936 413704 700942
rect 413652 700878 413704 700884
rect 429856 700874 429884 703520
rect 429844 700868 429896 700874
rect 429844 700810 429896 700816
rect 462332 700738 462360 703520
rect 462320 700732 462372 700738
rect 462320 700674 462372 700680
rect 478524 700670 478552 703520
rect 478512 700664 478564 700670
rect 478512 700606 478564 700612
rect 494808 700602 494836 703520
rect 494796 700596 494848 700602
rect 494796 700538 494848 700544
rect 527192 700466 527220 703520
rect 527180 700460 527232 700466
rect 527180 700402 527232 700408
rect 543476 700398 543504 703520
rect 543464 700392 543516 700398
rect 543464 700334 543516 700340
rect 559668 700330 559696 703520
rect 559656 700324 559708 700330
rect 559656 700266 559708 700272
rect 364984 700188 365036 700194
rect 364984 700130 365036 700136
rect 348792 700120 348844 700126
rect 348792 700062 348844 700068
rect 332508 700052 332560 700058
rect 332508 699994 332560 700000
rect 580170 698048 580226 698057
rect 580170 697983 580226 697992
rect 580184 696998 580212 697983
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 299664 688628 299716 688634
rect 299664 688570 299716 688576
rect 300124 688628 300176 688634
rect 300124 688570 300176 688576
rect 299676 685930 299704 688570
rect 580170 686352 580226 686361
rect 580170 686287 580226 686296
rect 299584 685902 299704 685930
rect 580184 685914 580212 686287
rect 580172 685908 580224 685914
rect 299584 684486 299612 685902
rect 580172 685850 580224 685856
rect 299572 684480 299624 684486
rect 299572 684422 299624 684428
rect 580170 674656 580226 674665
rect 580170 674591 580226 674600
rect 580184 673538 580212 674591
rect 580172 673532 580224 673538
rect 580172 673474 580224 673480
rect 299940 666596 299992 666602
rect 299940 666538 299992 666544
rect 299952 659682 299980 666538
rect 299768 659654 299980 659682
rect 267832 652792 267884 652798
rect 267832 652734 267884 652740
rect 267004 495508 267056 495514
rect 267004 495450 267056 495456
rect 267016 402626 267044 495450
rect 267004 402620 267056 402626
rect 267004 402562 267056 402568
rect 267556 402552 267608 402558
rect 267556 402494 267608 402500
rect 266556 399894 267030 399922
rect 267568 399908 267596 402494
rect 267844 402234 267872 652734
rect 299768 647290 299796 659654
rect 580170 651128 580226 651137
rect 580170 651063 580226 651072
rect 580184 650078 580212 651063
rect 580172 650072 580224 650078
rect 580172 650014 580224 650020
rect 299664 647284 299716 647290
rect 299664 647226 299716 647232
rect 299756 647284 299808 647290
rect 299756 647226 299808 647232
rect 299676 640422 299704 647226
rect 299664 640416 299716 640422
rect 299664 640358 299716 640364
rect 299756 640416 299808 640422
rect 299756 640358 299808 640364
rect 299768 630698 299796 640358
rect 580170 639432 580226 639441
rect 580170 639367 580226 639376
rect 580184 638994 580212 639367
rect 580172 638988 580224 638994
rect 580172 638930 580224 638936
rect 299572 630692 299624 630698
rect 299572 630634 299624 630640
rect 299756 630692 299808 630698
rect 299756 630634 299808 630640
rect 299584 630578 299612 630634
rect 299584 630550 299704 630578
rect 299676 621058 299704 630550
rect 580170 627736 580226 627745
rect 580170 627671 580226 627680
rect 580184 626618 580212 627671
rect 580172 626612 580224 626618
rect 580172 626554 580224 626560
rect 299676 621030 299796 621058
rect 299768 611386 299796 621030
rect 299572 611380 299624 611386
rect 299572 611322 299624 611328
rect 299756 611380 299808 611386
rect 299756 611322 299808 611328
rect 299584 611266 299612 611322
rect 299584 611238 299704 611266
rect 299676 608598 299704 611238
rect 299664 608592 299716 608598
rect 299664 608534 299716 608540
rect 580170 604208 580226 604217
rect 580170 604143 580226 604152
rect 580184 603158 580212 604143
rect 580172 603152 580224 603158
rect 580172 603094 580224 603100
rect 299848 601724 299900 601730
rect 299848 601666 299900 601672
rect 299860 598942 299888 601666
rect 299848 598936 299900 598942
rect 299848 598878 299900 598884
rect 269304 594856 269356 594862
rect 269304 594798 269356 594804
rect 269212 402960 269264 402966
rect 269212 402902 269264 402908
rect 269120 402484 269172 402490
rect 269120 402426 269172 402432
rect 267844 402206 268148 402234
rect 268016 402076 268068 402082
rect 268016 402018 268068 402024
rect 268028 399908 268056 402018
rect 227168 399774 227220 399780
rect 227180 295322 227208 399774
rect 251758 399758 252232 399786
rect 268120 399786 268148 402206
rect 269132 399908 269160 402426
rect 269224 399922 269252 402902
rect 269316 400058 269344 594798
rect 580170 592512 580226 592521
rect 580170 592447 580226 592456
rect 580184 592074 580212 592447
rect 580172 592068 580224 592074
rect 580172 592010 580224 592016
rect 299940 589348 299992 589354
rect 299940 589290 299992 589296
rect 299952 582486 299980 589290
rect 299940 582480 299992 582486
rect 299940 582422 299992 582428
rect 299848 582344 299900 582350
rect 299848 582286 299900 582292
rect 299860 572642 299888 582286
rect 580170 580816 580226 580825
rect 580170 580751 580226 580760
rect 580184 579698 580212 580751
rect 580172 579692 580224 579698
rect 580172 579634 580224 579640
rect 299676 572614 299888 572642
rect 299676 569922 299704 572614
rect 299584 569894 299704 569922
rect 299584 563174 299612 569894
rect 299572 563168 299624 563174
rect 299572 563110 299624 563116
rect 299572 563032 299624 563038
rect 299572 562974 299624 562980
rect 299584 560561 299612 562974
rect 299570 560552 299626 560561
rect 299570 560487 299626 560496
rect 299570 560416 299626 560425
rect 299570 560351 299626 560360
rect 299584 553518 299612 560351
rect 580170 557288 580226 557297
rect 580170 557223 580226 557232
rect 580184 556238 580212 557223
rect 580172 556232 580224 556238
rect 580172 556174 580224 556180
rect 299572 553512 299624 553518
rect 299572 553454 299624 553460
rect 299480 553376 299532 553382
rect 299480 553318 299532 553324
rect 299492 549273 299520 553318
rect 299294 549264 299350 549273
rect 299294 549199 299350 549208
rect 299478 549264 299534 549273
rect 299478 549199 299534 549208
rect 299308 543726 299336 549199
rect 580170 545592 580226 545601
rect 580170 545527 580226 545536
rect 580184 545154 580212 545527
rect 580172 545148 580224 545154
rect 580172 545090 580224 545096
rect 299296 543720 299348 543726
rect 299296 543662 299348 543668
rect 299480 543720 299532 543726
rect 299480 543662 299532 543668
rect 299492 539594 299520 543662
rect 299492 539566 299612 539594
rect 270776 538280 270828 538286
rect 270776 538222 270828 538228
rect 269764 437504 269816 437510
rect 269764 437446 269816 437452
rect 269776 402218 269804 437446
rect 270684 402824 270736 402830
rect 270684 402766 270736 402772
rect 269764 402212 269816 402218
rect 269764 402154 269816 402160
rect 269316 400030 269896 400058
rect 269868 399922 269896 400030
rect 269224 399894 269606 399922
rect 269868 399894 270158 399922
rect 270696 399908 270724 402766
rect 270788 402506 270816 538222
rect 299584 531350 299612 539566
rect 580170 533896 580226 533905
rect 580170 533831 580226 533840
rect 580184 532778 580212 533831
rect 580172 532772 580224 532778
rect 580172 532714 580224 532720
rect 299572 531344 299624 531350
rect 299572 531286 299624 531292
rect 299756 531344 299808 531350
rect 299756 531286 299808 531292
rect 299768 524482 299796 531286
rect 299756 524476 299808 524482
rect 299756 524418 299808 524424
rect 299848 524408 299900 524414
rect 299848 524350 299900 524356
rect 299860 521665 299888 524350
rect 299662 521656 299718 521665
rect 299662 521591 299718 521600
rect 299846 521656 299902 521665
rect 299846 521591 299902 521600
rect 299676 512038 299704 521591
rect 299664 512032 299716 512038
rect 299664 511974 299716 511980
rect 299940 512032 299992 512038
rect 299940 511974 299992 511980
rect 299952 502382 299980 511974
rect 580170 510368 580226 510377
rect 580170 510303 580226 510312
rect 580184 509318 580212 510303
rect 580172 509312 580224 509318
rect 580172 509254 580224 509260
rect 299756 502376 299808 502382
rect 299478 502344 299534 502353
rect 299478 502279 299534 502288
rect 299754 502344 299756 502353
rect 299940 502376 299992 502382
rect 299808 502344 299810 502353
rect 299940 502318 299992 502324
rect 299754 502279 299810 502288
rect 299492 492697 299520 502279
rect 580170 498672 580226 498681
rect 580170 498607 580226 498616
rect 580184 498234 580212 498607
rect 580172 498228 580224 498234
rect 580172 498170 580224 498176
rect 299478 492688 299534 492697
rect 299478 492623 299534 492632
rect 299662 492688 299718 492697
rect 299662 492623 299664 492632
rect 299716 492623 299718 492632
rect 299664 492594 299716 492600
rect 580170 486840 580226 486849
rect 580170 486775 580226 486784
rect 580184 485858 580212 486775
rect 580172 485852 580224 485858
rect 580172 485794 580224 485800
rect 299664 485784 299716 485790
rect 299664 485726 299716 485732
rect 299676 483018 299704 485726
rect 299676 482990 299796 483018
rect 272524 480276 272576 480282
rect 272524 480218 272576 480224
rect 272248 402756 272300 402762
rect 272248 402698 272300 402704
rect 270788 402478 271552 402506
rect 271236 402416 271288 402422
rect 271236 402358 271288 402364
rect 271248 399908 271276 402358
rect 271524 399922 271552 402478
rect 271524 399894 271722 399922
rect 272260 399908 272288 402698
rect 272536 402082 272564 480218
rect 299768 476134 299796 482990
rect 299572 476128 299624 476134
rect 299756 476128 299808 476134
rect 299624 476076 299704 476082
rect 299572 476070 299704 476076
rect 299756 476070 299808 476076
rect 299584 476054 299704 476070
rect 299676 473346 299704 476054
rect 299664 473340 299716 473346
rect 299664 473282 299716 473288
rect 299664 466404 299716 466410
rect 299664 466346 299716 466352
rect 299676 463706 299704 466346
rect 299676 463678 299796 463706
rect 299768 460902 299796 463678
rect 580170 463448 580226 463457
rect 580170 463383 580226 463392
rect 580184 462398 580212 463383
rect 580172 462392 580224 462398
rect 580172 462334 580224 462340
rect 299388 460896 299440 460902
rect 299388 460838 299440 460844
rect 299756 460896 299808 460902
rect 299756 460838 299808 460844
rect 299400 451330 299428 460838
rect 580170 451752 580226 451761
rect 580170 451687 580226 451696
rect 299400 451302 299520 451330
rect 580184 451314 580212 451687
rect 299492 449886 299520 451302
rect 580172 451308 580224 451314
rect 580172 451250 580224 451256
rect 299480 449880 299532 449886
rect 299480 449822 299532 449828
rect 299572 440292 299624 440298
rect 299572 440234 299624 440240
rect 299584 436830 299612 440234
rect 580170 439920 580226 439929
rect 580170 439855 580226 439864
rect 580184 438938 580212 439855
rect 580172 438932 580224 438938
rect 580172 438874 580224 438880
rect 299572 436824 299624 436830
rect 299572 436766 299624 436772
rect 299572 427780 299624 427786
rect 299572 427722 299624 427728
rect 273904 423700 273956 423706
rect 273904 423642 273956 423648
rect 273812 402620 273864 402626
rect 273812 402562 273864 402568
rect 272800 402348 272852 402354
rect 272800 402290 272852 402296
rect 272524 402076 272576 402082
rect 272524 402018 272576 402024
rect 272812 399908 272840 402290
rect 273260 402076 273312 402082
rect 273260 402018 273312 402024
rect 273272 399908 273300 402018
rect 273824 399908 273852 402562
rect 273916 402082 273944 423642
rect 299584 418146 299612 427722
rect 299584 418118 299796 418146
rect 299768 415410 299796 418118
rect 580170 416528 580226 416537
rect 580170 416463 580226 416472
rect 580184 415478 580212 416463
rect 580172 415472 580224 415478
rect 580172 415414 580224 415420
rect 299756 415404 299808 415410
rect 299756 415346 299808 415352
rect 299664 405748 299716 405754
rect 299664 405690 299716 405696
rect 274364 402280 274416 402286
rect 274364 402222 274416 402228
rect 273904 402076 273956 402082
rect 273904 402018 273956 402024
rect 274376 399908 274404 402222
rect 275376 402212 275428 402218
rect 275376 402154 275428 402160
rect 274916 402076 274968 402082
rect 274916 402018 274968 402024
rect 274928 399908 274956 402018
rect 275388 399908 275416 402154
rect 299676 402150 299704 405690
rect 580170 404832 580226 404841
rect 580170 404767 580226 404776
rect 580184 404394 580212 404767
rect 580172 404388 580224 404394
rect 580172 404330 580224 404336
rect 299664 402144 299716 402150
rect 299664 402086 299716 402092
rect 493324 402008 493376 402014
rect 493324 401950 493376 401956
rect 278596 401804 278648 401810
rect 278596 401746 278648 401752
rect 277492 401328 277544 401334
rect 277492 401270 277544 401276
rect 276480 401260 276532 401266
rect 276480 401202 276532 401208
rect 275652 399968 275704 399974
rect 275704 399916 275954 399922
rect 275652 399910 275954 399916
rect 275664 399894 275954 399910
rect 276492 399908 276520 401202
rect 277504 399908 277532 401270
rect 278044 400716 278096 400722
rect 278044 400658 278096 400664
rect 278056 399908 278084 400658
rect 278608 399908 278636 401746
rect 280160 401736 280212 401742
rect 280160 401678 280212 401684
rect 280172 399908 280200 401678
rect 281724 401668 281776 401674
rect 281724 401610 281776 401616
rect 280712 401124 280764 401130
rect 280712 401066 280764 401072
rect 280724 399908 280752 401066
rect 281172 400580 281224 400586
rect 281172 400522 281224 400528
rect 281184 399908 281212 400522
rect 281736 399908 281764 401610
rect 290464 401192 290516 401198
rect 290464 401134 290516 401140
rect 284852 401056 284904 401062
rect 284852 400998 284904 401004
rect 283840 400784 283892 400790
rect 283840 400726 283892 400732
rect 283852 399908 283880 400726
rect 284864 399908 284892 400998
rect 286968 400648 287020 400654
rect 286968 400590 287020 400596
rect 285956 400376 286008 400382
rect 285956 400318 286008 400324
rect 285968 399908 285996 400318
rect 286980 399908 287008 400590
rect 278780 399832 278832 399838
rect 268120 399758 268594 399786
rect 278832 399780 279082 399786
rect 278780 399774 279082 399780
rect 278792 399758 279082 399774
rect 281920 399770 282302 399786
rect 281908 399764 282302 399770
rect 281960 399758 282302 399764
rect 281908 399706 281960 399712
rect 233608 399696 233660 399702
rect 233358 399644 233608 399650
rect 233358 399638 233660 399644
rect 233358 399622 233648 399638
rect 236486 399634 236776 399650
rect 236486 399628 236788 399634
rect 236486 399622 236736 399628
rect 236736 399570 236788 399576
rect 289268 399560 289320 399566
rect 232254 399498 232544 399514
rect 239614 399498 239904 399514
rect 289320 399508 289662 399514
rect 289268 399502 289662 399508
rect 232254 399492 232556 399498
rect 232254 399486 232504 399492
rect 239614 399492 239916 399498
rect 239614 399486 239864 399492
rect 232504 399434 232556 399440
rect 289280 399486 289662 399502
rect 239864 399434 239916 399440
rect 285036 399424 285088 399430
rect 231582 399392 231638 399401
rect 231242 399350 231582 399378
rect 232962 399392 233018 399401
rect 232806 399350 232962 399378
rect 231582 399327 231638 399336
rect 237194 399392 237250 399401
rect 233910 399350 234200 399378
rect 234370 399350 234568 399378
rect 237038 399350 237194 399378
rect 232962 399327 233018 399336
rect 234172 399294 234200 399350
rect 234540 399294 234568 399350
rect 237194 399327 237250 399336
rect 238298 399392 238354 399401
rect 242530 399392 242586 399401
rect 238354 399350 238602 399378
rect 242282 399350 242530 399378
rect 238298 399327 238354 399336
rect 242530 399327 242586 399336
rect 276846 399392 276902 399401
rect 283010 399392 283066 399401
rect 276902 399350 277058 399378
rect 279344 399362 279634 399378
rect 282472 399362 282762 399378
rect 279332 399356 279634 399362
rect 276846 399327 276902 399336
rect 279384 399350 279634 399356
rect 282460 399356 282762 399362
rect 279332 399298 279384 399304
rect 282512 399350 282762 399356
rect 284482 399392 284538 399401
rect 283066 399350 283314 399378
rect 284418 399350 284482 399378
rect 283010 399327 283066 399336
rect 286138 399392 286194 399401
rect 285088 399372 285430 399378
rect 285036 399366 285430 399372
rect 285048 399350 285430 399366
rect 284482 399327 284538 399336
rect 287334 399392 287390 399401
rect 286194 399350 286442 399378
rect 286138 399327 286194 399336
rect 287886 399392 287942 399401
rect 287390 399350 287546 399378
rect 287334 399327 287390 399336
rect 287942 399350 288098 399378
rect 288360 399362 288558 399378
rect 288728 399362 289110 399378
rect 288348 399356 288558 399362
rect 287886 399327 287942 399336
rect 282460 399298 282512 399304
rect 288400 399350 288558 399356
rect 288716 399356 289110 399362
rect 288348 399298 288400 399304
rect 288768 399350 289110 399356
rect 288716 399298 288768 399304
rect 234160 399288 234212 399294
rect 229112 399214 230230 399242
rect 234160 399230 234212 399236
rect 234528 399288 234580 399294
rect 234528 399230 234580 399236
rect 228364 337136 228416 337142
rect 228364 337078 228416 337084
rect 227628 335368 227680 335374
rect 227628 335310 227680 335316
rect 227168 295316 227220 295322
rect 227168 295258 227220 295264
rect 227076 151768 227128 151774
rect 227076 151710 227128 151716
rect 226984 11756 227036 11762
rect 226984 11698 227036 11704
rect 227640 3874 227668 335310
rect 228376 14482 228404 337078
rect 229008 330880 229060 330886
rect 229008 330822 229060 330828
rect 228364 14476 228416 14482
rect 228364 14418 228416 14424
rect 228916 11756 228968 11762
rect 228916 11698 228968 11704
rect 225328 3868 225380 3874
rect 225328 3810 225380 3816
rect 226248 3868 226300 3874
rect 226248 3810 226300 3816
rect 226524 3868 226576 3874
rect 226524 3810 226576 3816
rect 227628 3868 227680 3874
rect 227628 3810 227680 3816
rect 227720 3868 227772 3874
rect 227720 3810 227772 3816
rect 224960 3460 225012 3466
rect 224960 3402 225012 3408
rect 220556 3318 220768 3346
rect 221752 3318 222148 3346
rect 222948 3318 223528 3346
rect 224144 3318 224908 3346
rect 220556 480 220584 3318
rect 221752 480 221780 3318
rect 222948 480 222976 3318
rect 224144 480 224172 3318
rect 224972 3233 225000 3402
rect 224958 3224 225014 3233
rect 224958 3159 225014 3168
rect 225340 480 225368 3810
rect 226536 480 226564 3810
rect 227732 480 227760 3810
rect 228928 480 228956 11698
rect 229020 3874 229048 330822
rect 229112 17950 229140 399214
rect 290476 346390 290504 401134
rect 297456 400988 297508 400994
rect 297456 400930 297508 400936
rect 294604 400920 294656 400926
rect 294604 400862 294656 400868
rect 290556 400240 290608 400246
rect 290556 400182 290608 400188
rect 290464 346384 290516 346390
rect 290464 346326 290516 346332
rect 229296 340054 230046 340082
rect 229192 335640 229244 335646
rect 229192 335582 229244 335588
rect 229100 17944 229152 17950
rect 229100 17886 229152 17892
rect 229204 4962 229232 335582
rect 229296 5030 229324 340054
rect 230124 335594 230152 340068
rect 230216 335646 230244 340068
rect 229388 335566 230152 335594
rect 230204 335640 230256 335646
rect 230204 335582 230256 335588
rect 229284 5024 229336 5030
rect 229284 4966 229336 4972
rect 229192 4956 229244 4962
rect 229192 4898 229244 4904
rect 229388 4826 229416 335566
rect 230308 335442 230336 340068
rect 230492 337414 230520 340068
rect 230480 337408 230532 337414
rect 230480 337350 230532 337356
rect 230388 336796 230440 336802
rect 230388 336738 230440 336744
rect 230296 335436 230348 335442
rect 230296 335378 230348 335384
rect 230400 335322 230428 336738
rect 230480 336524 230532 336530
rect 230480 336466 230532 336472
rect 229756 335294 230428 335322
rect 229560 328500 229612 328506
rect 229560 328442 229612 328448
rect 229572 318782 229600 328442
rect 229756 319462 229784 335294
rect 230492 335186 230520 336466
rect 230584 335510 230612 340068
rect 230690 340054 230796 340082
rect 230664 335640 230716 335646
rect 230664 335582 230716 335588
rect 230572 335504 230624 335510
rect 230572 335446 230624 335452
rect 230400 335158 230520 335186
rect 229744 319456 229796 319462
rect 229744 319398 229796 319404
rect 229560 318776 229612 318782
rect 229560 318718 229612 318724
rect 229468 310820 229520 310826
rect 229468 310762 229520 310768
rect 229480 309126 229508 310762
rect 229468 309120 229520 309126
rect 229468 309062 229520 309068
rect 229560 299532 229612 299538
rect 229560 299474 229612 299480
rect 229572 294522 229600 299474
rect 229572 294494 229692 294522
rect 229664 282826 229692 294494
rect 229572 282798 229692 282826
rect 229572 280158 229600 282798
rect 229560 280152 229612 280158
rect 229560 280094 229612 280100
rect 229652 270564 229704 270570
rect 229652 270506 229704 270512
rect 229664 263514 229692 270506
rect 229572 263486 229692 263514
rect 229572 260846 229600 263486
rect 229560 260840 229612 260846
rect 229560 260782 229612 260788
rect 229652 251252 229704 251258
rect 229652 251194 229704 251200
rect 229664 244202 229692 251194
rect 229572 244174 229692 244202
rect 229572 241505 229600 244174
rect 229558 241496 229614 241505
rect 229558 241431 229614 241440
rect 229834 241496 229890 241505
rect 229834 241431 229890 241440
rect 229848 231878 229876 241431
rect 229652 231872 229704 231878
rect 229652 231814 229704 231820
rect 229836 231872 229888 231878
rect 229836 231814 229888 231820
rect 229664 224890 229692 231814
rect 229572 224862 229692 224890
rect 229572 222193 229600 224862
rect 229558 222184 229614 222193
rect 229558 222119 229614 222128
rect 229834 222184 229890 222193
rect 229834 222119 229890 222128
rect 229848 212566 229876 222119
rect 229652 212560 229704 212566
rect 229652 212502 229704 212508
rect 229836 212560 229888 212566
rect 229836 212502 229888 212508
rect 229664 205578 229692 212502
rect 229572 205550 229692 205578
rect 229572 202881 229600 205550
rect 229558 202872 229614 202881
rect 229558 202807 229614 202816
rect 229834 202872 229890 202881
rect 229834 202807 229890 202816
rect 229848 193254 229876 202807
rect 229652 193248 229704 193254
rect 229652 193190 229704 193196
rect 229836 193248 229888 193254
rect 229836 193190 229888 193196
rect 229664 186266 229692 193190
rect 229572 186238 229692 186266
rect 229572 183569 229600 186238
rect 229558 183560 229614 183569
rect 229558 183495 229614 183504
rect 229834 183560 229890 183569
rect 229834 183495 229890 183504
rect 229848 173942 229876 183495
rect 229652 173936 229704 173942
rect 229652 173878 229704 173884
rect 229836 173936 229888 173942
rect 229836 173878 229888 173884
rect 229664 166954 229692 173878
rect 229572 166926 229692 166954
rect 229572 164218 229600 166926
rect 229560 164212 229612 164218
rect 229560 164154 229612 164160
rect 229836 164212 229888 164218
rect 229836 164154 229888 164160
rect 229848 154601 229876 164154
rect 229650 154592 229706 154601
rect 229650 154527 229706 154536
rect 229834 154592 229890 154601
rect 229834 154527 229890 154536
rect 229664 147642 229692 154527
rect 229572 147614 229692 147642
rect 229572 138038 229600 147614
rect 229560 138032 229612 138038
rect 229560 137974 229612 137980
rect 229468 137964 229520 137970
rect 229468 137906 229520 137912
rect 229480 135289 229508 137906
rect 229466 135280 229522 135289
rect 229466 135215 229522 135224
rect 229650 135280 229706 135289
rect 229650 135215 229706 135224
rect 229664 128330 229692 135215
rect 229572 128302 229692 128330
rect 229572 118726 229600 128302
rect 229560 118720 229612 118726
rect 229560 118662 229612 118668
rect 229468 118652 229520 118658
rect 229468 118594 229520 118600
rect 229480 115977 229508 118594
rect 229466 115968 229522 115977
rect 229466 115903 229522 115912
rect 229650 115968 229706 115977
rect 229650 115903 229706 115912
rect 229664 109018 229692 115903
rect 229572 108990 229692 109018
rect 229572 99414 229600 108990
rect 229560 99408 229612 99414
rect 229560 99350 229612 99356
rect 229468 99340 229520 99346
rect 229468 99282 229520 99288
rect 229480 96665 229508 99282
rect 229466 96656 229522 96665
rect 229466 96591 229522 96600
rect 229650 96656 229706 96665
rect 229650 96591 229706 96600
rect 229664 89706 229692 96591
rect 229572 89678 229692 89706
rect 229572 80102 229600 89678
rect 229560 80096 229612 80102
rect 229560 80038 229612 80044
rect 229652 80028 229704 80034
rect 229652 79970 229704 79976
rect 229664 77246 229692 79970
rect 229652 77240 229704 77246
rect 229652 77182 229704 77188
rect 229560 67652 229612 67658
rect 229560 67594 229612 67600
rect 229572 60738 229600 67594
rect 229480 60722 229600 60738
rect 229468 60716 229600 60722
rect 229520 60710 229600 60716
rect 229652 60716 229704 60722
rect 229468 60658 229520 60664
rect 229652 60658 229704 60664
rect 229664 57934 229692 60658
rect 229652 57928 229704 57934
rect 229652 57870 229704 57876
rect 229560 48340 229612 48346
rect 229560 48282 229612 48288
rect 229572 41426 229600 48282
rect 229480 41410 229600 41426
rect 229468 41404 229600 41410
rect 229520 41398 229600 41404
rect 229652 41404 229704 41410
rect 229468 41346 229520 41352
rect 229652 41346 229704 41352
rect 229664 38622 229692 41346
rect 229652 38616 229704 38622
rect 229652 38558 229704 38564
rect 229560 29028 229612 29034
rect 229560 28970 229612 28976
rect 229572 22166 229600 28970
rect 229560 22160 229612 22166
rect 229560 22102 229612 22108
rect 229560 22024 229612 22030
rect 229560 21966 229612 21972
rect 229572 10334 229600 21966
rect 229560 10328 229612 10334
rect 229560 10270 229612 10276
rect 229376 4820 229428 4826
rect 229376 4762 229428 4768
rect 229008 3868 229060 3874
rect 229008 3810 229060 3816
rect 229744 3528 229796 3534
rect 229744 3470 229796 3476
rect 229756 3346 229784 3470
rect 229664 3318 229784 3346
rect 229836 3324 229888 3330
rect 229664 3058 229692 3318
rect 229836 3266 229888 3272
rect 229848 3233 229876 3266
rect 229834 3224 229890 3233
rect 229834 3159 229890 3168
rect 229652 3052 229704 3058
rect 229652 2994 229704 3000
rect 230400 610 230428 335158
rect 230676 6186 230704 335582
rect 230664 6180 230716 6186
rect 230664 6122 230716 6128
rect 230768 4622 230796 340054
rect 230860 10402 230888 340068
rect 230952 337550 230980 340068
rect 230940 337544 230992 337550
rect 230940 337486 230992 337492
rect 231044 337482 231072 340068
rect 231136 340054 231242 340082
rect 231032 337476 231084 337482
rect 231032 337418 231084 337424
rect 231136 335646 231164 340054
rect 231320 336802 231348 340068
rect 231308 336796 231360 336802
rect 231308 336738 231360 336744
rect 231124 335640 231176 335646
rect 231124 335582 231176 335588
rect 231124 335504 231176 335510
rect 231124 335446 231176 335452
rect 230848 10396 230900 10402
rect 230848 10338 230900 10344
rect 230756 4616 230808 4622
rect 230756 4558 230808 4564
rect 231136 3369 231164 335446
rect 231308 10328 231360 10334
rect 231308 10270 231360 10276
rect 231122 3360 231178 3369
rect 231122 3295 231178 3304
rect 230112 604 230164 610
rect 230112 546 230164 552
rect 230388 604 230440 610
rect 230388 546 230440 552
rect 230124 480 230152 546
rect 231320 480 231348 10270
rect 231412 3505 231440 340068
rect 231492 332648 231544 332654
rect 231492 332590 231544 332596
rect 231504 326398 231532 332590
rect 231492 326392 231544 326398
rect 231492 326334 231544 326340
rect 231596 3641 231624 340068
rect 231688 8974 231716 340068
rect 231780 332654 231808 340068
rect 231964 337686 231992 340068
rect 231952 337680 232004 337686
rect 231952 337622 232004 337628
rect 232056 337618 232084 340068
rect 232044 337612 232096 337618
rect 232044 337554 232096 337560
rect 231860 337476 231912 337482
rect 231860 337418 231912 337424
rect 231872 334626 231900 337418
rect 231952 337408 232004 337414
rect 231952 337350 232004 337356
rect 231964 335374 231992 337350
rect 232044 335844 232096 335850
rect 232044 335786 232096 335792
rect 231952 335368 232004 335374
rect 231952 335310 232004 335316
rect 231860 334620 231912 334626
rect 231860 334562 231912 334568
rect 231768 332648 231820 332654
rect 231768 332590 231820 332596
rect 232056 313954 232084 335786
rect 232044 313948 232096 313954
rect 232044 313890 232096 313896
rect 232148 10470 232176 340068
rect 232240 340054 232346 340082
rect 232240 335918 232268 340054
rect 232424 339946 232452 340068
rect 232332 339918 232452 339946
rect 232228 335912 232280 335918
rect 232228 335854 232280 335860
rect 232228 335708 232280 335714
rect 232228 335650 232280 335656
rect 232240 10538 232268 335650
rect 232332 335646 232360 339918
rect 232516 335782 232544 340068
rect 232608 340054 232714 340082
rect 232504 335776 232556 335782
rect 232504 335718 232556 335724
rect 232608 335714 232636 340054
rect 232688 335912 232740 335918
rect 232688 335854 232740 335860
rect 232596 335708 232648 335714
rect 232596 335650 232648 335656
rect 232320 335640 232372 335646
rect 232320 335582 232372 335588
rect 232700 315314 232728 335854
rect 232792 335850 232820 340068
rect 232884 337822 232912 340068
rect 232872 337816 232924 337822
rect 232872 337758 232924 337764
rect 232780 335844 232832 335850
rect 232780 335786 232832 335792
rect 232964 335776 233016 335782
rect 232964 335718 233016 335724
rect 232780 335640 232832 335646
rect 232780 335582 232832 335588
rect 232688 315308 232740 315314
rect 232688 315250 232740 315256
rect 232228 10532 232280 10538
rect 232228 10474 232280 10480
rect 232136 10464 232188 10470
rect 232136 10406 232188 10412
rect 232504 10396 232556 10402
rect 232504 10338 232556 10344
rect 231676 8968 231728 8974
rect 231676 8910 231728 8916
rect 231582 3632 231638 3641
rect 231582 3567 231638 3576
rect 231398 3496 231454 3505
rect 231398 3431 231454 3440
rect 232516 480 232544 10338
rect 232792 3777 232820 335582
rect 232976 3913 233004 335718
rect 233068 10606 233096 340068
rect 233160 312594 233188 340068
rect 233266 340054 233372 340082
rect 233240 335980 233292 335986
rect 233240 335922 233292 335928
rect 233252 334234 233280 335922
rect 233344 334354 233372 340054
rect 233436 335850 233464 340068
rect 233424 335844 233476 335850
rect 233424 335786 233476 335792
rect 233424 335708 233476 335714
rect 233424 335650 233476 335656
rect 233332 334348 233384 334354
rect 233332 334290 233384 334296
rect 233252 334206 233372 334234
rect 233344 324970 233372 334206
rect 233436 329118 233464 335650
rect 233528 333962 233556 340068
rect 233620 337754 233648 340068
rect 233712 340054 233818 340082
rect 233608 337748 233660 337754
rect 233608 337690 233660 337696
rect 233608 337612 233660 337618
rect 233608 337554 233660 337560
rect 233620 336054 233648 337554
rect 233608 336048 233660 336054
rect 233608 335990 233660 335996
rect 233712 335714 233740 340054
rect 233792 336660 233844 336666
rect 233792 336602 233844 336608
rect 233700 335708 233752 335714
rect 233700 335650 233752 335656
rect 233804 334098 233832 336602
rect 233896 334506 233924 340068
rect 234002 340054 234108 340082
rect 234080 335714 234108 340054
rect 234172 335986 234200 340068
rect 234160 335980 234212 335986
rect 234160 335922 234212 335928
rect 234160 335844 234212 335850
rect 234160 335786 234212 335792
rect 234068 335708 234120 335714
rect 234068 335650 234120 335656
rect 233896 334478 234108 334506
rect 233804 334070 233924 334098
rect 233528 333934 233740 333962
rect 233608 333872 233660 333878
rect 233608 333814 233660 333820
rect 233516 331220 233568 331226
rect 233516 331162 233568 331168
rect 233424 329112 233476 329118
rect 233424 329054 233476 329060
rect 233332 324964 233384 324970
rect 233332 324906 233384 324912
rect 233528 321638 233556 331162
rect 233516 321632 233568 321638
rect 233516 321574 233568 321580
rect 233148 312588 233200 312594
rect 233148 312530 233200 312536
rect 233620 305658 233648 333814
rect 233712 331226 233740 333934
rect 233700 331220 233752 331226
rect 233700 331162 233752 331168
rect 233896 322250 233924 334070
rect 234080 333878 234108 334478
rect 234068 333872 234120 333878
rect 234068 333814 234120 333820
rect 234068 331832 234120 331838
rect 234068 331774 234120 331780
rect 233976 327140 234028 327146
rect 233976 327082 234028 327088
rect 233884 322244 233936 322250
rect 233884 322186 233936 322192
rect 233700 321632 233752 321638
rect 233700 321574 233752 321580
rect 233712 307086 233740 321574
rect 233988 318918 234016 327082
rect 233976 318912 234028 318918
rect 233976 318854 234028 318860
rect 233976 318776 234028 318782
rect 233976 318718 234028 318724
rect 233988 307766 234016 318718
rect 233976 307760 234028 307766
rect 233976 307702 234028 307708
rect 233792 307692 233844 307698
rect 233792 307634 233844 307640
rect 233700 307080 233752 307086
rect 233700 307022 233752 307028
rect 233608 305652 233660 305658
rect 233608 305594 233660 305600
rect 233804 294658 233832 307634
rect 233804 294630 233924 294658
rect 233896 282946 233924 294630
rect 233700 282940 233752 282946
rect 233700 282882 233752 282888
rect 233884 282940 233936 282946
rect 233884 282882 233936 282888
rect 233712 282826 233740 282882
rect 233712 282798 233832 282826
rect 233804 273306 233832 282798
rect 233804 273278 233924 273306
rect 233896 263634 233924 273278
rect 233700 263628 233752 263634
rect 233700 263570 233752 263576
rect 233884 263628 233936 263634
rect 233884 263570 233936 263576
rect 233712 263514 233740 263570
rect 233712 263486 233832 263514
rect 233804 253994 233832 263486
rect 233804 253966 233924 253994
rect 233896 244322 233924 253966
rect 233700 244316 233752 244322
rect 233700 244258 233752 244264
rect 233884 244316 233936 244322
rect 233884 244258 233936 244264
rect 233712 244202 233740 244258
rect 233712 244174 233832 244202
rect 233804 234682 233832 244174
rect 233804 234654 233924 234682
rect 233896 225010 233924 234654
rect 233700 225004 233752 225010
rect 233700 224946 233752 224952
rect 233884 225004 233936 225010
rect 233884 224946 233936 224952
rect 233712 224890 233740 224946
rect 233712 224862 233832 224890
rect 233804 215370 233832 224862
rect 233804 215342 233924 215370
rect 233896 205698 233924 215342
rect 233700 205692 233752 205698
rect 233700 205634 233752 205640
rect 233884 205692 233936 205698
rect 233884 205634 233936 205640
rect 233712 205578 233740 205634
rect 233712 205550 233832 205578
rect 233804 196058 233832 205550
rect 233804 196030 233924 196058
rect 233896 186386 233924 196030
rect 233700 186380 233752 186386
rect 233700 186322 233752 186328
rect 233884 186380 233936 186386
rect 233884 186322 233936 186328
rect 233712 186266 233740 186322
rect 233712 186238 233832 186266
rect 233804 179194 233832 186238
rect 233804 179166 233924 179194
rect 233896 167074 233924 179166
rect 233700 167068 233752 167074
rect 233700 167010 233752 167016
rect 233884 167068 233936 167074
rect 233884 167010 233936 167016
rect 233712 166954 233740 167010
rect 233712 166926 233832 166954
rect 233804 154442 233832 166926
rect 233804 154414 234016 154442
rect 233988 144945 234016 154414
rect 233790 144936 233846 144945
rect 233790 144871 233846 144880
rect 233974 144936 234030 144945
rect 233974 144871 234030 144880
rect 233804 140026 233832 144871
rect 233804 139998 233924 140026
rect 233896 128382 233924 139998
rect 233700 128376 233752 128382
rect 233884 128376 233936 128382
rect 233752 128324 233832 128330
rect 233700 128318 233832 128324
rect 233884 128318 233936 128324
rect 233712 128302 233832 128318
rect 233804 120714 233832 128302
rect 233804 120686 233924 120714
rect 233896 109070 233924 120686
rect 233700 109064 233752 109070
rect 233884 109064 233936 109070
rect 233752 109012 233832 109018
rect 233700 109006 233832 109012
rect 233884 109006 233936 109012
rect 233712 108990 233832 109006
rect 233804 104854 233832 108990
rect 233792 104848 233844 104854
rect 233792 104790 233844 104796
rect 233976 95260 234028 95266
rect 233976 95202 234028 95208
rect 233988 87009 234016 95202
rect 233790 87000 233846 87009
rect 233790 86935 233846 86944
rect 233974 87000 234030 87009
rect 233974 86935 234030 86944
rect 233804 77314 233832 86935
rect 233792 77308 233844 77314
rect 233792 77250 233844 77256
rect 233884 77308 233936 77314
rect 233884 77250 233936 77256
rect 233896 67658 233924 77250
rect 233792 67652 233844 67658
rect 233792 67594 233844 67600
rect 233884 67652 233936 67658
rect 233884 67594 233936 67600
rect 233804 60738 233832 67594
rect 233804 60710 233924 60738
rect 233896 50946 233924 60710
rect 233804 50918 233924 50946
rect 233804 41426 233832 50918
rect 233804 41398 233924 41426
rect 233896 31770 233924 41398
rect 233712 31742 233924 31770
rect 233712 31634 233740 31742
rect 233712 31606 233832 31634
rect 233804 12594 233832 31606
rect 233712 12566 233832 12594
rect 233056 10600 233108 10606
rect 233056 10542 233108 10548
rect 233712 4978 233740 12566
rect 233620 4950 233740 4978
rect 233620 4049 233648 4950
rect 233700 4820 233752 4826
rect 233700 4762 233752 4768
rect 233606 4040 233662 4049
rect 233606 3975 233662 3984
rect 232962 3904 233018 3913
rect 232962 3839 233018 3848
rect 232778 3768 232834 3777
rect 232778 3703 232834 3712
rect 233712 480 233740 4762
rect 234080 3534 234108 331774
rect 234172 330546 234200 335786
rect 234160 330540 234212 330546
rect 234160 330482 234212 330488
rect 234264 304298 234292 340068
rect 234356 331838 234384 340068
rect 234436 335708 234488 335714
rect 234436 335650 234488 335656
rect 234344 331832 234396 331838
rect 234344 331774 234396 331780
rect 234252 304292 234304 304298
rect 234252 304234 234304 304240
rect 234068 3528 234120 3534
rect 234068 3470 234120 3476
rect 234448 3330 234476 335650
rect 234540 323610 234568 340068
rect 234632 335646 234660 340068
rect 234738 340054 234844 340082
rect 234620 335640 234672 335646
rect 234620 335582 234672 335588
rect 234816 331702 234844 340054
rect 234908 337618 234936 340068
rect 234896 337612 234948 337618
rect 234896 337554 234948 337560
rect 235000 331906 235028 340068
rect 234988 331900 235040 331906
rect 234988 331842 235040 331848
rect 235092 331786 235120 340068
rect 235276 337482 235304 340068
rect 235264 337476 235316 337482
rect 235264 337418 235316 337424
rect 234908 331758 235120 331786
rect 234804 331696 234856 331702
rect 234804 331638 234856 331644
rect 234528 323604 234580 323610
rect 234528 323546 234580 323552
rect 234908 318102 234936 331758
rect 235080 331696 235132 331702
rect 235080 331638 235132 331644
rect 234896 318096 234948 318102
rect 234896 318038 234948 318044
rect 234986 241496 235042 241505
rect 234986 241431 235042 241440
rect 235000 231878 235028 241431
rect 234988 231872 235040 231878
rect 234988 231814 235040 231820
rect 234986 220824 235042 220833
rect 234986 220759 235042 220768
rect 235000 211177 235028 220759
rect 234986 211168 235042 211177
rect 234986 211103 235042 211112
rect 234988 201408 235040 201414
rect 234988 201350 235040 201356
rect 235000 183598 235028 201350
rect 234988 183592 235040 183598
rect 234986 183560 234988 183569
rect 235040 183560 235042 183569
rect 234986 183495 235042 183504
rect 235000 173942 235028 183495
rect 234988 173936 235040 173942
rect 234988 173878 235040 173884
rect 234988 172508 235040 172514
rect 234988 172450 235040 172456
rect 235000 162897 235028 172450
rect 234986 162888 235042 162897
rect 234986 162823 235042 162832
rect 234804 6180 234856 6186
rect 234804 6122 234856 6128
rect 234436 3324 234488 3330
rect 234436 3266 234488 3272
rect 234816 480 234844 6122
rect 235092 3466 235120 331638
rect 235368 327758 235396 340068
rect 235356 327752 235408 327758
rect 235356 327694 235408 327700
rect 235460 327570 235488 340068
rect 235644 333266 235672 340068
rect 235632 333260 235684 333266
rect 235632 333202 235684 333208
rect 235540 331628 235592 331634
rect 235540 331570 235592 331576
rect 235184 327542 235488 327570
rect 235184 317422 235212 327542
rect 235172 317416 235224 317422
rect 235172 317358 235224 317364
rect 235356 301980 235408 301986
rect 235356 301922 235408 301928
rect 235368 298110 235396 301922
rect 235356 298104 235408 298110
rect 235356 298046 235408 298052
rect 235356 289808 235408 289814
rect 235356 289750 235408 289756
rect 235184 278798 235212 278829
rect 235368 278798 235396 289750
rect 235552 280158 235580 331570
rect 235736 331294 235764 340068
rect 235828 331634 235856 340068
rect 235908 335640 235960 335646
rect 235908 335582 235960 335588
rect 235816 331628 235868 331634
rect 235816 331570 235868 331576
rect 235724 331288 235776 331294
rect 235724 331230 235776 331236
rect 235724 331152 235776 331158
rect 235724 331094 235776 331100
rect 235736 326466 235764 331094
rect 235724 326460 235776 326466
rect 235724 326402 235776 326408
rect 235920 311166 235948 335582
rect 236012 335170 236040 340068
rect 236104 335714 236132 340068
rect 236092 335708 236144 335714
rect 236092 335650 236144 335656
rect 236196 335458 236224 340068
rect 236380 335714 236408 340068
rect 236472 335968 236500 340068
rect 236564 336122 236592 340068
rect 236656 340054 236762 340082
rect 236552 336116 236604 336122
rect 236552 336058 236604 336064
rect 236472 335940 236592 335968
rect 236460 335844 236512 335850
rect 236460 335786 236512 335792
rect 236368 335708 236420 335714
rect 236368 335650 236420 335656
rect 236104 335430 236224 335458
rect 236276 335504 236328 335510
rect 236276 335446 236328 335452
rect 236000 335164 236052 335170
rect 236000 335106 236052 335112
rect 235908 311160 235960 311166
rect 235908 311102 235960 311108
rect 235540 280152 235592 280158
rect 235540 280094 235592 280100
rect 235172 278792 235224 278798
rect 235356 278792 235408 278798
rect 235224 278740 235304 278746
rect 235172 278734 235304 278740
rect 235356 278734 235408 278740
rect 235184 278718 235304 278734
rect 235276 273970 235304 278718
rect 235264 273964 235316 273970
rect 235264 273906 235316 273912
rect 235540 270564 235592 270570
rect 235540 270506 235592 270512
rect 235172 260908 235224 260914
rect 235172 260850 235224 260856
rect 235184 259418 235212 260850
rect 235172 259412 235224 259418
rect 235172 259354 235224 259360
rect 235172 244044 235224 244050
rect 235172 243986 235224 243992
rect 235184 241505 235212 243986
rect 235552 241505 235580 270506
rect 235170 241496 235226 241505
rect 235170 241431 235226 241440
rect 235538 241496 235594 241505
rect 235538 241431 235594 241440
rect 235722 241496 235778 241505
rect 235722 241431 235778 241440
rect 235264 231872 235316 231878
rect 235264 231814 235316 231820
rect 235276 225026 235304 231814
rect 235736 230518 235764 241431
rect 235540 230512 235592 230518
rect 235540 230454 235592 230460
rect 235724 230512 235776 230518
rect 235724 230454 235776 230460
rect 235276 224998 235396 225026
rect 235368 222222 235396 224998
rect 235172 222216 235224 222222
rect 235172 222158 235224 222164
rect 235356 222216 235408 222222
rect 235356 222158 235408 222164
rect 235184 220833 235212 222158
rect 235552 220833 235580 230454
rect 235170 220824 235226 220833
rect 235170 220759 235226 220768
rect 235538 220824 235594 220833
rect 235538 220759 235594 220768
rect 235722 220824 235778 220833
rect 235722 220759 235778 220768
rect 235736 211177 235764 220759
rect 235170 211168 235226 211177
rect 235170 211103 235226 211112
rect 235538 211168 235594 211177
rect 235538 211103 235594 211112
rect 235722 211168 235778 211177
rect 235722 211103 235778 211112
rect 235184 202842 235212 211103
rect 235552 202910 235580 211103
rect 235540 202904 235592 202910
rect 235540 202846 235592 202852
rect 235632 202904 235684 202910
rect 235632 202846 235684 202852
rect 235172 202836 235224 202842
rect 235172 202778 235224 202784
rect 235264 202836 235316 202842
rect 235264 202778 235316 202784
rect 235276 201482 235304 202778
rect 235264 201476 235316 201482
rect 235264 201418 235316 201424
rect 235644 193254 235672 202846
rect 235540 193248 235592 193254
rect 235540 193190 235592 193196
rect 235632 193248 235684 193254
rect 235632 193190 235684 193196
rect 235552 188442 235580 193190
rect 235460 188414 235580 188442
rect 235172 183592 235224 183598
rect 235170 183560 235172 183569
rect 235224 183560 235226 183569
rect 235170 183495 235226 183504
rect 235460 173942 235488 188414
rect 235264 173936 235316 173942
rect 235264 173878 235316 173884
rect 235448 173936 235500 173942
rect 235448 173878 235500 173884
rect 235540 173936 235592 173942
rect 235540 173878 235592 173884
rect 235276 172514 235304 173878
rect 235264 172508 235316 172514
rect 235264 172450 235316 172456
rect 235170 162888 235226 162897
rect 235170 162823 235226 162832
rect 235184 162790 235212 162823
rect 235172 162784 235224 162790
rect 235172 162726 235224 162732
rect 235172 157412 235224 157418
rect 235172 157354 235224 157360
rect 235184 144906 235212 157354
rect 235552 144906 235580 173878
rect 235172 144900 235224 144906
rect 235172 144842 235224 144848
rect 235540 144900 235592 144906
rect 235540 144842 235592 144848
rect 235264 144832 235316 144838
rect 235264 144774 235316 144780
rect 235276 143546 235304 144774
rect 235264 143540 235316 143546
rect 235264 143482 235316 143488
rect 235540 135312 235592 135318
rect 235540 135254 235592 135260
rect 235264 133952 235316 133958
rect 235264 133894 235316 133900
rect 235276 124234 235304 133894
rect 235552 125594 235580 135254
rect 235540 125588 235592 125594
rect 235540 125530 235592 125536
rect 235264 124228 235316 124234
rect 235264 124170 235316 124176
rect 235264 122868 235316 122874
rect 235264 122810 235316 122816
rect 235276 114510 235304 122810
rect 235540 116000 235592 116006
rect 235540 115942 235592 115948
rect 235264 114504 235316 114510
rect 235264 114446 235316 114452
rect 235356 114504 235408 114510
rect 235356 114446 235408 114452
rect 235368 99550 235396 114446
rect 235356 99544 235408 99550
rect 235356 99486 235408 99492
rect 235172 99408 235224 99414
rect 235172 99350 235224 99356
rect 235184 86970 235212 99350
rect 235552 87145 235580 115942
rect 235538 87136 235594 87145
rect 235538 87071 235594 87080
rect 235446 87000 235502 87009
rect 235172 86964 235224 86970
rect 235172 86906 235224 86912
rect 235264 86964 235316 86970
rect 235446 86935 235502 86944
rect 235264 86906 235316 86912
rect 235276 85542 235304 86906
rect 235264 85536 235316 85542
rect 235264 85478 235316 85484
rect 235460 77314 235488 86935
rect 235448 77308 235500 77314
rect 235448 77250 235500 77256
rect 235540 77308 235592 77314
rect 235540 77250 235592 77256
rect 235264 75948 235316 75954
rect 235264 75890 235316 75896
rect 235276 70514 235304 75890
rect 235264 70508 235316 70514
rect 235264 70450 235316 70456
rect 235172 70372 235224 70378
rect 235172 70314 235224 70320
rect 235184 58002 235212 70314
rect 235552 67590 235580 77250
rect 235540 67584 235592 67590
rect 235540 67526 235592 67532
rect 235172 57996 235224 58002
rect 235172 57938 235224 57944
rect 235264 57996 235316 58002
rect 235264 57938 235316 57944
rect 235540 57996 235592 58002
rect 235540 57938 235592 57944
rect 235276 48414 235304 57938
rect 235172 48408 235224 48414
rect 235172 48350 235224 48356
rect 235264 48408 235316 48414
rect 235264 48350 235316 48356
rect 235184 46918 235212 48350
rect 235172 46912 235224 46918
rect 235172 46854 235224 46860
rect 235172 37324 235224 37330
rect 235172 37266 235224 37272
rect 235184 19378 235212 37266
rect 235552 28966 235580 57938
rect 235540 28960 235592 28966
rect 235540 28902 235592 28908
rect 235172 19372 235224 19378
rect 235172 19314 235224 19320
rect 235264 19372 235316 19378
rect 235264 19314 235316 19320
rect 235540 19372 235592 19378
rect 235540 19314 235592 19320
rect 235276 14498 235304 19314
rect 235184 14470 235304 14498
rect 235184 3670 235212 14470
rect 235552 3874 235580 19314
rect 236000 10464 236052 10470
rect 236000 10406 236052 10412
rect 235540 3868 235592 3874
rect 235540 3810 235592 3816
rect 235172 3664 235224 3670
rect 235172 3606 235224 3612
rect 235080 3460 235132 3466
rect 235080 3402 235132 3408
rect 236012 480 236040 10406
rect 236104 3806 236132 335430
rect 236184 335368 236236 335374
rect 236184 335310 236236 335316
rect 236196 3942 236224 335310
rect 236288 4010 236316 335446
rect 236368 335164 236420 335170
rect 236368 335106 236420 335112
rect 236380 9042 236408 335106
rect 236472 9178 236500 335786
rect 236564 335730 236592 335940
rect 236656 335850 236684 340054
rect 236840 336666 236868 340068
rect 236828 336660 236880 336666
rect 236828 336602 236880 336608
rect 236932 336274 236960 340068
rect 236840 336246 236960 336274
rect 237024 340054 237130 340082
rect 236644 335844 236696 335850
rect 236644 335786 236696 335792
rect 236564 335702 236776 335730
rect 236552 335640 236604 335646
rect 236552 335582 236604 335588
rect 236644 335640 236696 335646
rect 236644 335582 236696 335588
rect 236460 9172 236512 9178
rect 236460 9114 236512 9120
rect 236564 9110 236592 335582
rect 236656 9246 236684 335582
rect 236748 10742 236776 335702
rect 236840 335374 236868 336246
rect 236920 336116 236972 336122
rect 236920 336058 236972 336064
rect 236932 335492 236960 336058
rect 237024 335646 237052 340054
rect 237104 336796 237156 336802
rect 237104 336738 237156 336744
rect 237012 335640 237064 335646
rect 237012 335582 237064 335588
rect 236932 335464 237052 335492
rect 236828 335368 236880 335374
rect 236828 335310 236880 335316
rect 236828 335232 236880 335238
rect 236828 335174 236880 335180
rect 236736 10736 236788 10742
rect 236736 10678 236788 10684
rect 236840 10674 236868 335174
rect 237024 328438 237052 335464
rect 237116 331974 237144 336738
rect 237208 336190 237236 340068
rect 237196 336184 237248 336190
rect 237196 336126 237248 336132
rect 237300 335510 237328 340068
rect 237288 335504 237340 335510
rect 237288 335446 237340 335452
rect 237484 334506 237512 340068
rect 237576 334694 237604 340068
rect 237668 335714 237696 340068
rect 237760 340054 237866 340082
rect 237656 335708 237708 335714
rect 237656 335650 237708 335656
rect 237564 334688 237616 334694
rect 237564 334630 237616 334636
rect 237484 334478 237696 334506
rect 237104 331968 237156 331974
rect 237104 331910 237156 331916
rect 237012 328432 237064 328438
rect 237012 328374 237064 328380
rect 237104 318844 237156 318850
rect 237104 318786 237156 318792
rect 237116 312576 237144 318786
rect 237116 312548 237328 312576
rect 237300 307766 237328 312548
rect 237288 307760 237340 307766
rect 237288 307702 237340 307708
rect 237196 298172 237248 298178
rect 237196 298114 237248 298120
rect 237208 282826 237236 298114
rect 237116 282798 237236 282826
rect 237116 280158 237144 282798
rect 237104 280152 237156 280158
rect 237104 280094 237156 280100
rect 237196 280152 237248 280158
rect 237196 280094 237248 280100
rect 237208 263514 237236 280094
rect 237116 263486 237236 263514
rect 237116 253994 237144 263486
rect 237024 253966 237144 253994
rect 237024 253910 237052 253966
rect 237012 253904 237064 253910
rect 237012 253846 237064 253852
rect 237196 253904 237248 253910
rect 237196 253846 237248 253852
rect 237208 251190 237236 253846
rect 237196 251184 237248 251190
rect 237196 251126 237248 251132
rect 237104 241528 237156 241534
rect 237104 241470 237156 241476
rect 237116 220810 237144 241470
rect 237024 220782 237144 220810
rect 237024 212566 237052 220782
rect 237012 212560 237064 212566
rect 237012 212502 237064 212508
rect 237012 212424 237064 212430
rect 237012 212366 237064 212372
rect 237024 205578 237052 212366
rect 237024 205550 237144 205578
rect 237116 202842 237144 205550
rect 237104 202836 237156 202842
rect 237104 202778 237156 202784
rect 237196 202836 237248 202842
rect 237196 202778 237248 202784
rect 237208 186266 237236 202778
rect 237116 186238 237236 186266
rect 237116 183530 237144 186238
rect 237104 183524 237156 183530
rect 237104 183466 237156 183472
rect 237196 183524 237248 183530
rect 237196 183466 237248 183472
rect 237208 166954 237236 183466
rect 237116 166926 237236 166954
rect 237116 157434 237144 166926
rect 237024 157406 237144 157434
rect 237024 157350 237052 157406
rect 237012 157344 237064 157350
rect 237012 157286 237064 157292
rect 237196 157344 237248 157350
rect 237196 157286 237248 157292
rect 237208 144974 237236 157286
rect 237104 144968 237156 144974
rect 237104 144910 237156 144916
rect 237196 144968 237248 144974
rect 237196 144910 237248 144916
rect 237116 138038 237144 144910
rect 237104 138032 237156 138038
rect 237104 137974 237156 137980
rect 237196 137964 237248 137970
rect 237196 137906 237248 137912
rect 237208 128330 237236 137906
rect 237116 128302 237236 128330
rect 237116 118726 237144 128302
rect 237104 118720 237156 118726
rect 237104 118662 237156 118668
rect 237196 118652 237248 118658
rect 237196 118594 237248 118600
rect 237208 109018 237236 118594
rect 237116 108990 237236 109018
rect 237116 100042 237144 108990
rect 237116 100014 237236 100042
rect 237208 85542 237236 100014
rect 237196 85536 237248 85542
rect 237196 85478 237248 85484
rect 237012 76016 237064 76022
rect 237012 75958 237064 75964
rect 237024 75886 237052 75958
rect 237012 75880 237064 75886
rect 237012 75822 237064 75828
rect 237196 57996 237248 58002
rect 237196 57938 237248 57944
rect 237208 51134 237236 57938
rect 237196 51128 237248 51134
rect 237196 51070 237248 51076
rect 237104 51060 237156 51066
rect 237104 51002 237156 51008
rect 237116 41426 237144 51002
rect 237024 41410 237144 41426
rect 237012 41404 237144 41410
rect 237064 41398 237144 41404
rect 237196 41404 237248 41410
rect 237012 41346 237064 41352
rect 237196 41346 237248 41352
rect 237208 31822 237236 41346
rect 237196 31816 237248 31822
rect 237196 31758 237248 31764
rect 237012 31748 237064 31754
rect 237012 31690 237064 31696
rect 237024 19378 237052 31690
rect 237012 19372 237064 19378
rect 237012 19314 237064 19320
rect 237104 19372 237156 19378
rect 237104 19314 237156 19320
rect 237116 14498 237144 19314
rect 237024 14470 237144 14498
rect 236828 10668 236880 10674
rect 236828 10610 236880 10616
rect 236644 9240 236696 9246
rect 236644 9182 236696 9188
rect 236552 9104 236604 9110
rect 236552 9046 236604 9052
rect 236368 9036 236420 9042
rect 236368 8978 236420 8984
rect 236276 4004 236328 4010
rect 236276 3946 236328 3952
rect 236184 3936 236236 3942
rect 236184 3878 236236 3884
rect 236092 3800 236144 3806
rect 236092 3742 236144 3748
rect 237024 3398 237052 14470
rect 237668 9314 237696 334478
rect 237760 9382 237788 340054
rect 237944 330614 237972 340068
rect 237932 330608 237984 330614
rect 237932 330550 237984 330556
rect 237748 9376 237800 9382
rect 237748 9318 237800 9324
rect 237656 9308 237708 9314
rect 237656 9250 237708 9256
rect 237288 4888 237340 4894
rect 237288 4830 237340 4836
rect 237012 3392 237064 3398
rect 237012 3334 237064 3340
rect 237300 2530 237328 4830
rect 238036 4146 238064 340068
rect 238116 335640 238168 335646
rect 238116 335582 238168 335588
rect 238024 4140 238076 4146
rect 238024 4082 238076 4088
rect 238128 3262 238156 335582
rect 238220 9450 238248 340068
rect 238312 320890 238340 340068
rect 238404 335646 238432 340068
rect 238484 335708 238536 335714
rect 238484 335650 238536 335656
rect 238392 335640 238444 335646
rect 238392 335582 238444 335588
rect 238300 320884 238352 320890
rect 238300 320826 238352 320832
rect 238208 9444 238260 9450
rect 238208 9386 238260 9392
rect 238392 6044 238444 6050
rect 238392 5986 238444 5992
rect 238116 3256 238168 3262
rect 238116 3198 238168 3204
rect 237208 2502 237328 2530
rect 237208 480 237236 2502
rect 238404 480 238432 5986
rect 238496 4078 238524 335650
rect 238588 9518 238616 340068
rect 238680 329186 238708 340068
rect 238786 340054 238892 340082
rect 238864 333826 238892 340054
rect 238956 335696 238984 340068
rect 239048 336802 239076 340068
rect 239036 336796 239088 336802
rect 239036 336738 239088 336744
rect 239140 335714 239168 340068
rect 239232 340054 239338 340082
rect 239128 335708 239180 335714
rect 238956 335668 239076 335696
rect 238864 333798 238984 333826
rect 238668 329180 238720 329186
rect 238668 329122 238720 329128
rect 238956 280106 238984 333798
rect 238864 280078 238984 280106
rect 238864 270638 238892 280078
rect 238852 270632 238904 270638
rect 238852 270574 238904 270580
rect 238944 270564 238996 270570
rect 238944 270506 238996 270512
rect 238956 241466 238984 270506
rect 238944 241460 238996 241466
rect 238944 241402 238996 241408
rect 238944 231872 238996 231878
rect 238944 231814 238996 231820
rect 238956 202842 238984 231814
rect 238944 202836 238996 202842
rect 238944 202778 238996 202784
rect 238944 191888 238996 191894
rect 238944 191830 238996 191836
rect 238956 162858 238984 191830
rect 238760 162852 238812 162858
rect 238760 162794 238812 162800
rect 238944 162852 238996 162858
rect 238944 162794 238996 162800
rect 238772 153241 238800 162794
rect 238758 153232 238814 153241
rect 238758 153167 238814 153176
rect 238942 153232 238998 153241
rect 238942 153167 238998 153176
rect 238956 145081 238984 153167
rect 238942 145072 238998 145081
rect 238942 145007 238998 145016
rect 238758 144800 238814 144809
rect 238758 144735 238814 144744
rect 238772 135289 238800 144735
rect 238758 135280 238814 135289
rect 238758 135215 238814 135224
rect 238942 135280 238998 135289
rect 238942 135215 238998 135224
rect 238956 125769 238984 135215
rect 238942 125760 238998 125769
rect 238942 125695 238998 125704
rect 238758 125352 238814 125361
rect 238758 125287 238814 125296
rect 238772 115977 238800 125287
rect 238758 115968 238814 115977
rect 238758 115903 238814 115912
rect 238942 115968 238998 115977
rect 238942 115903 238998 115912
rect 238576 9512 238628 9518
rect 238576 9454 238628 9460
rect 238484 4072 238536 4078
rect 238484 4014 238536 4020
rect 238956 3602 238984 115903
rect 239048 9586 239076 335668
rect 239128 335650 239180 335656
rect 239128 335572 239180 335578
rect 239128 335514 239180 335520
rect 239036 9580 239088 9586
rect 239036 9522 239088 9528
rect 239140 8838 239168 335514
rect 239232 9654 239260 340054
rect 239416 333334 239444 340068
rect 239404 333328 239456 333334
rect 239404 333270 239456 333276
rect 239220 9648 239272 9654
rect 239220 9590 239272 9596
rect 239128 8832 239180 8838
rect 239128 8774 239180 8780
rect 238944 3596 238996 3602
rect 238944 3538 238996 3544
rect 239508 3194 239536 340068
rect 239588 335640 239640 335646
rect 239588 335582 239640 335588
rect 239600 4298 239628 335582
rect 239692 8906 239720 340068
rect 239784 327826 239812 340068
rect 239876 335646 239904 340068
rect 239956 335708 240008 335714
rect 239956 335650 240008 335656
rect 239864 335640 239916 335646
rect 239864 335582 239916 335588
rect 239772 327820 239824 327826
rect 239772 327762 239824 327768
rect 239680 8900 239732 8906
rect 239680 8842 239732 8848
rect 239600 4270 239720 4298
rect 239588 4140 239640 4146
rect 239588 4082 239640 4088
rect 239496 3188 239548 3194
rect 239496 3130 239548 3136
rect 239600 480 239628 4082
rect 239692 3126 239720 4270
rect 239680 3120 239732 3126
rect 239680 3062 239732 3068
rect 239968 3058 239996 335650
rect 240060 335578 240088 340068
rect 240048 335572 240100 335578
rect 240048 335514 240100 335520
rect 240048 335436 240100 335442
rect 240048 335378 240100 335384
rect 240060 4146 240088 335378
rect 240152 318170 240180 340068
rect 240244 338026 240272 340068
rect 240232 338020 240284 338026
rect 240232 337962 240284 337968
rect 240232 337884 240284 337890
rect 240232 337826 240284 337832
rect 240244 334830 240272 337826
rect 240324 337544 240376 337550
rect 240324 337486 240376 337492
rect 240336 336598 240364 337486
rect 240324 336592 240376 336598
rect 240324 336534 240376 336540
rect 240324 335708 240376 335714
rect 240324 335650 240376 335656
rect 240232 334824 240284 334830
rect 240232 334766 240284 334772
rect 240232 334620 240284 334626
rect 240232 334562 240284 334568
rect 240244 325038 240272 334562
rect 240232 325032 240284 325038
rect 240232 324974 240284 324980
rect 240140 318164 240192 318170
rect 240140 318106 240192 318112
rect 240336 8702 240364 335650
rect 240428 8770 240456 340068
rect 240520 334626 240548 340068
rect 240626 340054 240732 340082
rect 240704 335646 240732 340054
rect 240796 335714 240824 340068
rect 240784 335708 240836 335714
rect 240784 335650 240836 335656
rect 240692 335640 240744 335646
rect 240692 335582 240744 335588
rect 240508 334620 240560 334626
rect 240508 334562 240560 334568
rect 240888 334506 240916 340068
rect 240980 338094 241008 340068
rect 240968 338088 241020 338094
rect 240968 338030 241020 338036
rect 240968 336796 241020 336802
rect 240968 336738 241020 336744
rect 240520 334478 240916 334506
rect 240520 309806 240548 334478
rect 240692 334416 240744 334422
rect 240980 334370 241008 336738
rect 241060 335640 241112 335646
rect 241060 335582 241112 335588
rect 240692 334358 240744 334364
rect 240704 316742 240732 334358
rect 240796 334342 241008 334370
rect 240796 323678 240824 334342
rect 240784 323672 240836 323678
rect 240784 323614 240836 323620
rect 240692 316736 240744 316742
rect 240692 316678 240744 316684
rect 240508 309800 240560 309806
rect 240508 309742 240560 309748
rect 240416 8764 240468 8770
rect 240416 8706 240468 8712
rect 240324 8696 240376 8702
rect 240324 8638 240376 8644
rect 240784 4956 240836 4962
rect 240784 4898 240836 4904
rect 240048 4140 240100 4146
rect 240048 4082 240100 4088
rect 239956 3052 240008 3058
rect 239956 2994 240008 3000
rect 240796 480 240824 4898
rect 241072 2990 241100 335582
rect 241164 8634 241192 340068
rect 241256 334422 241284 340068
rect 241244 334416 241296 334422
rect 241244 334358 241296 334364
rect 241152 8628 241204 8634
rect 241152 8570 241204 8576
rect 241348 3738 241376 340068
rect 241532 333810 241560 340068
rect 241624 336802 241652 340068
rect 241716 337822 241744 340068
rect 241808 340054 241914 340082
rect 241704 337816 241756 337822
rect 241704 337758 241756 337764
rect 241612 336796 241664 336802
rect 241612 336738 241664 336744
rect 241520 333804 241572 333810
rect 241520 333746 241572 333752
rect 241808 8498 241836 340054
rect 241992 337278 242020 340068
rect 241980 337272 242032 337278
rect 241980 337214 242032 337220
rect 241888 333804 241940 333810
rect 241888 333746 241940 333752
rect 241900 8566 241928 333746
rect 241980 8968 242032 8974
rect 241980 8910 242032 8916
rect 241888 8560 241940 8566
rect 241888 8502 241940 8508
rect 241796 8492 241848 8498
rect 241796 8434 241848 8440
rect 241336 3732 241388 3738
rect 241336 3674 241388 3680
rect 241060 2984 241112 2990
rect 241060 2926 241112 2932
rect 241992 480 242020 8910
rect 242084 2922 242112 340068
rect 242164 335640 242216 335646
rect 242164 335582 242216 335588
rect 242072 2916 242124 2922
rect 242072 2858 242124 2864
rect 242176 2854 242204 335582
rect 242268 8430 242296 340068
rect 242360 322318 242388 340068
rect 242452 335646 242480 340068
rect 242440 335640 242492 335646
rect 242440 335582 242492 335588
rect 242532 335640 242584 335646
rect 242532 335582 242584 335588
rect 242348 322312 242400 322318
rect 242348 322254 242400 322260
rect 242544 320958 242572 335582
rect 242532 320952 242584 320958
rect 242532 320894 242584 320900
rect 242256 8424 242308 8430
rect 242256 8366 242308 8372
rect 242636 8362 242664 340068
rect 242728 335646 242756 340068
rect 242820 337754 242848 340068
rect 242808 337748 242860 337754
rect 242808 337690 242860 337696
rect 243004 337550 243032 340068
rect 242992 337544 243044 337550
rect 242992 337486 243044 337492
rect 242900 337476 242952 337482
rect 242900 337418 242952 337424
rect 242912 336394 242940 337418
rect 242992 337272 243044 337278
rect 242992 337214 243044 337220
rect 242900 336388 242952 336394
rect 242900 336330 242952 336336
rect 242900 335844 242952 335850
rect 242900 335786 242952 335792
rect 242716 335640 242768 335646
rect 242716 335582 242768 335588
rect 242912 333402 242940 335786
rect 243004 334762 243032 337214
rect 242992 334756 243044 334762
rect 242992 334698 243044 334704
rect 242900 333396 242952 333402
rect 242900 333338 242952 333344
rect 243096 330682 243124 340068
rect 243188 335850 243216 340068
rect 243176 335844 243228 335850
rect 243176 335786 243228 335792
rect 243176 335708 243228 335714
rect 243176 335650 243228 335656
rect 243084 330676 243136 330682
rect 243084 330618 243136 330624
rect 242624 8356 242676 8362
rect 242624 8298 242676 8304
rect 243188 6322 243216 335650
rect 243268 335640 243320 335646
rect 243268 335582 243320 335588
rect 243176 6316 243228 6322
rect 243176 6258 243228 6264
rect 243280 6254 243308 335582
rect 243372 335458 243400 340068
rect 243464 335646 243492 340068
rect 243452 335640 243504 335646
rect 243452 335582 243504 335588
rect 243372 335430 243492 335458
rect 243360 292596 243412 292602
rect 243360 292538 243412 292544
rect 243372 234598 243400 292538
rect 243360 234592 243412 234598
rect 243360 234534 243412 234540
rect 243360 215348 243412 215354
rect 243360 215290 243412 215296
rect 243372 99346 243400 215290
rect 243360 99340 243412 99346
rect 243360 99282 243412 99288
rect 243360 70440 243412 70446
rect 243360 70382 243412 70388
rect 243372 7614 243400 70382
rect 243360 7608 243412 7614
rect 243360 7550 243412 7556
rect 243268 6248 243320 6254
rect 243268 6190 243320 6196
rect 243464 5098 243492 335430
rect 243556 292670 243584 340068
rect 243544 292664 243596 292670
rect 243544 292606 243596 292612
rect 243544 234592 243596 234598
rect 243544 234534 243596 234540
rect 243556 215422 243584 234534
rect 243544 215416 243596 215422
rect 243544 215358 243596 215364
rect 243544 99340 243596 99346
rect 243544 99282 243596 99288
rect 243556 70446 243584 99282
rect 243544 70440 243596 70446
rect 243544 70382 243596 70388
rect 243740 5166 243768 340068
rect 243832 335714 243860 340068
rect 243820 335708 243872 335714
rect 243820 335650 243872 335656
rect 243924 318238 243952 340068
rect 244016 340054 244122 340082
rect 243912 318232 243964 318238
rect 243912 318174 243964 318180
rect 244016 5234 244044 340054
rect 244200 327894 244228 340068
rect 244306 340054 244412 340082
rect 244280 336796 244332 336802
rect 244280 336738 244332 336744
rect 244292 329254 244320 336738
rect 244384 332738 244412 340054
rect 244476 333470 244504 340068
rect 244464 333464 244516 333470
rect 244464 333406 244516 333412
rect 244568 332874 244596 340068
rect 244674 340054 244780 340082
rect 244752 335594 244780 340054
rect 244844 335714 244872 340068
rect 244832 335708 244884 335714
rect 244832 335650 244884 335656
rect 244936 335646 244964 340068
rect 244924 335640 244976 335646
rect 244752 335566 244872 335594
rect 244924 335582 244976 335588
rect 244568 332846 244780 332874
rect 244384 332710 244596 332738
rect 244372 332648 244424 332654
rect 244372 332590 244424 332596
rect 244384 330750 244412 332590
rect 244372 330744 244424 330750
rect 244372 330686 244424 330692
rect 244280 329248 244332 329254
rect 244280 329190 244332 329196
rect 244188 327888 244240 327894
rect 244188 327830 244240 327836
rect 244568 316810 244596 332710
rect 244752 325106 244780 332846
rect 244740 325100 244792 325106
rect 244740 325042 244792 325048
rect 244556 316804 244608 316810
rect 244556 316746 244608 316752
rect 244844 315382 244872 335566
rect 244832 315376 244884 315382
rect 244832 315318 244884 315324
rect 245028 314022 245056 340068
rect 245120 337210 245148 340068
rect 245108 337204 245160 337210
rect 245108 337146 245160 337152
rect 245108 335708 245160 335714
rect 245108 335650 245160 335656
rect 245120 332042 245148 335650
rect 245108 332036 245160 332042
rect 245108 331978 245160 331984
rect 245304 323354 245332 340068
rect 245396 328438 245424 340068
rect 245488 332654 245516 340068
rect 245568 335640 245620 335646
rect 245568 335582 245620 335588
rect 245476 332648 245528 332654
rect 245476 332590 245528 332596
rect 245384 328432 245436 328438
rect 245384 328374 245436 328380
rect 245212 323326 245332 323354
rect 245212 321026 245240 323326
rect 245580 322386 245608 335582
rect 245672 332110 245700 340068
rect 245764 334150 245792 340068
rect 245856 336802 245884 340068
rect 245844 336796 245896 336802
rect 245844 336738 245896 336744
rect 245936 335640 245988 335646
rect 245936 335582 245988 335588
rect 245752 334144 245804 334150
rect 245752 334086 245804 334092
rect 245660 332104 245712 332110
rect 245660 332046 245712 332052
rect 245948 323746 245976 335582
rect 246040 329322 246068 340068
rect 246028 329316 246080 329322
rect 246028 329258 246080 329264
rect 245936 323740 245988 323746
rect 245936 323682 245988 323688
rect 245568 322380 245620 322386
rect 245568 322322 245620 322328
rect 245200 321020 245252 321026
rect 245200 320962 245252 320968
rect 245200 320340 245252 320346
rect 245200 320282 245252 320288
rect 245212 318782 245240 320282
rect 245200 318776 245252 318782
rect 245200 318718 245252 318724
rect 245016 314016 245068 314022
rect 245016 313958 245068 313964
rect 246132 312662 246160 340068
rect 246224 337278 246252 340068
rect 246212 337272 246264 337278
rect 246212 337214 246264 337220
rect 246212 334144 246264 334150
rect 246212 334086 246264 334092
rect 246224 319530 246252 334086
rect 246408 326534 246436 340068
rect 246396 326528 246448 326534
rect 246396 326470 246448 326476
rect 246212 319524 246264 319530
rect 246212 319466 246264 319472
rect 246120 312656 246172 312662
rect 246120 312598 246172 312604
rect 245200 311840 245252 311846
rect 245200 311782 245252 311788
rect 245212 225026 245240 311782
rect 246500 311234 246528 340068
rect 246592 337890 246620 340068
rect 246580 337884 246632 337890
rect 246580 337826 246632 337832
rect 246776 337074 246804 340068
rect 246764 337068 246816 337074
rect 246764 337010 246816 337016
rect 246868 335646 246896 340068
rect 246960 337618 246988 340068
rect 246948 337612 247000 337618
rect 246948 337554 247000 337560
rect 246948 337068 247000 337074
rect 246948 337010 247000 337016
rect 246856 335640 246908 335646
rect 246856 335582 246908 335588
rect 246960 335102 246988 337010
rect 246948 335096 247000 335102
rect 246948 335038 247000 335044
rect 247144 327962 247172 340068
rect 247236 333554 247264 340068
rect 247328 336258 247356 340068
rect 247408 338224 247460 338230
rect 247408 338166 247460 338172
rect 247316 336252 247368 336258
rect 247316 336194 247368 336200
rect 247420 333674 247448 338166
rect 247512 333690 247540 340068
rect 247604 335646 247632 340068
rect 247696 338230 247724 340068
rect 247788 340054 247894 340082
rect 247684 338224 247736 338230
rect 247684 338166 247736 338172
rect 247684 338088 247736 338094
rect 247684 338030 247736 338036
rect 247592 335640 247644 335646
rect 247592 335582 247644 335588
rect 247408 333668 247460 333674
rect 247512 333662 247632 333690
rect 247408 333610 247460 333616
rect 247236 333526 247540 333554
rect 247316 333464 247368 333470
rect 247316 333406 247368 333412
rect 247132 327956 247184 327962
rect 247132 327898 247184 327904
rect 246488 311228 246540 311234
rect 246488 311170 246540 311176
rect 245120 224998 245240 225026
rect 245120 224890 245148 224998
rect 245120 224862 245240 224890
rect 245212 222193 245240 224862
rect 245014 222184 245070 222193
rect 245014 222119 245070 222128
rect 245198 222184 245254 222193
rect 245198 222119 245254 222128
rect 245028 212566 245056 222119
rect 245016 212560 245068 212566
rect 245016 212502 245068 212508
rect 245200 212560 245252 212566
rect 245200 212502 245252 212508
rect 245212 202881 245240 212502
rect 245014 202872 245070 202881
rect 245014 202807 245070 202816
rect 245198 202872 245254 202881
rect 245198 202807 245254 202816
rect 245028 193254 245056 202807
rect 245016 193248 245068 193254
rect 245016 193190 245068 193196
rect 245200 193248 245252 193254
rect 245200 193190 245252 193196
rect 245212 183569 245240 193190
rect 245014 183560 245070 183569
rect 245014 183495 245070 183504
rect 245198 183560 245254 183569
rect 245198 183495 245254 183504
rect 245028 180810 245056 183495
rect 245016 180804 245068 180810
rect 245016 180746 245068 180752
rect 245292 171148 245344 171154
rect 245292 171090 245344 171096
rect 245304 161430 245332 171090
rect 245292 161424 245344 161430
rect 245292 161366 245344 161372
rect 245016 151836 245068 151842
rect 245016 151778 245068 151784
rect 245028 143585 245056 151778
rect 245014 143576 245070 143585
rect 245014 143511 245070 143520
rect 245198 143576 245254 143585
rect 245198 143511 245254 143520
rect 245212 138718 245240 143511
rect 245200 138712 245252 138718
rect 245200 138654 245252 138660
rect 245384 135176 245436 135182
rect 245384 135118 245436 135124
rect 245396 133906 245424 135118
rect 245396 133878 245516 133906
rect 245488 128330 245516 133878
rect 245396 128302 245516 128330
rect 245396 125526 245424 128302
rect 245108 125520 245160 125526
rect 245108 125462 245160 125468
rect 245384 125520 245436 125526
rect 245384 125462 245436 125468
rect 245120 124166 245148 125462
rect 245108 124160 245160 124166
rect 245108 124102 245160 124108
rect 245108 114572 245160 114578
rect 245108 114514 245160 114520
rect 245120 109070 245148 114514
rect 245108 109064 245160 109070
rect 245108 109006 245160 109012
rect 245200 108996 245252 109002
rect 245200 108938 245252 108944
rect 245212 106162 245240 108938
rect 245212 106134 245332 106162
rect 245304 89706 245332 106134
rect 245212 89678 245332 89706
rect 245212 85542 245240 89678
rect 245200 85536 245252 85542
rect 245200 85478 245252 85484
rect 245200 75948 245252 75954
rect 245200 75890 245252 75896
rect 245212 70514 245240 75890
rect 245200 70508 245252 70514
rect 245200 70450 245252 70456
rect 245108 67652 245160 67658
rect 245108 67594 245160 67600
rect 245120 64954 245148 67594
rect 245120 64926 245332 64954
rect 245304 57934 245332 64926
rect 245292 57928 245344 57934
rect 245292 57870 245344 57876
rect 245200 48340 245252 48346
rect 245200 48282 245252 48288
rect 245212 41426 245240 48282
rect 245212 41398 245332 41426
rect 245304 15910 245332 41398
rect 245292 15904 245344 15910
rect 245292 15846 245344 15852
rect 247328 7818 247356 333406
rect 247408 333396 247460 333402
rect 247408 333338 247460 333344
rect 247420 7886 247448 333338
rect 247408 7880 247460 7886
rect 247408 7822 247460 7828
rect 247316 7812 247368 7818
rect 247316 7754 247368 7760
rect 247512 7682 247540 333526
rect 247604 326602 247632 333662
rect 247592 326596 247644 326602
rect 247592 326538 247644 326544
rect 247500 7676 247552 7682
rect 247500 7618 247552 7624
rect 244004 5228 244056 5234
rect 244004 5170 244056 5176
rect 247696 5166 247724 338030
rect 247788 6390 247816 340054
rect 247868 335640 247920 335646
rect 247868 335582 247920 335588
rect 247880 7750 247908 335582
rect 247972 333470 248000 340068
rect 248064 334898 248092 340068
rect 248156 340054 248262 340082
rect 248052 334892 248104 334898
rect 248052 334834 248104 334840
rect 247960 333464 248012 333470
rect 247960 333406 248012 333412
rect 247868 7744 247920 7750
rect 247868 7686 247920 7692
rect 248156 6458 248184 340054
rect 248340 333402 248368 340068
rect 248432 336326 248460 340068
rect 248512 337000 248564 337006
rect 248512 336942 248564 336948
rect 248420 336320 248472 336326
rect 248420 336262 248472 336268
rect 248524 335594 248552 336942
rect 248432 335566 248552 335594
rect 248328 333396 248380 333402
rect 248328 333338 248380 333344
rect 248432 330818 248460 335566
rect 248420 330812 248472 330818
rect 248420 330754 248472 330760
rect 248418 228032 248474 228041
rect 248418 227967 248474 227976
rect 248432 227905 248460 227967
rect 248418 227896 248474 227905
rect 248418 227831 248474 227840
rect 248616 6526 248644 340068
rect 248708 335594 248736 340068
rect 248800 335714 248828 340068
rect 248892 340054 248998 340082
rect 248892 335782 248920 340054
rect 248880 335776 248932 335782
rect 248880 335718 248932 335724
rect 248788 335708 248840 335714
rect 248788 335650 248840 335656
rect 248880 335640 248932 335646
rect 248708 335566 248828 335594
rect 248880 335582 248932 335588
rect 248696 335504 248748 335510
rect 248696 335446 248748 335452
rect 248708 8022 248736 335446
rect 248696 8016 248748 8022
rect 248696 7958 248748 7964
rect 248800 7954 248828 335566
rect 248788 7948 248840 7954
rect 248788 7890 248840 7896
rect 248892 6594 248920 335582
rect 249076 335510 249104 340068
rect 249182 340054 249288 340082
rect 249260 335646 249288 340054
rect 249248 335640 249300 335646
rect 249248 335582 249300 335588
rect 249064 335504 249116 335510
rect 249064 335446 249116 335452
rect 249352 6662 249380 340068
rect 249444 8090 249472 340068
rect 249432 8084 249484 8090
rect 249432 8026 249484 8032
rect 249340 6656 249392 6662
rect 249340 6598 249392 6604
rect 248880 6588 248932 6594
rect 248880 6530 248932 6536
rect 248604 6520 248656 6526
rect 248604 6462 248656 6468
rect 248144 6452 248196 6458
rect 248144 6394 248196 6400
rect 247776 6384 247828 6390
rect 247776 6326 247828 6332
rect 249536 5370 249564 340068
rect 249616 335640 249668 335646
rect 249616 335582 249668 335588
rect 249524 5364 249576 5370
rect 249524 5306 249576 5312
rect 249628 5302 249656 335582
rect 249720 6730 249748 340068
rect 249812 335594 249840 340068
rect 249918 340054 250024 340082
rect 249812 335566 249932 335594
rect 249800 335504 249852 335510
rect 249800 335446 249852 335452
rect 249708 6724 249760 6730
rect 249708 6666 249760 6672
rect 249812 5438 249840 335446
rect 249904 8158 249932 335566
rect 249892 8152 249944 8158
rect 249892 8094 249944 8100
rect 249800 5432 249852 5438
rect 249800 5374 249852 5380
rect 249616 5296 249668 5302
rect 249616 5238 249668 5244
rect 249996 5234 250024 340054
rect 250088 6798 250116 340068
rect 250180 8226 250208 340068
rect 250272 335510 250300 340068
rect 250364 340054 250470 340082
rect 250260 335504 250312 335510
rect 250260 335446 250312 335452
rect 250258 280120 250314 280129
rect 250258 280055 250314 280064
rect 250272 273154 250300 280055
rect 250260 273148 250312 273154
rect 250260 273090 250312 273096
rect 250168 8220 250220 8226
rect 250168 8162 250220 8168
rect 250364 6866 250392 340054
rect 250548 333334 250576 340068
rect 250654 340054 250760 340082
rect 250732 335646 250760 340054
rect 250720 335640 250772 335646
rect 250720 335582 250772 335588
rect 250536 333328 250588 333334
rect 250536 333270 250588 333276
rect 250628 328500 250680 328506
rect 250628 328442 250680 328448
rect 250640 311794 250668 328442
rect 250640 311766 250760 311794
rect 250732 280226 250760 311766
rect 250536 280220 250588 280226
rect 250536 280162 250588 280168
rect 250720 280220 250772 280226
rect 250720 280162 250772 280168
rect 250442 280120 250498 280129
rect 250548 280106 250576 280162
rect 250498 280078 250576 280106
rect 250442 280055 250498 280064
rect 250720 273148 250772 273154
rect 250720 273090 250772 273096
rect 250732 261089 250760 273090
rect 250718 261080 250774 261089
rect 250718 261015 250774 261024
rect 250442 260944 250498 260953
rect 250442 260879 250498 260888
rect 250456 260846 250484 260879
rect 250444 260840 250496 260846
rect 250444 260782 250496 260788
rect 250720 253836 250772 253842
rect 250720 253778 250772 253784
rect 250732 234666 250760 253778
rect 250720 234660 250772 234666
rect 250720 234602 250772 234608
rect 250720 234524 250772 234530
rect 250720 234466 250772 234472
rect 250732 225026 250760 234466
rect 250640 224998 250760 225026
rect 250640 224890 250668 224998
rect 250640 224862 250760 224890
rect 250732 205714 250760 224862
rect 250640 205686 250760 205714
rect 250640 205578 250668 205686
rect 250640 205550 250760 205578
rect 250732 186402 250760 205550
rect 250640 186374 250760 186402
rect 250640 186266 250668 186374
rect 250640 186238 250760 186266
rect 250732 167090 250760 186238
rect 250640 167062 250760 167090
rect 250640 166954 250668 167062
rect 250640 166926 250760 166954
rect 250732 142361 250760 166926
rect 250718 142352 250774 142361
rect 250718 142287 250774 142296
rect 250626 142216 250682 142225
rect 250626 142151 250682 142160
rect 250640 140758 250668 142151
rect 250628 140752 250680 140758
rect 250628 140694 250680 140700
rect 250536 128308 250588 128314
rect 250536 128250 250588 128256
rect 250548 125610 250576 128250
rect 250548 125582 250668 125610
rect 250640 125526 250668 125582
rect 250628 125520 250680 125526
rect 250628 125462 250680 125468
rect 250720 125520 250772 125526
rect 250720 125462 250772 125468
rect 250732 111790 250760 125462
rect 250720 111784 250772 111790
rect 250720 111726 250772 111732
rect 250628 102196 250680 102202
rect 250628 102138 250680 102144
rect 250640 82822 250668 102138
rect 250628 82816 250680 82822
rect 250628 82758 250680 82764
rect 250444 68332 250496 68338
rect 250444 68274 250496 68280
rect 250456 58018 250484 68274
rect 250456 57990 250576 58018
rect 250548 48362 250576 57990
rect 250456 48334 250576 48362
rect 250456 44169 250484 48334
rect 250442 44160 250498 44169
rect 250442 44095 250498 44104
rect 250718 44160 250774 44169
rect 250718 44095 250774 44104
rect 250732 19394 250760 44095
rect 250548 19366 250760 19394
rect 250548 19310 250576 19366
rect 250536 19304 250588 19310
rect 250536 19246 250588 19252
rect 250444 9716 250496 9722
rect 250444 9658 250496 9664
rect 250456 9602 250484 9658
rect 250456 9574 250576 9602
rect 250548 8294 250576 9574
rect 250536 8288 250588 8294
rect 250536 8230 250588 8236
rect 250352 6860 250404 6866
rect 250352 6802 250404 6808
rect 250076 6792 250128 6798
rect 250076 6734 250128 6740
rect 250824 6118 250852 340068
rect 250916 77246 250944 340068
rect 250904 77240 250956 77246
rect 250904 77182 250956 77188
rect 251008 77178 251036 340068
rect 251192 335646 251220 340068
rect 251284 337006 251312 340068
rect 251376 337482 251404 340068
rect 251468 340054 251574 340082
rect 251364 337476 251416 337482
rect 251364 337418 251416 337424
rect 251272 337000 251324 337006
rect 251272 336942 251324 336948
rect 251272 336864 251324 336870
rect 251272 336806 251324 336812
rect 251088 335640 251140 335646
rect 251088 335582 251140 335588
rect 251180 335640 251232 335646
rect 251180 335582 251232 335588
rect 251100 77246 251128 335582
rect 251284 335458 251312 336806
rect 251468 335730 251496 340054
rect 251192 335430 251312 335458
rect 251376 335702 251496 335730
rect 251088 77240 251140 77246
rect 251088 77182 251140 77188
rect 250996 77172 251048 77178
rect 250996 77114 251048 77120
rect 250904 72480 250956 72486
rect 250904 72422 250956 72428
rect 250916 7546 250944 72422
rect 250996 71732 251048 71738
rect 250996 71674 251048 71680
rect 250904 7540 250956 7546
rect 250904 7482 250956 7488
rect 250812 6112 250864 6118
rect 250812 6054 250864 6060
rect 249984 5228 250036 5234
rect 249984 5170 250036 5176
rect 243728 5160 243780 5166
rect 243728 5102 243780 5108
rect 244372 5160 244424 5166
rect 244372 5102 244424 5108
rect 247684 5160 247736 5166
rect 247684 5102 247736 5108
rect 243452 5092 243504 5098
rect 243452 5034 243504 5040
rect 243176 4072 243228 4078
rect 243176 4014 243228 4020
rect 242164 2848 242216 2854
rect 242164 2790 242216 2796
rect 243188 480 243216 4014
rect 244384 480 244412 5102
rect 251008 4690 251036 71674
rect 251088 70440 251140 70446
rect 251088 70382 251140 70388
rect 251100 4758 251128 70382
rect 251192 10334 251220 335430
rect 251376 332246 251404 335702
rect 251548 335640 251600 335646
rect 251548 335582 251600 335588
rect 251456 335504 251508 335510
rect 251456 335446 251508 335452
rect 251364 332240 251416 332246
rect 251364 332182 251416 332188
rect 251468 325174 251496 335446
rect 251560 329390 251588 335582
rect 251652 335306 251680 340068
rect 251744 335986 251772 340068
rect 251836 340054 251942 340082
rect 251732 335980 251784 335986
rect 251732 335922 251784 335928
rect 251836 335866 251864 340054
rect 251744 335838 251864 335866
rect 251744 335510 251772 335838
rect 251732 335504 251784 335510
rect 251732 335446 251784 335452
rect 251640 335300 251692 335306
rect 251640 335242 251692 335248
rect 252020 335186 252048 340068
rect 252126 340054 252232 340082
rect 252204 337006 252232 340054
rect 252192 337000 252244 337006
rect 252192 336942 252244 336948
rect 251652 335158 252048 335186
rect 251548 329384 251600 329390
rect 251548 329326 251600 329332
rect 251652 328030 251680 335158
rect 251732 335096 251784 335102
rect 251732 335038 251784 335044
rect 251640 328024 251692 328030
rect 251640 327966 251692 327972
rect 251456 325168 251508 325174
rect 251456 325110 251508 325116
rect 251744 319598 251772 335038
rect 251916 334008 251968 334014
rect 251916 333950 251968 333956
rect 251824 329044 251876 329050
rect 251824 328986 251876 328992
rect 251732 319592 251784 319598
rect 251732 319534 251784 319540
rect 251180 10328 251232 10334
rect 251180 10270 251232 10276
rect 251836 8974 251864 328986
rect 251928 326398 251956 333950
rect 252296 333826 252324 340068
rect 252388 334014 252416 340068
rect 252480 336462 252508 340068
rect 252560 337000 252612 337006
rect 252560 336942 252612 336948
rect 252468 336456 252520 336462
rect 252468 336398 252520 336404
rect 252572 336274 252600 336942
rect 252480 336246 252600 336274
rect 252376 334008 252428 334014
rect 252376 333950 252428 333956
rect 252296 333798 252416 333826
rect 252008 328500 252060 328506
rect 252008 328442 252060 328448
rect 251916 326392 251968 326398
rect 251916 326334 251968 326340
rect 252020 11762 252048 328442
rect 252100 326392 252152 326398
rect 252100 326334 252152 326340
rect 252112 311794 252140 326334
rect 252388 323814 252416 333798
rect 252480 333742 252508 336246
rect 252664 333810 252692 340068
rect 252652 333804 252704 333810
rect 252652 333746 252704 333752
rect 252468 333736 252520 333742
rect 252468 333678 252520 333684
rect 252756 326670 252784 340068
rect 252848 335034 252876 340068
rect 252940 340054 253046 340082
rect 252940 337074 252968 340054
rect 253020 338156 253072 338162
rect 253020 338098 253072 338104
rect 253032 337414 253060 338098
rect 253020 337408 253072 337414
rect 253020 337350 253072 337356
rect 252928 337068 252980 337074
rect 252928 337010 252980 337016
rect 252928 335640 252980 335646
rect 252928 335582 252980 335588
rect 252836 335028 252888 335034
rect 252836 334970 252888 334976
rect 252744 326664 252796 326670
rect 252744 326606 252796 326612
rect 252376 323808 252428 323814
rect 252376 323750 252428 323756
rect 252112 311766 252232 311794
rect 252204 296682 252232 311766
rect 252192 296676 252244 296682
rect 252192 296618 252244 296624
rect 252284 296676 252336 296682
rect 252284 296618 252336 296624
rect 252296 251326 252324 296618
rect 252284 251320 252336 251326
rect 252284 251262 252336 251268
rect 252192 249824 252244 249830
rect 252192 249766 252244 249772
rect 252204 244338 252232 249766
rect 252112 244310 252232 244338
rect 252112 244254 252140 244310
rect 252100 244248 252152 244254
rect 252100 244190 252152 244196
rect 252284 244248 252336 244254
rect 252284 244190 252336 244196
rect 252296 229106 252324 244190
rect 252204 229078 252324 229106
rect 252204 208350 252232 229078
rect 252192 208344 252244 208350
rect 252192 208286 252244 208292
rect 252284 198756 252336 198762
rect 252284 198698 252336 198704
rect 252296 189106 252324 198698
rect 252100 189100 252152 189106
rect 252100 189042 252152 189048
rect 252284 189100 252336 189106
rect 252284 189042 252336 189048
rect 252112 186318 252140 189042
rect 252100 186312 252152 186318
rect 252100 186254 252152 186260
rect 252192 176724 252244 176730
rect 252192 176666 252244 176672
rect 252204 174010 252232 176666
rect 252192 174004 252244 174010
rect 252192 173946 252244 173952
rect 252192 168360 252244 168366
rect 252192 168302 252244 168308
rect 252204 164898 252232 168302
rect 252192 164892 252244 164898
rect 252192 164834 252244 164840
rect 252008 11756 252060 11762
rect 252008 11698 252060 11704
rect 252940 10402 252968 335582
rect 253124 322454 253152 340068
rect 253216 338162 253244 340068
rect 253308 340054 253414 340082
rect 253204 338156 253256 338162
rect 253204 338098 253256 338104
rect 253204 337952 253256 337958
rect 253204 337894 253256 337900
rect 253112 322448 253164 322454
rect 253112 322390 253164 322396
rect 253216 10470 253244 337894
rect 253308 330886 253336 340054
rect 253296 330880 253348 330886
rect 253296 330822 253348 330828
rect 253492 328506 253520 340068
rect 253584 336530 253612 340068
rect 253768 336870 253796 340068
rect 253756 336864 253808 336870
rect 253756 336806 253808 336812
rect 253572 336524 253624 336530
rect 253572 336466 253624 336472
rect 253860 335646 253888 340068
rect 253966 340054 254072 340082
rect 253848 335640 253900 335646
rect 253848 335582 253900 335588
rect 254044 333538 254072 340054
rect 254136 335850 254164 340068
rect 254228 337958 254256 340068
rect 254216 337952 254268 337958
rect 254216 337894 254268 337900
rect 254124 335844 254176 335850
rect 254124 335786 254176 335792
rect 254320 335730 254348 340068
rect 254136 335702 254348 335730
rect 254412 340054 254518 340082
rect 254032 333532 254084 333538
rect 254032 333474 254084 333480
rect 253480 328500 253532 328506
rect 253480 328442 253532 328448
rect 253204 10464 253256 10470
rect 253204 10406 253256 10412
rect 252928 10396 252980 10402
rect 252928 10338 252980 10344
rect 251824 8968 251876 8974
rect 251824 8910 251876 8916
rect 253848 8288 253900 8294
rect 253848 8230 253900 8236
rect 251088 4752 251140 4758
rect 251088 4694 251140 4700
rect 250996 4684 251048 4690
rect 250996 4626 251048 4632
rect 250352 3868 250404 3874
rect 250352 3810 250404 3816
rect 247960 3664 248012 3670
rect 247960 3606 248012 3612
rect 245568 3596 245620 3602
rect 245568 3538 245620 3544
rect 245580 480 245608 3538
rect 246764 3392 246816 3398
rect 246764 3334 246816 3340
rect 246776 480 246804 3334
rect 247972 480 248000 3606
rect 249156 2984 249208 2990
rect 249156 2926 249208 2932
rect 249168 480 249196 2926
rect 250364 480 250392 3810
rect 252652 3460 252704 3466
rect 252652 3402 252704 3408
rect 251456 604 251508 610
rect 251456 546 251508 552
rect 251468 480 251496 546
rect 252664 480 252692 3402
rect 253860 480 253888 8230
rect 254136 4894 254164 335702
rect 254308 335640 254360 335646
rect 254308 335582 254360 335588
rect 254216 333532 254268 333538
rect 254216 333474 254268 333480
rect 254124 4888 254176 4894
rect 254124 4830 254176 4836
rect 254228 4826 254256 333474
rect 254320 4962 254348 335582
rect 254412 6050 254440 340054
rect 254596 337142 254624 340068
rect 254584 337136 254636 337142
rect 254584 337078 254636 337084
rect 254584 336796 254636 336802
rect 254584 336738 254636 336744
rect 254492 335844 254544 335850
rect 254492 335786 254544 335792
rect 254504 6186 254532 335786
rect 254492 6180 254544 6186
rect 254492 6122 254544 6128
rect 254400 6044 254452 6050
rect 254400 5986 254452 5992
rect 254308 4956 254360 4962
rect 254308 4898 254360 4904
rect 254216 4820 254268 4826
rect 254216 4762 254268 4768
rect 254596 3670 254624 336738
rect 254688 335646 254716 340068
rect 254676 335640 254728 335646
rect 254676 335582 254728 335588
rect 254872 329050 254900 340068
rect 254964 333946 254992 340068
rect 255056 338094 255084 340068
rect 255044 338088 255096 338094
rect 255044 338030 255096 338036
rect 254952 333940 255004 333946
rect 254952 333882 255004 333888
rect 254860 329044 254912 329050
rect 254860 328986 254912 328992
rect 254676 328500 254728 328506
rect 254676 328442 254728 328448
rect 254584 3664 254636 3670
rect 254584 3606 254636 3612
rect 254688 610 254716 328442
rect 254860 316124 254912 316130
rect 254860 316066 254912 316072
rect 254872 314673 254900 316066
rect 254858 314664 254914 314673
rect 254858 314599 254914 314608
rect 254766 305008 254822 305017
rect 254766 304943 254768 304952
rect 254820 304943 254822 304952
rect 255044 304972 255096 304978
rect 254768 304914 254820 304920
rect 255044 304914 255096 304920
rect 255056 295361 255084 304914
rect 254858 295352 254914 295361
rect 254858 295287 254860 295296
rect 254912 295287 254914 295296
rect 255042 295352 255098 295361
rect 255042 295287 255098 295296
rect 254860 295258 254912 295264
rect 254860 285728 254912 285734
rect 254860 285670 254912 285676
rect 254872 280786 254900 285670
rect 254872 280758 255084 280786
rect 255056 280106 255084 280758
rect 254964 280078 255084 280106
rect 254964 259434 254992 280078
rect 254872 259406 254992 259434
rect 254872 251258 254900 259406
rect 254860 251252 254912 251258
rect 254860 251194 254912 251200
rect 254860 249824 254912 249830
rect 254860 249766 254912 249772
rect 254872 231690 254900 249766
rect 254780 231662 254900 231690
rect 254780 222222 254808 231662
rect 254768 222216 254820 222222
rect 254768 222158 254820 222164
rect 254860 222148 254912 222154
rect 254860 222090 254912 222096
rect 254872 218226 254900 222090
rect 254872 218198 254992 218226
rect 254964 202910 254992 218198
rect 254860 202904 254912 202910
rect 254860 202846 254912 202852
rect 254952 202904 255004 202910
rect 254952 202846 255004 202852
rect 254872 189258 254900 202846
rect 254780 189230 254900 189258
rect 254780 189038 254808 189230
rect 254768 189032 254820 189038
rect 254768 188974 254820 188980
rect 254952 179444 255004 179450
rect 254952 179386 255004 179392
rect 254964 168366 254992 179386
rect 254952 168360 255004 168366
rect 254952 168302 255004 168308
rect 254860 158772 254912 158778
rect 254860 158714 254912 158720
rect 254872 150482 254900 158714
rect 254860 150476 254912 150482
rect 254860 150418 254912 150424
rect 255044 150476 255096 150482
rect 255044 150418 255096 150424
rect 255056 142066 255084 150418
rect 254964 142038 255084 142066
rect 254964 140758 254992 142038
rect 254952 140752 255004 140758
rect 254952 140694 255004 140700
rect 255044 140752 255096 140758
rect 255044 140694 255096 140700
rect 255056 135232 255084 140694
rect 254964 135204 255084 135232
rect 254964 125662 254992 135204
rect 254952 125656 255004 125662
rect 254952 125598 255004 125604
rect 254860 125588 254912 125594
rect 254860 125530 254912 125536
rect 254872 124166 254900 125530
rect 254860 124160 254912 124166
rect 254860 124102 254912 124108
rect 255136 124160 255188 124166
rect 255136 124102 255188 124108
rect 255148 122806 255176 124102
rect 255136 122800 255188 122806
rect 255136 122742 255188 122748
rect 255044 113212 255096 113218
rect 255044 113154 255096 113160
rect 255056 106162 255084 113154
rect 254872 106134 255084 106162
rect 254872 104854 254900 106134
rect 254860 104848 254912 104854
rect 254860 104790 254912 104796
rect 255044 95260 255096 95266
rect 255044 95202 255096 95208
rect 255056 91089 255084 95202
rect 254766 91080 254822 91089
rect 254766 91015 254822 91024
rect 255042 91080 255098 91089
rect 255042 91015 255098 91024
rect 254780 81462 254808 91015
rect 254964 81462 254992 81493
rect 254768 81456 254820 81462
rect 254952 81456 255004 81462
rect 254768 81398 254820 81404
rect 254872 81404 254952 81410
rect 254872 81398 255004 81404
rect 254872 81382 254992 81398
rect 254872 80073 254900 81382
rect 254858 80064 254914 80073
rect 254858 79999 254914 80008
rect 255042 80064 255098 80073
rect 255042 79999 255098 80008
rect 255056 70417 255084 79999
rect 254858 70408 254914 70417
rect 254858 70343 254914 70352
rect 255042 70408 255098 70417
rect 255042 70343 255098 70352
rect 254872 60654 254900 70343
rect 254860 60648 254912 60654
rect 254860 60590 254912 60596
rect 255044 51128 255096 51134
rect 255044 51070 255096 51076
rect 255056 42838 255084 51070
rect 254768 42832 254820 42838
rect 254768 42774 254820 42780
rect 255044 42832 255096 42838
rect 255044 42774 255096 42780
rect 254780 34542 254808 42774
rect 254768 34536 254820 34542
rect 254768 34478 254820 34484
rect 254860 34536 254912 34542
rect 254860 34478 254912 34484
rect 254872 13138 254900 34478
rect 254780 13110 254900 13138
rect 254780 8276 254808 13110
rect 254780 8248 254900 8276
rect 254872 4078 254900 8248
rect 255044 4140 255096 4146
rect 255044 4082 255096 4088
rect 254860 4072 254912 4078
rect 254860 4014 254912 4020
rect 254676 604 254728 610
rect 254676 546 254728 552
rect 255056 480 255084 4082
rect 255240 3602 255268 340068
rect 255332 335186 255360 340068
rect 255424 336802 255452 340068
rect 255412 336796 255464 336802
rect 255412 336738 255464 336744
rect 255608 335322 255636 340068
rect 255700 335458 255728 340068
rect 255792 335782 255820 340068
rect 255884 340054 255990 340082
rect 255780 335776 255832 335782
rect 255780 335718 255832 335724
rect 255884 335578 255912 340054
rect 256068 335714 256096 340068
rect 256056 335708 256108 335714
rect 256056 335650 256108 335656
rect 255872 335572 255924 335578
rect 255872 335514 255924 335520
rect 255700 335430 256004 335458
rect 255608 335294 255728 335322
rect 255332 335158 255636 335186
rect 255504 335096 255556 335102
rect 255504 335038 255556 335044
rect 255228 3596 255280 3602
rect 255228 3538 255280 3544
rect 255516 3466 255544 335038
rect 255504 3460 255556 3466
rect 255504 3402 255556 3408
rect 255608 3398 255636 335158
rect 255596 3392 255648 3398
rect 255596 3334 255648 3340
rect 255700 2990 255728 335294
rect 255872 328500 255924 328506
rect 255872 328442 255924 328448
rect 255884 297378 255912 328442
rect 255792 297350 255912 297378
rect 255792 296698 255820 297350
rect 255792 296670 255912 296698
rect 255884 295322 255912 296670
rect 255872 295316 255924 295322
rect 255872 295258 255924 295264
rect 255780 289128 255832 289134
rect 255778 289096 255780 289105
rect 255832 289096 255834 289105
rect 255778 289031 255834 289040
rect 255778 276040 255834 276049
rect 255778 275975 255834 275984
rect 255792 274650 255820 275975
rect 255780 274644 255832 274650
rect 255780 274586 255832 274592
rect 255780 264988 255832 264994
rect 255780 264930 255832 264936
rect 255792 255270 255820 264930
rect 255780 255264 255832 255270
rect 255780 255206 255832 255212
rect 255872 237448 255924 237454
rect 255872 237390 255924 237396
rect 255884 237266 255912 237390
rect 255792 237238 255912 237266
rect 255792 227769 255820 237238
rect 255778 227760 255834 227769
rect 255778 227695 255834 227704
rect 255872 219564 255924 219570
rect 255872 219506 255924 219512
rect 255884 218006 255912 219506
rect 255872 218000 255924 218006
rect 255872 217942 255924 217948
rect 255872 208412 255924 208418
rect 255872 208354 255924 208360
rect 255884 198694 255912 208354
rect 255872 198688 255924 198694
rect 255872 198630 255924 198636
rect 255780 191344 255832 191350
rect 255780 191286 255832 191292
rect 255792 189038 255820 191286
rect 255780 189032 255832 189038
rect 255780 188974 255832 188980
rect 255872 184204 255924 184210
rect 255872 184146 255924 184152
rect 255884 157418 255912 184146
rect 255976 157434 256004 335430
rect 256054 227760 256110 227769
rect 256054 227695 256110 227704
rect 256068 219570 256096 227695
rect 256056 219564 256108 219570
rect 256056 219506 256108 219512
rect 255872 157412 255924 157418
rect 255976 157406 256096 157434
rect 255872 157354 255924 157360
rect 256068 157026 256096 157406
rect 255976 156998 256096 157026
rect 255872 154556 255924 154562
rect 255872 154498 255924 154504
rect 255884 135250 255912 154498
rect 255872 135244 255924 135250
rect 255872 135186 255924 135192
rect 255870 125624 255926 125633
rect 255870 125559 255926 125568
rect 255884 124166 255912 125559
rect 255872 124160 255924 124166
rect 255872 124102 255924 124108
rect 255870 106312 255926 106321
rect 255870 106247 255926 106256
rect 255884 98734 255912 106247
rect 255872 98728 255924 98734
rect 255872 98670 255924 98676
rect 255780 81456 255832 81462
rect 255780 81398 255832 81404
rect 255792 73098 255820 81398
rect 255780 73092 255832 73098
rect 255780 73034 255832 73040
rect 255872 63572 255924 63578
rect 255872 63514 255924 63520
rect 255884 62098 255912 63514
rect 255792 62070 255912 62098
rect 255792 62014 255820 62070
rect 255780 62008 255832 62014
rect 255780 61950 255832 61956
rect 255780 52488 255832 52494
rect 255780 52430 255832 52436
rect 255792 44266 255820 52430
rect 255780 44260 255832 44266
rect 255780 44202 255832 44208
rect 255872 42832 255924 42838
rect 255792 42792 255872 42820
rect 255792 34610 255820 42792
rect 255872 42774 255924 42780
rect 255780 34604 255832 34610
rect 255780 34546 255832 34552
rect 255872 34536 255924 34542
rect 255872 34478 255924 34484
rect 255884 8294 255912 34478
rect 255872 8288 255924 8294
rect 255872 8230 255924 8236
rect 255976 3874 256004 156998
rect 256056 135244 256108 135250
rect 256056 135186 256108 135192
rect 256068 125633 256096 135186
rect 256054 125624 256110 125633
rect 256054 125559 256110 125568
rect 256056 124160 256108 124166
rect 256056 124102 256108 124108
rect 256068 106321 256096 124102
rect 256054 106312 256110 106321
rect 256054 106247 256110 106256
rect 256056 98728 256108 98734
rect 256056 98670 256108 98676
rect 256068 81462 256096 98670
rect 256056 81456 256108 81462
rect 256056 81398 256108 81404
rect 256160 4146 256188 340068
rect 256148 4140 256200 4146
rect 256148 4082 256200 4088
rect 255964 3868 256016 3874
rect 255964 3810 256016 3816
rect 255688 2984 255740 2990
rect 255688 2926 255740 2932
rect 256344 626 256372 340068
rect 256436 328166 256464 340068
rect 256528 336870 256556 340068
rect 256712 337074 256740 340068
rect 256700 337068 256752 337074
rect 256700 337010 256752 337016
rect 256804 336938 256832 340068
rect 256792 336932 256844 336938
rect 256792 336874 256844 336880
rect 256516 336864 256568 336870
rect 256516 336806 256568 336812
rect 256896 334694 256924 340068
rect 256884 334688 256936 334694
rect 256884 334630 256936 334636
rect 256424 328160 256476 328166
rect 256424 328102 256476 328108
rect 256700 328160 256752 328166
rect 256700 328102 256752 328108
rect 256712 316130 256740 328102
rect 256608 316124 256660 316130
rect 256608 316066 256660 316072
rect 256700 316124 256752 316130
rect 256700 316066 256752 316072
rect 256620 314673 256648 316066
rect 256422 314664 256478 314673
rect 256422 314599 256478 314608
rect 256606 314664 256662 314673
rect 256606 314599 256662 314608
rect 256436 305017 256464 314599
rect 256422 305008 256478 305017
rect 256422 304943 256478 304952
rect 256606 305008 256662 305017
rect 256606 304943 256662 304952
rect 256620 295322 256648 304943
rect 256424 295316 256476 295322
rect 256424 295258 256476 295264
rect 256608 295316 256660 295322
rect 256608 295258 256660 295264
rect 256436 285705 256464 295258
rect 256422 285696 256478 285705
rect 256422 285631 256478 285640
rect 256606 285696 256662 285705
rect 256606 285631 256662 285640
rect 256620 238762 256648 285631
rect 256974 259448 257030 259457
rect 256974 259383 257030 259392
rect 256988 249830 257016 259383
rect 256976 249824 257028 249830
rect 256976 249766 257028 249772
rect 256528 238746 256648 238762
rect 256516 238740 256660 238746
rect 256568 238734 256608 238740
rect 256516 238682 256568 238688
rect 256608 238682 256660 238688
rect 256620 220930 256648 238682
rect 256608 220924 256660 220930
rect 256608 220866 256660 220872
rect 256424 220788 256476 220794
rect 256424 220730 256476 220736
rect 256436 193225 256464 220730
rect 256422 193216 256478 193225
rect 256422 193151 256478 193160
rect 256606 193216 256662 193225
rect 256606 193151 256662 193160
rect 256620 106298 256648 193151
rect 256528 106270 256648 106298
rect 256528 104854 256556 106270
rect 256516 104848 256568 104854
rect 256516 104790 256568 104796
rect 256700 95260 256752 95266
rect 256700 95202 256752 95208
rect 256712 89026 256740 95202
rect 256620 88998 256740 89026
rect 256620 82822 256648 88998
rect 256424 82816 256476 82822
rect 256424 82758 256476 82764
rect 256608 82816 256660 82822
rect 256608 82758 256660 82764
rect 256436 73166 256464 82758
rect 256424 73160 256476 73166
rect 256424 73102 256476 73108
rect 256608 63572 256660 63578
rect 256608 63514 256660 63520
rect 256620 44130 256648 63514
rect 256974 62112 257030 62121
rect 256974 62047 257030 62056
rect 256988 52494 257016 62047
rect 256976 52488 257028 52494
rect 256976 52430 257028 52436
rect 256608 44124 256660 44130
rect 256608 44066 256660 44072
rect 256608 18012 256660 18018
rect 256608 17954 256660 17960
rect 256620 17898 256648 17954
rect 256528 17870 256648 17898
rect 256528 9722 256556 17870
rect 256516 9716 256568 9722
rect 256516 9658 256568 9664
rect 256516 8356 256568 8362
rect 256516 8298 256568 8304
rect 256528 1902 256556 8298
rect 257080 3874 257108 340068
rect 257172 337618 257200 340068
rect 257160 337612 257212 337618
rect 257160 337554 257212 337560
rect 257264 337482 257292 340068
rect 257252 337476 257304 337482
rect 257252 337418 257304 337424
rect 257448 337142 257476 340068
rect 257540 337550 257568 340068
rect 257528 337544 257580 337550
rect 257528 337486 257580 337492
rect 257436 337136 257488 337142
rect 257436 337078 257488 337084
rect 257344 336864 257396 336870
rect 257344 336806 257396 336812
rect 257160 334688 257212 334694
rect 257160 334630 257212 334636
rect 257172 328438 257200 334630
rect 257160 328432 257212 328438
rect 257160 328374 257212 328380
rect 257252 328432 257304 328438
rect 257252 328374 257304 328380
rect 257264 287094 257292 328374
rect 257160 287088 257212 287094
rect 257160 287030 257212 287036
rect 257252 287088 257304 287094
rect 257252 287030 257304 287036
rect 257172 266370 257200 287030
rect 257172 266342 257292 266370
rect 257264 260914 257292 266342
rect 257160 260908 257212 260914
rect 257160 260850 257212 260856
rect 257252 260908 257304 260914
rect 257252 260850 257304 260856
rect 257172 259457 257200 260850
rect 257158 259448 257214 259457
rect 257158 259383 257214 259392
rect 257252 249824 257304 249830
rect 257252 249766 257304 249772
rect 257264 229129 257292 249766
rect 257250 229120 257306 229129
rect 257250 229055 257306 229064
rect 257250 228984 257306 228993
rect 257250 228919 257306 228928
rect 257264 169114 257292 228919
rect 257252 169108 257304 169114
rect 257252 169050 257304 169056
rect 257250 164248 257306 164257
rect 257250 164183 257306 164192
rect 257264 154698 257292 164183
rect 257252 154692 257304 154698
rect 257252 154634 257304 154640
rect 257160 154556 257212 154562
rect 257160 154498 257212 154504
rect 257172 130422 257200 154498
rect 257160 130416 257212 130422
rect 257160 130358 257212 130364
rect 257252 130348 257304 130354
rect 257252 130290 257304 130296
rect 257264 124166 257292 130290
rect 257252 124160 257304 124166
rect 257252 124102 257304 124108
rect 257252 114572 257304 114578
rect 257252 114514 257304 114520
rect 257264 95266 257292 114514
rect 257252 95260 257304 95266
rect 257252 95202 257304 95208
rect 257252 93900 257304 93906
rect 257252 93842 257304 93848
rect 257264 84266 257292 93842
rect 257172 84238 257292 84266
rect 257172 77874 257200 84238
rect 257172 77846 257292 77874
rect 257264 68406 257292 77846
rect 257252 68400 257304 68406
rect 257252 68342 257304 68348
rect 257160 63572 257212 63578
rect 257160 63514 257212 63520
rect 257172 62121 257200 63514
rect 257158 62112 257214 62121
rect 257158 62047 257214 62056
rect 257252 52488 257304 52494
rect 257252 52430 257304 52436
rect 257264 48346 257292 52430
rect 257160 48340 257212 48346
rect 257160 48282 257212 48288
rect 257252 48340 257304 48346
rect 257252 48282 257304 48288
rect 257172 39370 257200 48282
rect 257160 39364 257212 39370
rect 257160 39306 257212 39312
rect 257252 34536 257304 34542
rect 257252 34478 257304 34484
rect 257264 27606 257292 34478
rect 257252 27600 257304 27606
rect 257252 27542 257304 27548
rect 257252 18012 257304 18018
rect 257252 17954 257304 17960
rect 257264 9722 257292 17954
rect 257160 9716 257212 9722
rect 257160 9658 257212 9664
rect 257252 9716 257304 9722
rect 257252 9658 257304 9664
rect 257172 3942 257200 9658
rect 257356 4078 257384 336806
rect 257436 336796 257488 336802
rect 257436 336738 257488 336744
rect 257448 318102 257476 336738
rect 257436 318096 257488 318102
rect 257436 318038 257488 318044
rect 257436 169108 257488 169114
rect 257436 169050 257488 169056
rect 257448 164257 257476 169050
rect 257434 164248 257490 164257
rect 257434 164183 257490 164192
rect 257632 4758 257660 340068
rect 257712 336932 257764 336938
rect 257712 336874 257764 336880
rect 257620 4752 257672 4758
rect 257620 4694 257672 4700
rect 257344 4072 257396 4078
rect 257344 4014 257396 4020
rect 257724 4010 257752 336874
rect 257816 5506 257844 340068
rect 257908 336802 257936 340068
rect 257896 336796 257948 336802
rect 257896 336738 257948 336744
rect 257804 5500 257856 5506
rect 257804 5442 257856 5448
rect 258000 5370 258028 340068
rect 258184 336802 258212 340068
rect 258276 337686 258304 340068
rect 258264 337680 258316 337686
rect 258264 337622 258316 337628
rect 258264 336932 258316 336938
rect 258264 336874 258316 336880
rect 258172 336796 258224 336802
rect 258172 336738 258224 336744
rect 258276 335628 258304 336874
rect 258368 335782 258396 340068
rect 258460 340054 258566 340082
rect 258356 335776 258408 335782
rect 258356 335718 258408 335724
rect 258276 335600 258396 335628
rect 258264 331220 258316 331226
rect 258264 331162 258316 331168
rect 258276 315518 258304 331162
rect 258264 315512 258316 315518
rect 258264 315454 258316 315460
rect 257988 5364 258040 5370
rect 257988 5306 258040 5312
rect 258368 4894 258396 335600
rect 258460 5234 258488 340054
rect 258644 337346 258672 340068
rect 258632 337340 258684 337346
rect 258632 337282 258684 337288
rect 258540 337068 258592 337074
rect 258540 337010 258592 337016
rect 258448 5228 258500 5234
rect 258448 5170 258500 5176
rect 258356 4888 258408 4894
rect 258356 4830 258408 4836
rect 258552 4146 258580 337010
rect 258736 336802 258764 340068
rect 258920 336870 258948 340068
rect 258908 336864 258960 336870
rect 258908 336806 258960 336812
rect 258632 336796 258684 336802
rect 258632 336738 258684 336744
rect 258724 336796 258776 336802
rect 258724 336738 258776 336744
rect 258644 5438 258672 336738
rect 258908 335776 258960 335782
rect 258908 335718 258960 335724
rect 258632 5432 258684 5438
rect 258632 5374 258684 5380
rect 258920 5302 258948 335718
rect 259012 327758 259040 340068
rect 259104 336938 259132 340068
rect 259196 340054 259302 340082
rect 259092 336932 259144 336938
rect 259092 336874 259144 336880
rect 259092 336796 259144 336802
rect 259092 336738 259144 336744
rect 259000 327752 259052 327758
rect 259000 327694 259052 327700
rect 258908 5296 258960 5302
rect 258908 5238 258960 5244
rect 259104 5166 259132 336738
rect 259092 5160 259144 5166
rect 259092 5102 259144 5108
rect 259196 5030 259224 340054
rect 259276 336864 259328 336870
rect 259276 336806 259328 336812
rect 259288 5098 259316 336806
rect 259380 331226 259408 340068
rect 259472 336802 259500 340068
rect 259656 337278 259684 340068
rect 259644 337272 259696 337278
rect 259644 337214 259696 337220
rect 259748 337142 259776 340068
rect 259736 337136 259788 337142
rect 259736 337078 259788 337084
rect 259460 336796 259512 336802
rect 259460 336738 259512 336744
rect 259840 333402 259868 340068
rect 259932 340054 260038 340082
rect 259828 333396 259880 333402
rect 259828 333338 259880 333344
rect 259932 331922 259960 340054
rect 260116 337210 260144 340068
rect 260104 337204 260156 337210
rect 260104 337146 260156 337152
rect 260208 337074 260236 340068
rect 260196 337068 260248 337074
rect 260196 337010 260248 337016
rect 260300 335628 260328 340068
rect 260380 336796 260432 336802
rect 260380 336738 260432 336744
rect 259840 331894 259960 331922
rect 260024 335600 260328 335628
rect 259368 331220 259420 331226
rect 259368 331162 259420 331168
rect 259840 301594 259868 331894
rect 259840 301566 259960 301594
rect 259932 270638 259960 301566
rect 259920 270632 259972 270638
rect 259920 270574 259972 270580
rect 259828 270496 259880 270502
rect 259828 270438 259880 270444
rect 259840 264330 259868 270438
rect 259840 264302 259960 264330
rect 259932 255270 259960 264302
rect 259920 255264 259972 255270
rect 259920 255206 259972 255212
rect 259920 245676 259972 245682
rect 259920 245618 259972 245624
rect 259932 217410 259960 245618
rect 259840 217382 259960 217410
rect 259840 205698 259868 217382
rect 259828 205692 259880 205698
rect 259828 205634 259880 205640
rect 259920 205624 259972 205630
rect 259920 205566 259972 205572
rect 259932 189145 259960 205566
rect 259918 189136 259974 189145
rect 259918 189071 259974 189080
rect 259734 189000 259790 189009
rect 259790 188958 259868 188986
rect 259734 188935 259790 188944
rect 259840 182050 259868 188958
rect 259840 182022 259960 182050
rect 259932 169794 259960 182022
rect 259920 169788 259972 169794
rect 259920 169730 259972 169736
rect 259736 169720 259788 169726
rect 259736 169662 259788 169668
rect 259748 160138 259776 169662
rect 259736 160132 259788 160138
rect 259736 160074 259788 160080
rect 259920 160132 259972 160138
rect 259920 160074 259972 160080
rect 259932 157434 259960 160074
rect 259840 157406 259960 157434
rect 259840 147694 259868 157406
rect 259828 147688 259880 147694
rect 259828 147630 259880 147636
rect 259920 147620 259972 147626
rect 259920 147562 259972 147568
rect 259932 138122 259960 147562
rect 259840 138094 259960 138122
rect 259840 128382 259868 138094
rect 259828 128376 259880 128382
rect 259828 128318 259880 128324
rect 259920 128308 259972 128314
rect 259920 128250 259972 128256
rect 259932 120714 259960 128250
rect 259840 120686 259960 120714
rect 259840 115938 259868 120686
rect 259828 115932 259880 115938
rect 259828 115874 259880 115880
rect 259920 115932 259972 115938
rect 259920 115874 259972 115880
rect 259932 95266 259960 115874
rect 259920 95260 259972 95266
rect 259920 95202 259972 95208
rect 259920 92540 259972 92546
rect 259920 92482 259972 92488
rect 259932 81462 259960 92482
rect 259828 81456 259880 81462
rect 259828 81398 259880 81404
rect 259920 81456 259972 81462
rect 259920 81398 259972 81404
rect 259840 73166 259868 81398
rect 259828 73160 259880 73166
rect 259828 73102 259880 73108
rect 259734 71768 259790 71777
rect 259734 71703 259790 71712
rect 259748 62150 259776 71703
rect 260024 63578 260052 335600
rect 260392 335458 260420 336738
rect 260300 335430 260420 335458
rect 260196 333396 260248 333402
rect 260196 333338 260248 333344
rect 260104 73160 260156 73166
rect 260104 73102 260156 73108
rect 260116 71777 260144 73102
rect 260102 71768 260158 71777
rect 260102 71703 260158 71712
rect 260012 63572 260064 63578
rect 260012 63514 260064 63520
rect 260012 63436 260064 63442
rect 260012 63378 260064 63384
rect 259736 62144 259788 62150
rect 259736 62086 259788 62092
rect 259828 62144 259880 62150
rect 259828 62086 259880 62092
rect 259840 51134 259868 62086
rect 259828 51128 259880 51134
rect 259828 51070 259880 51076
rect 259920 51060 259972 51066
rect 259920 51002 259972 51008
rect 259932 43466 259960 51002
rect 259840 43438 259960 43466
rect 259840 27606 259868 43438
rect 259828 27600 259880 27606
rect 259828 27542 259880 27548
rect 259920 27600 259972 27606
rect 259920 27542 259972 27548
rect 259932 9314 259960 27542
rect 259920 9308 259972 9314
rect 259920 9250 259972 9256
rect 260024 9246 260052 63378
rect 260012 9240 260064 9246
rect 260012 9182 260064 9188
rect 259276 5092 259328 5098
rect 259276 5034 259328 5040
rect 259184 5024 259236 5030
rect 259184 4966 259236 4972
rect 260208 4826 260236 333338
rect 260300 4962 260328 335430
rect 260484 332382 260512 340068
rect 260576 337414 260604 340068
rect 260564 337408 260616 337414
rect 260564 337350 260616 337356
rect 260472 332376 260524 332382
rect 260472 332318 260524 332324
rect 260668 324358 260696 340068
rect 260748 337204 260800 337210
rect 260748 337146 260800 337152
rect 260760 335102 260788 337146
rect 260748 335096 260800 335102
rect 260748 335038 260800 335044
rect 260852 333554 260880 340068
rect 260944 336530 260972 340068
rect 261036 336802 261064 340068
rect 261220 336938 261248 340068
rect 261312 338094 261340 340068
rect 261300 338088 261352 338094
rect 261300 338030 261352 338036
rect 261208 336932 261260 336938
rect 261208 336874 261260 336880
rect 261024 336796 261076 336802
rect 261024 336738 261076 336744
rect 261024 336660 261076 336666
rect 261024 336602 261076 336608
rect 260932 336524 260984 336530
rect 260932 336466 260984 336472
rect 261036 333606 261064 336602
rect 260760 333526 260880 333554
rect 261024 333600 261076 333606
rect 261024 333542 261076 333548
rect 260760 333282 260788 333526
rect 261300 333328 261352 333334
rect 260760 333254 260972 333282
rect 261300 333270 261352 333276
rect 260840 331220 260892 331226
rect 260840 331162 260892 331168
rect 260380 324352 260432 324358
rect 260378 324320 260380 324329
rect 260656 324352 260708 324358
rect 260432 324320 260434 324329
rect 260378 324255 260434 324264
rect 260654 324320 260656 324329
rect 260708 324320 260710 324329
rect 260654 324255 260710 324264
rect 260668 321910 260696 324255
rect 260656 321904 260708 321910
rect 260656 321846 260708 321852
rect 260656 314696 260708 314702
rect 260656 314638 260708 314644
rect 260668 266529 260696 314638
rect 260852 311370 260880 331162
rect 260944 328166 260972 333254
rect 261208 332988 261260 332994
rect 261208 332930 261260 332936
rect 260932 328160 260984 328166
rect 260932 328102 260984 328108
rect 260840 311364 260892 311370
rect 260840 311306 260892 311312
rect 260654 266520 260710 266529
rect 260654 266455 260710 266464
rect 260654 266384 260710 266393
rect 260654 266319 260710 266328
rect 260668 247042 260696 266319
rect 260656 247036 260708 247042
rect 260656 246978 260708 246984
rect 260564 237448 260616 237454
rect 260564 237390 260616 237396
rect 260576 227769 260604 237390
rect 260562 227760 260618 227769
rect 260562 227695 260618 227704
rect 260746 227760 260802 227769
rect 260746 227695 260802 227704
rect 260760 219502 260788 227695
rect 260748 219496 260800 219502
rect 260748 219438 260800 219444
rect 260656 219428 260708 219434
rect 260656 219370 260708 219376
rect 260668 218006 260696 219370
rect 260656 218000 260708 218006
rect 260656 217942 260708 217948
rect 260932 218000 260984 218006
rect 260932 217942 260984 217948
rect 260944 208457 260972 217942
rect 260930 208448 260986 208457
rect 260930 208383 260986 208392
rect 260746 208312 260802 208321
rect 260746 208247 260802 208256
rect 260760 198694 260788 208247
rect 260656 198688 260708 198694
rect 260656 198630 260708 198636
rect 260748 198688 260800 198694
rect 260748 198630 260800 198636
rect 260668 197334 260696 198630
rect 260656 197328 260708 197334
rect 260656 197270 260708 197276
rect 260656 187740 260708 187746
rect 260656 187682 260708 187688
rect 260668 179450 260696 187682
rect 260656 179444 260708 179450
rect 260656 179386 260708 179392
rect 260656 178084 260708 178090
rect 260656 178026 260708 178032
rect 260668 177993 260696 178026
rect 260654 177984 260710 177993
rect 260654 177919 260710 177928
rect 260838 177984 260894 177993
rect 260838 177919 260894 177928
rect 260852 168473 260880 177919
rect 260654 168464 260710 168473
rect 260654 168399 260710 168408
rect 260838 168464 260894 168473
rect 260838 168399 260894 168408
rect 260668 162874 260696 168399
rect 260576 162846 260696 162874
rect 260576 158710 260604 162846
rect 260564 158704 260616 158710
rect 260564 158646 260616 158652
rect 260656 149116 260708 149122
rect 260656 149058 260708 149064
rect 260668 140842 260696 149058
rect 260576 140814 260696 140842
rect 260576 140758 260604 140814
rect 260564 140752 260616 140758
rect 260564 140694 260616 140700
rect 260564 129804 260616 129810
rect 260564 129746 260616 129752
rect 260576 111790 260604 129746
rect 260472 111784 260524 111790
rect 260472 111726 260524 111732
rect 260564 111784 260616 111790
rect 260564 111726 260616 111732
rect 260484 110430 260512 111726
rect 260472 110424 260524 110430
rect 260472 110366 260524 110372
rect 260564 102128 260616 102134
rect 260564 102070 260616 102076
rect 260576 100745 260604 102070
rect 260562 100736 260618 100745
rect 260562 100671 260618 100680
rect 260654 100600 260710 100609
rect 260654 100535 260710 100544
rect 260668 78010 260696 100535
rect 260576 77982 260696 78010
rect 260576 45558 260604 77982
rect 260564 45552 260616 45558
rect 260564 45494 260616 45500
rect 260564 45416 260616 45422
rect 260564 45358 260616 45364
rect 260576 34678 260604 45358
rect 260564 34672 260616 34678
rect 260564 34614 260616 34620
rect 260656 34536 260708 34542
rect 260656 34478 260708 34484
rect 260668 29034 260696 34478
rect 260656 29028 260708 29034
rect 260656 28970 260708 28976
rect 260564 28960 260616 28966
rect 260564 28902 260616 28908
rect 260576 26194 260604 28902
rect 260576 26166 260696 26194
rect 260668 16590 260696 26166
rect 260656 16584 260708 16590
rect 260656 16526 260708 16532
rect 261220 9110 261248 332930
rect 261208 9104 261260 9110
rect 261208 9046 261260 9052
rect 261312 9042 261340 333270
rect 261404 332994 261432 340068
rect 261484 336796 261536 336802
rect 261484 336738 261536 336744
rect 261392 332988 261444 332994
rect 261392 332930 261444 332936
rect 261496 326482 261524 336738
rect 261588 333690 261616 340068
rect 261680 333810 261708 340068
rect 261668 333804 261720 333810
rect 261668 333746 261720 333752
rect 261588 333662 261708 333690
rect 261576 333600 261628 333606
rect 261576 333542 261628 333548
rect 261404 326454 261524 326482
rect 261300 9036 261352 9042
rect 261300 8978 261352 8984
rect 261404 8974 261432 326454
rect 261588 326346 261616 333542
rect 261496 326318 261616 326346
rect 261680 326330 261708 333662
rect 261772 333334 261800 340068
rect 261852 336932 261904 336938
rect 261852 336874 261904 336880
rect 261760 333328 261812 333334
rect 261760 333270 261812 333276
rect 261760 328500 261812 328506
rect 261760 328442 261812 328448
rect 261668 326324 261720 326330
rect 261392 8968 261444 8974
rect 261392 8910 261444 8916
rect 261496 8294 261524 326318
rect 261668 326266 261720 326272
rect 261668 326120 261720 326126
rect 261668 326062 261720 326068
rect 261680 319734 261708 326062
rect 261668 319728 261720 319734
rect 261668 319670 261720 319676
rect 261772 313954 261800 328442
rect 261864 325310 261892 336874
rect 261956 331294 261984 340068
rect 262048 335034 262076 340068
rect 262036 335028 262088 335034
rect 262036 334970 262088 334976
rect 261944 331288 261996 331294
rect 261944 331230 261996 331236
rect 262140 330886 262168 340068
rect 262220 337272 262272 337278
rect 262220 337214 262272 337220
rect 262232 334626 262260 337214
rect 262220 334620 262272 334626
rect 262220 334562 262272 334568
rect 262128 330880 262180 330886
rect 262128 330822 262180 330828
rect 261852 325304 261904 325310
rect 261852 325246 261904 325252
rect 262324 323950 262352 340068
rect 262416 337090 262444 340068
rect 262508 337210 262536 340068
rect 262496 337204 262548 337210
rect 262496 337146 262548 337152
rect 262416 337062 262536 337090
rect 262508 336462 262536 337062
rect 262496 336456 262548 336462
rect 262496 336398 262548 336404
rect 262496 336320 262548 336326
rect 262496 336262 262548 336268
rect 262508 333470 262536 336262
rect 262588 335776 262640 335782
rect 262588 335718 262640 335724
rect 262496 333464 262548 333470
rect 262496 333406 262548 333412
rect 262600 331922 262628 335718
rect 262508 331894 262628 331922
rect 262402 324320 262458 324329
rect 262402 324255 262458 324264
rect 262312 323944 262364 323950
rect 262312 323886 262364 323892
rect 262416 314702 262444 324255
rect 262404 314696 262456 314702
rect 262404 314638 262456 314644
rect 261760 313948 261812 313954
rect 261760 313890 261812 313896
rect 262508 293350 262536 331894
rect 262692 331362 262720 340068
rect 262784 338026 262812 340068
rect 262772 338020 262824 338026
rect 262772 337962 262824 337968
rect 262876 336870 262904 340068
rect 262956 337204 263008 337210
rect 262956 337146 263008 337152
rect 262864 336864 262916 336870
rect 262864 336806 262916 336812
rect 262772 336796 262824 336802
rect 262772 336738 262824 336744
rect 262680 331356 262732 331362
rect 262680 331298 262732 331304
rect 262680 324352 262732 324358
rect 262678 324320 262680 324329
rect 262732 324320 262734 324329
rect 262678 324255 262734 324264
rect 262588 314696 262640 314702
rect 262588 314638 262640 314644
rect 262600 306542 262628 314638
rect 262588 306536 262640 306542
rect 262588 306478 262640 306484
rect 262680 306400 262732 306406
rect 262680 306342 262732 306348
rect 262496 293344 262548 293350
rect 262496 293286 262548 293292
rect 262692 266506 262720 306342
rect 262600 266478 262720 266506
rect 262600 266370 262628 266478
rect 262600 266342 262720 266370
rect 262692 247042 262720 266342
rect 262496 247036 262548 247042
rect 262496 246978 262548 246984
rect 262680 247036 262732 247042
rect 262680 246978 262732 246984
rect 262508 237425 262536 246978
rect 262494 237416 262550 237425
rect 262494 237351 262550 237360
rect 262678 237416 262734 237425
rect 262678 237351 262734 237360
rect 262692 234734 262720 237351
rect 262680 234728 262732 234734
rect 262680 234670 262732 234676
rect 262496 229084 262548 229090
rect 262496 229026 262548 229032
rect 262508 219450 262536 229026
rect 262508 219422 262720 219450
rect 262692 218006 262720 219422
rect 262680 218000 262732 218006
rect 262680 217942 262732 217948
rect 262680 198756 262732 198762
rect 262680 198698 262732 198704
rect 262692 189038 262720 198698
rect 262680 189032 262732 189038
rect 262680 188974 262732 188980
rect 262680 179444 262732 179450
rect 262680 179386 262732 179392
rect 262692 169726 262720 179386
rect 262680 169720 262732 169726
rect 262680 169662 262732 169668
rect 262680 160132 262732 160138
rect 262680 160074 262732 160080
rect 262692 140758 262720 160074
rect 262680 140752 262732 140758
rect 262680 140694 262732 140700
rect 262680 131164 262732 131170
rect 262680 131106 262732 131112
rect 262692 111790 262720 131106
rect 262680 111784 262732 111790
rect 262680 111726 262732 111732
rect 262680 102264 262732 102270
rect 262680 102206 262732 102212
rect 262692 102134 262720 102206
rect 262680 102128 262732 102134
rect 262680 102070 262732 102076
rect 262588 91112 262640 91118
rect 262588 91054 262640 91060
rect 262600 81462 262628 91054
rect 262588 81456 262640 81462
rect 262588 81398 262640 81404
rect 262496 81388 262548 81394
rect 262496 81330 262548 81336
rect 262508 75290 262536 81330
rect 262416 75262 262536 75290
rect 262416 66858 262444 75262
rect 262416 66830 262628 66858
rect 262600 45558 262628 66830
rect 262588 45552 262640 45558
rect 262588 45494 262640 45500
rect 262680 45552 262732 45558
rect 262680 45494 262732 45500
rect 262692 16590 262720 45494
rect 262680 16584 262732 16590
rect 262680 16526 262732 16532
rect 261484 8288 261536 8294
rect 261484 8230 261536 8236
rect 262588 6996 262640 7002
rect 262588 6938 262640 6944
rect 262600 6848 262628 6938
rect 262600 6820 262720 6848
rect 262692 5642 262720 6820
rect 262680 5636 262732 5642
rect 262680 5578 262732 5584
rect 262784 5574 262812 336738
rect 262864 336728 262916 336734
rect 262864 336670 262916 336676
rect 262876 333554 262904 336670
rect 262968 333674 262996 337146
rect 262956 333668 263008 333674
rect 262956 333610 263008 333616
rect 262876 333526 262996 333554
rect 262864 333464 262916 333470
rect 262864 333406 262916 333412
rect 262772 5568 262824 5574
rect 262772 5510 262824 5516
rect 260288 4956 260340 4962
rect 260288 4898 260340 4904
rect 260196 4820 260248 4826
rect 260196 4762 260248 4768
rect 262876 4146 262904 333406
rect 262968 6934 262996 333526
rect 263060 322454 263088 340068
rect 263152 336802 263180 340068
rect 263258 340054 263364 340082
rect 263232 336864 263284 336870
rect 263232 336806 263284 336812
rect 263140 336796 263192 336802
rect 263140 336738 263192 336744
rect 263244 331378 263272 336806
rect 263336 335628 263364 340054
rect 263428 335782 263456 340068
rect 263520 338314 263548 340068
rect 263612 338434 263640 340068
rect 263600 338428 263652 338434
rect 263600 338370 263652 338376
rect 263520 338286 263640 338314
rect 263416 335776 263468 335782
rect 263416 335718 263468 335724
rect 263336 335600 263548 335628
rect 263244 331350 263364 331378
rect 263232 331288 263284 331294
rect 263232 331230 263284 331236
rect 263048 322448 263100 322454
rect 263048 322390 263100 322396
rect 263244 310010 263272 331230
rect 263336 326738 263364 331350
rect 263520 329458 263548 335600
rect 263508 329452 263560 329458
rect 263508 329394 263560 329400
rect 263324 326732 263376 326738
rect 263324 326674 263376 326680
rect 263612 324358 263640 338286
rect 263692 337136 263744 337142
rect 263690 337104 263692 337113
rect 263744 337104 263746 337113
rect 263690 337039 263746 337048
rect 263796 337006 263824 340068
rect 263784 337000 263836 337006
rect 263784 336942 263836 336948
rect 263888 327010 263916 340068
rect 263980 337958 264008 340068
rect 263968 337952 264020 337958
rect 263968 337894 264020 337900
rect 264164 337822 264192 340068
rect 264152 337816 264204 337822
rect 264152 337758 264204 337764
rect 263968 337136 264020 337142
rect 263968 337078 264020 337084
rect 263876 327004 263928 327010
rect 263876 326946 263928 326952
rect 263600 324352 263652 324358
rect 263600 324294 263652 324300
rect 263232 310004 263284 310010
rect 263232 309946 263284 309952
rect 263980 308582 264008 337078
rect 264152 336864 264204 336870
rect 264152 336806 264204 336812
rect 264060 326392 264112 326398
rect 264060 326334 264112 326340
rect 263968 308576 264020 308582
rect 263968 308518 264020 308524
rect 262956 6928 263008 6934
rect 262956 6870 263008 6876
rect 264072 5778 264100 326334
rect 264164 5846 264192 336806
rect 264256 326398 264284 340068
rect 264348 337346 264376 340068
rect 264336 337340 264388 337346
rect 264336 337282 264388 337288
rect 264428 337000 264480 337006
rect 264428 336942 264480 336948
rect 264440 328098 264468 336942
rect 264428 328092 264480 328098
rect 264428 328034 264480 328040
rect 264336 327004 264388 327010
rect 264336 326946 264388 326952
rect 264244 326392 264296 326398
rect 264244 326334 264296 326340
rect 264348 306406 264376 326946
rect 264532 318306 264560 340068
rect 264624 336870 264652 340068
rect 264612 336864 264664 336870
rect 264612 336806 264664 336812
rect 264716 333606 264744 340068
rect 264796 337340 264848 337346
rect 264796 337282 264848 337288
rect 264704 333600 264756 333606
rect 264704 333542 264756 333548
rect 264808 332450 264836 337282
rect 264900 337142 264928 340068
rect 264888 337136 264940 337142
rect 264888 337078 264940 337084
rect 264796 332444 264848 332450
rect 264796 332386 264848 332392
rect 264520 318300 264572 318306
rect 264520 318242 264572 318248
rect 264244 306400 264296 306406
rect 264242 306368 264244 306377
rect 264336 306400 264388 306406
rect 264296 306368 264298 306377
rect 264336 306342 264388 306348
rect 264426 306368 264482 306377
rect 264242 306303 264298 306312
rect 264426 306303 264482 306312
rect 264440 296750 264468 306303
rect 264244 296744 264296 296750
rect 264244 296686 264296 296692
rect 264428 296744 264480 296750
rect 264428 296686 264480 296692
rect 264256 237386 264284 296686
rect 264244 237380 264296 237386
rect 264244 237322 264296 237328
rect 264244 219496 264296 219502
rect 264244 219438 264296 219444
rect 264256 218006 264284 219438
rect 264244 218000 264296 218006
rect 264244 217942 264296 217948
rect 264428 208412 264480 208418
rect 264428 208354 264480 208360
rect 264440 198762 264468 208354
rect 264244 198756 264296 198762
rect 264244 198698 264296 198704
rect 264428 198756 264480 198762
rect 264428 198698 264480 198704
rect 264256 189038 264284 198698
rect 264244 189032 264296 189038
rect 264244 188974 264296 188980
rect 264244 179444 264296 179450
rect 264244 179386 264296 179392
rect 264256 169726 264284 179386
rect 264244 169720 264296 169726
rect 264244 169662 264296 169668
rect 264244 160132 264296 160138
rect 264244 160074 264296 160080
rect 264256 140758 264284 160074
rect 264244 140752 264296 140758
rect 264244 140694 264296 140700
rect 264244 131164 264296 131170
rect 264244 131106 264296 131112
rect 264256 102134 264284 131106
rect 264244 102128 264296 102134
rect 264244 102070 264296 102076
rect 264244 92540 264296 92546
rect 264244 92482 264296 92488
rect 264256 92426 264284 92482
rect 264256 92398 264376 92426
rect 264348 82906 264376 92398
rect 264256 82878 264376 82906
rect 264256 82822 264284 82878
rect 264244 82816 264296 82822
rect 264244 82758 264296 82764
rect 264336 75812 264388 75818
rect 264336 75754 264388 75760
rect 264348 66298 264376 75754
rect 264244 66292 264296 66298
rect 264244 66234 264296 66240
rect 264336 66292 264388 66298
rect 264336 66234 264388 66240
rect 264256 45558 264284 66234
rect 264244 45552 264296 45558
rect 264244 45494 264296 45500
rect 264244 35964 264296 35970
rect 264244 35906 264296 35912
rect 264256 26246 264284 35906
rect 264244 26240 264296 26246
rect 264244 26182 264296 26188
rect 264244 16652 264296 16658
rect 264244 16594 264296 16600
rect 264256 6866 264284 16594
rect 264244 6860 264296 6866
rect 264244 6802 264296 6808
rect 264992 5914 265020 340068
rect 265084 10062 265112 340068
rect 265268 337754 265296 340068
rect 265256 337748 265308 337754
rect 265256 337690 265308 337696
rect 265360 336870 265388 340068
rect 265348 336864 265400 336870
rect 265348 336806 265400 336812
rect 265452 335374 265480 340068
rect 265636 337482 265664 340068
rect 265624 337476 265676 337482
rect 265624 337418 265676 337424
rect 265624 336796 265676 336802
rect 265624 336738 265676 336744
rect 265164 335368 265216 335374
rect 265164 335310 265216 335316
rect 265440 335368 265492 335374
rect 265440 335310 265492 335316
rect 265532 335368 265584 335374
rect 265532 335310 265584 335316
rect 265176 327078 265204 335310
rect 265440 327412 265492 327418
rect 265440 327354 265492 327360
rect 265164 327072 265216 327078
rect 265164 327014 265216 327020
rect 265256 327072 265308 327078
rect 265256 327014 265308 327020
rect 265268 302954 265296 327014
rect 265268 302926 265388 302954
rect 265072 10056 265124 10062
rect 265072 9998 265124 10004
rect 264980 5908 265032 5914
rect 264980 5850 265032 5856
rect 264152 5840 264204 5846
rect 264152 5782 264204 5788
rect 264060 5772 264112 5778
rect 264060 5714 264112 5720
rect 265360 4214 265388 302926
rect 265452 6118 265480 327354
rect 265544 327078 265572 335310
rect 265636 329390 265664 336738
rect 265728 335510 265756 340068
rect 265716 335504 265768 335510
rect 265716 335446 265768 335452
rect 265624 329384 265676 329390
rect 265624 329326 265676 329332
rect 265532 327072 265584 327078
rect 265532 327014 265584 327020
rect 265624 327072 265676 327078
rect 265624 327014 265676 327020
rect 265636 302954 265664 327014
rect 265636 302926 265756 302954
rect 265728 10130 265756 302926
rect 265820 10198 265848 340068
rect 265900 338428 265952 338434
rect 265900 338370 265952 338376
rect 265912 334966 265940 338370
rect 266004 336326 266032 340068
rect 265992 336320 266044 336326
rect 265992 336262 266044 336268
rect 266096 335714 266124 340068
rect 266084 335708 266136 335714
rect 266084 335650 266136 335656
rect 266188 335594 266216 340068
rect 266372 337550 266400 340068
rect 266360 337544 266412 337550
rect 266360 337486 266412 337492
rect 266360 337000 266412 337006
rect 266360 336942 266412 336948
rect 266268 336864 266320 336870
rect 266268 336806 266320 336812
rect 266280 336734 266308 336806
rect 266268 336728 266320 336734
rect 266268 336670 266320 336676
rect 266004 335566 266216 335594
rect 265900 334960 265952 334966
rect 265900 334902 265952 334908
rect 266004 10266 266032 335566
rect 266084 335504 266136 335510
rect 266084 335446 266136 335452
rect 266372 335458 266400 336942
rect 266464 335594 266492 340068
rect 266556 335714 266584 340068
rect 266740 337550 266768 340068
rect 266636 337544 266688 337550
rect 266636 337486 266688 337492
rect 266728 337544 266780 337550
rect 266728 337486 266780 337492
rect 266648 336802 266676 337486
rect 266728 337272 266780 337278
rect 266728 337214 266780 337220
rect 266636 336796 266688 336802
rect 266636 336738 266688 336744
rect 266544 335708 266596 335714
rect 266544 335650 266596 335656
rect 266464 335566 266676 335594
rect 265992 10260 266044 10266
rect 265992 10202 266044 10208
rect 265808 10192 265860 10198
rect 265808 10134 265860 10140
rect 265716 10124 265768 10130
rect 265716 10066 265768 10072
rect 265440 6112 265492 6118
rect 265440 6054 265492 6060
rect 266096 6050 266124 335446
rect 266372 335430 266584 335458
rect 266360 335368 266412 335374
rect 266360 335310 266412 335316
rect 266268 327140 266320 327146
rect 266268 327082 266320 327088
rect 266280 299538 266308 327082
rect 266372 326670 266400 335310
rect 266452 332036 266504 332042
rect 266452 331978 266504 331984
rect 266360 326664 266412 326670
rect 266360 326606 266412 326612
rect 266176 299532 266228 299538
rect 266176 299474 266228 299480
rect 266268 299532 266320 299538
rect 266268 299474 266320 299480
rect 266084 6044 266136 6050
rect 266084 5986 266136 5992
rect 266188 5982 266216 299474
rect 266266 228032 266322 228041
rect 266266 227967 266322 227976
rect 266280 227769 266308 227967
rect 266266 227760 266322 227769
rect 266266 227695 266322 227704
rect 266464 6662 266492 331978
rect 266556 6730 266584 335430
rect 266648 326398 266676 335566
rect 266740 332042 266768 337214
rect 266728 332036 266780 332042
rect 266728 331978 266780 331984
rect 266832 331922 266860 340068
rect 266924 336802 266952 340068
rect 267016 340054 267122 340082
rect 266912 336796 266964 336802
rect 266912 336738 266964 336744
rect 267016 335374 267044 340054
rect 267200 337006 267228 340068
rect 267188 337000 267240 337006
rect 267188 336942 267240 336948
rect 267096 336864 267148 336870
rect 267096 336806 267148 336812
rect 267004 335368 267056 335374
rect 267004 335310 267056 335316
rect 266740 331894 266860 331922
rect 266636 326392 266688 326398
rect 266636 326334 266688 326340
rect 266740 6798 266768 331894
rect 266820 326392 266872 326398
rect 266820 326334 266872 326340
rect 266832 6866 266860 326334
rect 267108 319666 267136 336806
rect 267292 335594 267320 340068
rect 267476 336870 267504 340068
rect 267568 337278 267596 340068
rect 267556 337272 267608 337278
rect 267556 337214 267608 337220
rect 267464 336864 267516 336870
rect 267464 336806 267516 336812
rect 267372 336796 267424 336802
rect 267372 336738 267424 336744
rect 267200 335566 267320 335594
rect 267096 319660 267148 319666
rect 267096 319602 267148 319608
rect 267200 10878 267228 335566
rect 267384 331922 267412 336738
rect 267464 335708 267516 335714
rect 267464 335650 267516 335656
rect 267292 331894 267412 331922
rect 267292 10946 267320 331894
rect 267372 326392 267424 326398
rect 267372 326334 267424 326340
rect 267280 10940 267332 10946
rect 267280 10882 267332 10888
rect 267188 10872 267240 10878
rect 267188 10814 267240 10820
rect 267384 10810 267412 326334
rect 267476 318850 267504 335650
rect 267660 326398 267688 340068
rect 267740 337136 267792 337142
rect 267738 337104 267740 337113
rect 267792 337104 267794 337113
rect 267738 337039 267794 337048
rect 267844 336870 267872 340068
rect 267832 336864 267884 336870
rect 267832 336806 267884 336812
rect 267740 336796 267792 336802
rect 267740 336738 267792 336744
rect 267752 326398 267780 336738
rect 267832 336728 267884 336734
rect 267832 336670 267884 336676
rect 267648 326392 267700 326398
rect 267648 326334 267700 326340
rect 267740 326392 267792 326398
rect 267740 326334 267792 326340
rect 267464 318844 267516 318850
rect 267464 318786 267516 318792
rect 267464 317484 267516 317490
rect 267464 317426 267516 317432
rect 267476 75886 267504 317426
rect 267464 75880 267516 75886
rect 267464 75822 267516 75828
rect 267464 66292 267516 66298
rect 267464 66234 267516 66240
rect 267476 11014 267504 66234
rect 267464 11008 267516 11014
rect 267464 10950 267516 10956
rect 267372 10804 267424 10810
rect 267372 10746 267424 10752
rect 267004 8288 267056 8294
rect 267004 8230 267056 8236
rect 266820 6860 266872 6866
rect 266820 6802 266872 6808
rect 266728 6792 266780 6798
rect 266728 6734 266780 6740
rect 266544 6724 266596 6730
rect 266544 6666 266596 6672
rect 266452 6656 266504 6662
rect 266452 6598 266504 6604
rect 266176 5976 266228 5982
rect 266176 5918 266228 5924
rect 265348 4208 265400 4214
rect 265348 4150 265400 4156
rect 265808 4208 265860 4214
rect 265808 4150 265860 4156
rect 258540 4140 258592 4146
rect 258540 4082 258592 4088
rect 259828 4140 259880 4146
rect 259828 4082 259880 4088
rect 262864 4140 262916 4146
rect 262864 4082 262916 4088
rect 264612 4140 264664 4146
rect 264612 4082 264664 4088
rect 258632 4072 258684 4078
rect 258632 4014 258684 4020
rect 257712 4004 257764 4010
rect 257712 3946 257764 3952
rect 257160 3936 257212 3942
rect 257160 3878 257212 3884
rect 257068 3868 257120 3874
rect 257068 3810 257120 3816
rect 256516 1896 256568 1902
rect 256516 1838 256568 1844
rect 257436 1896 257488 1902
rect 257436 1838 257488 1844
rect 256252 598 256372 626
rect 256252 480 256280 598
rect 257448 480 257476 1838
rect 258644 480 258672 4014
rect 259840 480 259868 4082
rect 261024 4004 261076 4010
rect 261024 3946 261076 3952
rect 261036 480 261064 3946
rect 262220 3936 262272 3942
rect 262220 3878 262272 3884
rect 262232 480 262260 3878
rect 263416 3868 263468 3874
rect 263416 3810 263468 3816
rect 263428 480 263456 3810
rect 264624 480 264652 4082
rect 265820 480 265848 4150
rect 267016 480 267044 8230
rect 267844 6390 267872 336670
rect 267936 335594 267964 340068
rect 268028 337346 268056 340068
rect 268108 337952 268160 337958
rect 268108 337894 268160 337900
rect 268016 337340 268068 337346
rect 268016 337282 268068 337288
rect 268016 337204 268068 337210
rect 268016 337146 268068 337152
rect 268028 335714 268056 337146
rect 268120 336394 268148 337894
rect 268108 336388 268160 336394
rect 268108 336330 268160 336336
rect 268016 335708 268068 335714
rect 268016 335650 268068 335656
rect 267936 335566 268148 335594
rect 268016 335504 268068 335510
rect 268016 335446 268068 335452
rect 267924 326392 267976 326398
rect 267924 326334 267976 326340
rect 267936 6526 267964 326334
rect 267924 6520 267976 6526
rect 267924 6462 267976 6468
rect 268028 6458 268056 335446
rect 268120 33810 268148 335566
rect 268212 332228 268240 340068
rect 268304 336802 268332 340068
rect 268410 340054 268516 340082
rect 268384 336864 268436 336870
rect 268384 336806 268436 336812
rect 268292 336796 268344 336802
rect 268292 336738 268344 336744
rect 268212 332200 268332 332228
rect 268304 316946 268332 332200
rect 268396 325242 268424 336806
rect 268488 335594 268516 340054
rect 268580 335714 268608 340068
rect 268672 337210 268700 340068
rect 268660 337204 268712 337210
rect 268660 337146 268712 337152
rect 268568 335708 268620 335714
rect 268568 335650 268620 335656
rect 268488 335566 268700 335594
rect 268568 335504 268620 335510
rect 268568 335446 268620 335452
rect 268384 325236 268436 325242
rect 268384 325178 268436 325184
rect 268292 316940 268344 316946
rect 268292 316882 268344 316888
rect 268580 311302 268608 335446
rect 268568 311296 268620 311302
rect 268568 311238 268620 311244
rect 268120 33782 268332 33810
rect 268108 6928 268160 6934
rect 268108 6870 268160 6876
rect 268016 6452 268068 6458
rect 268016 6394 268068 6400
rect 267832 6384 267884 6390
rect 267832 6326 267884 6332
rect 268120 480 268148 6870
rect 268304 6594 268332 33782
rect 268672 10674 268700 335566
rect 268660 10668 268712 10674
rect 268660 10610 268712 10616
rect 268764 10606 268792 340068
rect 268856 340054 268962 340082
rect 268856 335510 268884 340054
rect 269040 337498 269068 340068
rect 269146 340054 269252 340082
rect 268948 337470 269068 337498
rect 268948 336802 268976 337470
rect 269028 337340 269080 337346
rect 269028 337282 269080 337288
rect 268936 336796 268988 336802
rect 268936 336738 268988 336744
rect 269040 336734 269068 337282
rect 269120 337068 269172 337074
rect 269120 337010 269172 337016
rect 269028 336728 269080 336734
rect 269028 336670 269080 336676
rect 268936 335708 268988 335714
rect 268936 335650 268988 335656
rect 268844 335504 268896 335510
rect 268844 335446 268896 335452
rect 268948 333538 268976 335650
rect 268936 333532 268988 333538
rect 268936 333474 268988 333480
rect 269028 327140 269080 327146
rect 269028 327082 269080 327088
rect 269040 306474 269068 327082
rect 268844 306468 268896 306474
rect 268844 306410 268896 306416
rect 269028 306468 269080 306474
rect 269028 306410 269080 306416
rect 268856 200122 268884 306410
rect 268844 200116 268896 200122
rect 268844 200058 268896 200064
rect 269028 200116 269080 200122
rect 269028 200058 269080 200064
rect 269040 190505 269068 200058
rect 268842 190496 268898 190505
rect 268842 190431 268898 190440
rect 269026 190496 269082 190505
rect 269026 190431 269082 190440
rect 268856 178022 268884 190431
rect 268844 178016 268896 178022
rect 268844 177958 268896 177964
rect 268936 168428 268988 168434
rect 268936 168370 268988 168376
rect 268948 161498 268976 168370
rect 268844 161492 268896 161498
rect 268844 161434 268896 161440
rect 268936 161492 268988 161498
rect 268936 161434 268988 161440
rect 268856 160070 268884 161434
rect 268844 160064 268896 160070
rect 268844 160006 268896 160012
rect 268936 150476 268988 150482
rect 268936 150418 268988 150424
rect 268948 142186 268976 150418
rect 268844 142180 268896 142186
rect 268844 142122 268896 142128
rect 268936 142180 268988 142186
rect 268936 142122 268988 142128
rect 268856 121446 268884 142122
rect 268844 121440 268896 121446
rect 268844 121382 268896 121388
rect 268844 111920 268896 111926
rect 268844 111862 268896 111868
rect 268856 111790 268884 111862
rect 268844 111784 268896 111790
rect 268844 111726 268896 111732
rect 268844 100768 268896 100774
rect 268844 100710 268896 100716
rect 268856 92478 268884 100710
rect 268844 92472 268896 92478
rect 268844 92414 268896 92420
rect 268936 87100 268988 87106
rect 268936 87042 268988 87048
rect 268948 76634 268976 87042
rect 268936 76628 268988 76634
rect 268936 76570 268988 76576
rect 269028 71800 269080 71806
rect 269028 71742 269080 71748
rect 269040 68542 269068 71742
rect 268844 68536 268896 68542
rect 268844 68478 268896 68484
rect 269028 68536 269080 68542
rect 269028 68478 269080 68484
rect 268856 26246 268884 68478
rect 268844 26240 268896 26246
rect 268844 26182 268896 26188
rect 268844 16652 268896 16658
rect 268844 16594 268896 16600
rect 268856 10742 268884 16594
rect 268844 10736 268896 10742
rect 268844 10678 268896 10684
rect 268752 10600 268804 10606
rect 268752 10542 268804 10548
rect 269132 10402 269160 337010
rect 269224 10538 269252 340054
rect 269316 328030 269344 340068
rect 269408 337006 269436 340068
rect 269396 337000 269448 337006
rect 269396 336942 269448 336948
rect 269500 336938 269528 340068
rect 269488 336932 269540 336938
rect 269488 336874 269540 336880
rect 269580 336864 269632 336870
rect 269580 336806 269632 336812
rect 269396 336796 269448 336802
rect 269396 336738 269448 336744
rect 269304 328024 269356 328030
rect 269304 327966 269356 327972
rect 269212 10532 269264 10538
rect 269212 10474 269264 10480
rect 269120 10396 269172 10402
rect 269120 10338 269172 10344
rect 268292 6588 268344 6594
rect 268292 6530 268344 6536
rect 269408 6254 269436 336738
rect 269488 335640 269540 335646
rect 269488 335582 269540 335588
rect 269500 326890 269528 335582
rect 269592 327010 269620 336806
rect 269684 327026 269712 340068
rect 269776 336802 269804 340068
rect 269868 337074 269896 340068
rect 269960 340054 270066 340082
rect 269856 337068 269908 337074
rect 269856 337010 269908 337016
rect 269764 336796 269816 336802
rect 269764 336738 269816 336744
rect 269580 327004 269632 327010
rect 269684 326998 269804 327026
rect 269580 326946 269632 326952
rect 269500 326862 269712 326890
rect 269488 326800 269540 326806
rect 269488 326742 269540 326748
rect 269396 6248 269448 6254
rect 269396 6190 269448 6196
rect 269500 6186 269528 326742
rect 269684 307902 269712 326862
rect 269776 323882 269804 326998
rect 269764 323876 269816 323882
rect 269764 323818 269816 323824
rect 269960 309942 269988 340054
rect 270040 336932 270092 336938
rect 270040 336874 270092 336880
rect 269948 309936 270000 309942
rect 269948 309878 270000 309884
rect 269672 307896 269724 307902
rect 269672 307838 269724 307844
rect 269580 307692 269632 307698
rect 269580 307634 269632 307640
rect 269592 56574 269620 307634
rect 269580 56568 269632 56574
rect 269580 56510 269632 56516
rect 269672 53644 269724 53650
rect 269672 53586 269724 53592
rect 269684 37262 269712 53586
rect 269580 37256 269632 37262
rect 269580 37198 269632 37204
rect 269672 37256 269724 37262
rect 269672 37198 269724 37204
rect 269592 27554 269620 37198
rect 269592 27526 269712 27554
rect 269684 18086 269712 27526
rect 269672 18080 269724 18086
rect 269672 18022 269724 18028
rect 269580 18012 269632 18018
rect 269580 17954 269632 17960
rect 269592 17898 269620 17954
rect 269592 17870 269712 17898
rect 269684 8430 269712 17870
rect 270052 10470 270080 336874
rect 270144 336870 270172 340068
rect 270132 336864 270184 336870
rect 270132 336806 270184 336812
rect 270132 336728 270184 336734
rect 270132 336670 270184 336676
rect 270040 10464 270092 10470
rect 270040 10406 270092 10412
rect 269672 8424 269724 8430
rect 269672 8366 269724 8372
rect 269580 8356 269632 8362
rect 269580 8298 269632 8304
rect 269488 6180 269540 6186
rect 269488 6122 269540 6128
rect 269304 4752 269356 4758
rect 269304 4694 269356 4700
rect 269316 480 269344 4694
rect 269592 2854 269620 8298
rect 270144 6322 270172 336670
rect 270236 10334 270264 340068
rect 270328 340054 270434 340082
rect 270328 335646 270356 340054
rect 270316 335640 270368 335646
rect 270316 335582 270368 335588
rect 270512 330818 270540 340068
rect 270500 330812 270552 330818
rect 270500 330754 270552 330760
rect 270604 321094 270632 340068
rect 270788 334150 270816 340068
rect 270880 338162 270908 340068
rect 270868 338156 270920 338162
rect 270868 338098 270920 338104
rect 270776 334144 270828 334150
rect 270776 334086 270828 334092
rect 270972 332330 271000 340068
rect 270788 332302 271000 332330
rect 271064 340054 271170 340082
rect 270788 325174 270816 332302
rect 270868 332240 270920 332246
rect 270868 332182 270920 332188
rect 270776 325168 270828 325174
rect 270776 325110 270828 325116
rect 270592 321088 270644 321094
rect 270592 321030 270644 321036
rect 270880 318238 270908 332182
rect 270960 332172 271012 332178
rect 270960 332114 271012 332120
rect 270868 318232 270920 318238
rect 270868 318174 270920 318180
rect 270500 318096 270552 318102
rect 270500 318038 270552 318044
rect 270224 10328 270276 10334
rect 270224 10270 270276 10276
rect 270132 6316 270184 6322
rect 270132 6258 270184 6264
rect 269580 2848 269632 2854
rect 269580 2790 269632 2796
rect 270512 1426 270540 318038
rect 270972 307154 271000 332114
rect 270960 307148 271012 307154
rect 270960 307090 271012 307096
rect 270592 5500 270644 5506
rect 270592 5442 270644 5448
rect 270500 1420 270552 1426
rect 270500 1362 270552 1368
rect 270604 1034 270632 5442
rect 271064 2990 271092 340054
rect 271248 333470 271276 340068
rect 271236 333464 271288 333470
rect 271236 333406 271288 333412
rect 271340 332246 271368 340068
rect 271328 332240 271380 332246
rect 271328 332182 271380 332188
rect 271524 299538 271552 340068
rect 271616 332110 271644 340068
rect 271708 332178 271736 340068
rect 271788 334144 271840 334150
rect 271788 334086 271840 334092
rect 271696 332172 271748 332178
rect 271696 332114 271748 332120
rect 271604 332104 271656 332110
rect 271604 332046 271656 332052
rect 271144 299532 271196 299538
rect 271144 299474 271196 299480
rect 271512 299532 271564 299538
rect 271512 299474 271564 299480
rect 271156 66230 271184 299474
rect 271800 295361 271828 334086
rect 271892 333334 271920 340068
rect 271984 338094 272012 340068
rect 271972 338088 272024 338094
rect 271972 338030 272024 338036
rect 271972 336796 272024 336802
rect 271972 336738 272024 336744
rect 271880 333328 271932 333334
rect 271880 333270 271932 333276
rect 271602 295352 271658 295361
rect 271602 295287 271658 295296
rect 271786 295352 271842 295361
rect 271786 295287 271842 295296
rect 271616 250458 271644 295287
rect 271524 250430 271644 250458
rect 271524 245682 271552 250430
rect 271512 245676 271564 245682
rect 271512 245618 271564 245624
rect 271788 245676 271840 245682
rect 271788 245618 271840 245624
rect 271800 237454 271828 245618
rect 271604 237448 271656 237454
rect 271604 237390 271656 237396
rect 271788 237448 271840 237454
rect 271788 237390 271840 237396
rect 271616 195974 271644 237390
rect 271604 195968 271656 195974
rect 271604 195910 271656 195916
rect 271696 186380 271748 186386
rect 271696 186322 271748 186328
rect 271708 178090 271736 186322
rect 271604 178084 271656 178090
rect 271604 178026 271656 178032
rect 271696 178084 271748 178090
rect 271696 178026 271748 178032
rect 271616 160070 271644 178026
rect 271604 160064 271656 160070
rect 271604 160006 271656 160012
rect 271696 149184 271748 149190
rect 271616 149132 271696 149138
rect 271616 149126 271748 149132
rect 271616 149110 271736 149126
rect 271616 149054 271644 149110
rect 271604 149048 271656 149054
rect 271604 148990 271656 148996
rect 271604 139528 271656 139534
rect 271604 139470 271656 139476
rect 271616 139398 271644 139470
rect 271604 139392 271656 139398
rect 271604 139334 271656 139340
rect 271512 129804 271564 129810
rect 271512 129746 271564 129752
rect 271524 126290 271552 129746
rect 271524 126262 271644 126290
rect 271144 66224 271196 66230
rect 271144 66166 271196 66172
rect 271236 66224 271288 66230
rect 271236 66166 271288 66172
rect 271248 48346 271276 66166
rect 271144 48340 271196 48346
rect 271144 48282 271196 48288
rect 271236 48340 271288 48346
rect 271236 48282 271288 48288
rect 271156 3058 271184 48282
rect 271616 37262 271644 126262
rect 271604 37256 271656 37262
rect 271604 37198 271656 37204
rect 271604 18012 271656 18018
rect 271604 17954 271656 17960
rect 271144 3052 271196 3058
rect 271144 2994 271196 3000
rect 271052 2984 271104 2990
rect 271052 2926 271104 2932
rect 271616 2922 271644 17954
rect 271984 3194 272012 336738
rect 272076 316878 272104 340068
rect 272260 336802 272288 340068
rect 272352 336802 272380 340068
rect 272248 336796 272300 336802
rect 272248 336738 272300 336744
rect 272340 336796 272392 336802
rect 272340 336738 272392 336744
rect 272340 335640 272392 335646
rect 272340 335582 272392 335588
rect 272248 333328 272300 333334
rect 272248 333270 272300 333276
rect 272156 326392 272208 326398
rect 272156 326334 272208 326340
rect 272064 316872 272116 316878
rect 272064 316814 272116 316820
rect 272168 3330 272196 326334
rect 272156 3324 272208 3330
rect 272156 3266 272208 3272
rect 271972 3188 272024 3194
rect 271972 3130 272024 3136
rect 272260 3126 272288 333270
rect 272352 3262 272380 335582
rect 272444 305726 272472 340068
rect 272536 340054 272642 340082
rect 272536 335646 272564 340054
rect 272720 336802 272748 340068
rect 272616 336796 272668 336802
rect 272616 336738 272668 336744
rect 272708 336796 272760 336802
rect 272708 336738 272760 336744
rect 272524 335640 272576 335646
rect 272524 335582 272576 335588
rect 272524 335504 272576 335510
rect 272524 335446 272576 335452
rect 272432 305720 272484 305726
rect 272432 305662 272484 305668
rect 272536 8294 272564 335446
rect 272628 330750 272656 336738
rect 272616 330744 272668 330750
rect 272616 330686 272668 330692
rect 272812 291922 272840 340068
rect 272892 336796 272944 336802
rect 272892 336738 272944 336744
rect 272904 325106 272932 336738
rect 272996 326398 273024 340068
rect 273088 336802 273116 340068
rect 273076 336796 273128 336802
rect 273076 336738 273128 336744
rect 273180 336734 273208 340068
rect 273260 337408 273312 337414
rect 273260 337350 273312 337356
rect 273168 336728 273220 336734
rect 273168 336670 273220 336676
rect 273076 336660 273128 336666
rect 273076 336602 273128 336608
rect 273088 326602 273116 336602
rect 273272 334830 273300 337350
rect 273364 337074 273392 340068
rect 273456 337414 273484 340068
rect 273444 337408 273496 337414
rect 273444 337350 273496 337356
rect 273352 337068 273404 337074
rect 273352 337010 273404 337016
rect 273548 337006 273576 340068
rect 273640 340054 273746 340082
rect 273536 337000 273588 337006
rect 273640 336977 273668 340054
rect 273536 336942 273588 336948
rect 273626 336968 273682 336977
rect 273352 336932 273404 336938
rect 273824 336938 273852 340068
rect 273626 336903 273682 336912
rect 273812 336932 273864 336938
rect 273352 336874 273404 336880
rect 273812 336874 273864 336880
rect 273260 334824 273312 334830
rect 273260 334766 273312 334772
rect 273364 329254 273392 336874
rect 273628 336864 273680 336870
rect 273628 336806 273680 336812
rect 273810 336832 273866 336841
rect 273444 336796 273496 336802
rect 273444 336738 273496 336744
rect 273352 329248 273404 329254
rect 273352 329190 273404 329196
rect 273168 327140 273220 327146
rect 273168 327082 273220 327088
rect 273076 326596 273128 326602
rect 273076 326538 273128 326544
rect 272984 326392 273036 326398
rect 272984 326334 273036 326340
rect 272892 325100 272944 325106
rect 272892 325042 272944 325048
rect 273180 304366 273208 327082
rect 273168 304360 273220 304366
rect 273168 304302 273220 304308
rect 273456 303006 273484 336738
rect 273536 336728 273588 336734
rect 273536 336670 273588 336676
rect 273444 303000 273496 303006
rect 273444 302942 273496 302948
rect 272800 291916 272852 291922
rect 272800 291858 272852 291864
rect 272524 8288 272576 8294
rect 272524 8230 272576 8236
rect 272892 5364 272944 5370
rect 272892 5306 272944 5312
rect 272340 3256 272392 3262
rect 272340 3198 272392 3204
rect 272248 3120 272300 3126
rect 272248 3062 272300 3068
rect 271604 2916 271656 2922
rect 271604 2858 271656 2864
rect 271696 1420 271748 1426
rect 271696 1362 271748 1368
rect 270512 1006 270632 1034
rect 270512 480 270540 1006
rect 271708 480 271736 1362
rect 272904 480 272932 5306
rect 273548 4010 273576 336670
rect 273640 327894 273668 336806
rect 273916 336802 273944 340068
rect 274008 340054 274114 340082
rect 273810 336767 273866 336776
rect 273904 336796 273956 336802
rect 273628 327888 273680 327894
rect 273628 327830 273680 327836
rect 273628 311228 273680 311234
rect 273628 311170 273680 311176
rect 273640 309126 273668 311170
rect 273628 309120 273680 309126
rect 273628 309062 273680 309068
rect 273628 296744 273680 296750
rect 273628 296686 273680 296692
rect 273640 263634 273668 296686
rect 273824 289814 273852 336767
rect 273904 336738 273956 336744
rect 274008 311234 274036 340054
rect 274088 337000 274140 337006
rect 274088 336942 274140 336948
rect 274100 315450 274128 336942
rect 274192 336870 274220 340068
rect 274180 336864 274232 336870
rect 274180 336806 274232 336812
rect 274284 326380 274312 340068
rect 274364 337068 274416 337074
rect 274364 337010 274416 337016
rect 274376 336734 274404 337010
rect 274468 336802 274496 340068
rect 274456 336796 274508 336802
rect 274456 336738 274508 336744
rect 274364 336728 274416 336734
rect 274364 336670 274416 336676
rect 274364 327140 274416 327146
rect 274364 327082 274416 327088
rect 274192 326352 274312 326380
rect 274088 315444 274140 315450
rect 274088 315386 274140 315392
rect 273996 311228 274048 311234
rect 273996 311170 274048 311176
rect 274192 290562 274220 326352
rect 274376 325650 274404 327082
rect 274364 325644 274416 325650
rect 274364 325586 274416 325592
rect 274560 319598 274588 340068
rect 274666 340054 274772 340082
rect 274744 326806 274772 340054
rect 274836 333062 274864 340068
rect 274928 337074 274956 340068
rect 274916 337068 274968 337074
rect 274916 337010 274968 337016
rect 275020 336802 275048 340068
rect 275008 336796 275060 336802
rect 275008 336738 275060 336744
rect 274824 333056 274876 333062
rect 274824 332998 274876 333004
rect 275008 331220 275060 331226
rect 275008 331162 275060 331168
rect 274732 326800 274784 326806
rect 274732 326742 274784 326748
rect 274548 319592 274600 319598
rect 274548 319534 274600 319540
rect 274364 316056 274416 316062
rect 274364 315998 274416 316004
rect 274376 311216 274404 315998
rect 274376 311188 274496 311216
rect 274468 299606 274496 311188
rect 274456 299600 274508 299606
rect 274456 299542 274508 299548
rect 274364 299464 274416 299470
rect 274364 299406 274416 299412
rect 274180 290556 274232 290562
rect 274180 290498 274232 290504
rect 273812 289808 273864 289814
rect 273812 289750 273864 289756
rect 273904 289808 273956 289814
rect 273904 289750 273956 289756
rect 273628 263628 273680 263634
rect 273628 263570 273680 263576
rect 273720 263560 273772 263566
rect 273720 263502 273772 263508
rect 273732 251258 273760 263502
rect 273720 251252 273772 251258
rect 273720 251194 273772 251200
rect 273812 251116 273864 251122
rect 273812 251058 273864 251064
rect 273824 241534 273852 251058
rect 273720 241528 273772 241534
rect 273720 241470 273772 241476
rect 273812 241528 273864 241534
rect 273812 241470 273864 241476
rect 273732 195242 273760 241470
rect 273916 214554 273944 289750
rect 274376 284968 274404 299406
rect 274284 284940 274404 284968
rect 274284 272626 274312 284940
rect 274192 272598 274312 272626
rect 274192 249830 274220 272598
rect 274180 249824 274232 249830
rect 274180 249766 274232 249772
rect 274272 249824 274324 249830
rect 274272 249766 274324 249772
rect 274284 247042 274312 249766
rect 274272 247036 274324 247042
rect 274272 246978 274324 246984
rect 274180 237448 274232 237454
rect 274180 237390 274232 237396
rect 274192 229090 274220 237390
rect 274180 229084 274232 229090
rect 274180 229026 274232 229032
rect 274364 229016 274416 229022
rect 274364 228958 274416 228964
rect 273916 214526 274036 214554
rect 274008 202910 274036 214526
rect 274376 213994 274404 228958
rect 274180 213988 274232 213994
rect 274180 213930 274232 213936
rect 274364 213988 274416 213994
rect 274364 213930 274416 213936
rect 273904 202904 273956 202910
rect 273904 202846 273956 202852
rect 273996 202904 274048 202910
rect 273996 202846 274048 202852
rect 273732 195214 273852 195242
rect 273824 183598 273852 195214
rect 273916 184278 273944 202846
rect 274192 200122 274220 213930
rect 274180 200116 274232 200122
rect 274180 200058 274232 200064
rect 274272 200048 274324 200054
rect 274272 199990 274324 199996
rect 273904 184272 273956 184278
rect 274284 184226 274312 199990
rect 273904 184214 273956 184220
rect 274192 184198 274312 184226
rect 273720 183592 273772 183598
rect 273720 183534 273772 183540
rect 273812 183592 273864 183598
rect 273812 183534 273864 183540
rect 273732 175930 273760 183534
rect 273812 180804 273864 180810
rect 273812 180746 273864 180752
rect 273640 175902 273760 175930
rect 273640 164286 273668 175902
rect 273824 171086 273852 180746
rect 273812 171080 273864 171086
rect 273812 171022 273864 171028
rect 273904 171080 273956 171086
rect 273904 171022 273956 171028
rect 273628 164280 273680 164286
rect 273628 164222 273680 164228
rect 273720 164144 273772 164150
rect 273720 164086 273772 164092
rect 273732 142186 273760 164086
rect 273916 142186 273944 171022
rect 274192 160070 274220 184198
rect 274180 160064 274232 160070
rect 274180 160006 274232 160012
rect 274180 159928 274232 159934
rect 274180 159870 274232 159876
rect 273628 142180 273680 142186
rect 273628 142122 273680 142128
rect 273720 142180 273772 142186
rect 273720 142122 273772 142128
rect 273812 142180 273864 142186
rect 273812 142122 273864 142128
rect 273904 142180 273956 142186
rect 273904 142122 273956 142128
rect 273640 111874 273668 142122
rect 273824 133890 273852 142122
rect 273812 133884 273864 133890
rect 273812 133826 273864 133832
rect 273996 133884 274048 133890
rect 273996 133826 274048 133832
rect 274008 128874 274036 133826
rect 274192 131102 274220 159870
rect 274180 131096 274232 131102
rect 274180 131038 274232 131044
rect 273916 128846 274036 128874
rect 273916 120086 273944 128846
rect 274088 121508 274140 121514
rect 274088 121450 274140 121456
rect 273904 120080 273956 120086
rect 273904 120022 273956 120028
rect 273640 111846 273760 111874
rect 274100 111858 274128 121450
rect 273732 74594 273760 111846
rect 274088 111852 274140 111858
rect 274088 111794 274140 111800
rect 274272 111852 274324 111858
rect 274272 111794 274324 111800
rect 273996 110492 274048 110498
rect 273996 110434 274048 110440
rect 274008 92478 274036 110434
rect 274284 102218 274312 111794
rect 274192 102190 274312 102218
rect 274192 99346 274220 102190
rect 274180 99340 274232 99346
rect 274180 99282 274232 99288
rect 273812 92472 273864 92478
rect 273812 92414 273864 92420
rect 273996 92472 274048 92478
rect 273996 92414 274048 92420
rect 273824 91089 273852 92414
rect 273810 91080 273866 91089
rect 273810 91015 273866 91024
rect 274086 91080 274142 91089
rect 274086 91015 274142 91024
rect 274100 76634 274128 91015
rect 274180 82884 274232 82890
rect 274180 82826 274232 82832
rect 274192 76634 274220 82826
rect 274088 76628 274140 76634
rect 274088 76570 274140 76576
rect 274180 76628 274232 76634
rect 274180 76570 274232 76576
rect 274456 76628 274508 76634
rect 274456 76570 274508 76576
rect 273628 74588 273680 74594
rect 273628 74530 273680 74536
rect 273720 74588 273772 74594
rect 273720 74530 273772 74536
rect 273640 66366 273668 74530
rect 274468 71754 274496 76570
rect 274376 71726 274496 71754
rect 273628 66360 273680 66366
rect 273628 66302 273680 66308
rect 273628 66224 273680 66230
rect 273628 66166 273680 66172
rect 273640 58682 273668 66166
rect 274376 63578 274404 71726
rect 273904 63572 273956 63578
rect 273904 63514 273956 63520
rect 274364 63572 274416 63578
rect 274364 63514 274416 63520
rect 273916 63458 273944 63514
rect 273916 63430 274036 63458
rect 273628 58676 273680 58682
rect 273628 58618 273680 58624
rect 273904 58676 273956 58682
rect 273904 58618 273956 58624
rect 273916 50402 273944 58618
rect 273824 50374 273944 50402
rect 273824 48362 273852 50374
rect 273732 48334 273852 48362
rect 274008 48346 274036 63430
rect 274272 63436 274324 63442
rect 274272 63378 274324 63384
rect 273904 48340 273956 48346
rect 273732 37262 273760 48334
rect 273904 48282 273956 48288
rect 273996 48340 274048 48346
rect 273996 48282 274048 48288
rect 273628 37256 273680 37262
rect 273628 37198 273680 37204
rect 273720 37256 273772 37262
rect 273720 37198 273772 37204
rect 273640 4078 273668 37198
rect 273916 33810 273944 48282
rect 273824 33782 273944 33810
rect 273824 4146 273852 33782
rect 274284 27606 274312 63378
rect 274272 27600 274324 27606
rect 274272 27542 274324 27548
rect 274272 18012 274324 18018
rect 274272 17954 274324 17960
rect 274088 5432 274140 5438
rect 274088 5374 274140 5380
rect 273812 4140 273864 4146
rect 273812 4082 273864 4088
rect 273628 4072 273680 4078
rect 273628 4014 273680 4020
rect 273536 4004 273588 4010
rect 273536 3946 273588 3952
rect 274100 480 274128 5374
rect 274284 3398 274312 17954
rect 275020 3738 275048 331162
rect 275112 3874 275140 340068
rect 275296 337006 275324 340068
rect 275284 337000 275336 337006
rect 275284 336942 275336 336948
rect 275192 336796 275244 336802
rect 275192 336738 275244 336744
rect 275284 336796 275336 336802
rect 275284 336738 275336 336744
rect 275204 323746 275232 336738
rect 275192 323740 275244 323746
rect 275192 323682 275244 323688
rect 275296 8378 275324 336738
rect 275388 314090 275416 340068
rect 275480 336802 275508 340068
rect 275560 337000 275612 337006
rect 275560 336942 275612 336948
rect 275468 336796 275520 336802
rect 275468 336738 275520 336744
rect 275572 333402 275600 336942
rect 275664 336258 275692 340068
rect 275652 336252 275704 336258
rect 275652 336194 275704 336200
rect 275560 333396 275612 333402
rect 275560 333338 275612 333344
rect 275756 333146 275784 340068
rect 275572 333118 275784 333146
rect 275376 314084 275428 314090
rect 275376 314026 275428 314032
rect 275572 301578 275600 333118
rect 275744 333056 275796 333062
rect 275744 332998 275796 333004
rect 275560 301572 275612 301578
rect 275560 301514 275612 301520
rect 275296 8350 275416 8378
rect 275284 8288 275336 8294
rect 275284 8230 275336 8236
rect 275100 3868 275152 3874
rect 275100 3810 275152 3816
rect 275008 3732 275060 3738
rect 275008 3674 275060 3680
rect 274272 3392 274324 3398
rect 274272 3334 274324 3340
rect 275296 480 275324 8230
rect 275388 3806 275416 8350
rect 275756 3942 275784 332998
rect 275848 331362 275876 340068
rect 276032 337822 276060 340068
rect 276020 337816 276072 337822
rect 276020 337758 276072 337764
rect 276020 337000 276072 337006
rect 276020 336942 276072 336948
rect 275836 331356 275888 331362
rect 275836 331298 275888 331304
rect 276032 300218 276060 336942
rect 276124 333334 276152 340068
rect 276230 340054 276336 340082
rect 276204 336864 276256 336870
rect 276204 336806 276256 336812
rect 276112 333328 276164 333334
rect 276112 333270 276164 333276
rect 276216 333282 276244 336806
rect 276308 334150 276336 340054
rect 276400 335714 276428 340068
rect 276492 336802 276520 340068
rect 276480 336796 276532 336802
rect 276480 336738 276532 336744
rect 276388 335708 276440 335714
rect 276388 335650 276440 335656
rect 276584 334234 276612 340068
rect 276400 334206 276612 334234
rect 276296 334144 276348 334150
rect 276296 334086 276348 334092
rect 276216 333254 276336 333282
rect 276308 316810 276336 333254
rect 276296 316804 276348 316810
rect 276296 316746 276348 316752
rect 276020 300212 276072 300218
rect 276020 300154 276072 300160
rect 275744 3936 275796 3942
rect 275744 3878 275796 3884
rect 275376 3800 275428 3806
rect 275376 3742 275428 3748
rect 276400 3602 276428 334206
rect 276480 334144 276532 334150
rect 276480 334086 276532 334092
rect 276492 8106 276520 334086
rect 276572 333328 276624 333334
rect 276572 333270 276624 333276
rect 276584 321026 276612 333270
rect 276768 322386 276796 340068
rect 276860 337006 276888 340068
rect 276966 340054 277072 340082
rect 277044 338570 277072 340054
rect 277032 338564 277084 338570
rect 277032 338506 277084 338512
rect 276940 337408 276992 337414
rect 276940 337350 276992 337356
rect 276848 337000 276900 337006
rect 276848 336942 276900 336948
rect 276848 336796 276900 336802
rect 276848 336738 276900 336744
rect 276756 322380 276808 322386
rect 276756 322322 276808 322328
rect 276572 321020 276624 321026
rect 276572 320962 276624 320968
rect 276860 289202 276888 336738
rect 276848 289196 276900 289202
rect 276848 289138 276900 289144
rect 276952 287706 276980 337350
rect 277032 337272 277084 337278
rect 277032 337214 277084 337220
rect 277044 335617 277072 337214
rect 277136 336870 277164 340068
rect 277228 337414 277256 340068
rect 277334 340054 277440 340082
rect 277216 337408 277268 337414
rect 277216 337350 277268 337356
rect 277412 337278 277440 340054
rect 277504 337890 277532 340068
rect 277492 337884 277544 337890
rect 277492 337826 277544 337832
rect 277400 337272 277452 337278
rect 277400 337214 277452 337220
rect 277400 337136 277452 337142
rect 277400 337078 277452 337084
rect 277124 336864 277176 336870
rect 277124 336806 277176 336812
rect 277216 335708 277268 335714
rect 277216 335650 277268 335656
rect 277030 335608 277086 335617
rect 277030 335543 277086 335552
rect 277032 335436 277084 335442
rect 277032 335378 277084 335384
rect 277044 327078 277072 335378
rect 277228 330682 277256 335650
rect 277306 335370 277362 335379
rect 277306 335305 277362 335314
rect 277320 331294 277348 335305
rect 277308 331288 277360 331294
rect 277308 331230 277360 331236
rect 277216 330676 277268 330682
rect 277216 330618 277268 330624
rect 277412 329186 277440 337078
rect 277596 337006 277624 340068
rect 277702 340054 277808 340082
rect 277584 337000 277636 337006
rect 277584 336942 277636 336948
rect 277492 336864 277544 336870
rect 277492 336806 277544 336812
rect 277400 329180 277452 329186
rect 277400 329122 277452 329128
rect 277032 327072 277084 327078
rect 277032 327014 277084 327020
rect 277124 327072 277176 327078
rect 277124 327014 277176 327020
rect 277030 324320 277086 324329
rect 277030 324255 277086 324264
rect 277044 297378 277072 324255
rect 277136 312610 277164 327014
rect 277400 324352 277452 324358
rect 277398 324320 277400 324329
rect 277452 324320 277454 324329
rect 277398 324255 277454 324264
rect 277504 322318 277532 336806
rect 277584 336796 277636 336802
rect 277584 336738 277636 336744
rect 277492 322312 277544 322318
rect 277492 322254 277544 322260
rect 277136 312582 277348 312610
rect 277044 297350 277256 297378
rect 277124 290488 277176 290494
rect 277124 290430 277176 290436
rect 277136 289814 277164 290430
rect 277124 289808 277176 289814
rect 277124 289750 277176 289756
rect 276940 287700 276992 287706
rect 276940 287642 276992 287648
rect 277228 283626 277256 297350
rect 277320 290494 277348 312582
rect 277596 298790 277624 336738
rect 277780 333418 277808 340054
rect 277872 337210 277900 340068
rect 277860 337204 277912 337210
rect 277860 337146 277912 337152
rect 277860 337068 277912 337074
rect 277860 337010 277912 337016
rect 277872 336802 277900 337010
rect 277964 336802 277992 340068
rect 277860 336796 277912 336802
rect 277860 336738 277912 336744
rect 277952 336796 278004 336802
rect 277952 336738 278004 336744
rect 277780 333390 277992 333418
rect 277860 333328 277912 333334
rect 277860 333270 277912 333276
rect 277768 310140 277820 310146
rect 277768 310082 277820 310088
rect 277780 302190 277808 310082
rect 277768 302184 277820 302190
rect 277768 302126 277820 302132
rect 277584 298784 277636 298790
rect 277584 298726 277636 298732
rect 277308 290488 277360 290494
rect 277308 290430 277360 290436
rect 277308 289808 277360 289814
rect 277308 289750 277360 289756
rect 277032 283620 277084 283626
rect 277032 283562 277084 283568
rect 277216 283620 277268 283626
rect 277216 283562 277268 283568
rect 277044 276049 277072 283562
rect 277320 283506 277348 289750
rect 277228 283478 277348 283506
rect 276846 276040 276902 276049
rect 276846 275975 276902 275984
rect 277030 276040 277086 276049
rect 277030 275975 277086 275984
rect 276860 271130 276888 275975
rect 277228 274650 277256 283478
rect 277216 274644 277268 274650
rect 277216 274586 277268 274592
rect 276860 271102 276980 271130
rect 276952 266354 276980 271102
rect 276940 266348 276992 266354
rect 276940 266290 276992 266296
rect 277216 264988 277268 264994
rect 277216 264930 277268 264936
rect 277032 256760 277084 256766
rect 276952 256708 277032 256714
rect 276952 256702 277084 256708
rect 276952 256698 277072 256702
rect 276940 256692 277072 256698
rect 276992 256686 277072 256692
rect 276940 256634 276992 256640
rect 277228 255270 277256 264930
rect 277216 255264 277268 255270
rect 277216 255206 277268 255212
rect 276940 249756 276992 249762
rect 276940 249698 276992 249704
rect 276952 247058 276980 249698
rect 276952 247030 277072 247058
rect 277044 229090 277072 247030
rect 277216 247036 277268 247042
rect 277216 246978 277268 246984
rect 277228 241534 277256 246978
rect 277216 241528 277268 241534
rect 277216 241470 277268 241476
rect 277216 237448 277268 237454
rect 277216 237390 277268 237396
rect 276940 229084 276992 229090
rect 276940 229026 276992 229032
rect 277032 229084 277084 229090
rect 277032 229026 277084 229032
rect 276952 200002 276980 229026
rect 277228 209778 277256 237390
rect 277584 212764 277636 212770
rect 277584 212706 277636 212712
rect 277596 212537 277624 212706
rect 277582 212528 277638 212537
rect 277582 212463 277638 212472
rect 277766 212528 277822 212537
rect 277766 212463 277822 212472
rect 277124 209772 277176 209778
rect 277124 209714 277176 209720
rect 277216 209772 277268 209778
rect 277216 209714 277268 209720
rect 277136 208350 277164 209714
rect 277124 208344 277176 208350
rect 277124 208286 277176 208292
rect 277216 208344 277268 208350
rect 277216 208286 277268 208292
rect 276952 199974 277072 200002
rect 277044 195242 277072 199974
rect 277228 198778 277256 208286
rect 277136 198750 277256 198778
rect 277136 197334 277164 198750
rect 277124 197328 277176 197334
rect 277124 197270 277176 197276
rect 277780 195974 277808 212463
rect 277768 195968 277820 195974
rect 277768 195910 277820 195916
rect 276860 195214 277072 195242
rect 276860 190482 276888 195214
rect 276860 190454 276980 190482
rect 276952 183598 276980 190454
rect 277124 187740 277176 187746
rect 277124 187682 277176 187688
rect 277136 183598 277164 187682
rect 276940 183592 276992 183598
rect 276940 183534 276992 183540
rect 277032 183592 277084 183598
rect 277032 183534 277084 183540
rect 277124 183592 277176 183598
rect 277124 183534 277176 183540
rect 277044 175930 277072 183534
rect 277216 183456 277268 183462
rect 277216 183398 277268 183404
rect 277228 178022 277256 183398
rect 277216 178016 277268 178022
rect 277216 177958 277268 177964
rect 277400 178016 277452 178022
rect 277400 177958 277452 177964
rect 276952 175902 277072 175930
rect 276952 164914 276980 175902
rect 276860 164886 276980 164914
rect 276860 160138 276888 164886
rect 277412 160138 277440 177958
rect 276848 160132 276900 160138
rect 276848 160074 276900 160080
rect 277032 160132 277084 160138
rect 277032 160074 277084 160080
rect 277124 160132 277176 160138
rect 277124 160074 277176 160080
rect 277400 160132 277452 160138
rect 277400 160074 277452 160080
rect 277044 132530 277072 160074
rect 277136 158710 277164 160074
rect 277124 158704 277176 158710
rect 277124 158646 277176 158652
rect 277216 158704 277268 158710
rect 277216 158646 277268 158652
rect 277228 149138 277256 158646
rect 277136 149110 277256 149138
rect 277136 149054 277164 149110
rect 277124 149048 277176 149054
rect 277124 148990 277176 148996
rect 277216 139460 277268 139466
rect 277216 139402 277268 139408
rect 276940 132524 276992 132530
rect 276940 132466 276992 132472
rect 277032 132524 277084 132530
rect 277032 132466 277084 132472
rect 276952 111790 276980 132466
rect 277228 116006 277256 139402
rect 277216 116000 277268 116006
rect 277216 115942 277268 115948
rect 276940 111784 276992 111790
rect 276940 111726 276992 111732
rect 277216 102264 277268 102270
rect 277216 102206 277268 102212
rect 277032 102196 277084 102202
rect 277032 102138 277084 102144
rect 276938 100736 276994 100745
rect 276938 100671 276994 100680
rect 276952 91118 276980 100671
rect 276940 91112 276992 91118
rect 276940 91054 276992 91060
rect 277044 68490 277072 102138
rect 277228 100745 277256 102206
rect 277214 100736 277270 100745
rect 277214 100671 277270 100680
rect 277124 91112 277176 91118
rect 277124 91054 277176 91060
rect 277136 84182 277164 91054
rect 277124 84176 277176 84182
rect 277124 84118 277176 84124
rect 277124 74588 277176 74594
rect 277124 74530 277176 74536
rect 277136 73098 277164 74530
rect 277124 73092 277176 73098
rect 277124 73034 277176 73040
rect 276952 68462 277072 68490
rect 276952 68218 276980 68462
rect 276952 68190 277072 68218
rect 277044 53854 277072 68190
rect 277216 63572 277268 63578
rect 277216 63514 277268 63520
rect 276940 53848 276992 53854
rect 276940 53790 276992 53796
rect 277032 53848 277084 53854
rect 277032 53790 277084 53796
rect 276952 45014 276980 53790
rect 277228 48346 277256 63514
rect 277584 60444 277636 60450
rect 277584 60386 277636 60392
rect 277596 53122 277624 60386
rect 277596 53094 277808 53122
rect 277124 48340 277176 48346
rect 277124 48282 277176 48288
rect 277216 48340 277268 48346
rect 277216 48282 277268 48288
rect 276940 45008 276992 45014
rect 276940 44950 276992 44956
rect 276848 37324 276900 37330
rect 276848 37266 276900 37272
rect 276860 33130 276888 37266
rect 276860 33102 276980 33130
rect 276952 19802 276980 33102
rect 276768 19774 276980 19802
rect 276768 19258 276796 19774
rect 276768 19230 276888 19258
rect 276492 8078 276612 8106
rect 276480 5296 276532 5302
rect 276480 5238 276532 5244
rect 276388 3596 276440 3602
rect 276388 3538 276440 3544
rect 276492 480 276520 5238
rect 276584 3670 276612 8078
rect 276572 3664 276624 3670
rect 276572 3606 276624 3612
rect 276860 3466 276888 19230
rect 277136 3534 277164 48282
rect 277780 41410 277808 53094
rect 277768 41404 277820 41410
rect 277768 41346 277820 41352
rect 277768 22160 277820 22166
rect 277768 22102 277820 22108
rect 277780 17270 277808 22102
rect 277768 17264 277820 17270
rect 277768 17206 277820 17212
rect 277676 5228 277728 5234
rect 277676 5170 277728 5176
rect 277124 3528 277176 3534
rect 277124 3470 277176 3476
rect 276848 3460 276900 3466
rect 276848 3402 276900 3408
rect 277688 480 277716 5170
rect 277872 3777 277900 333270
rect 277964 310146 277992 333390
rect 277952 310140 278004 310146
rect 277952 310082 278004 310088
rect 277952 302184 278004 302190
rect 277952 302126 278004 302132
rect 277964 212770 277992 302126
rect 277952 212764 278004 212770
rect 277952 212706 278004 212712
rect 277952 195900 278004 195906
rect 277952 195842 278004 195848
rect 277964 60450 277992 195842
rect 277952 60444 278004 60450
rect 277952 60386 278004 60392
rect 277952 41336 278004 41342
rect 277952 41278 278004 41284
rect 277964 22166 277992 41278
rect 277952 22160 278004 22166
rect 277952 22102 278004 22108
rect 278056 3913 278084 340068
rect 278240 332042 278268 340068
rect 278332 336870 278360 340068
rect 278424 336920 278452 340068
rect 278608 337142 278636 340068
rect 278596 337136 278648 337142
rect 278596 337078 278648 337084
rect 278700 337074 278728 340068
rect 278806 340054 278912 340082
rect 278688 337068 278740 337074
rect 278688 337010 278740 337016
rect 278596 337000 278648 337006
rect 278596 336942 278648 336948
rect 278424 336892 278544 336920
rect 278320 336864 278372 336870
rect 278320 336806 278372 336812
rect 278412 336796 278464 336802
rect 278412 336738 278464 336744
rect 278228 332036 278280 332042
rect 278228 331978 278280 331984
rect 278424 312730 278452 336738
rect 278516 333334 278544 336892
rect 278504 333328 278556 333334
rect 278504 333270 278556 333276
rect 278608 330614 278636 336942
rect 278688 336728 278740 336734
rect 278688 336670 278740 336676
rect 278700 336410 278728 336670
rect 278700 336382 278820 336410
rect 278792 335238 278820 336382
rect 278780 335232 278832 335238
rect 278780 335174 278832 335180
rect 278884 333282 278912 340054
rect 278976 335442 279004 340068
rect 279068 335510 279096 340068
rect 279160 336870 279188 340068
rect 279240 337204 279292 337210
rect 279240 337146 279292 337152
rect 279148 336864 279200 336870
rect 279148 336806 279200 336812
rect 279056 335504 279108 335510
rect 279056 335446 279108 335452
rect 278964 335436 279016 335442
rect 278964 335378 279016 335384
rect 279148 335232 279200 335238
rect 279148 335174 279200 335180
rect 278884 333254 279004 333282
rect 278596 330608 278648 330614
rect 278596 330550 278648 330556
rect 278976 326126 279004 333254
rect 278964 326120 279016 326126
rect 278964 326062 279016 326068
rect 279160 323814 279188 335174
rect 279252 326194 279280 337146
rect 279344 333282 279372 340068
rect 279436 335594 279464 340068
rect 279528 336802 279556 340068
rect 279712 338094 279740 340068
rect 279700 338088 279752 338094
rect 279700 338030 279752 338036
rect 279516 336796 279568 336802
rect 279516 336738 279568 336744
rect 279436 335566 279740 335594
rect 279608 335504 279660 335510
rect 279608 335446 279660 335452
rect 279516 335436 279568 335442
rect 279516 335378 279568 335384
rect 279344 333254 279464 333282
rect 279332 326392 279384 326398
rect 279332 326334 279384 326340
rect 279240 326188 279292 326194
rect 279240 326130 279292 326136
rect 279148 323808 279200 323814
rect 279148 323750 279200 323756
rect 279344 320958 279372 326334
rect 279332 320952 279384 320958
rect 279332 320894 279384 320900
rect 279332 316736 279384 316742
rect 279332 316678 279384 316684
rect 278780 313948 278832 313954
rect 278780 313890 278832 313896
rect 278412 312724 278464 312730
rect 278412 312666 278464 312672
rect 278688 227792 278740 227798
rect 278686 227760 278688 227769
rect 278740 227760 278742 227769
rect 278686 227695 278742 227704
rect 278136 17264 278188 17270
rect 278136 17206 278188 17212
rect 278148 4049 278176 17206
rect 278134 4040 278190 4049
rect 278134 3975 278190 3984
rect 278042 3904 278098 3913
rect 278042 3839 278098 3848
rect 277858 3768 277914 3777
rect 277858 3703 277914 3712
rect 278792 626 278820 313890
rect 279344 307086 279372 316678
rect 279436 314022 279464 333254
rect 279528 326398 279556 335378
rect 279516 326392 279568 326398
rect 279516 326334 279568 326340
rect 279516 326256 279568 326262
rect 279516 326198 279568 326204
rect 279424 314016 279476 314022
rect 279424 313958 279476 313964
rect 279528 312662 279556 326198
rect 279516 312656 279568 312662
rect 279516 312598 279568 312604
rect 279332 307080 279384 307086
rect 279332 307022 279384 307028
rect 279620 286346 279648 335446
rect 279608 286340 279660 286346
rect 279608 286282 279660 286288
rect 279712 284986 279740 335566
rect 279804 326534 279832 340068
rect 279792 326528 279844 326534
rect 279792 326470 279844 326476
rect 279896 326380 279924 340068
rect 280080 337822 280108 340068
rect 280068 337816 280120 337822
rect 280068 337758 280120 337764
rect 280068 336864 280120 336870
rect 280068 336806 280120 336812
rect 279976 336796 280028 336802
rect 279976 336738 280028 336744
rect 279804 326352 279924 326380
rect 279804 316742 279832 326352
rect 279988 326210 280016 336738
rect 279896 326182 280016 326210
rect 279792 316736 279844 316742
rect 279792 316678 279844 316684
rect 279896 316554 279924 326182
rect 279976 326120 280028 326126
rect 279976 326062 280028 326068
rect 279804 316526 279924 316554
rect 279804 307170 279832 316526
rect 279804 307142 279924 307170
rect 279792 307080 279844 307086
rect 279792 307022 279844 307028
rect 279700 284980 279752 284986
rect 279700 284922 279752 284928
rect 279804 283626 279832 307022
rect 279792 283620 279844 283626
rect 279792 283562 279844 283568
rect 279896 8106 279924 307142
rect 279804 8078 279924 8106
rect 279988 8090 280016 326062
rect 279976 8084 280028 8090
rect 279804 3369 279832 8078
rect 279976 8026 280028 8032
rect 279976 7880 280028 7886
rect 279976 7822 280028 7828
rect 279884 6928 279936 6934
rect 279884 6870 279936 6876
rect 279896 3505 279924 6870
rect 279988 3641 280016 7822
rect 280080 6934 280108 336806
rect 280172 336802 280200 340068
rect 280160 336796 280212 336802
rect 280160 336738 280212 336744
rect 280264 335594 280292 340068
rect 280344 337612 280396 337618
rect 280344 337554 280396 337560
rect 280356 336666 280384 337554
rect 280448 337414 280476 340068
rect 280436 337408 280488 337414
rect 280436 337350 280488 337356
rect 280436 336796 280488 336802
rect 280436 336738 280488 336744
rect 280344 336660 280396 336666
rect 280344 336602 280396 336608
rect 280344 335708 280396 335714
rect 280344 335650 280396 335656
rect 280172 335566 280292 335594
rect 280172 282198 280200 335566
rect 280356 335458 280384 335650
rect 280264 335430 280384 335458
rect 280448 335458 280476 336738
rect 280540 335594 280568 340068
rect 280632 336870 280660 340068
rect 280712 338020 280764 338026
rect 280712 337962 280764 337968
rect 280724 337210 280752 337962
rect 280816 337929 280844 340068
rect 280802 337920 280858 337929
rect 280802 337855 280858 337864
rect 280804 337612 280856 337618
rect 280804 337554 280856 337560
rect 280712 337204 280764 337210
rect 280712 337146 280764 337152
rect 280712 337000 280764 337006
rect 280712 336942 280764 336948
rect 280620 336864 280672 336870
rect 280620 336806 280672 336812
rect 280724 335714 280752 336942
rect 280816 335714 280844 337554
rect 280712 335708 280764 335714
rect 280712 335650 280764 335656
rect 280804 335708 280856 335714
rect 280804 335650 280856 335656
rect 280540 335566 280844 335594
rect 280712 335504 280764 335510
rect 280448 335430 280660 335458
rect 280712 335446 280764 335452
rect 280264 326126 280292 335430
rect 280344 335368 280396 335374
rect 280344 335310 280396 335316
rect 280528 335368 280580 335374
rect 280528 335310 280580 335316
rect 280356 329322 280384 335310
rect 280344 329316 280396 329322
rect 280344 329258 280396 329264
rect 280252 326120 280304 326126
rect 280252 326062 280304 326068
rect 280540 318170 280568 335310
rect 280632 326210 280660 335430
rect 280724 326346 280752 335446
rect 280816 326482 280844 335566
rect 280908 335050 280936 340068
rect 281000 336802 281028 340068
rect 281184 338026 281212 340068
rect 281172 338020 281224 338026
rect 281172 337962 281224 337968
rect 281080 337340 281132 337346
rect 281080 337282 281132 337288
rect 280988 336796 281040 336802
rect 280988 336738 281040 336744
rect 281092 335170 281120 337282
rect 281172 337204 281224 337210
rect 281172 337146 281224 337152
rect 281080 335164 281132 335170
rect 281080 335106 281132 335112
rect 280908 335022 281028 335050
rect 280816 326454 280936 326482
rect 280724 326318 280844 326346
rect 280632 326182 280752 326210
rect 280724 319530 280752 326182
rect 280712 319524 280764 319530
rect 280712 319466 280764 319472
rect 280528 318164 280580 318170
rect 280528 318106 280580 318112
rect 280160 282192 280212 282198
rect 280160 282134 280212 282140
rect 280252 29096 280304 29102
rect 280250 29064 280252 29073
rect 280304 29064 280306 29073
rect 280250 28999 280306 29008
rect 280816 6934 280844 326318
rect 280908 311234 280936 326454
rect 280896 311228 280948 311234
rect 280896 311170 280948 311176
rect 281000 309874 281028 335022
rect 281184 332314 281212 337146
rect 281172 332308 281224 332314
rect 281172 332250 281224 332256
rect 281276 332194 281304 340068
rect 281368 337006 281396 340068
rect 281552 337210 281580 340068
rect 281540 337204 281592 337210
rect 281540 337146 281592 337152
rect 281356 337000 281408 337006
rect 281356 336942 281408 336948
rect 281356 336864 281408 336870
rect 281356 336806 281408 336812
rect 281092 332166 281304 332194
rect 280988 309868 281040 309874
rect 280988 309810 281040 309816
rect 281092 308514 281120 332166
rect 281368 326380 281396 336806
rect 281448 336796 281500 336802
rect 281448 336738 281500 336744
rect 281276 326352 281396 326380
rect 281080 308508 281132 308514
rect 281080 308450 281132 308456
rect 281276 280838 281304 326352
rect 281460 326210 281488 336738
rect 281644 331242 281672 340068
rect 281736 331362 281764 340068
rect 281920 337793 281948 340068
rect 281906 337784 281962 337793
rect 281906 337719 281962 337728
rect 281816 337068 281868 337074
rect 281816 337010 281868 337016
rect 281828 333418 281856 337010
rect 281908 336864 281960 336870
rect 281908 336806 281960 336812
rect 281920 333554 281948 336806
rect 282012 333690 282040 340068
rect 282104 337006 282132 340068
rect 282288 338094 282316 340068
rect 282276 338088 282328 338094
rect 282276 338030 282328 338036
rect 282380 337074 282408 340068
rect 282368 337068 282420 337074
rect 282368 337010 282420 337016
rect 282092 337000 282144 337006
rect 282092 336942 282144 336948
rect 282276 336932 282328 336938
rect 282276 336874 282328 336880
rect 282184 336796 282236 336802
rect 282184 336738 282236 336744
rect 282012 333662 282132 333690
rect 281920 333526 282040 333554
rect 281828 333390 281948 333418
rect 281724 331356 281776 331362
rect 281724 331298 281776 331304
rect 281644 331214 281856 331242
rect 281540 327752 281592 327758
rect 281540 327694 281592 327700
rect 281368 326182 281488 326210
rect 281264 280832 281316 280838
rect 281264 280774 281316 280780
rect 281368 279478 281396 326182
rect 281448 326120 281500 326126
rect 281448 326062 281500 326068
rect 281356 279472 281408 279478
rect 281356 279414 281408 279420
rect 281460 180130 281488 326062
rect 281448 180124 281500 180130
rect 281448 180066 281500 180072
rect 280068 6928 280120 6934
rect 280068 6870 280120 6876
rect 280804 6928 280856 6934
rect 280804 6870 280856 6876
rect 280068 5160 280120 5166
rect 280068 5102 280120 5108
rect 279974 3632 280030 3641
rect 279974 3567 280030 3576
rect 279882 3496 279938 3505
rect 279882 3431 279938 3440
rect 279790 3360 279846 3369
rect 279790 3295 279846 3304
rect 278792 598 278912 626
rect 278884 480 278912 598
rect 280080 480 280108 5102
rect 281264 5092 281316 5098
rect 281264 5034 281316 5040
rect 281276 480 281304 5034
rect 281552 610 281580 327694
rect 281828 325038 281856 331214
rect 281920 327826 281948 333390
rect 281908 327820 281960 327826
rect 281908 327762 281960 327768
rect 281816 325032 281868 325038
rect 281816 324974 281868 324980
rect 282012 276690 282040 333526
rect 282104 326398 282132 333662
rect 282092 326392 282144 326398
rect 282092 326334 282144 326340
rect 282196 307086 282224 336738
rect 282184 307080 282236 307086
rect 282184 307022 282236 307028
rect 282000 276684 282052 276690
rect 282000 276626 282052 276632
rect 282288 273970 282316 336874
rect 282472 336870 282500 340068
rect 282656 338065 282684 340068
rect 282642 338056 282698 338065
rect 282642 337991 282698 338000
rect 282644 337000 282696 337006
rect 282644 336942 282696 336948
rect 282460 336864 282512 336870
rect 282460 336806 282512 336812
rect 282368 326392 282420 326398
rect 282368 326334 282420 326340
rect 282380 318102 282408 326334
rect 282368 318096 282420 318102
rect 282368 318038 282420 318044
rect 282656 291854 282684 336942
rect 282748 336802 282776 340068
rect 282840 336938 282868 340068
rect 283024 337958 283052 340068
rect 283012 337952 283064 337958
rect 283012 337894 283064 337900
rect 283012 337544 283064 337550
rect 283012 337486 283064 337492
rect 282920 337204 282972 337210
rect 282920 337146 282972 337152
rect 282828 336932 282880 336938
rect 282828 336874 282880 336880
rect 282932 336870 282960 337146
rect 282920 336864 282972 336870
rect 282920 336806 282972 336812
rect 282736 336796 282788 336802
rect 282736 336738 282788 336744
rect 283024 336682 283052 337486
rect 283116 336802 283144 340068
rect 283104 336796 283156 336802
rect 283104 336738 283156 336744
rect 282932 336654 283052 336682
rect 282932 335374 282960 336654
rect 283208 335594 283236 340068
rect 283392 337210 283420 340068
rect 283288 337204 283340 337210
rect 283288 337146 283340 337152
rect 283380 337204 283432 337210
rect 283380 337146 283432 337152
rect 283300 337090 283328 337146
rect 283300 337062 283420 337090
rect 283288 336864 283340 336870
rect 283288 336806 283340 336812
rect 283024 335566 283236 335594
rect 282920 335368 282972 335374
rect 282920 335310 282972 335316
rect 282644 291848 282696 291854
rect 282644 291790 282696 291796
rect 282276 273964 282328 273970
rect 282276 273906 282328 273912
rect 283024 272542 283052 335566
rect 283300 335458 283328 336806
rect 283208 335430 283328 335458
rect 283012 272536 283064 272542
rect 283012 272478 283064 272484
rect 283208 269822 283236 335430
rect 283288 335368 283340 335374
rect 283288 335310 283340 335316
rect 283392 335322 283420 337062
rect 283484 335510 283512 340068
rect 283472 335504 283524 335510
rect 283472 335446 283524 335452
rect 283576 335442 283604 340068
rect 283760 337550 283788 340068
rect 283748 337544 283800 337550
rect 283748 337486 283800 337492
rect 283656 336796 283708 336802
rect 283656 336738 283708 336744
rect 283564 335436 283616 335442
rect 283564 335378 283616 335384
rect 283300 327962 283328 335310
rect 283392 335294 283604 335322
rect 283472 335232 283524 335238
rect 283472 335174 283524 335180
rect 283288 327956 283340 327962
rect 283288 327898 283340 327904
rect 283484 315382 283512 335174
rect 283472 315376 283524 315382
rect 283472 315318 283524 315324
rect 283196 269816 283248 269822
rect 283196 269758 283248 269764
rect 283576 4962 283604 335294
rect 283668 316742 283696 336738
rect 283656 316736 283708 316742
rect 283656 316678 283708 316684
rect 283852 304298 283880 340068
rect 283944 336870 283972 340068
rect 284128 337890 284156 340068
rect 284116 337884 284168 337890
rect 284116 337826 284168 337832
rect 284116 337544 284168 337550
rect 284116 337486 284168 337492
rect 284024 337204 284076 337210
rect 284024 337146 284076 337152
rect 283932 336864 283984 336870
rect 283932 336806 283984 336812
rect 284036 335714 284064 337146
rect 284128 336122 284156 337486
rect 284116 336116 284168 336122
rect 284116 336058 284168 336064
rect 284024 335708 284076 335714
rect 284024 335650 284076 335656
rect 284220 335594 284248 340068
rect 284312 336802 284340 340068
rect 284496 337686 284524 340068
rect 284484 337680 284536 337686
rect 284484 337622 284536 337628
rect 284392 337204 284444 337210
rect 284392 337146 284444 337152
rect 284300 336796 284352 336802
rect 284300 336738 284352 336744
rect 283944 335566 284248 335594
rect 283840 304292 283892 304298
rect 283840 304234 283892 304240
rect 283944 302938 283972 335566
rect 284024 335504 284076 335510
rect 284024 335446 284076 335452
rect 284208 335504 284260 335510
rect 284208 335446 284260 335452
rect 284036 305658 284064 335446
rect 284116 335436 284168 335442
rect 284116 335378 284168 335384
rect 284024 305652 284076 305658
rect 284024 305594 284076 305600
rect 283932 302932 283984 302938
rect 283932 302874 283984 302880
rect 284128 271182 284156 335378
rect 284220 333334 284248 335446
rect 284208 333328 284260 333334
rect 284208 333270 284260 333276
rect 284404 326330 284432 337146
rect 284484 337068 284536 337074
rect 284484 337010 284536 337016
rect 284392 326324 284444 326330
rect 284392 326266 284444 326272
rect 284496 300150 284524 337010
rect 284588 336870 284616 340068
rect 284694 340054 284800 340082
rect 284576 336864 284628 336870
rect 284576 336806 284628 336812
rect 284772 326482 284800 340054
rect 284864 337618 284892 340068
rect 284852 337612 284904 337618
rect 284852 337554 284904 337560
rect 284956 336802 284984 340068
rect 284944 336796 284996 336802
rect 284944 336738 284996 336744
rect 284944 331152 284996 331158
rect 284944 331094 284996 331100
rect 284680 326454 284800 326482
rect 284484 300144 284536 300150
rect 284484 300086 284536 300092
rect 284680 298110 284708 326454
rect 284760 326392 284812 326398
rect 284760 326334 284812 326340
rect 284668 298104 284720 298110
rect 284668 298046 284720 298052
rect 284576 288448 284628 288454
rect 284576 288390 284628 288396
rect 284588 282962 284616 288390
rect 284496 282934 284616 282962
rect 284496 282826 284524 282934
rect 284496 282798 284616 282826
rect 284588 273306 284616 282798
rect 284588 273278 284708 273306
rect 284116 271176 284168 271182
rect 284116 271118 284168 271124
rect 284680 267034 284708 273278
rect 284668 267028 284720 267034
rect 284668 266970 284720 266976
rect 284772 265674 284800 326334
rect 284852 326324 284904 326330
rect 284852 326266 284904 326272
rect 284760 265668 284812 265674
rect 284760 265610 284812 265616
rect 284864 182850 284892 326266
rect 284956 278050 284984 331094
rect 285048 326398 285076 340068
rect 285232 336977 285260 340068
rect 285324 337074 285352 340068
rect 285416 337210 285444 340068
rect 285496 337612 285548 337618
rect 285496 337554 285548 337560
rect 285404 337204 285456 337210
rect 285404 337146 285456 337152
rect 285312 337068 285364 337074
rect 285312 337010 285364 337016
rect 285218 336968 285274 336977
rect 285218 336903 285274 336912
rect 285128 336864 285180 336870
rect 285128 336806 285180 336812
rect 285404 336864 285456 336870
rect 285404 336806 285456 336812
rect 285036 326392 285088 326398
rect 285036 326334 285088 326340
rect 285140 301510 285168 336806
rect 285220 336796 285272 336802
rect 285220 336738 285272 336744
rect 285232 315314 285260 336738
rect 285312 336728 285364 336734
rect 285312 336670 285364 336676
rect 285220 315308 285272 315314
rect 285220 315250 285272 315256
rect 285128 301504 285180 301510
rect 285128 301446 285180 301452
rect 284944 278044 284996 278050
rect 284944 277986 284996 277992
rect 285324 268394 285352 336670
rect 285416 331974 285444 336806
rect 285508 334694 285536 337554
rect 285600 337074 285628 340068
rect 285588 337068 285640 337074
rect 285588 337010 285640 337016
rect 285586 336968 285642 336977
rect 285586 336903 285642 336912
rect 285496 334688 285548 334694
rect 285496 334630 285548 334636
rect 285404 331968 285456 331974
rect 285404 331910 285456 331916
rect 285600 330546 285628 336903
rect 285588 330540 285640 330546
rect 285588 330482 285640 330488
rect 285692 323678 285720 340068
rect 285680 323672 285732 323678
rect 285680 323614 285732 323620
rect 285680 315512 285732 315518
rect 285680 315454 285732 315460
rect 285312 268388 285364 268394
rect 285312 268330 285364 268336
rect 284852 182844 284904 182850
rect 284852 182786 284904 182792
rect 284760 5024 284812 5030
rect 284760 4966 284812 4972
rect 283564 4956 283616 4962
rect 283564 4898 283616 4904
rect 283656 4888 283708 4894
rect 283656 4830 283708 4836
rect 281540 604 281592 610
rect 281540 546 281592 552
rect 282460 604 282512 610
rect 282460 546 282512 552
rect 282472 480 282500 546
rect 283668 480 283696 4830
rect 284772 480 284800 4966
rect 285692 610 285720 315454
rect 285784 290494 285812 340068
rect 285968 337414 285996 340068
rect 285956 337408 286008 337414
rect 285956 337350 286008 337356
rect 286060 335714 286088 340068
rect 286048 335708 286100 335714
rect 286048 335650 286100 335656
rect 286152 335594 286180 340068
rect 286336 337074 286364 340068
rect 286324 337068 286376 337074
rect 286324 337010 286376 337016
rect 286232 336864 286284 336870
rect 286232 336806 286284 336812
rect 285968 335566 286180 335594
rect 285772 290488 285824 290494
rect 285772 290430 285824 290436
rect 285968 262886 285996 335566
rect 286244 335458 286272 336806
rect 286324 335708 286376 335714
rect 286324 335650 286376 335656
rect 286060 335430 286272 335458
rect 285956 262880 286008 262886
rect 285956 262822 286008 262828
rect 286060 261526 286088 335430
rect 286140 335368 286192 335374
rect 286140 335310 286192 335316
rect 286048 261520 286100 261526
rect 286048 261462 286100 261468
rect 286152 260166 286180 335310
rect 286336 332874 286364 335650
rect 286428 333010 286456 340068
rect 286520 336870 286548 340068
rect 286508 336864 286560 336870
rect 286508 336806 286560 336812
rect 286428 332982 286640 333010
rect 286336 332846 286456 332874
rect 286428 313954 286456 332846
rect 286416 313948 286468 313954
rect 286416 313890 286468 313896
rect 286612 297498 286640 332982
rect 286704 327758 286732 340068
rect 286692 327752 286744 327758
rect 286692 327694 286744 327700
rect 286796 312594 286824 340068
rect 286888 335374 286916 340068
rect 287072 338026 287100 340068
rect 287060 338020 287112 338026
rect 287060 337962 287112 337968
rect 286968 337068 287020 337074
rect 286968 337010 287020 337016
rect 286876 335368 286928 335374
rect 286876 335310 286928 335316
rect 286980 333266 287008 337010
rect 287060 334620 287112 334626
rect 287060 334562 287112 334568
rect 286968 333260 287020 333266
rect 286968 333202 287020 333208
rect 286784 312588 286836 312594
rect 286784 312530 286836 312536
rect 286600 297492 286652 297498
rect 286600 297434 286652 297440
rect 286140 260160 286192 260166
rect 286140 260102 286192 260108
rect 287072 4214 287100 334562
rect 287164 331158 287192 340068
rect 287256 336954 287284 340068
rect 287440 337210 287468 340068
rect 287428 337204 287480 337210
rect 287428 337146 287480 337152
rect 287256 336926 287468 336954
rect 287336 336864 287388 336870
rect 287336 336806 287388 336812
rect 287244 336796 287296 336802
rect 287244 336738 287296 336744
rect 287152 331152 287204 331158
rect 287152 331094 287204 331100
rect 287256 258738 287284 336738
rect 287244 258732 287296 258738
rect 287244 258674 287296 258680
rect 287348 257378 287376 336806
rect 287440 331294 287468 336926
rect 287532 332738 287560 340068
rect 287624 336802 287652 340068
rect 287704 337816 287756 337822
rect 287702 337784 287704 337793
rect 287756 337784 287758 337793
rect 287702 337719 287758 337728
rect 287808 337686 287836 340068
rect 287796 337680 287848 337686
rect 287796 337622 287848 337628
rect 287796 337204 287848 337210
rect 287796 337146 287848 337152
rect 287612 336796 287664 336802
rect 287612 336738 287664 336744
rect 287808 336054 287836 337146
rect 287796 336048 287848 336054
rect 287796 335990 287848 335996
rect 287532 332710 287836 332738
rect 287428 331288 287480 331294
rect 287428 331230 287480 331236
rect 287704 331152 287756 331158
rect 287704 331094 287756 331100
rect 287428 326392 287480 326398
rect 287428 326334 287480 326340
rect 287440 309806 287468 326334
rect 287612 326324 287664 326330
rect 287612 326266 287664 326272
rect 287428 309800 287480 309806
rect 287428 309742 287480 309748
rect 287336 257372 287388 257378
rect 287336 257314 287388 257320
rect 287624 28286 287652 326266
rect 287716 319462 287744 331094
rect 287808 326398 287836 332710
rect 287796 326392 287848 326398
rect 287796 326334 287848 326340
rect 287704 319456 287756 319462
rect 287704 319398 287756 319404
rect 287900 296002 287928 340068
rect 287992 336870 288020 340068
rect 288070 338056 288126 338065
rect 288070 337991 288126 338000
rect 288084 337890 288112 337991
rect 288072 337884 288124 337890
rect 288072 337826 288124 337832
rect 287980 336864 288032 336870
rect 287980 336806 288032 336812
rect 287980 331220 288032 331226
rect 287980 331162 288032 331168
rect 287992 324850 288020 331162
rect 288176 324970 288204 340068
rect 288164 324964 288216 324970
rect 288164 324906 288216 324912
rect 287992 324822 288204 324850
rect 287980 322924 288032 322930
rect 287980 322866 288032 322872
rect 287888 295996 287940 296002
rect 287888 295938 287940 295944
rect 287992 294642 288020 322866
rect 288176 313970 288204 324822
rect 288268 322930 288296 340068
rect 288360 326330 288388 340068
rect 288544 337006 288572 340068
rect 288532 337000 288584 337006
rect 288532 336942 288584 336948
rect 288636 335510 288664 340068
rect 288624 335504 288676 335510
rect 288624 335446 288676 335452
rect 288624 329588 288676 329594
rect 288624 329530 288676 329536
rect 288348 326324 288400 326330
rect 288348 326266 288400 326272
rect 288256 322924 288308 322930
rect 288256 322866 288308 322872
rect 288176 313942 288388 313970
rect 288360 298110 288388 313942
rect 288636 308446 288664 329530
rect 288624 308440 288676 308446
rect 288624 308382 288676 308388
rect 288348 298104 288400 298110
rect 288348 298046 288400 298052
rect 288728 297430 288756 340068
rect 288912 336870 288940 340068
rect 289004 336938 289032 340068
rect 288992 336932 289044 336938
rect 288992 336874 289044 336880
rect 288900 336864 288952 336870
rect 288900 336806 288952 336812
rect 289096 321706 289124 340068
rect 289280 337142 289308 340068
rect 289268 337136 289320 337142
rect 289268 337078 289320 337084
rect 289372 335714 289400 340068
rect 289360 335708 289412 335714
rect 289360 335650 289412 335656
rect 289464 335594 289492 340068
rect 289542 337920 289598 337929
rect 289542 337855 289598 337864
rect 289556 337754 289584 337855
rect 289544 337748 289596 337754
rect 289544 337690 289596 337696
rect 289544 337136 289596 337142
rect 289544 337078 289596 337084
rect 289188 335566 289492 335594
rect 289188 323610 289216 335566
rect 289268 335504 289320 335510
rect 289268 335446 289320 335452
rect 289176 323604 289228 323610
rect 289176 323546 289228 323552
rect 289280 322250 289308 335446
rect 289556 331906 289584 337078
rect 289648 334626 289676 340068
rect 289636 334620 289688 334626
rect 289636 334562 289688 334568
rect 289544 331900 289596 331906
rect 289544 331842 289596 331848
rect 289740 328522 289768 340068
rect 289832 337929 289860 340068
rect 289818 337920 289874 337929
rect 289818 337855 289874 337864
rect 290464 337272 290516 337278
rect 290464 337214 290516 337220
rect 289648 328494 289768 328522
rect 289648 323490 289676 328494
rect 289464 323462 289676 323490
rect 289268 322244 289320 322250
rect 289268 322186 289320 322192
rect 289084 321700 289136 321706
rect 289084 321642 289136 321648
rect 288992 321564 289044 321570
rect 288992 321506 289044 321512
rect 288716 297424 288768 297430
rect 288716 297366 288768 297372
rect 289004 296070 289032 321506
rect 289268 318844 289320 318850
rect 289268 318786 289320 318792
rect 289280 298110 289308 318786
rect 289464 311166 289492 323462
rect 289452 311160 289504 311166
rect 289452 311102 289504 311108
rect 289268 298104 289320 298110
rect 289268 298046 289320 298052
rect 288992 296064 289044 296070
rect 288992 296006 289044 296012
rect 287980 294636 288032 294642
rect 287980 294578 288032 294584
rect 289084 288448 289136 288454
rect 289084 288390 289136 288396
rect 289096 282962 289124 288390
rect 288912 282934 289124 282962
rect 288912 264246 288940 282934
rect 288900 264240 288952 264246
rect 288900 264182 288952 264188
rect 289728 227792 289780 227798
rect 289726 227760 289728 227769
rect 289780 227760 289782 227769
rect 289726 227695 289782 227704
rect 289728 29096 289780 29102
rect 289726 29064 289728 29073
rect 289780 29064 289782 29073
rect 289726 28999 289782 29008
rect 287612 28280 287664 28286
rect 287612 28222 287664 28228
rect 290476 15910 290504 337214
rect 290568 322930 290596 400182
rect 290648 399900 290700 399906
rect 290648 399842 290700 399848
rect 290660 393310 290688 399842
rect 291936 399696 291988 399702
rect 291936 399638 291988 399644
rect 291844 398880 291896 398886
rect 291844 398822 291896 398828
rect 290648 393304 290700 393310
rect 290648 393246 290700 393252
rect 291856 369850 291884 398822
rect 291844 369844 291896 369850
rect 291844 369786 291896 369792
rect 291200 338088 291252 338094
rect 291200 338030 291252 338036
rect 290832 337952 290884 337958
rect 290832 337894 290884 337900
rect 291106 337920 291162 337929
rect 290740 337000 290792 337006
rect 290740 336942 290792 336948
rect 290648 336864 290700 336870
rect 290648 336806 290700 336812
rect 290556 322924 290608 322930
rect 290556 322866 290608 322872
rect 290660 320890 290688 336806
rect 290752 323610 290780 336942
rect 290844 326398 290872 337894
rect 291106 337855 291162 337864
rect 290832 326392 290884 326398
rect 290832 326334 290884 326340
rect 290740 323604 290792 323610
rect 290740 323546 290792 323552
rect 290648 320884 290700 320890
rect 290648 320826 290700 320832
rect 291120 256018 291148 337855
rect 291212 336190 291240 338030
rect 291844 337204 291896 337210
rect 291844 337146 291896 337152
rect 291200 336184 291252 336190
rect 291200 336126 291252 336132
rect 291108 256012 291160 256018
rect 291108 255954 291160 255960
rect 290464 15904 290516 15910
rect 290464 15846 290516 15852
rect 291856 13122 291884 337146
rect 291948 111790 291976 399638
rect 292028 336932 292080 336938
rect 292028 336874 292080 336880
rect 292040 293282 292068 336874
rect 293960 336660 294012 336666
rect 293960 336602 294012 336608
rect 292580 335096 292632 335102
rect 292580 335038 292632 335044
rect 292028 293276 292080 293282
rect 292028 293218 292080 293224
rect 291936 111784 291988 111790
rect 291936 111726 291988 111732
rect 291844 13116 291896 13122
rect 291844 13058 291896 13064
rect 291936 9308 291988 9314
rect 291936 9250 291988 9256
rect 289544 6928 289596 6934
rect 289544 6870 289596 6876
rect 287152 4752 287204 4758
rect 287152 4694 287204 4700
rect 287060 4208 287112 4214
rect 287060 4150 287112 4156
rect 285680 604 285732 610
rect 285680 546 285732 552
rect 285956 604 286008 610
rect 285956 546 286008 552
rect 285968 480 285996 546
rect 287164 480 287192 4694
rect 288348 4208 288400 4214
rect 288348 4150 288400 4156
rect 288360 480 288388 4150
rect 289556 480 289584 6870
rect 290740 4820 290792 4826
rect 290740 4762 290792 4768
rect 290752 480 290780 4762
rect 291948 480 291976 9250
rect 292592 3482 292620 335038
rect 293972 3482 294000 336602
rect 294616 64870 294644 400862
rect 297364 338020 297416 338026
rect 297364 337962 297416 337968
rect 294696 336728 294748 336734
rect 294696 336670 294748 336676
rect 294604 64864 294656 64870
rect 294604 64806 294656 64812
rect 294708 19990 294736 336670
rect 296720 336592 296772 336598
rect 296720 336534 296772 336540
rect 294696 19984 294748 19990
rect 294696 19926 294748 19932
rect 295524 9240 295576 9246
rect 295524 9182 295576 9188
rect 292592 3454 293172 3482
rect 293972 3454 294368 3482
rect 293144 480 293172 3454
rect 294340 480 294368 3454
rect 295536 480 295564 9182
rect 296732 4214 296760 336534
rect 296812 332376 296864 332382
rect 296812 332318 296864 332324
rect 296720 4208 296772 4214
rect 296720 4150 296772 4156
rect 296824 1442 296852 332318
rect 297376 18630 297404 337962
rect 297468 158710 297496 400930
rect 301596 400852 301648 400858
rect 301596 400794 301648 400800
rect 298836 399628 298888 399634
rect 298836 399570 298888 399576
rect 298744 337884 298796 337890
rect 298744 337826 298796 337832
rect 297456 158704 297508 158710
rect 297456 158646 297508 158652
rect 297364 18624 297416 18630
rect 297364 18566 297416 18572
rect 298756 14482 298784 337826
rect 298848 205630 298876 399570
rect 301504 337816 301556 337822
rect 301504 337758 301556 337764
rect 300860 335980 300912 335986
rect 300860 335922 300912 335928
rect 299480 328160 299532 328166
rect 299480 328102 299532 328108
rect 298836 205624 298888 205630
rect 298836 205566 298888 205572
rect 298744 14476 298796 14482
rect 298744 14418 298796 14424
rect 299112 9172 299164 9178
rect 299112 9114 299164 9120
rect 297916 4208 297968 4214
rect 297916 4150 297968 4156
rect 296732 1414 296852 1442
rect 296732 480 296760 1414
rect 297928 480 297956 4150
rect 299124 480 299152 9114
rect 299492 610 299520 328102
rect 300872 610 300900 335922
rect 301516 11762 301544 337758
rect 301608 252550 301636 400794
rect 304264 400512 304316 400518
rect 304264 400454 304316 400460
rect 302976 399492 303028 399498
rect 302976 399434 303028 399440
rect 302884 337884 302936 337890
rect 302884 337826 302936 337832
rect 301596 252544 301648 252550
rect 301596 252486 301648 252492
rect 302146 227896 302202 227905
rect 302146 227831 302202 227840
rect 302160 227497 302188 227831
rect 302146 227488 302202 227497
rect 302146 227423 302202 227432
rect 302146 76120 302202 76129
rect 302146 76055 302202 76064
rect 302160 75721 302188 76055
rect 302146 75712 302202 75721
rect 302146 75647 302202 75656
rect 301504 11756 301556 11762
rect 301504 11698 301556 11704
rect 302896 8974 302924 337826
rect 302988 299470 303016 399434
rect 303620 325304 303672 325310
rect 303620 325246 303672 325252
rect 302976 299464 303028 299470
rect 302976 299406 303028 299412
rect 302608 8968 302660 8974
rect 302608 8910 302660 8916
rect 302884 8968 302936 8974
rect 302884 8910 302936 8916
rect 299480 604 299532 610
rect 299480 546 299532 552
rect 300308 604 300360 610
rect 300308 546 300360 552
rect 300860 604 300912 610
rect 300860 546 300912 552
rect 301412 604 301464 610
rect 301412 546 301464 552
rect 300320 480 300348 546
rect 301424 480 301452 546
rect 302620 480 302648 8910
rect 303632 610 303660 325246
rect 304276 41410 304304 400454
rect 308404 400444 308456 400450
rect 308404 400386 308456 400392
rect 305644 399288 305696 399294
rect 305644 399230 305696 399236
rect 305000 335164 305052 335170
rect 305000 335106 305052 335112
rect 304264 41404 304316 41410
rect 304264 41346 304316 41352
rect 303620 604 303672 610
rect 303620 546 303672 552
rect 303804 604 303856 610
rect 303804 546 303856 552
rect 303816 480 303844 546
rect 305012 480 305040 335106
rect 305656 88330 305684 399230
rect 307758 333806 307814 333815
rect 307758 333741 307814 333750
rect 307758 333568 307814 333577
rect 307758 333503 307814 333512
rect 306380 319728 306432 319734
rect 306380 319670 306432 319676
rect 305644 88324 305696 88330
rect 305644 88266 305696 88272
rect 306196 9104 306248 9110
rect 306196 9046 306248 9052
rect 306208 480 306236 9046
rect 306392 3482 306420 319670
rect 307772 3482 307800 333503
rect 308416 182170 308444 400386
rect 413284 400308 413336 400314
rect 413284 400250 413336 400256
rect 312544 399084 312596 399090
rect 312544 399026 312596 399032
rect 309782 398576 309838 398585
rect 309782 398511 309838 398520
rect 309796 276010 309824 398511
rect 311900 335028 311952 335034
rect 311900 334970 311952 334976
rect 310520 311364 310572 311370
rect 310520 311306 310572 311312
rect 309784 276004 309836 276010
rect 309784 275946 309836 275952
rect 309140 227792 309192 227798
rect 309138 227760 309140 227769
rect 309192 227760 309194 227769
rect 309138 227695 309194 227704
rect 308404 182164 308456 182170
rect 308404 182106 308456 182112
rect 309140 76016 309192 76022
rect 309138 75984 309140 75993
rect 309192 75984 309194 75993
rect 309138 75919 309194 75928
rect 309784 9036 309836 9042
rect 309784 8978 309836 8984
rect 306392 3454 307432 3482
rect 307772 3454 308628 3482
rect 307404 480 307432 3454
rect 308600 480 308628 3454
rect 309796 480 309824 8978
rect 310532 3482 310560 311306
rect 311912 3482 311940 334970
rect 312556 124166 312584 399026
rect 319444 399016 319496 399022
rect 319444 398958 319496 398964
rect 316684 337612 316736 337618
rect 316684 337554 316736 337560
rect 315304 337544 315356 337550
rect 315304 337486 315356 337492
rect 314660 336456 314712 336462
rect 314660 336398 314712 336404
rect 313280 330880 313332 330886
rect 313280 330822 313332 330828
rect 312634 227896 312690 227905
rect 312634 227831 312690 227840
rect 312648 227798 312676 227831
rect 312636 227792 312688 227798
rect 312636 227734 312688 227740
rect 312544 124160 312596 124166
rect 312544 124102 312596 124108
rect 313292 3482 313320 330822
rect 313372 323944 313424 323950
rect 313372 323886 313424 323892
rect 313384 4214 313412 323886
rect 313922 76120 313978 76129
rect 313922 76055 313978 76064
rect 313936 76022 313964 76055
rect 313924 76016 313976 76022
rect 313924 75958 313976 75964
rect 313372 4208 313424 4214
rect 313372 4150 313424 4156
rect 314568 4208 314620 4214
rect 314568 4150 314620 4156
rect 310532 3454 311020 3482
rect 311912 3454 312216 3482
rect 313292 3454 313412 3482
rect 310992 480 311020 3454
rect 312188 480 312216 3454
rect 313384 480 313412 3454
rect 314580 480 314608 4150
rect 314672 3618 314700 336398
rect 315316 4826 315344 337486
rect 316040 333668 316092 333674
rect 316040 333610 316092 333616
rect 315304 4820 315356 4826
rect 315304 4762 315356 4768
rect 314672 3590 315804 3618
rect 315776 480 315804 3590
rect 316052 3482 316080 333610
rect 316696 7614 316724 337554
rect 318800 332308 318852 332314
rect 318800 332250 318852 332256
rect 317420 310004 317472 310010
rect 317420 309946 317472 309952
rect 316684 7608 316736 7614
rect 316684 7550 316736 7556
rect 317432 3482 317460 309946
rect 318812 3482 318840 332250
rect 319456 135250 319484 398958
rect 326342 398440 326398 398449
rect 326342 398375 326398 398384
rect 326356 358766 326384 398375
rect 326344 358760 326396 358766
rect 326344 358702 326396 358708
rect 320824 337680 320876 337686
rect 320824 337622 320876 337628
rect 320180 326732 320232 326738
rect 320180 326674 320232 326680
rect 319444 135244 319496 135250
rect 319444 135186 319496 135192
rect 320192 3482 320220 326674
rect 320836 21418 320864 337622
rect 346400 337476 346452 337482
rect 346400 337418 346452 337424
rect 331220 336388 331272 336394
rect 331220 336330 331272 336336
rect 327080 334960 327132 334966
rect 327080 334902 327132 334908
rect 322940 329452 322992 329458
rect 322940 329394 322992 329400
rect 321560 322448 321612 322454
rect 321560 322390 321612 322396
rect 320824 21412 320876 21418
rect 320824 21354 320876 21360
rect 321572 3482 321600 322390
rect 322848 5568 322900 5574
rect 322848 5510 322900 5516
rect 316052 3454 317000 3482
rect 317432 3454 318104 3482
rect 318812 3454 319300 3482
rect 320192 3454 320496 3482
rect 321572 3454 321692 3482
rect 316972 480 317000 3454
rect 318076 480 318104 3454
rect 319272 480 319300 3454
rect 320468 480 320496 3454
rect 321664 480 321692 3454
rect 322860 480 322888 5510
rect 322952 3482 322980 329394
rect 324320 293344 324372 293350
rect 324320 293286 324372 293292
rect 323582 227896 323638 227905
rect 323582 227831 323638 227840
rect 323596 227633 323624 227831
rect 323582 227624 323638 227633
rect 323582 227559 323638 227568
rect 323582 76120 323638 76129
rect 323582 76055 323638 76064
rect 323596 75857 323624 76055
rect 323582 75848 323638 75857
rect 323582 75783 323638 75792
rect 324332 3482 324360 293286
rect 326436 5636 326488 5642
rect 326436 5578 326488 5584
rect 322952 3454 324084 3482
rect 324332 3454 325280 3482
rect 324056 480 324084 3454
rect 325252 480 325280 3454
rect 326448 480 326476 5578
rect 327092 3482 327120 334902
rect 328460 328092 328512 328098
rect 328460 328034 328512 328040
rect 328472 228138 328500 328034
rect 328460 228132 328512 228138
rect 328460 228074 328512 228080
rect 328458 228032 328514 228041
rect 328514 227990 328592 228018
rect 328458 227967 328514 227976
rect 328460 227928 328512 227934
rect 328460 227870 328512 227876
rect 328472 76362 328500 227870
rect 328564 227633 328592 227990
rect 328550 227624 328606 227633
rect 328550 227559 328606 227568
rect 328460 76356 328512 76362
rect 328460 76298 328512 76304
rect 328458 76256 328514 76265
rect 328514 76214 328592 76242
rect 328458 76191 328514 76200
rect 328460 76152 328512 76158
rect 328460 76094 328512 76100
rect 328472 3482 328500 76094
rect 328564 75857 328592 76214
rect 328550 75848 328606 75857
rect 328550 75783 328606 75792
rect 330024 5704 330076 5710
rect 330024 5646 330076 5652
rect 327092 3454 327672 3482
rect 328472 3454 328868 3482
rect 327644 480 327672 3454
rect 328840 480 328868 3454
rect 330036 480 330064 5646
rect 331232 480 331260 336330
rect 338120 333600 338172 333606
rect 338120 333542 338172 333548
rect 333980 332240 334032 332246
rect 333980 332182 334032 332188
rect 333612 5772 333664 5778
rect 333612 5714 333664 5720
rect 332416 4888 332468 4894
rect 332416 4830 332468 4836
rect 332428 480 332456 4830
rect 333624 480 333652 5714
rect 333992 3482 334020 332182
rect 335360 318300 335412 318306
rect 335360 318242 335412 318248
rect 335372 3482 335400 318242
rect 337108 5840 337160 5846
rect 337108 5782 337160 5788
rect 333992 3454 334756 3482
rect 335372 3454 335952 3482
rect 334728 480 334756 3454
rect 335924 480 335952 3454
rect 337120 480 337148 5782
rect 338132 3482 338160 333542
rect 342260 329384 342312 329390
rect 342260 329326 342312 329332
rect 339500 308576 339552 308582
rect 339500 308518 339552 308524
rect 338132 3454 338344 3482
rect 338316 480 338344 3454
rect 339512 480 339540 308518
rect 340880 10056 340932 10062
rect 340880 9998 340932 10004
rect 340696 5908 340748 5914
rect 340696 5850 340748 5856
rect 340708 480 340736 5850
rect 340892 3482 340920 9998
rect 342272 3482 342300 329326
rect 345020 10124 345072 10130
rect 345020 10066 345072 10072
rect 344284 5976 344336 5982
rect 344284 5918 344336 5924
rect 340892 3454 341932 3482
rect 342272 3454 343128 3482
rect 341904 480 341932 3454
rect 343100 480 343128 3454
rect 344296 480 344324 5918
rect 345032 3482 345060 10066
rect 346412 3482 346440 337418
rect 349160 336320 349212 336326
rect 349160 336262 349212 336268
rect 347780 326800 347832 326806
rect 347780 326742 347832 326748
rect 347792 326466 347820 326742
rect 347780 326460 347832 326466
rect 347780 326402 347832 326408
rect 347780 10192 347832 10198
rect 347780 10134 347832 10140
rect 347792 4214 347820 10134
rect 347872 6044 347924 6050
rect 347872 5986 347924 5992
rect 347780 4208 347832 4214
rect 347780 4150 347832 4156
rect 345032 3454 345520 3482
rect 346412 3454 346716 3482
rect 345492 480 345520 3454
rect 346688 480 346716 3454
rect 347884 480 347912 5986
rect 349068 4208 349120 4214
rect 349068 4150 349120 4156
rect 349080 480 349108 4150
rect 349172 3482 349200 336262
rect 353300 334892 353352 334898
rect 353300 334834 353352 334840
rect 351920 10260 351972 10266
rect 351920 10202 351972 10208
rect 351368 6112 351420 6118
rect 351368 6054 351420 6060
rect 349172 3454 350304 3482
rect 350276 480 350304 3454
rect 351380 480 351408 6054
rect 351932 3482 351960 10202
rect 351932 3454 352604 3482
rect 352576 480 352604 3454
rect 353312 1306 353340 334834
rect 374000 333532 374052 333538
rect 374000 333474 374052 333480
rect 356060 332172 356112 332178
rect 356060 332114 356112 332120
rect 354956 6860 355008 6866
rect 354956 6802 355008 6808
rect 353312 1278 353800 1306
rect 353772 480 353800 1278
rect 354968 480 354996 6802
rect 356072 4214 356100 332114
rect 360200 326664 360252 326670
rect 360200 326606 360252 326612
rect 356152 11008 356204 11014
rect 356152 10950 356204 10956
rect 356060 4208 356112 4214
rect 356060 4150 356112 4156
rect 356164 480 356192 10950
rect 358820 10940 358872 10946
rect 358820 10882 358872 10888
rect 358544 6792 358596 6798
rect 358544 6734 358596 6740
rect 357348 4208 357400 4214
rect 357348 4150 357400 4156
rect 357360 480 357388 4150
rect 358556 480 358584 6734
rect 358832 3482 358860 10882
rect 360212 3482 360240 326606
rect 367100 325236 367152 325242
rect 367100 325178 367152 325184
rect 364340 319660 364392 319666
rect 364340 319602 364392 319608
rect 362960 10872 363012 10878
rect 362960 10814 363012 10820
rect 362132 6724 362184 6730
rect 362132 6666 362184 6672
rect 358832 3454 359780 3482
rect 360212 3454 360976 3482
rect 359752 480 359780 3454
rect 360948 480 360976 3454
rect 362144 480 362172 6666
rect 362972 3482 363000 10814
rect 364352 3482 364380 319602
rect 365720 10804 365772 10810
rect 365720 10746 365772 10752
rect 365732 4214 365760 10746
rect 365812 6656 365864 6662
rect 365812 6598 365864 6604
rect 365720 4208 365772 4214
rect 365720 4150 365772 4156
rect 362972 3454 363368 3482
rect 364352 3454 364564 3482
rect 363340 480 363368 3454
rect 364536 480 364564 3454
rect 365824 3346 365852 6598
rect 366916 4208 366968 4214
rect 366916 4150 366968 4156
rect 365732 3318 365852 3346
rect 365732 480 365760 3318
rect 366928 480 366956 4150
rect 367112 3482 367140 325178
rect 371240 316940 371292 316946
rect 371240 316882 371292 316888
rect 369860 10736 369912 10742
rect 369860 10678 369912 10684
rect 369216 6588 369268 6594
rect 369216 6530 369268 6536
rect 367112 3454 368060 3482
rect 368032 480 368060 3454
rect 369228 480 369256 6530
rect 369872 3482 369900 10678
rect 371252 3482 371280 316882
rect 372804 6520 372856 6526
rect 372804 6462 372856 6468
rect 369872 3454 370452 3482
rect 371252 3454 371648 3482
rect 370424 480 370452 3454
rect 371620 480 371648 3454
rect 372816 480 372844 6462
rect 374012 4214 374040 333474
rect 400312 333464 400364 333470
rect 400312 333406 400364 333412
rect 393320 330812 393372 330818
rect 393320 330754 393372 330760
rect 382280 328024 382332 328030
rect 382280 327966 382332 327972
rect 378140 311296 378192 311302
rect 378140 311238 378192 311244
rect 374092 10668 374144 10674
rect 374092 10610 374144 10616
rect 374000 4208 374052 4214
rect 374000 4150 374052 4156
rect 374104 1442 374132 10610
rect 376760 10600 376812 10606
rect 376760 10542 376812 10548
rect 376392 6452 376444 6458
rect 376392 6394 376444 6400
rect 375196 4208 375248 4214
rect 375196 4150 375248 4156
rect 374012 1414 374132 1442
rect 374012 480 374040 1414
rect 375208 480 375236 4150
rect 376404 480 376432 6394
rect 376772 3482 376800 10542
rect 378152 3482 378180 311238
rect 380900 10532 380952 10538
rect 380900 10474 380952 10480
rect 379980 6384 380032 6390
rect 379980 6326 380032 6332
rect 376772 3454 377628 3482
rect 378152 3454 378824 3482
rect 377600 480 377628 3454
rect 378796 480 378824 3454
rect 379992 480 380020 6326
rect 380912 3482 380940 10474
rect 382292 3482 382320 327966
rect 385040 323876 385092 323882
rect 385040 323818 385092 323824
rect 383660 10464 383712 10470
rect 383660 10406 383712 10412
rect 383568 6316 383620 6322
rect 383568 6258 383620 6264
rect 380912 3454 381216 3482
rect 382292 3454 382412 3482
rect 381188 480 381216 3454
rect 382384 480 382412 3454
rect 383580 480 383608 6258
rect 383672 3482 383700 10406
rect 385052 3482 385080 323818
rect 389180 309936 389232 309942
rect 389180 309878 389232 309884
rect 387800 10396 387852 10402
rect 387800 10338 387852 10344
rect 387064 6248 387116 6254
rect 387064 6190 387116 6196
rect 383672 3454 384712 3482
rect 385052 3454 385908 3482
rect 384684 480 384712 3454
rect 385880 480 385908 3454
rect 387076 480 387104 6190
rect 387812 3482 387840 10338
rect 389192 3482 389220 309878
rect 390560 10328 390612 10334
rect 390560 10270 390612 10276
rect 387812 3454 388300 3482
rect 389192 3454 389496 3482
rect 388272 480 388300 3454
rect 389468 480 389496 3454
rect 390572 2854 390600 10270
rect 390652 6180 390704 6186
rect 390652 6122 390704 6128
rect 390560 2848 390612 2854
rect 390560 2790 390612 2796
rect 390664 480 390692 6122
rect 393332 3482 393360 330754
rect 397460 329316 397512 329322
rect 397460 329258 397512 329264
rect 394700 321088 394752 321094
rect 394700 321030 394752 321036
rect 394712 3482 394740 321030
rect 397472 3482 397500 329258
rect 398840 325168 398892 325174
rect 398840 325110 398892 325116
rect 398104 29300 398156 29306
rect 398104 29242 398156 29248
rect 398116 29209 398144 29242
rect 398102 29200 398158 29209
rect 398102 29135 398158 29144
rect 398852 3482 398880 325110
rect 400324 3482 400352 333406
rect 404360 332104 404412 332110
rect 404360 332046 404412 332052
rect 401600 318232 401652 318238
rect 401600 318174 401652 318180
rect 401612 3482 401640 318174
rect 404372 3482 404400 332046
rect 411260 330744 411312 330750
rect 411260 330686 411312 330692
rect 408500 327956 408552 327962
rect 408500 327898 408552 327904
rect 405740 307148 405792 307154
rect 405740 307090 405792 307096
rect 405646 29336 405702 29345
rect 405646 29271 405648 29280
rect 405700 29271 405702 29280
rect 405648 29242 405700 29248
rect 405752 3482 405780 307090
rect 393332 3454 394280 3482
rect 394712 3454 395476 3482
rect 397472 3454 397868 3482
rect 398852 3454 399064 3482
rect 400324 3454 401364 3482
rect 401612 3454 402560 3482
rect 404372 3454 404952 3482
rect 405752 3454 406148 3482
rect 391848 2848 391900 2854
rect 391848 2790 391900 2796
rect 393044 2848 393096 2854
rect 393044 2790 393096 2796
rect 391860 480 391888 2790
rect 393056 480 393084 2790
rect 394252 480 394280 3454
rect 395448 480 395476 3454
rect 396632 2916 396684 2922
rect 396632 2858 396684 2864
rect 396644 480 396672 2858
rect 397840 480 397868 3454
rect 399036 480 399064 3454
rect 400220 2984 400272 2990
rect 400220 2926 400272 2932
rect 400232 480 400260 2926
rect 401336 480 401364 3454
rect 402532 480 402560 3454
rect 403716 3052 403768 3058
rect 403716 2994 403768 3000
rect 403728 480 403756 2994
rect 404924 480 404952 3454
rect 406120 480 406148 3454
rect 407304 3120 407356 3126
rect 407304 3062 407356 3068
rect 407316 480 407344 3062
rect 408512 480 408540 327898
rect 408592 316872 408644 316878
rect 408592 316814 408644 316820
rect 408604 3482 408632 316814
rect 411272 3482 411300 330686
rect 412640 305720 412692 305726
rect 412640 305662 412692 305668
rect 412652 3482 412680 305662
rect 413296 218006 413324 400250
rect 489184 336728 489236 336734
rect 489184 336670 489236 336676
rect 443092 336252 443144 336258
rect 443092 336194 443144 336200
rect 422300 334824 422352 334830
rect 422300 334766 422352 334772
rect 415400 326596 415452 326602
rect 415400 326538 415452 326544
rect 413284 218000 413336 218006
rect 413284 217942 413336 217948
rect 415306 76120 415362 76129
rect 415306 76055 415362 76064
rect 415320 75993 415348 76055
rect 415306 75984 415362 75993
rect 415306 75919 415362 75928
rect 415412 3482 415440 326538
rect 418160 325100 418212 325106
rect 418160 325042 418212 325048
rect 416872 291916 416924 291922
rect 416872 291858 416924 291864
rect 408604 3454 409736 3482
rect 411272 3454 412128 3482
rect 412652 3454 413324 3482
rect 415412 3454 415716 3482
rect 409708 480 409736 3454
rect 410892 3188 410944 3194
rect 410892 3130 410944 3136
rect 410904 480 410932 3130
rect 412100 480 412128 3454
rect 413296 480 413324 3454
rect 414480 3256 414532 3262
rect 414480 3198 414532 3204
rect 414492 480 414520 3198
rect 415688 480 415716 3454
rect 416884 480 416912 291858
rect 418066 228032 418122 228041
rect 418066 227967 418068 227976
rect 418120 227967 418122 227976
rect 418068 227938 418120 227944
rect 417332 29232 417384 29238
rect 417330 29200 417332 29209
rect 417384 29200 417386 29209
rect 417330 29135 417386 29144
rect 418172 3482 418200 325042
rect 419540 304360 419592 304366
rect 419540 304302 419592 304308
rect 419552 3482 419580 304302
rect 422312 3482 422340 334766
rect 440240 333396 440292 333402
rect 440240 333338 440292 333344
rect 425152 329248 425204 329254
rect 425152 329190 425204 329196
rect 423680 315444 423732 315450
rect 423680 315386 423732 315392
rect 423692 3482 423720 315386
rect 424966 228032 425022 228041
rect 424966 227967 424968 227976
rect 425020 227967 425022 227976
rect 424968 227938 425020 227944
rect 424966 29336 425022 29345
rect 424966 29271 425022 29280
rect 424980 29238 425008 29271
rect 424968 29232 425020 29238
rect 424968 29174 425020 29180
rect 425060 4140 425112 4146
rect 425060 4082 425112 4088
rect 418172 3454 419212 3482
rect 419552 3454 420408 3482
rect 422312 3454 422800 3482
rect 423692 3454 423996 3482
rect 417976 3324 418028 3330
rect 417976 3266 418028 3272
rect 417988 480 418016 3266
rect 419184 480 419212 3454
rect 420380 480 420408 3454
rect 421564 3392 421616 3398
rect 421564 3334 421616 3340
rect 421576 480 421604 3334
rect 422772 480 422800 3454
rect 423968 480 423996 3454
rect 425072 2802 425100 4082
rect 425164 2922 425192 329190
rect 429200 327888 429252 327894
rect 429200 327830 429252 327836
rect 426440 303000 426492 303006
rect 426440 302942 426492 302948
rect 426452 3482 426480 302942
rect 428740 4072 428792 4078
rect 428740 4014 428792 4020
rect 426452 3454 427584 3482
rect 425152 2916 425204 2922
rect 425152 2858 425204 2864
rect 426348 2916 426400 2922
rect 426348 2858 426400 2864
rect 425072 2774 425192 2802
rect 425164 480 425192 2774
rect 426360 480 426388 2858
rect 427556 480 427584 3454
rect 428752 480 428780 4014
rect 429212 3482 429240 327830
rect 433340 326528 433392 326534
rect 433340 326470 433392 326476
rect 430580 290556 430632 290562
rect 430580 290498 430632 290504
rect 430592 3482 430620 290498
rect 432328 4004 432380 4010
rect 432328 3946 432380 3952
rect 429212 3454 429976 3482
rect 430592 3454 431172 3482
rect 429948 480 429976 3454
rect 431144 480 431172 3454
rect 432340 480 432368 3946
rect 433352 3398 433380 326470
rect 436100 323808 436152 323814
rect 436100 323750 436152 323756
rect 433432 319592 433484 319598
rect 433432 319534 433484 319540
rect 433444 3482 433472 319534
rect 435824 3936 435876 3942
rect 435824 3878 435876 3884
rect 433444 3454 433564 3482
rect 433340 3392 433392 3398
rect 433340 3334 433392 3340
rect 433536 480 433564 3454
rect 434628 3392 434680 3398
rect 434628 3334 434680 3340
rect 434640 480 434668 3334
rect 435836 480 435864 3878
rect 436112 3482 436140 323750
rect 437480 323740 437532 323746
rect 437480 323682 437532 323688
rect 437386 227896 437442 227905
rect 437386 227831 437388 227840
rect 437440 227831 437442 227840
rect 437388 227802 437440 227808
rect 437386 76120 437442 76129
rect 437386 76055 437388 76064
rect 437440 76055 437442 76064
rect 437388 76026 437440 76032
rect 436744 29300 436796 29306
rect 436744 29242 436796 29248
rect 436756 29209 436784 29242
rect 436742 29200 436798 29209
rect 436742 29135 436798 29144
rect 437492 3482 437520 323682
rect 439412 3868 439464 3874
rect 439412 3810 439464 3816
rect 436112 3454 437060 3482
rect 437492 3454 438256 3482
rect 437032 480 437060 3454
rect 438228 480 438256 3454
rect 439424 480 439452 3810
rect 440252 3482 440280 333338
rect 441620 314084 441672 314090
rect 441620 314026 441672 314032
rect 441632 3482 441660 314026
rect 443000 3800 443052 3806
rect 443000 3742 443052 3748
rect 440252 3454 440648 3482
rect 441632 3454 441844 3482
rect 440620 480 440648 3454
rect 441816 480 441844 3454
rect 443012 480 443040 3742
rect 443104 3482 443132 336194
rect 483020 336184 483072 336190
rect 483020 336126 483072 336132
rect 467840 332036 467892 332042
rect 467840 331978 467892 331984
rect 451280 330676 451332 330682
rect 451280 330618 451332 330624
rect 448520 321020 448572 321026
rect 448520 320962 448572 320968
rect 447140 318164 447192 318170
rect 447140 318106 447192 318112
rect 444380 301572 444432 301578
rect 444380 301514 444432 301520
rect 444288 227860 444340 227866
rect 444288 227802 444340 227808
rect 444300 227769 444328 227802
rect 444286 227760 444342 227769
rect 444286 227695 444342 227704
rect 444288 76084 444340 76090
rect 444288 76026 444340 76032
rect 444300 75993 444328 76026
rect 444286 75984 444342 75993
rect 444286 75919 444342 75928
rect 444286 29336 444342 29345
rect 444286 29271 444288 29280
rect 444340 29271 444342 29280
rect 444288 29242 444340 29248
rect 444392 3482 444420 301514
rect 446588 3732 446640 3738
rect 446588 3674 446640 3680
rect 443104 3454 444236 3482
rect 444392 3454 445432 3482
rect 444208 480 444236 3454
rect 445404 480 445432 3454
rect 446600 480 446628 3674
rect 447152 3482 447180 318106
rect 448532 3482 448560 320962
rect 450176 3664 450228 3670
rect 450176 3606 450228 3612
rect 447152 3454 447824 3482
rect 448532 3454 449020 3482
rect 447796 480 447824 3454
rect 448992 480 449020 3454
rect 450188 480 450216 3606
rect 451292 480 451320 330618
rect 462320 330608 462372 330614
rect 462320 330550 462372 330556
rect 454040 322380 454092 322386
rect 454040 322322 454092 322328
rect 451372 289196 451424 289202
rect 451372 289138 451424 289144
rect 451384 3482 451412 289138
rect 453672 3596 453724 3602
rect 453672 3538 453724 3544
rect 451384 3454 452516 3482
rect 452488 480 452516 3454
rect 453684 480 453712 3538
rect 454052 3482 454080 322322
rect 458180 316804 458232 316810
rect 458180 316746 458232 316752
rect 455420 300212 455472 300218
rect 455420 300154 455472 300160
rect 455432 3482 455460 300154
rect 456706 227896 456762 227905
rect 456890 227896 456946 227905
rect 456762 227854 456890 227882
rect 456706 227831 456762 227840
rect 456890 227831 456946 227840
rect 456706 76120 456762 76129
rect 456890 76120 456946 76129
rect 456762 76078 456890 76106
rect 456706 76055 456762 76064
rect 456890 76055 456946 76064
rect 456708 29232 456760 29238
rect 456706 29200 456708 29209
rect 456760 29200 456762 29209
rect 456706 29135 456762 29144
rect 457260 3528 457312 3534
rect 454052 3454 454908 3482
rect 455432 3454 456104 3482
rect 457260 3470 457312 3476
rect 458192 3482 458220 316746
rect 460940 315376 460992 315382
rect 460940 315318 460992 315324
rect 459652 287700 459704 287706
rect 459652 287642 459704 287648
rect 454880 480 454908 3454
rect 456076 480 456104 3454
rect 457272 480 457300 3470
rect 458192 3454 458496 3482
rect 458468 480 458496 3454
rect 459664 480 459692 287642
rect 460952 3482 460980 315318
rect 462332 3482 462360 330550
rect 465080 326460 465132 326466
rect 465080 326402 465132 326408
rect 463606 29336 463662 29345
rect 463606 29271 463662 29280
rect 463620 29238 463648 29271
rect 463608 29232 463660 29238
rect 463608 29174 463660 29180
rect 464434 4040 464490 4049
rect 464434 3975 464490 3984
rect 460848 3460 460900 3466
rect 460952 3454 462084 3482
rect 462332 3454 463280 3482
rect 460848 3402 460900 3408
rect 460860 480 460888 3402
rect 462056 480 462084 3454
rect 463252 480 463280 3454
rect 464448 480 464476 3975
rect 465092 3482 465120 326402
rect 466460 312724 466512 312730
rect 466460 312666 466512 312672
rect 466472 3482 466500 312666
rect 467852 3534 467880 331978
rect 471980 329180 472032 329186
rect 471980 329122 472032 329128
rect 469220 322312 469272 322318
rect 469220 322254 469272 322260
rect 467930 3904 467986 3913
rect 467930 3839 467986 3848
rect 467840 3528 467892 3534
rect 465092 3454 465672 3482
rect 466472 3454 466868 3482
rect 467840 3470 467892 3476
rect 465644 480 465672 3454
rect 466840 480 466868 3454
rect 467944 480 467972 3839
rect 469128 3528 469180 3534
rect 469128 3470 469180 3476
rect 469232 3482 469260 322254
rect 471244 256012 471296 256018
rect 471244 255954 471296 255960
rect 469140 480 469168 3470
rect 469232 3454 470364 3482
rect 471256 3466 471284 255954
rect 471518 3768 471574 3777
rect 471518 3703 471574 3712
rect 470336 480 470364 3454
rect 471244 3460 471296 3466
rect 471244 3402 471296 3408
rect 471532 480 471560 3703
rect 471992 3346 472020 329122
rect 476120 320952 476172 320958
rect 476120 320894 476172 320900
rect 473360 298784 473412 298790
rect 473360 298726 473412 298732
rect 473372 3346 473400 298726
rect 475384 264240 475436 264246
rect 475384 264182 475436 264188
rect 475292 29232 475344 29238
rect 475290 29200 475292 29209
rect 475344 29200 475346 29209
rect 475290 29135 475346 29144
rect 475106 3632 475162 3641
rect 475106 3567 475162 3576
rect 471992 3318 472756 3346
rect 473372 3318 473952 3346
rect 472728 480 472756 3318
rect 473924 480 473952 3318
rect 475120 480 475148 3567
rect 475396 3534 475424 264182
rect 476026 227896 476082 227905
rect 476026 227831 476028 227840
rect 476080 227831 476082 227840
rect 476028 227802 476080 227808
rect 475384 3528 475436 3534
rect 475384 3470 475436 3476
rect 476132 3346 476160 320894
rect 478880 314016 478932 314022
rect 478880 313958 478932 313964
rect 477500 286340 477552 286346
rect 477500 286282 477552 286288
rect 476132 3318 476344 3346
rect 476316 480 476344 3318
rect 477512 480 477540 286282
rect 478694 3496 478750 3505
rect 478694 3431 478750 3440
rect 478708 480 478736 3431
rect 478892 3346 478920 313958
rect 482284 296064 482336 296070
rect 482284 296006 482336 296012
rect 480260 284980 480312 284986
rect 480260 284922 480312 284928
rect 480272 3482 480300 284922
rect 482296 3602 482324 296006
rect 482928 227860 482980 227866
rect 482928 227802 482980 227808
rect 482940 227769 482968 227802
rect 482926 227760 482982 227769
rect 482926 227695 482982 227704
rect 482926 76120 482982 76129
rect 482926 76055 482982 76064
rect 482940 75993 482968 76055
rect 482926 75984 482982 75993
rect 482926 75919 482982 75928
rect 482926 29336 482982 29345
rect 482926 29271 482982 29280
rect 482940 29238 482968 29271
rect 482928 29232 482980 29238
rect 482928 29174 482980 29180
rect 482284 3596 482336 3602
rect 482284 3538 482336 3544
rect 483032 3482 483060 336126
rect 487160 319524 487212 319530
rect 487160 319466 487212 319472
rect 484400 312656 484452 312662
rect 484400 312598 484452 312604
rect 484412 3482 484440 312598
rect 485780 283620 485832 283626
rect 485780 283562 485832 283568
rect 480272 3454 481128 3482
rect 483032 3454 483520 3482
rect 484412 3454 484624 3482
rect 478892 3318 479932 3346
rect 479904 480 479932 3318
rect 481100 480 481128 3454
rect 482282 3360 482338 3369
rect 482282 3295 482338 3304
rect 482296 480 482324 3295
rect 483492 480 483520 3454
rect 484596 480 484624 3454
rect 485792 480 485820 283562
rect 486976 4820 487028 4826
rect 486976 4762 487028 4768
rect 486988 480 487016 4762
rect 487172 3482 487200 319466
rect 488540 282192 488592 282198
rect 488540 282134 488592 282140
rect 488552 3618 488580 282134
rect 489196 4826 489224 336670
rect 491300 311228 491352 311234
rect 491300 311170 491352 311176
rect 490564 7608 490616 7614
rect 490564 7550 490616 7556
rect 489184 4820 489236 4826
rect 489184 4762 489236 4768
rect 488552 3590 489408 3618
rect 487172 3454 488212 3482
rect 488184 480 488212 3454
rect 489380 480 489408 3590
rect 490576 480 490604 7550
rect 491312 626 491340 311170
rect 492680 280832 492732 280838
rect 492680 280774 492732 280780
rect 491312 598 491800 626
rect 492692 610 492720 280774
rect 493336 171086 493364 401950
rect 500224 401940 500276 401946
rect 500224 401882 500276 401888
rect 498844 401872 498896 401878
rect 498844 401814 498896 401820
rect 494060 309868 494112 309874
rect 494060 309810 494112 309816
rect 493324 171080 493376 171086
rect 493324 171022 493376 171028
rect 494072 3398 494100 309810
rect 498200 308508 498252 308514
rect 498200 308450 498252 308456
rect 495440 279472 495492 279478
rect 495440 279414 495492 279420
rect 495348 227928 495400 227934
rect 495346 227896 495348 227905
rect 495400 227896 495402 227905
rect 495346 227831 495402 227840
rect 495164 29232 495216 29238
rect 495162 29200 495164 29209
rect 495216 29200 495218 29209
rect 495162 29135 495218 29144
rect 494152 8968 494204 8974
rect 494152 8910 494204 8916
rect 494060 3392 494112 3398
rect 494060 3334 494112 3340
rect 491772 480 491800 598
rect 492680 604 492732 610
rect 492680 546 492732 552
rect 492956 604 493008 610
rect 492956 546 493008 552
rect 492968 480 492996 546
rect 494164 480 494192 8910
rect 495348 3392 495400 3398
rect 495348 3334 495400 3340
rect 495360 480 495388 3334
rect 495452 610 495480 279414
rect 497004 227928 497056 227934
rect 497002 227896 497004 227905
rect 497056 227896 497058 227905
rect 497002 227831 497058 227840
rect 497740 4820 497792 4826
rect 497740 4762 497792 4768
rect 495440 604 495492 610
rect 495440 546 495492 552
rect 496544 604 496596 610
rect 496544 546 496596 552
rect 496556 480 496584 546
rect 497752 480 497780 4762
rect 498212 610 498240 308450
rect 498856 264926 498884 401814
rect 500236 311846 500264 401882
rect 579804 393304 579856 393310
rect 579804 393246 579856 393252
rect 579816 393009 579844 393246
rect 579802 393000 579858 393009
rect 579802 392935 579858 392944
rect 580172 369844 580224 369850
rect 580172 369786 580224 369792
rect 580184 369617 580212 369786
rect 580170 369608 580226 369617
rect 580170 369543 580226 369552
rect 580080 358760 580132 358766
rect 580080 358702 580132 358708
rect 580092 357921 580120 358702
rect 580078 357912 580134 357921
rect 580078 357847 580134 357856
rect 579804 346384 579856 346390
rect 579804 346326 579856 346332
rect 579816 346089 579844 346326
rect 579802 346080 579858 346089
rect 579802 346015 579858 346024
rect 521660 336116 521712 336122
rect 521660 336058 521712 336064
rect 500960 334756 501012 334762
rect 500960 334698 501012 334704
rect 500224 311840 500276 311846
rect 500224 311782 500276 311788
rect 498844 264920 498896 264926
rect 498844 264862 498896 264868
rect 499580 180124 499632 180130
rect 499580 180066 499632 180072
rect 499592 3482 499620 180066
rect 500972 3482 501000 334698
rect 518900 333328 518952 333334
rect 518900 333270 518952 333276
rect 509240 327820 509292 327826
rect 509240 327762 509292 327768
rect 502340 325032 502392 325038
rect 502340 324974 502392 324980
rect 502248 76084 502300 76090
rect 502248 76026 502300 76032
rect 502260 75857 502288 76026
rect 502246 75848 502302 75857
rect 502246 75783 502302 75792
rect 502246 29336 502302 29345
rect 502246 29271 502302 29280
rect 502260 29238 502288 29271
rect 502248 29232 502300 29238
rect 502248 29174 502300 29180
rect 502352 3482 502380 324974
rect 505100 318096 505152 318102
rect 505100 318038 505152 318044
rect 502432 278044 502484 278050
rect 502432 277986 502484 277992
rect 502444 3670 502472 277986
rect 503720 11756 503772 11762
rect 503720 11698 503772 11704
rect 502432 3664 502484 3670
rect 502432 3606 502484 3612
rect 503628 3664 503680 3670
rect 503628 3606 503680 3612
rect 499592 3454 500172 3482
rect 500972 3454 501276 3482
rect 502352 3454 502472 3482
rect 498200 604 498252 610
rect 498200 546 498252 552
rect 498936 604 498988 610
rect 498936 546 498988 552
rect 498948 480 498976 546
rect 500144 480 500172 3454
rect 501248 480 501276 3454
rect 502444 480 502472 3454
rect 503640 480 503668 3606
rect 503732 3482 503760 11698
rect 505112 3482 505140 318038
rect 506480 291848 506532 291854
rect 506480 291790 506532 291796
rect 506492 3482 506520 291790
rect 507860 13116 507912 13122
rect 507860 13058 507912 13064
rect 507872 3482 507900 13058
rect 509252 3482 509280 327762
rect 516140 316736 516192 316742
rect 516140 316678 516192 316684
rect 512000 307080 512052 307086
rect 512000 307022 512052 307028
rect 510620 276684 510672 276690
rect 510620 276626 510672 276632
rect 510526 76256 510582 76265
rect 510526 76191 510582 76200
rect 510540 76090 510568 76191
rect 510528 76084 510580 76090
rect 510528 76026 510580 76032
rect 510632 3482 510660 276626
rect 503732 3454 504864 3482
rect 505112 3454 506060 3482
rect 506492 3454 507256 3482
rect 507872 3454 508452 3482
rect 509252 3454 509648 3482
rect 510632 3454 510844 3482
rect 504836 480 504864 3454
rect 506032 480 506060 3454
rect 507228 480 507256 3454
rect 508424 480 508452 3454
rect 509620 480 509648 3454
rect 510816 480 510844 3454
rect 512012 3398 512040 307022
rect 513380 273964 513432 273970
rect 513380 273906 513432 273912
rect 512092 14476 512144 14482
rect 512092 14418 512144 14424
rect 512000 3392 512052 3398
rect 512000 3334 512052 3340
rect 512104 1442 512132 14418
rect 513392 3482 513420 273906
rect 514666 227896 514722 227905
rect 514666 227831 514668 227840
rect 514720 227831 514722 227840
rect 514668 227802 514720 227808
rect 513564 29232 513616 29238
rect 513562 29200 513564 29209
rect 513616 29200 513618 29209
rect 513562 29135 513618 29144
rect 514760 15904 514812 15910
rect 514760 15846 514812 15852
rect 514772 3482 514800 15846
rect 516152 3482 516180 316678
rect 517520 272536 517572 272542
rect 517520 272478 517572 272484
rect 517532 3482 517560 272478
rect 518912 3482 518940 333270
rect 520280 305652 520332 305658
rect 520280 305594 520332 305600
rect 513392 3454 514432 3482
rect 514772 3454 515628 3482
rect 516152 3454 516824 3482
rect 517532 3454 517928 3482
rect 518912 3454 519124 3482
rect 513196 3392 513248 3398
rect 513196 3334 513248 3340
rect 512012 1414 512132 1442
rect 512012 480 512040 1414
rect 513208 480 513236 3334
rect 514404 480 514432 3454
rect 515600 480 515628 3454
rect 516796 480 516824 3454
rect 517900 480 517928 3454
rect 519096 480 519124 3454
rect 520292 480 520320 305594
rect 520372 271176 520424 271182
rect 520372 271118 520424 271124
rect 520384 3482 520412 271118
rect 521568 227860 521620 227866
rect 521568 227802 521620 227808
rect 521580 227769 521608 227802
rect 521566 227760 521622 227769
rect 521566 227695 521622 227704
rect 521566 76528 521622 76537
rect 521566 76463 521622 76472
rect 521580 75993 521608 76463
rect 521566 75984 521622 75993
rect 521566 75919 521622 75928
rect 521566 29336 521622 29345
rect 521566 29271 521622 29280
rect 521580 29238 521608 29271
rect 521568 29232 521620 29238
rect 521568 29174 521620 29180
rect 521672 3482 521700 336058
rect 557540 336048 557592 336054
rect 557540 335990 557592 335996
rect 532700 334688 532752 334694
rect 532700 334630 532752 334636
rect 528560 331968 528612 331974
rect 528560 331910 528612 331916
rect 523040 304292 523092 304298
rect 523040 304234 523092 304240
rect 523052 3482 523080 304234
rect 527180 302932 527232 302938
rect 527180 302874 527232 302880
rect 524420 269816 524472 269822
rect 524420 269758 524472 269764
rect 524432 3482 524460 269758
rect 525800 18624 525852 18630
rect 525800 18566 525852 18572
rect 525812 3482 525840 18566
rect 527192 3482 527220 302874
rect 520384 3454 521516 3482
rect 521672 3454 522712 3482
rect 523052 3454 523908 3482
rect 524432 3454 525104 3482
rect 525812 3454 526300 3482
rect 527192 3454 527496 3482
rect 521488 480 521516 3454
rect 522684 480 522712 3454
rect 523880 480 523908 3454
rect 525076 480 525104 3454
rect 526272 480 526300 3454
rect 527468 480 527496 3454
rect 528572 3398 528600 331910
rect 529940 301504 529992 301510
rect 529940 301446 529992 301452
rect 528652 268388 528704 268394
rect 528652 268330 528704 268336
rect 528560 3392 528612 3398
rect 528560 3334 528612 3340
rect 528664 480 528692 268330
rect 529952 3482 529980 301446
rect 531320 267028 531372 267034
rect 531320 266970 531372 266976
rect 531332 3482 531360 266970
rect 532712 3482 532740 334630
rect 546500 333260 546552 333266
rect 546500 333202 546552 333208
rect 536840 330540 536892 330546
rect 536840 330482 536892 330488
rect 534080 315308 534132 315314
rect 534080 315250 534132 315256
rect 533986 227896 534042 227905
rect 533986 227831 534042 227840
rect 534000 227798 534028 227831
rect 533988 227792 534040 227798
rect 533988 227734 534040 227740
rect 533986 76120 534042 76129
rect 533986 76055 533988 76064
rect 534040 76055 534042 76064
rect 533988 76026 534040 76032
rect 533804 29232 533856 29238
rect 533802 29200 533804 29209
rect 533856 29200 533858 29209
rect 533802 29135 533858 29144
rect 534092 3482 534120 315250
rect 535460 265668 535512 265674
rect 535460 265610 535512 265616
rect 535472 3482 535500 265610
rect 536852 3482 536880 330482
rect 539600 329112 539652 329118
rect 539600 329054 539652 329060
rect 536932 300144 536984 300150
rect 536932 300086 536984 300092
rect 536944 3670 536972 300086
rect 538220 182844 538272 182850
rect 538220 182786 538272 182792
rect 536932 3664 536984 3670
rect 536932 3606 536984 3612
rect 538128 3664 538180 3670
rect 538128 3606 538180 3612
rect 529952 3454 531084 3482
rect 531332 3454 532280 3482
rect 532712 3454 533476 3482
rect 534092 3454 534580 3482
rect 535472 3454 535776 3482
rect 536852 3454 536972 3482
rect 529848 3392 529900 3398
rect 529848 3334 529900 3340
rect 529860 480 529888 3334
rect 531056 480 531084 3454
rect 532252 480 532280 3454
rect 533448 480 533476 3454
rect 534552 480 534580 3454
rect 535748 480 535776 3454
rect 536944 480 536972 3454
rect 538140 480 538168 3606
rect 538232 3482 538260 182786
rect 539612 3482 539640 329054
rect 540980 323672 541032 323678
rect 540980 323614 541032 323620
rect 540888 227792 540940 227798
rect 540886 227760 540888 227769
rect 540940 227760 540942 227769
rect 540886 227695 540942 227704
rect 540888 76084 540940 76090
rect 540888 76026 540940 76032
rect 540900 75993 540928 76026
rect 540886 75984 540942 75993
rect 540886 75919 540942 75928
rect 540886 29336 540942 29345
rect 540886 29271 540942 29280
rect 540900 29238 540928 29271
rect 540888 29232 540940 29238
rect 540888 29174 540940 29180
rect 540992 3482 541020 323614
rect 545120 313948 545172 313954
rect 545120 313890 545172 313896
rect 542360 290488 542412 290494
rect 542360 290430 542412 290436
rect 542372 3482 542400 290430
rect 543740 19984 543792 19990
rect 543740 19926 543792 19932
rect 543752 3482 543780 19926
rect 545132 3482 545160 313890
rect 546512 3670 546540 333202
rect 550640 327752 550692 327758
rect 550640 327694 550692 327700
rect 547880 297492 547932 297498
rect 547880 297434 547932 297440
rect 546592 262880 546644 262886
rect 546592 262822 546644 262828
rect 546500 3664 546552 3670
rect 546500 3606 546552 3612
rect 546604 3482 546632 262822
rect 547696 3664 547748 3670
rect 547696 3606 547748 3612
rect 538232 3454 539364 3482
rect 539612 3454 540560 3482
rect 540992 3454 541756 3482
rect 542372 3454 542952 3482
rect 543752 3454 544148 3482
rect 545132 3454 545344 3482
rect 539336 480 539364 3454
rect 540532 480 540560 3454
rect 541728 480 541756 3454
rect 542924 480 542952 3454
rect 544120 480 544148 3454
rect 545316 480 545344 3454
rect 546512 3454 546632 3482
rect 546512 480 546540 3454
rect 547708 480 547736 3606
rect 547892 3482 547920 297434
rect 549260 261520 549312 261526
rect 549260 261462 549312 261468
rect 549272 3482 549300 261462
rect 550652 3482 550680 327694
rect 554780 326392 554832 326398
rect 554780 326334 554832 326340
rect 552020 312588 552072 312594
rect 552020 312530 552072 312536
rect 552032 3482 552060 312530
rect 553400 260160 553452 260166
rect 553400 260102 553452 260108
rect 553308 227928 553360 227934
rect 553306 227896 553308 227905
rect 553360 227896 553362 227905
rect 553306 227831 553362 227840
rect 553308 76152 553360 76158
rect 553306 76120 553308 76129
rect 553360 76120 553362 76129
rect 553306 76055 553362 76064
rect 552480 29232 552532 29238
rect 552478 29200 552480 29209
rect 552532 29200 552534 29209
rect 552478 29135 552534 29144
rect 553412 3482 553440 260102
rect 554596 227928 554648 227934
rect 554594 227896 554596 227905
rect 554648 227896 554650 227905
rect 554594 227831 554650 227840
rect 554596 76152 554648 76158
rect 554594 76120 554596 76129
rect 554648 76120 554650 76129
rect 554594 76055 554650 76064
rect 547892 3454 548932 3482
rect 549272 3454 550128 3482
rect 550652 3454 551232 3482
rect 552032 3454 552428 3482
rect 553412 3454 553624 3482
rect 548904 480 548932 3454
rect 550100 480 550128 3454
rect 551204 480 551232 3454
rect 552400 480 552428 3454
rect 553596 480 553624 3454
rect 554792 480 554820 326334
rect 554872 319456 554924 319462
rect 554872 319398 554924 319404
rect 554884 3482 554912 319398
rect 556804 309800 556856 309806
rect 556804 309742 556856 309748
rect 556160 289128 556212 289134
rect 556160 289070 556212 289076
rect 556172 3618 556200 289070
rect 556816 4146 556844 309742
rect 556804 4140 556856 4146
rect 556804 4082 556856 4088
rect 556172 3590 557212 3618
rect 554884 3454 556016 3482
rect 555988 480 556016 3454
rect 557184 480 557212 3590
rect 557552 3482 557580 335990
rect 573364 334620 573416 334626
rect 573364 334562 573416 334568
rect 564440 324964 564492 324970
rect 564440 324906 564492 324912
rect 563060 295996 563112 296002
rect 563060 295938 563112 295944
rect 560944 294636 560996 294642
rect 560944 294578 560996 294584
rect 560300 258732 560352 258738
rect 560300 258674 560352 258680
rect 560206 29336 560262 29345
rect 560206 29271 560262 29280
rect 560220 29238 560248 29271
rect 560208 29232 560260 29238
rect 560208 29174 560260 29180
rect 559564 4140 559616 4146
rect 559564 4082 559616 4088
rect 557552 3454 558408 3482
rect 558380 480 558408 3454
rect 559576 480 559604 4082
rect 560312 3482 560340 258674
rect 560312 3454 560800 3482
rect 560772 480 560800 3454
rect 560956 3058 560984 294578
rect 561680 21412 561732 21418
rect 561680 21354 561732 21360
rect 561692 3482 561720 21354
rect 563072 3482 563100 295938
rect 563152 257372 563204 257378
rect 563152 257314 563204 257320
rect 563164 3670 563192 257314
rect 563152 3664 563204 3670
rect 563152 3606 563204 3612
rect 564348 3664 564400 3670
rect 564348 3606 564400 3612
rect 561692 3454 561996 3482
rect 563072 3454 563192 3482
rect 560944 3052 560996 3058
rect 560944 2994 560996 3000
rect 561968 480 561996 3454
rect 563164 480 563192 3454
rect 564360 480 564388 3606
rect 564452 3482 564480 324906
rect 568580 323604 568632 323610
rect 568580 323546 568632 323552
rect 567844 322244 567896 322250
rect 567844 322186 567896 322192
rect 567200 28280 567252 28286
rect 567200 28222 567252 28228
rect 564452 3454 565584 3482
rect 565556 480 565584 3454
rect 567212 3346 567240 28222
rect 567856 3602 567884 322186
rect 567844 3596 567896 3602
rect 567844 3538 567896 3544
rect 568592 3346 568620 323546
rect 571432 320884 571484 320890
rect 571432 320826 571484 320832
rect 570604 297424 570656 297430
rect 570604 297366 570656 297372
rect 570616 3602 570644 297366
rect 571444 3738 571472 320826
rect 571984 311160 572036 311166
rect 571984 311102 572036 311108
rect 571432 3732 571484 3738
rect 571432 3674 571484 3680
rect 571996 3670 572024 311102
rect 572720 293276 572772 293282
rect 572720 293218 572772 293224
rect 572628 3732 572680 3738
rect 572628 3674 572680 3680
rect 571984 3664 572036 3670
rect 571984 3606 572036 3612
rect 570236 3596 570288 3602
rect 570236 3538 570288 3544
rect 570604 3596 570656 3602
rect 570604 3538 570656 3544
rect 571432 3596 571484 3602
rect 571432 3538 571484 3544
rect 567212 3318 567884 3346
rect 568592 3318 569080 3346
rect 566740 3052 566792 3058
rect 566740 2994 566792 3000
rect 566752 480 566780 2994
rect 567856 480 567884 3318
rect 569052 480 569080 3318
rect 570248 480 570276 3538
rect 571444 480 571472 3538
rect 572640 480 572668 3674
rect 572732 3346 572760 293218
rect 573376 3738 573404 334562
rect 574744 331900 574796 331906
rect 574744 331842 574796 331848
rect 573364 3732 573416 3738
rect 573364 3674 573416 3680
rect 574756 3602 574784 331842
rect 580172 322924 580224 322930
rect 580172 322866 580224 322872
rect 580184 322697 580212 322866
rect 580170 322688 580226 322697
rect 580170 322623 580226 322632
rect 580172 311840 580224 311846
rect 580172 311782 580224 311788
rect 580184 310865 580212 311782
rect 580170 310856 580226 310865
rect 580170 310791 580226 310800
rect 574836 308440 574888 308446
rect 574836 308382 574888 308388
rect 574744 3596 574796 3602
rect 574744 3538 574796 3544
rect 572732 3318 573864 3346
rect 574848 3330 574876 308382
rect 579804 299464 579856 299470
rect 579804 299406 579856 299412
rect 579816 299169 579844 299406
rect 579802 299160 579858 299169
rect 579802 299095 579858 299104
rect 580172 276004 580224 276010
rect 580172 275946 580224 275952
rect 580184 275777 580212 275946
rect 580170 275768 580226 275777
rect 580170 275703 580226 275712
rect 580172 264920 580224 264926
rect 580172 264862 580224 264868
rect 580184 263945 580212 264862
rect 580170 263936 580226 263945
rect 580170 263871 580226 263880
rect 579804 252544 579856 252550
rect 579804 252486 579856 252492
rect 579816 252249 579844 252486
rect 579802 252240 579858 252249
rect 579802 252175 579858 252184
rect 580172 218000 580224 218006
rect 580172 217942 580224 217948
rect 580184 217025 580212 217942
rect 580170 217016 580226 217025
rect 580170 216951 580226 216960
rect 579804 205624 579856 205630
rect 579804 205566 579856 205572
rect 579816 205329 579844 205566
rect 579802 205320 579858 205329
rect 579802 205255 579858 205264
rect 580172 182164 580224 182170
rect 580172 182106 580224 182112
rect 580184 181937 580212 182106
rect 580170 181928 580226 181937
rect 580170 181863 580226 181872
rect 580172 171080 580224 171086
rect 580172 171022 580224 171028
rect 580184 170105 580212 171022
rect 580170 170096 580226 170105
rect 580170 170031 580226 170040
rect 579804 158704 579856 158710
rect 579804 158646 579856 158652
rect 579816 158409 579844 158646
rect 579802 158400 579858 158409
rect 579802 158335 579858 158344
rect 580172 135244 580224 135250
rect 580172 135186 580224 135192
rect 580184 134881 580212 135186
rect 580170 134872 580226 134881
rect 580170 134807 580226 134816
rect 580172 124160 580224 124166
rect 580172 124102 580224 124108
rect 580184 123185 580212 124102
rect 580170 123176 580226 123185
rect 580170 123111 580226 123120
rect 579804 111784 579856 111790
rect 579804 111726 579856 111732
rect 579816 111489 579844 111726
rect 579802 111480 579858 111489
rect 579802 111415 579858 111424
rect 580172 88324 580224 88330
rect 580172 88266 580224 88272
rect 580184 87961 580212 88266
rect 580170 87952 580226 87961
rect 580170 87887 580226 87896
rect 579804 64864 579856 64870
rect 579804 64806 579856 64812
rect 579816 64569 579844 64806
rect 579802 64560 579858 64569
rect 579802 64495 579858 64504
rect 580172 41404 580224 41410
rect 580172 41346 580224 41352
rect 580184 41041 580212 41346
rect 580170 41032 580226 41041
rect 580170 40967 580226 40976
rect 579804 17944 579856 17950
rect 579804 17886 579856 17892
rect 579816 17649 579844 17886
rect 579802 17640 579858 17649
rect 579802 17575 579858 17584
rect 579804 3732 579856 3738
rect 579804 3674 579856 3680
rect 576216 3596 576268 3602
rect 576216 3538 576268 3544
rect 575020 3392 575072 3398
rect 575020 3334 575072 3340
rect 573836 480 573864 3318
rect 574836 3324 574888 3330
rect 574836 3266 574888 3272
rect 575032 480 575060 3334
rect 576228 480 576256 3538
rect 578608 3528 578660 3534
rect 578608 3470 578660 3476
rect 577412 3324 577464 3330
rect 577412 3266 577464 3272
rect 577424 480 577452 3266
rect 578620 480 578648 3470
rect 579816 480 579844 3674
rect 581000 3664 581052 3670
rect 581000 3606 581052 3612
rect 581012 480 581040 3606
rect 582196 3460 582248 3466
rect 582196 3402 582248 3408
rect 582208 480 582236 3402
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8822 -960 8934 480
rect 10018 -960 10130 480
rect 11214 -960 11326 480
rect 12410 -960 12522 480
rect 13606 -960 13718 480
rect 14802 -960 14914 480
rect 15998 -960 16110 480
rect 17194 -960 17306 480
rect 18298 -960 18410 480
rect 19494 -960 19606 480
rect 20690 -960 20802 480
rect 21886 -960 21998 480
rect 23082 -960 23194 480
rect 24278 -960 24390 480
rect 25474 -960 25586 480
rect 26670 -960 26782 480
rect 27866 -960 27978 480
rect 29062 -960 29174 480
rect 30258 -960 30370 480
rect 31454 -960 31566 480
rect 32650 -960 32762 480
rect 33846 -960 33958 480
rect 34950 -960 35062 480
rect 36146 -960 36258 480
rect 37342 -960 37454 480
rect 38538 -960 38650 480
rect 39734 -960 39846 480
rect 40930 -960 41042 480
rect 42126 -960 42238 480
rect 43322 -960 43434 480
rect 44518 -960 44630 480
rect 45714 -960 45826 480
rect 46910 -960 47022 480
rect 48106 -960 48218 480
rect 49302 -960 49414 480
rect 50498 -960 50610 480
rect 51602 -960 51714 480
rect 52798 -960 52910 480
rect 53994 -960 54106 480
rect 55190 -960 55302 480
rect 56386 -960 56498 480
rect 57582 -960 57694 480
rect 58778 -960 58890 480
rect 59974 -960 60086 480
rect 61170 -960 61282 480
rect 62366 -960 62478 480
rect 63562 -960 63674 480
rect 64758 -960 64870 480
rect 65954 -960 66066 480
rect 67150 -960 67262 480
rect 68254 -960 68366 480
rect 69450 -960 69562 480
rect 70646 -960 70758 480
rect 71842 -960 71954 480
rect 73038 -960 73150 480
rect 74234 -960 74346 480
rect 75430 -960 75542 480
rect 76626 -960 76738 480
rect 77822 -960 77934 480
rect 79018 -960 79130 480
rect 80214 -960 80326 480
rect 81410 -960 81522 480
rect 82606 -960 82718 480
rect 83802 -960 83914 480
rect 84906 -960 85018 480
rect 86102 -960 86214 480
rect 87298 -960 87410 480
rect 88494 -960 88606 480
rect 89690 -960 89802 480
rect 90886 -960 90998 480
rect 92082 -960 92194 480
rect 93278 -960 93390 480
rect 94474 -960 94586 480
rect 95670 -960 95782 480
rect 96866 -960 96978 480
rect 98062 -960 98174 480
rect 99258 -960 99370 480
rect 100454 -960 100566 480
rect 101558 -960 101670 480
rect 102754 -960 102866 480
rect 103950 -960 104062 480
rect 105146 -960 105258 480
rect 106342 -960 106454 480
rect 107538 -960 107650 480
rect 108734 -960 108846 480
rect 109930 -960 110042 480
rect 111126 -960 111238 480
rect 112322 -960 112434 480
rect 113518 -960 113630 480
rect 114714 -960 114826 480
rect 115910 -960 116022 480
rect 117106 -960 117218 480
rect 118210 -960 118322 480
rect 119406 -960 119518 480
rect 120602 -960 120714 480
rect 121798 -960 121910 480
rect 122994 -960 123106 480
rect 124190 -960 124302 480
rect 125386 -960 125498 480
rect 126582 -960 126694 480
rect 127778 -960 127890 480
rect 128974 -960 129086 480
rect 130170 -960 130282 480
rect 131366 -960 131478 480
rect 132562 -960 132674 480
rect 133758 -960 133870 480
rect 134862 -960 134974 480
rect 136058 -960 136170 480
rect 137254 -960 137366 480
rect 138450 -960 138562 480
rect 139646 -960 139758 480
rect 140842 -960 140954 480
rect 142038 -960 142150 480
rect 143234 -960 143346 480
rect 144430 -960 144542 480
rect 145626 -960 145738 480
rect 146822 -960 146934 480
rect 148018 -960 148130 480
rect 149214 -960 149326 480
rect 150410 -960 150522 480
rect 151514 -960 151626 480
rect 152710 -960 152822 480
rect 153906 -960 154018 480
rect 155102 -960 155214 480
rect 156298 -960 156410 480
rect 157494 -960 157606 480
rect 158690 -960 158802 480
rect 159886 -960 159998 480
rect 161082 -960 161194 480
rect 162278 -960 162390 480
rect 163474 -960 163586 480
rect 164670 -960 164782 480
rect 165866 -960 165978 480
rect 167062 -960 167174 480
rect 168166 -960 168278 480
rect 169362 -960 169474 480
rect 170558 -960 170670 480
rect 171754 -960 171866 480
rect 172950 -960 173062 480
rect 174146 -960 174258 480
rect 175342 -960 175454 480
rect 176538 -960 176650 480
rect 177734 -960 177846 480
rect 178930 -960 179042 480
rect 180126 -960 180238 480
rect 181322 -960 181434 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184818 -960 184930 480
rect 186014 -960 186126 480
rect 187210 -960 187322 480
rect 188406 -960 188518 480
rect 189602 -960 189714 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197974 -960 198086 480
rect 199170 -960 199282 480
rect 200366 -960 200478 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206254 -960 206366 480
rect 207450 -960 207562 480
rect 208646 -960 208758 480
rect 209842 -960 209954 480
rect 211038 -960 211150 480
rect 212234 -960 212346 480
rect 213430 -960 213542 480
rect 214626 -960 214738 480
rect 215822 -960 215934 480
rect 217018 -960 217130 480
rect 218122 -960 218234 480
rect 219318 -960 219430 480
rect 220514 -960 220626 480
rect 221710 -960 221822 480
rect 222906 -960 223018 480
rect 224102 -960 224214 480
rect 225298 -960 225410 480
rect 226494 -960 226606 480
rect 227690 -960 227802 480
rect 228886 -960 228998 480
rect 230082 -960 230194 480
rect 231278 -960 231390 480
rect 232474 -960 232586 480
rect 233670 -960 233782 480
rect 234774 -960 234886 480
rect 235970 -960 236082 480
rect 237166 -960 237278 480
rect 238362 -960 238474 480
rect 239558 -960 239670 480
rect 240754 -960 240866 480
rect 241950 -960 242062 480
rect 243146 -960 243258 480
rect 244342 -960 244454 480
rect 245538 -960 245650 480
rect 246734 -960 246846 480
rect 247930 -960 248042 480
rect 249126 -960 249238 480
rect 250322 -960 250434 480
rect 251426 -960 251538 480
rect 252622 -960 252734 480
rect 253818 -960 253930 480
rect 255014 -960 255126 480
rect 256210 -960 256322 480
rect 257406 -960 257518 480
rect 258602 -960 258714 480
rect 259798 -960 259910 480
rect 260994 -960 261106 480
rect 262190 -960 262302 480
rect 263386 -960 263498 480
rect 264582 -960 264694 480
rect 265778 -960 265890 480
rect 266974 -960 267086 480
rect 268078 -960 268190 480
rect 269274 -960 269386 480
rect 270470 -960 270582 480
rect 271666 -960 271778 480
rect 272862 -960 272974 480
rect 274058 -960 274170 480
rect 275254 -960 275366 480
rect 276450 -960 276562 480
rect 277646 -960 277758 480
rect 278842 -960 278954 480
rect 280038 -960 280150 480
rect 281234 -960 281346 480
rect 282430 -960 282542 480
rect 283626 -960 283738 480
rect 284730 -960 284842 480
rect 285926 -960 286038 480
rect 287122 -960 287234 480
rect 288318 -960 288430 480
rect 289514 -960 289626 480
rect 290710 -960 290822 480
rect 291906 -960 292018 480
rect 293102 -960 293214 480
rect 294298 -960 294410 480
rect 295494 -960 295606 480
rect 296690 -960 296802 480
rect 297886 -960 297998 480
rect 299082 -960 299194 480
rect 300278 -960 300390 480
rect 301382 -960 301494 480
rect 302578 -960 302690 480
rect 303774 -960 303886 480
rect 304970 -960 305082 480
rect 306166 -960 306278 480
rect 307362 -960 307474 480
rect 308558 -960 308670 480
rect 309754 -960 309866 480
rect 310950 -960 311062 480
rect 312146 -960 312258 480
rect 313342 -960 313454 480
rect 314538 -960 314650 480
rect 315734 -960 315846 480
rect 316930 -960 317042 480
rect 318034 -960 318146 480
rect 319230 -960 319342 480
rect 320426 -960 320538 480
rect 321622 -960 321734 480
rect 322818 -960 322930 480
rect 324014 -960 324126 480
rect 325210 -960 325322 480
rect 326406 -960 326518 480
rect 327602 -960 327714 480
rect 328798 -960 328910 480
rect 329994 -960 330106 480
rect 331190 -960 331302 480
rect 332386 -960 332498 480
rect 333582 -960 333694 480
rect 334686 -960 334798 480
rect 335882 -960 335994 480
rect 337078 -960 337190 480
rect 338274 -960 338386 480
rect 339470 -960 339582 480
rect 340666 -960 340778 480
rect 341862 -960 341974 480
rect 343058 -960 343170 480
rect 344254 -960 344366 480
rect 345450 -960 345562 480
rect 346646 -960 346758 480
rect 347842 -960 347954 480
rect 349038 -960 349150 480
rect 350234 -960 350346 480
rect 351338 -960 351450 480
rect 352534 -960 352646 480
rect 353730 -960 353842 480
rect 354926 -960 355038 480
rect 356122 -960 356234 480
rect 357318 -960 357430 480
rect 358514 -960 358626 480
rect 359710 -960 359822 480
rect 360906 -960 361018 480
rect 362102 -960 362214 480
rect 363298 -960 363410 480
rect 364494 -960 364606 480
rect 365690 -960 365802 480
rect 366886 -960 366998 480
rect 367990 -960 368102 480
rect 369186 -960 369298 480
rect 370382 -960 370494 480
rect 371578 -960 371690 480
rect 372774 -960 372886 480
rect 373970 -960 374082 480
rect 375166 -960 375278 480
rect 376362 -960 376474 480
rect 377558 -960 377670 480
rect 378754 -960 378866 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384642 -960 384754 480
rect 385838 -960 385950 480
rect 387034 -960 387146 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395406 -960 395518 480
rect 396602 -960 396714 480
rect 397798 -960 397910 480
rect 398994 -960 399106 480
rect 400190 -960 400302 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403686 -960 403798 480
rect 404882 -960 404994 480
rect 406078 -960 406190 480
rect 407274 -960 407386 480
rect 408470 -960 408582 480
rect 409666 -960 409778 480
rect 410862 -960 410974 480
rect 412058 -960 412170 480
rect 413254 -960 413366 480
rect 414450 -960 414562 480
rect 415646 -960 415758 480
rect 416842 -960 416954 480
rect 417946 -960 418058 480
rect 419142 -960 419254 480
rect 420338 -960 420450 480
rect 421534 -960 421646 480
rect 422730 -960 422842 480
rect 423926 -960 424038 480
rect 425122 -960 425234 480
rect 426318 -960 426430 480
rect 427514 -960 427626 480
rect 428710 -960 428822 480
rect 429906 -960 430018 480
rect 431102 -960 431214 480
rect 432298 -960 432410 480
rect 433494 -960 433606 480
rect 434598 -960 434710 480
rect 435794 -960 435906 480
rect 436990 -960 437102 480
rect 438186 -960 438298 480
rect 439382 -960 439494 480
rect 440578 -960 440690 480
rect 441774 -960 441886 480
rect 442970 -960 443082 480
rect 444166 -960 444278 480
rect 445362 -960 445474 480
rect 446558 -960 446670 480
rect 447754 -960 447866 480
rect 448950 -960 449062 480
rect 450146 -960 450258 480
rect 451250 -960 451362 480
rect 452446 -960 452558 480
rect 453642 -960 453754 480
rect 454838 -960 454950 480
rect 456034 -960 456146 480
rect 457230 -960 457342 480
rect 458426 -960 458538 480
rect 459622 -960 459734 480
rect 460818 -960 460930 480
rect 462014 -960 462126 480
rect 463210 -960 463322 480
rect 464406 -960 464518 480
rect 465602 -960 465714 480
rect 466798 -960 466910 480
rect 467902 -960 468014 480
rect 469098 -960 469210 480
rect 470294 -960 470406 480
rect 471490 -960 471602 480
rect 472686 -960 472798 480
rect 473882 -960 473994 480
rect 475078 -960 475190 480
rect 476274 -960 476386 480
rect 477470 -960 477582 480
rect 478666 -960 478778 480
rect 479862 -960 479974 480
rect 481058 -960 481170 480
rect 482254 -960 482366 480
rect 483450 -960 483562 480
rect 484554 -960 484666 480
rect 485750 -960 485862 480
rect 486946 -960 487058 480
rect 488142 -960 488254 480
rect 489338 -960 489450 480
rect 490534 -960 490646 480
rect 491730 -960 491842 480
rect 492926 -960 493038 480
rect 494122 -960 494234 480
rect 495318 -960 495430 480
rect 496514 -960 496626 480
rect 497710 -960 497822 480
rect 498906 -960 499018 480
rect 500102 -960 500214 480
rect 501206 -960 501318 480
rect 502402 -960 502514 480
rect 503598 -960 503710 480
rect 504794 -960 504906 480
rect 505990 -960 506102 480
rect 507186 -960 507298 480
rect 508382 -960 508494 480
rect 509578 -960 509690 480
rect 510774 -960 510886 480
rect 511970 -960 512082 480
rect 513166 -960 513278 480
rect 514362 -960 514474 480
rect 515558 -960 515670 480
rect 516754 -960 516866 480
rect 517858 -960 517970 480
rect 519054 -960 519166 480
rect 520250 -960 520362 480
rect 521446 -960 521558 480
rect 522642 -960 522754 480
rect 523838 -960 523950 480
rect 525034 -960 525146 480
rect 526230 -960 526342 480
rect 527426 -960 527538 480
rect 528622 -960 528734 480
rect 529818 -960 529930 480
rect 531014 -960 531126 480
rect 532210 -960 532322 480
rect 533406 -960 533518 480
rect 534510 -960 534622 480
rect 535706 -960 535818 480
rect 536902 -960 537014 480
rect 538098 -960 538210 480
rect 539294 -960 539406 480
rect 540490 -960 540602 480
rect 541686 -960 541798 480
rect 542882 -960 542994 480
rect 544078 -960 544190 480
rect 545274 -960 545386 480
rect 546470 -960 546582 480
rect 547666 -960 547778 480
rect 548862 -960 548974 480
rect 550058 -960 550170 480
rect 551162 -960 551274 480
rect 552358 -960 552470 480
rect 553554 -960 553666 480
rect 554750 -960 554862 480
rect 555946 -960 556058 480
rect 557142 -960 557254 480
rect 558338 -960 558450 480
rect 559534 -960 559646 480
rect 560730 -960 560842 480
rect 561926 -960 562038 480
rect 563122 -960 563234 480
rect 564318 -960 564430 480
rect 565514 -960 565626 480
rect 566710 -960 566822 480
rect 567814 -960 567926 480
rect 569010 -960 569122 480
rect 570206 -960 570318 480
rect 571402 -960 571514 480
rect 572598 -960 572710 480
rect 573794 -960 573906 480
rect 574990 -960 575102 480
rect 576186 -960 576298 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3422 682216 3478 682272
rect 3054 653520 3110 653576
rect 3330 595992 3386 596048
rect 3330 553016 3386 553072
rect 3238 538600 3294 538656
rect 3330 495508 3386 495544
rect 3330 495488 3332 495508
rect 3332 495488 3384 495508
rect 3384 495488 3386 495508
rect 2962 481072 3018 481128
rect 3330 437960 3386 438016
rect 3330 423700 3386 423736
rect 3330 423680 3332 423700
rect 3332 423680 3384 423700
rect 3384 423680 3386 423700
rect 3514 667956 3570 667992
rect 3514 667936 3516 667956
rect 3516 667936 3568 667956
rect 3568 667936 3570 667956
rect 3514 624824 3570 624880
rect 3606 610408 3662 610464
rect 3698 567296 3754 567352
rect 3882 509904 3938 509960
rect 4066 452376 4122 452432
rect 154210 482976 154266 483032
rect 154486 482976 154542 483032
rect 218886 695680 218942 695736
rect 219254 695544 219310 695600
rect 218978 540912 219034 540968
rect 219162 540912 219218 540968
rect 218978 531256 219034 531312
rect 219162 531256 219218 531312
rect 218794 521600 218850 521656
rect 218978 521600 219034 521656
rect 218978 473320 219034 473376
rect 219254 473320 219310 473376
rect 218978 425040 219034 425096
rect 219346 425040 219402 425096
rect 3146 394984 3202 395040
rect 3422 380568 3478 380624
rect 2962 366152 3018 366208
rect 3422 337456 3478 337512
rect 3422 308760 3478 308816
rect 3054 294344 3110 294400
rect 2870 265648 2926 265704
rect 3422 251232 3478 251288
rect 17222 397976 17278 398032
rect 3974 323040 4030 323096
rect 3790 280064 3846 280120
rect 3606 236952 3662 237008
rect 3146 222536 3202 222592
rect 3422 208120 3478 208176
rect 3330 194520 3386 194576
rect 3330 193840 3386 193896
rect 3238 179424 3294 179480
rect 3514 165008 3570 165064
rect 3146 150728 3202 150784
rect 3238 136312 3294 136368
rect 3422 122032 3478 122088
rect 3422 108976 3478 109032
rect 3422 107616 3478 107672
rect 3422 93200 3478 93256
rect 3422 78920 3478 78976
rect 3330 64504 3386 64560
rect 3422 50088 3478 50144
rect 3422 35844 3424 35864
rect 3424 35844 3476 35864
rect 3476 35844 3478 35864
rect 3422 35808 3478 35844
rect 3146 21392 3202 21448
rect 3422 7112 3478 7168
rect 6458 3304 6514 3360
rect 14830 3440 14886 3496
rect 16026 3576 16082 3632
rect 25502 3848 25558 3904
rect 24306 3712 24362 3768
rect 32678 3984 32734 4040
rect 200762 398248 200818 398304
rect 198002 398112 198058 398168
rect 225694 398656 225750 398712
rect 258078 402464 258134 402520
rect 261206 402484 261262 402520
rect 261206 402464 261208 402484
rect 261208 402464 261260 402484
rect 261260 402464 261262 402484
rect 580170 697992 580226 698048
rect 580170 686296 580226 686352
rect 580170 674600 580226 674656
rect 580170 651072 580226 651128
rect 580170 639376 580226 639432
rect 580170 627680 580226 627736
rect 580170 604152 580226 604208
rect 580170 592456 580226 592512
rect 580170 580760 580226 580816
rect 299570 560496 299626 560552
rect 299570 560360 299626 560416
rect 580170 557232 580226 557288
rect 299294 549208 299350 549264
rect 299478 549208 299534 549264
rect 580170 545536 580226 545592
rect 580170 533840 580226 533896
rect 299662 521600 299718 521656
rect 299846 521600 299902 521656
rect 580170 510312 580226 510368
rect 299478 502288 299534 502344
rect 299754 502324 299756 502344
rect 299756 502324 299808 502344
rect 299808 502324 299810 502344
rect 299754 502288 299810 502324
rect 580170 498616 580226 498672
rect 299478 492632 299534 492688
rect 299662 492652 299718 492688
rect 299662 492632 299664 492652
rect 299664 492632 299716 492652
rect 299716 492632 299718 492652
rect 580170 486784 580226 486840
rect 580170 463392 580226 463448
rect 580170 451696 580226 451752
rect 580170 439864 580226 439920
rect 580170 416472 580226 416528
rect 580170 404776 580226 404832
rect 231582 399336 231638 399392
rect 232962 399336 233018 399392
rect 237194 399336 237250 399392
rect 238298 399336 238354 399392
rect 242530 399336 242586 399392
rect 276846 399336 276902 399392
rect 283010 399336 283066 399392
rect 284482 399336 284538 399392
rect 286138 399336 286194 399392
rect 287334 399336 287390 399392
rect 287886 399336 287942 399392
rect 224958 3168 225014 3224
rect 229558 241440 229614 241496
rect 229834 241440 229890 241496
rect 229558 222128 229614 222184
rect 229834 222128 229890 222184
rect 229558 202816 229614 202872
rect 229834 202816 229890 202872
rect 229558 183504 229614 183560
rect 229834 183504 229890 183560
rect 229650 154536 229706 154592
rect 229834 154536 229890 154592
rect 229466 135224 229522 135280
rect 229650 135224 229706 135280
rect 229466 115912 229522 115968
rect 229650 115912 229706 115968
rect 229466 96600 229522 96656
rect 229650 96600 229706 96656
rect 229834 3168 229890 3224
rect 231122 3304 231178 3360
rect 231582 3576 231638 3632
rect 231398 3440 231454 3496
rect 233790 144880 233846 144936
rect 233974 144880 234030 144936
rect 233790 86944 233846 87000
rect 233974 86944 234030 87000
rect 233606 3984 233662 4040
rect 232962 3848 233018 3904
rect 232778 3712 232834 3768
rect 234986 241440 235042 241496
rect 234986 220768 235042 220824
rect 234986 211112 235042 211168
rect 234986 183540 234988 183560
rect 234988 183540 235040 183560
rect 235040 183540 235042 183560
rect 234986 183504 235042 183540
rect 234986 162832 235042 162888
rect 235170 241440 235226 241496
rect 235538 241440 235594 241496
rect 235722 241440 235778 241496
rect 235170 220768 235226 220824
rect 235538 220768 235594 220824
rect 235722 220768 235778 220824
rect 235170 211112 235226 211168
rect 235538 211112 235594 211168
rect 235722 211112 235778 211168
rect 235170 183540 235172 183560
rect 235172 183540 235224 183560
rect 235224 183540 235226 183560
rect 235170 183504 235226 183540
rect 235170 162832 235226 162888
rect 235538 87080 235594 87136
rect 235446 86944 235502 87000
rect 238758 153176 238814 153232
rect 238942 153176 238998 153232
rect 238942 145016 238998 145072
rect 238758 144744 238814 144800
rect 238758 135224 238814 135280
rect 238942 135224 238998 135280
rect 238942 125704 238998 125760
rect 238758 125296 238814 125352
rect 238758 115912 238814 115968
rect 238942 115912 238998 115968
rect 245014 222128 245070 222184
rect 245198 222128 245254 222184
rect 245014 202816 245070 202872
rect 245198 202816 245254 202872
rect 245014 183504 245070 183560
rect 245198 183504 245254 183560
rect 245014 143520 245070 143576
rect 245198 143520 245254 143576
rect 248418 227976 248474 228032
rect 248418 227840 248474 227896
rect 250258 280064 250314 280120
rect 250442 280064 250498 280120
rect 250718 261024 250774 261080
rect 250442 260888 250498 260944
rect 250718 142296 250774 142352
rect 250626 142160 250682 142216
rect 250442 44104 250498 44160
rect 250718 44104 250774 44160
rect 254858 314608 254914 314664
rect 254766 304972 254822 305008
rect 254766 304952 254768 304972
rect 254768 304952 254820 304972
rect 254820 304952 254822 304972
rect 254858 295316 254914 295352
rect 254858 295296 254860 295316
rect 254860 295296 254912 295316
rect 254912 295296 254914 295316
rect 255042 295296 255098 295352
rect 254766 91024 254822 91080
rect 255042 91024 255098 91080
rect 254858 80008 254914 80064
rect 255042 80008 255098 80064
rect 254858 70352 254914 70408
rect 255042 70352 255098 70408
rect 255778 289076 255780 289096
rect 255780 289076 255832 289096
rect 255832 289076 255834 289096
rect 255778 289040 255834 289076
rect 255778 275984 255834 276040
rect 255778 227704 255834 227760
rect 256054 227704 256110 227760
rect 255870 125568 255926 125624
rect 255870 106256 255926 106312
rect 256054 125568 256110 125624
rect 256054 106256 256110 106312
rect 256422 314608 256478 314664
rect 256606 314608 256662 314664
rect 256422 304952 256478 305008
rect 256606 304952 256662 305008
rect 256422 285640 256478 285696
rect 256606 285640 256662 285696
rect 256974 259392 257030 259448
rect 256422 193160 256478 193216
rect 256606 193160 256662 193216
rect 256974 62056 257030 62112
rect 257158 259392 257214 259448
rect 257250 229064 257306 229120
rect 257250 228928 257306 228984
rect 257250 164192 257306 164248
rect 257158 62056 257214 62112
rect 257434 164192 257490 164248
rect 259918 189080 259974 189136
rect 259734 188944 259790 189000
rect 259734 71712 259790 71768
rect 260102 71712 260158 71768
rect 260378 324300 260380 324320
rect 260380 324300 260432 324320
rect 260432 324300 260434 324320
rect 260378 324264 260434 324300
rect 260654 324300 260656 324320
rect 260656 324300 260708 324320
rect 260708 324300 260710 324320
rect 260654 324264 260710 324300
rect 260654 266464 260710 266520
rect 260654 266328 260710 266384
rect 260562 227704 260618 227760
rect 260746 227704 260802 227760
rect 260930 208392 260986 208448
rect 260746 208256 260802 208312
rect 260654 177928 260710 177984
rect 260838 177928 260894 177984
rect 260654 168408 260710 168464
rect 260838 168408 260894 168464
rect 260562 100680 260618 100736
rect 260654 100544 260710 100600
rect 262402 324264 262458 324320
rect 262678 324300 262680 324320
rect 262680 324300 262732 324320
rect 262732 324300 262734 324320
rect 262678 324264 262734 324300
rect 262494 237360 262550 237416
rect 262678 237360 262734 237416
rect 263690 337084 263692 337104
rect 263692 337084 263744 337104
rect 263744 337084 263746 337104
rect 263690 337048 263746 337084
rect 264242 306348 264244 306368
rect 264244 306348 264296 306368
rect 264296 306348 264298 306368
rect 264242 306312 264298 306348
rect 264426 306312 264482 306368
rect 266266 227976 266322 228032
rect 266266 227704 266322 227760
rect 267738 337084 267740 337104
rect 267740 337084 267792 337104
rect 267792 337084 267794 337104
rect 267738 337048 267794 337084
rect 268842 190440 268898 190496
rect 269026 190440 269082 190496
rect 271602 295296 271658 295352
rect 271786 295296 271842 295352
rect 273626 336912 273682 336968
rect 273810 336776 273866 336832
rect 273810 91024 273866 91080
rect 274086 91024 274142 91080
rect 277030 335552 277086 335608
rect 277306 335314 277362 335370
rect 277030 324264 277086 324320
rect 277398 324300 277400 324320
rect 277400 324300 277452 324320
rect 277452 324300 277454 324320
rect 277398 324264 277454 324300
rect 276846 275984 276902 276040
rect 277030 275984 277086 276040
rect 277582 212472 277638 212528
rect 277766 212472 277822 212528
rect 276938 100680 276994 100736
rect 277214 100680 277270 100736
rect 278686 227740 278688 227760
rect 278688 227740 278740 227760
rect 278740 227740 278742 227760
rect 278686 227704 278742 227740
rect 278134 3984 278190 4040
rect 278042 3848 278098 3904
rect 277858 3712 277914 3768
rect 280802 337864 280858 337920
rect 280250 29044 280252 29064
rect 280252 29044 280304 29064
rect 280304 29044 280306 29064
rect 280250 29008 280306 29044
rect 281906 337728 281962 337784
rect 279974 3576 280030 3632
rect 279882 3440 279938 3496
rect 279790 3304 279846 3360
rect 282642 338000 282698 338056
rect 285218 336912 285274 336968
rect 285586 336912 285642 336968
rect 287702 337764 287704 337784
rect 287704 337764 287756 337784
rect 287756 337764 287758 337784
rect 287702 337728 287758 337764
rect 288070 338000 288126 338056
rect 289542 337864 289598 337920
rect 289818 337864 289874 337920
rect 289726 227740 289728 227760
rect 289728 227740 289780 227760
rect 289780 227740 289782 227760
rect 289726 227704 289782 227740
rect 289726 29044 289728 29064
rect 289728 29044 289780 29064
rect 289780 29044 289782 29064
rect 289726 29008 289782 29044
rect 291106 337864 291162 337920
rect 302146 227840 302202 227896
rect 302146 227432 302202 227488
rect 302146 76064 302202 76120
rect 302146 75656 302202 75712
rect 307758 333804 307814 333806
rect 307758 333752 307760 333804
rect 307760 333752 307812 333804
rect 307812 333752 307814 333804
rect 307758 333750 307814 333752
rect 307758 333512 307814 333568
rect 309782 398520 309838 398576
rect 309138 227740 309140 227760
rect 309140 227740 309192 227760
rect 309192 227740 309194 227760
rect 309138 227704 309194 227740
rect 309138 75964 309140 75984
rect 309140 75964 309192 75984
rect 309192 75964 309194 75984
rect 309138 75928 309194 75964
rect 312634 227840 312690 227896
rect 313922 76064 313978 76120
rect 326342 398384 326398 398440
rect 323582 227840 323638 227896
rect 323582 227568 323638 227624
rect 323582 76064 323638 76120
rect 323582 75792 323638 75848
rect 328458 227976 328514 228032
rect 328550 227568 328606 227624
rect 328458 76200 328514 76256
rect 328550 75792 328606 75848
rect 398102 29144 398158 29200
rect 405646 29300 405702 29336
rect 405646 29280 405648 29300
rect 405648 29280 405700 29300
rect 405700 29280 405702 29300
rect 415306 76064 415362 76120
rect 415306 75928 415362 75984
rect 418066 227996 418122 228032
rect 418066 227976 418068 227996
rect 418068 227976 418120 227996
rect 418120 227976 418122 227996
rect 417330 29180 417332 29200
rect 417332 29180 417384 29200
rect 417384 29180 417386 29200
rect 417330 29144 417386 29180
rect 424966 227996 425022 228032
rect 424966 227976 424968 227996
rect 424968 227976 425020 227996
rect 425020 227976 425022 227996
rect 424966 29280 425022 29336
rect 437386 227860 437442 227896
rect 437386 227840 437388 227860
rect 437388 227840 437440 227860
rect 437440 227840 437442 227860
rect 437386 76084 437442 76120
rect 437386 76064 437388 76084
rect 437388 76064 437440 76084
rect 437440 76064 437442 76084
rect 436742 29144 436798 29200
rect 444286 227704 444342 227760
rect 444286 75928 444342 75984
rect 444286 29300 444342 29336
rect 444286 29280 444288 29300
rect 444288 29280 444340 29300
rect 444340 29280 444342 29300
rect 456706 227840 456762 227896
rect 456890 227840 456946 227896
rect 456706 76064 456762 76120
rect 456890 76064 456946 76120
rect 456706 29180 456708 29200
rect 456708 29180 456760 29200
rect 456760 29180 456762 29200
rect 456706 29144 456762 29180
rect 463606 29280 463662 29336
rect 464434 3984 464490 4040
rect 467930 3848 467986 3904
rect 471518 3712 471574 3768
rect 475290 29180 475292 29200
rect 475292 29180 475344 29200
rect 475344 29180 475346 29200
rect 475290 29144 475346 29180
rect 475106 3576 475162 3632
rect 476026 227860 476082 227896
rect 476026 227840 476028 227860
rect 476028 227840 476080 227860
rect 476080 227840 476082 227860
rect 478694 3440 478750 3496
rect 482926 227704 482982 227760
rect 482926 76064 482982 76120
rect 482926 75928 482982 75984
rect 482926 29280 482982 29336
rect 482282 3304 482338 3360
rect 495346 227876 495348 227896
rect 495348 227876 495400 227896
rect 495400 227876 495402 227896
rect 495346 227840 495402 227876
rect 495162 29180 495164 29200
rect 495164 29180 495216 29200
rect 495216 29180 495218 29200
rect 495162 29144 495218 29180
rect 497002 227876 497004 227896
rect 497004 227876 497056 227896
rect 497056 227876 497058 227896
rect 497002 227840 497058 227876
rect 579802 392944 579858 393000
rect 580170 369552 580226 369608
rect 580078 357856 580134 357912
rect 579802 346024 579858 346080
rect 502246 75792 502302 75848
rect 502246 29280 502302 29336
rect 510526 76200 510582 76256
rect 514666 227860 514722 227896
rect 514666 227840 514668 227860
rect 514668 227840 514720 227860
rect 514720 227840 514722 227860
rect 513562 29180 513564 29200
rect 513564 29180 513616 29200
rect 513616 29180 513618 29200
rect 513562 29144 513618 29180
rect 521566 227704 521622 227760
rect 521566 76472 521622 76528
rect 521566 75928 521622 75984
rect 521566 29280 521622 29336
rect 533986 227840 534042 227896
rect 533986 76084 534042 76120
rect 533986 76064 533988 76084
rect 533988 76064 534040 76084
rect 534040 76064 534042 76084
rect 533802 29180 533804 29200
rect 533804 29180 533856 29200
rect 533856 29180 533858 29200
rect 533802 29144 533858 29180
rect 540886 227740 540888 227760
rect 540888 227740 540940 227760
rect 540940 227740 540942 227760
rect 540886 227704 540942 227740
rect 540886 75928 540942 75984
rect 540886 29280 540942 29336
rect 553306 227876 553308 227896
rect 553308 227876 553360 227896
rect 553360 227876 553362 227896
rect 553306 227840 553362 227876
rect 553306 76100 553308 76120
rect 553308 76100 553360 76120
rect 553360 76100 553362 76120
rect 553306 76064 553362 76100
rect 552478 29180 552480 29200
rect 552480 29180 552532 29200
rect 552532 29180 552534 29200
rect 552478 29144 552534 29180
rect 554594 227876 554596 227896
rect 554596 227876 554648 227896
rect 554648 227876 554650 227896
rect 554594 227840 554650 227876
rect 554594 76100 554596 76120
rect 554596 76100 554648 76120
rect 554648 76100 554650 76120
rect 554594 76064 554650 76100
rect 560206 29280 560262 29336
rect 580170 322632 580226 322688
rect 580170 310800 580226 310856
rect 579802 299104 579858 299160
rect 580170 275712 580226 275768
rect 580170 263880 580226 263936
rect 579802 252184 579858 252240
rect 580170 216960 580226 217016
rect 579802 205264 579858 205320
rect 580170 181872 580226 181928
rect 580170 170040 580226 170096
rect 579802 158344 579858 158400
rect 580170 134816 580226 134872
rect 580170 123120 580226 123176
rect 579802 111424 579858 111480
rect 580170 87896 580226 87952
rect 579802 64504 579858 64560
rect 580170 40976 580226 41032
rect 579802 17584 579858 17640
<< metal3 >>
rect 580165 698050 580231 698053
rect 583520 698050 584960 698140
rect 580165 698048 584960 698050
rect 580165 697992 580170 698048
rect 580226 697992 584960 698048
rect 580165 697990 584960 697992
rect 580165 697987 580231 697990
rect 583520 697900 584960 697990
rect -960 696540 480 696780
rect 218881 695738 218947 695741
rect 218881 695736 219450 695738
rect 218881 695680 218886 695736
rect 218942 695680 219450 695736
rect 218881 695678 219450 695680
rect 218881 695675 218947 695678
rect 219249 695602 219315 695605
rect 219390 695602 219450 695678
rect 219249 695600 219450 695602
rect 219249 695544 219254 695600
rect 219310 695544 219450 695600
rect 219249 695542 219450 695544
rect 219249 695539 219315 695542
rect 580165 686354 580231 686357
rect 583520 686354 584960 686444
rect 580165 686352 584960 686354
rect 580165 686296 580170 686352
rect 580226 686296 584960 686352
rect 580165 686294 584960 686296
rect 580165 686291 580231 686294
rect 583520 686204 584960 686294
rect -960 682274 480 682364
rect 3417 682274 3483 682277
rect -960 682272 3483 682274
rect -960 682216 3422 682272
rect 3478 682216 3483 682272
rect -960 682214 3483 682216
rect -960 682124 480 682214
rect 3417 682211 3483 682214
rect 580165 674658 580231 674661
rect 583520 674658 584960 674748
rect 580165 674656 584960 674658
rect 580165 674600 580170 674656
rect 580226 674600 584960 674656
rect 580165 674598 584960 674600
rect 580165 674595 580231 674598
rect 583520 674508 584960 674598
rect -960 667994 480 668084
rect 3509 667994 3575 667997
rect -960 667992 3575 667994
rect -960 667936 3514 667992
rect 3570 667936 3575 667992
rect -960 667934 3575 667936
rect -960 667844 480 667934
rect 3509 667931 3575 667934
rect 583520 662676 584960 662916
rect -960 653578 480 653668
rect 3049 653578 3115 653581
rect -960 653576 3115 653578
rect -960 653520 3054 653576
rect 3110 653520 3115 653576
rect -960 653518 3115 653520
rect -960 653428 480 653518
rect 3049 653515 3115 653518
rect 580165 651130 580231 651133
rect 583520 651130 584960 651220
rect 580165 651128 584960 651130
rect 580165 651072 580170 651128
rect 580226 651072 584960 651128
rect 580165 651070 584960 651072
rect 580165 651067 580231 651070
rect 583520 650980 584960 651070
rect 580165 639434 580231 639437
rect 583520 639434 584960 639524
rect 580165 639432 584960 639434
rect 580165 639376 580170 639432
rect 580226 639376 584960 639432
rect 580165 639374 584960 639376
rect 580165 639371 580231 639374
rect 583520 639284 584960 639374
rect -960 639012 480 639252
rect 580165 627738 580231 627741
rect 583520 627738 584960 627828
rect 580165 627736 584960 627738
rect 580165 627680 580170 627736
rect 580226 627680 584960 627736
rect 580165 627678 584960 627680
rect 580165 627675 580231 627678
rect 583520 627588 584960 627678
rect -960 624882 480 624972
rect 3509 624882 3575 624885
rect -960 624880 3575 624882
rect -960 624824 3514 624880
rect 3570 624824 3575 624880
rect -960 624822 3575 624824
rect -960 624732 480 624822
rect 3509 624819 3575 624822
rect 583520 615756 584960 615996
rect -960 610466 480 610556
rect 3601 610466 3667 610469
rect -960 610464 3667 610466
rect -960 610408 3606 610464
rect 3662 610408 3667 610464
rect -960 610406 3667 610408
rect -960 610316 480 610406
rect 3601 610403 3667 610406
rect 580165 604210 580231 604213
rect 583520 604210 584960 604300
rect 580165 604208 584960 604210
rect 580165 604152 580170 604208
rect 580226 604152 584960 604208
rect 580165 604150 584960 604152
rect 580165 604147 580231 604150
rect 583520 604060 584960 604150
rect -960 596050 480 596140
rect 3325 596050 3391 596053
rect -960 596048 3391 596050
rect -960 595992 3330 596048
rect 3386 595992 3391 596048
rect -960 595990 3391 595992
rect -960 595900 480 595990
rect 3325 595987 3391 595990
rect 580165 592514 580231 592517
rect 583520 592514 584960 592604
rect 580165 592512 584960 592514
rect 580165 592456 580170 592512
rect 580226 592456 584960 592512
rect 580165 592454 584960 592456
rect 580165 592451 580231 592454
rect 583520 592364 584960 592454
rect -960 581620 480 581860
rect 580165 580818 580231 580821
rect 583520 580818 584960 580908
rect 580165 580816 584960 580818
rect 580165 580760 580170 580816
rect 580226 580760 584960 580816
rect 580165 580758 584960 580760
rect 580165 580755 580231 580758
rect 583520 580668 584960 580758
rect 583520 568836 584960 569076
rect -960 567354 480 567444
rect 3693 567354 3759 567357
rect -960 567352 3759 567354
rect -960 567296 3698 567352
rect 3754 567296 3759 567352
rect -960 567294 3759 567296
rect -960 567204 480 567294
rect 3693 567291 3759 567294
rect 299565 560554 299631 560557
rect 299430 560552 299631 560554
rect 299430 560496 299570 560552
rect 299626 560496 299631 560552
rect 299430 560494 299631 560496
rect 299430 560418 299490 560494
rect 299565 560491 299631 560494
rect 299565 560418 299631 560421
rect 299430 560416 299631 560418
rect 299430 560360 299570 560416
rect 299626 560360 299631 560416
rect 299430 560358 299631 560360
rect 299565 560355 299631 560358
rect 580165 557290 580231 557293
rect 583520 557290 584960 557380
rect 580165 557288 584960 557290
rect 580165 557232 580170 557288
rect 580226 557232 584960 557288
rect 580165 557230 584960 557232
rect 580165 557227 580231 557230
rect 583520 557140 584960 557230
rect -960 553074 480 553164
rect 3325 553074 3391 553077
rect -960 553072 3391 553074
rect -960 553016 3330 553072
rect 3386 553016 3391 553072
rect -960 553014 3391 553016
rect -960 552924 480 553014
rect 3325 553011 3391 553014
rect 299289 549266 299355 549269
rect 299473 549266 299539 549269
rect 299289 549264 299539 549266
rect 299289 549208 299294 549264
rect 299350 549208 299478 549264
rect 299534 549208 299539 549264
rect 299289 549206 299539 549208
rect 299289 549203 299355 549206
rect 299473 549203 299539 549206
rect 580165 545594 580231 545597
rect 583520 545594 584960 545684
rect 580165 545592 584960 545594
rect 580165 545536 580170 545592
rect 580226 545536 584960 545592
rect 580165 545534 584960 545536
rect 580165 545531 580231 545534
rect 583520 545444 584960 545534
rect 218973 540970 219039 540973
rect 219157 540970 219223 540973
rect 218973 540968 219223 540970
rect 218973 540912 218978 540968
rect 219034 540912 219162 540968
rect 219218 540912 219223 540968
rect 218973 540910 219223 540912
rect 218973 540907 219039 540910
rect 219157 540907 219223 540910
rect -960 538658 480 538748
rect 3233 538658 3299 538661
rect -960 538656 3299 538658
rect -960 538600 3238 538656
rect 3294 538600 3299 538656
rect -960 538598 3299 538600
rect -960 538508 480 538598
rect 3233 538595 3299 538598
rect 580165 533898 580231 533901
rect 583520 533898 584960 533988
rect 580165 533896 584960 533898
rect 580165 533840 580170 533896
rect 580226 533840 584960 533896
rect 580165 533838 584960 533840
rect 580165 533835 580231 533838
rect 583520 533748 584960 533838
rect 218973 531314 219039 531317
rect 219157 531314 219223 531317
rect 218973 531312 219223 531314
rect 218973 531256 218978 531312
rect 219034 531256 219162 531312
rect 219218 531256 219223 531312
rect 218973 531254 219223 531256
rect 218973 531251 219039 531254
rect 219157 531251 219223 531254
rect -960 524092 480 524332
rect 583520 521916 584960 522156
rect 218789 521658 218855 521661
rect 218973 521658 219039 521661
rect 218789 521656 219039 521658
rect 218789 521600 218794 521656
rect 218850 521600 218978 521656
rect 219034 521600 219039 521656
rect 218789 521598 219039 521600
rect 218789 521595 218855 521598
rect 218973 521595 219039 521598
rect 299657 521658 299723 521661
rect 299841 521658 299907 521661
rect 299657 521656 299907 521658
rect 299657 521600 299662 521656
rect 299718 521600 299846 521656
rect 299902 521600 299907 521656
rect 299657 521598 299907 521600
rect 299657 521595 299723 521598
rect 299841 521595 299907 521598
rect 580165 510370 580231 510373
rect 583520 510370 584960 510460
rect 580165 510368 584960 510370
rect 580165 510312 580170 510368
rect 580226 510312 584960 510368
rect 580165 510310 584960 510312
rect 580165 510307 580231 510310
rect 583520 510220 584960 510310
rect -960 509962 480 510052
rect 3877 509962 3943 509965
rect -960 509960 3943 509962
rect -960 509904 3882 509960
rect 3938 509904 3943 509960
rect -960 509902 3943 509904
rect -960 509812 480 509902
rect 3877 509899 3943 509902
rect 299473 502346 299539 502349
rect 299749 502346 299815 502349
rect 299473 502344 299815 502346
rect 299473 502288 299478 502344
rect 299534 502288 299754 502344
rect 299810 502288 299815 502344
rect 299473 502286 299815 502288
rect 299473 502283 299539 502286
rect 299749 502283 299815 502286
rect 580165 498674 580231 498677
rect 583520 498674 584960 498764
rect 580165 498672 584960 498674
rect 580165 498616 580170 498672
rect 580226 498616 584960 498672
rect 580165 498614 584960 498616
rect 580165 498611 580231 498614
rect 583520 498524 584960 498614
rect -960 495546 480 495636
rect 3325 495546 3391 495549
rect -960 495544 3391 495546
rect -960 495488 3330 495544
rect 3386 495488 3391 495544
rect -960 495486 3391 495488
rect -960 495396 480 495486
rect 3325 495483 3391 495486
rect 299473 492690 299539 492693
rect 299657 492690 299723 492693
rect 299473 492688 299723 492690
rect 299473 492632 299478 492688
rect 299534 492632 299662 492688
rect 299718 492632 299723 492688
rect 299473 492630 299723 492632
rect 299473 492627 299539 492630
rect 299657 492627 299723 492630
rect 580165 486842 580231 486845
rect 583520 486842 584960 486932
rect 580165 486840 584960 486842
rect 580165 486784 580170 486840
rect 580226 486784 584960 486840
rect 580165 486782 584960 486784
rect 580165 486779 580231 486782
rect 583520 486692 584960 486782
rect 154205 483034 154271 483037
rect 154481 483034 154547 483037
rect 154205 483032 154547 483034
rect 154205 482976 154210 483032
rect 154266 482976 154486 483032
rect 154542 482976 154547 483032
rect 154205 482974 154547 482976
rect 154205 482971 154271 482974
rect 154481 482971 154547 482974
rect -960 481130 480 481220
rect 2957 481130 3023 481133
rect -960 481128 3023 481130
rect -960 481072 2962 481128
rect 3018 481072 3023 481128
rect -960 481070 3023 481072
rect -960 480980 480 481070
rect 2957 481067 3023 481070
rect 583520 474996 584960 475236
rect 218973 473378 219039 473381
rect 219249 473378 219315 473381
rect 218973 473376 219315 473378
rect 218973 473320 218978 473376
rect 219034 473320 219254 473376
rect 219310 473320 219315 473376
rect 218973 473318 219315 473320
rect 218973 473315 219039 473318
rect 219249 473315 219315 473318
rect -960 466700 480 466940
rect 580165 463450 580231 463453
rect 583520 463450 584960 463540
rect 580165 463448 584960 463450
rect 580165 463392 580170 463448
rect 580226 463392 584960 463448
rect 580165 463390 584960 463392
rect 580165 463387 580231 463390
rect 583520 463300 584960 463390
rect -960 452434 480 452524
rect 4061 452434 4127 452437
rect -960 452432 4127 452434
rect -960 452376 4066 452432
rect 4122 452376 4127 452432
rect -960 452374 4127 452376
rect -960 452284 480 452374
rect 4061 452371 4127 452374
rect 580165 451754 580231 451757
rect 583520 451754 584960 451844
rect 580165 451752 584960 451754
rect 580165 451696 580170 451752
rect 580226 451696 584960 451752
rect 580165 451694 584960 451696
rect 580165 451691 580231 451694
rect 583520 451604 584960 451694
rect 580165 439922 580231 439925
rect 583520 439922 584960 440012
rect 580165 439920 584960 439922
rect 580165 439864 580170 439920
rect 580226 439864 584960 439920
rect 580165 439862 584960 439864
rect 580165 439859 580231 439862
rect 583520 439772 584960 439862
rect -960 438018 480 438108
rect 3325 438018 3391 438021
rect -960 438016 3391 438018
rect -960 437960 3330 438016
rect 3386 437960 3391 438016
rect -960 437958 3391 437960
rect -960 437868 480 437958
rect 3325 437955 3391 437958
rect 583520 428076 584960 428316
rect 218973 425098 219039 425101
rect 219341 425098 219407 425101
rect 218973 425096 219407 425098
rect 218973 425040 218978 425096
rect 219034 425040 219346 425096
rect 219402 425040 219407 425096
rect 218973 425038 219407 425040
rect 218973 425035 219039 425038
rect 219341 425035 219407 425038
rect -960 423738 480 423828
rect 3325 423738 3391 423741
rect -960 423736 3391 423738
rect -960 423680 3330 423736
rect 3386 423680 3391 423736
rect -960 423678 3391 423680
rect -960 423588 480 423678
rect 3325 423675 3391 423678
rect 580165 416530 580231 416533
rect 583520 416530 584960 416620
rect 580165 416528 584960 416530
rect 580165 416472 580170 416528
rect 580226 416472 584960 416528
rect 580165 416470 584960 416472
rect 580165 416467 580231 416470
rect 583520 416380 584960 416470
rect -960 409172 480 409412
rect 580165 404834 580231 404837
rect 583520 404834 584960 404924
rect 580165 404832 584960 404834
rect 580165 404776 580170 404832
rect 580226 404776 584960 404832
rect 580165 404774 584960 404776
rect 580165 404771 580231 404774
rect 583520 404684 584960 404774
rect 258073 402522 258139 402525
rect 261201 402522 261267 402525
rect 258073 402520 261267 402522
rect 258073 402464 258078 402520
rect 258134 402464 261206 402520
rect 261262 402464 261267 402520
rect 258073 402462 261267 402464
rect 258073 402459 258139 402462
rect 261201 402459 261267 402462
rect 231577 399394 231643 399397
rect 232957 399396 233023 399397
rect 237189 399396 237255 399397
rect 231710 399394 231716 399396
rect 231577 399392 231716 399394
rect 231577 399336 231582 399392
rect 231638 399336 231716 399392
rect 231577 399334 231716 399336
rect 231577 399331 231643 399334
rect 231710 399332 231716 399334
rect 231780 399332 231786 399396
rect 232957 399392 233004 399396
rect 233068 399394 233074 399396
rect 232957 399336 232962 399392
rect 232957 399332 233004 399336
rect 233068 399334 233114 399394
rect 237189 399392 237236 399396
rect 237300 399394 237306 399396
rect 237189 399336 237194 399392
rect 233068 399332 233074 399334
rect 237189 399332 237236 399336
rect 237300 399334 237346 399394
rect 237300 399332 237306 399334
rect 238150 399332 238156 399396
rect 238220 399394 238226 399396
rect 238293 399394 238359 399397
rect 238220 399392 238359 399394
rect 238220 399336 238298 399392
rect 238354 399336 238359 399392
rect 238220 399334 238359 399336
rect 238220 399332 238226 399334
rect 232957 399331 233023 399332
rect 237189 399331 237255 399332
rect 238293 399331 238359 399334
rect 242525 399394 242591 399397
rect 276841 399396 276907 399397
rect 242750 399394 242756 399396
rect 242525 399392 242756 399394
rect 242525 399336 242530 399392
rect 242586 399336 242756 399392
rect 242525 399334 242756 399336
rect 242525 399331 242591 399334
rect 242750 399332 242756 399334
rect 242820 399332 242826 399396
rect 276790 399394 276796 399396
rect 276750 399334 276796 399394
rect 276860 399392 276907 399396
rect 276902 399336 276907 399392
rect 276790 399332 276796 399334
rect 276860 399332 276907 399336
rect 282862 399332 282868 399396
rect 282932 399394 282938 399396
rect 283005 399394 283071 399397
rect 282932 399392 283071 399394
rect 282932 399336 283010 399392
rect 283066 399336 283071 399392
rect 282932 399334 283071 399336
rect 282932 399332 282938 399334
rect 276841 399331 276907 399332
rect 283005 399331 283071 399334
rect 284334 399332 284340 399396
rect 284404 399394 284410 399396
rect 284477 399394 284543 399397
rect 284404 399392 284543 399394
rect 284404 399336 284482 399392
rect 284538 399336 284543 399392
rect 284404 399334 284543 399336
rect 284404 399332 284410 399334
rect 284477 399331 284543 399334
rect 285622 399332 285628 399396
rect 285692 399394 285698 399396
rect 286133 399394 286199 399397
rect 287329 399396 287395 399397
rect 287881 399396 287947 399397
rect 287278 399394 287284 399396
rect 285692 399392 286199 399394
rect 285692 399336 286138 399392
rect 286194 399336 286199 399392
rect 285692 399334 286199 399336
rect 287238 399334 287284 399394
rect 287348 399392 287395 399396
rect 287830 399394 287836 399396
rect 287390 399336 287395 399392
rect 285692 399332 285698 399334
rect 286133 399331 286199 399334
rect 287278 399332 287284 399334
rect 287348 399332 287395 399336
rect 287790 399334 287836 399394
rect 287900 399392 287947 399396
rect 287942 399336 287947 399392
rect 287830 399332 287836 399334
rect 287900 399332 287947 399336
rect 287329 399331 287395 399332
rect 287881 399331 287947 399332
rect 225689 398714 225755 398717
rect 276790 398714 276796 398716
rect 225689 398712 276796 398714
rect 225689 398656 225694 398712
rect 225750 398656 276796 398712
rect 225689 398654 276796 398656
rect 225689 398651 225755 398654
rect 276790 398652 276796 398654
rect 276860 398652 276866 398716
rect 238150 398516 238156 398580
rect 238220 398578 238226 398580
rect 309777 398578 309843 398581
rect 238220 398576 309843 398578
rect 238220 398520 309782 398576
rect 309838 398520 309843 398576
rect 238220 398518 309843 398520
rect 238220 398516 238226 398518
rect 309777 398515 309843 398518
rect 242750 398380 242756 398444
rect 242820 398442 242826 398444
rect 326337 398442 326403 398445
rect 242820 398440 326403 398442
rect 242820 398384 326342 398440
rect 326398 398384 326403 398440
rect 242820 398382 326403 398384
rect 242820 398380 242826 398382
rect 326337 398379 326403 398382
rect 200757 398306 200823 398309
rect 287278 398306 287284 398308
rect 200757 398304 287284 398306
rect 200757 398248 200762 398304
rect 200818 398248 287284 398304
rect 200757 398246 287284 398248
rect 200757 398243 200823 398246
rect 287278 398244 287284 398246
rect 287348 398244 287354 398308
rect 197997 398170 198063 398173
rect 287830 398170 287836 398172
rect 197997 398168 287836 398170
rect 197997 398112 198002 398168
rect 198058 398112 287836 398168
rect 197997 398110 287836 398112
rect 197997 398107 198063 398110
rect 287830 398108 287836 398110
rect 287900 398108 287906 398172
rect 17217 398034 17283 398037
rect 284334 398034 284340 398036
rect 17217 398032 284340 398034
rect 17217 397976 17222 398032
rect 17278 397976 284340 398032
rect 17217 397974 284340 397976
rect 17217 397971 17283 397974
rect 284334 397972 284340 397974
rect 284404 397972 284410 398036
rect -960 395042 480 395132
rect 3141 395042 3207 395045
rect -960 395040 3207 395042
rect -960 394984 3146 395040
rect 3202 394984 3207 395040
rect -960 394982 3207 394984
rect -960 394892 480 394982
rect 3141 394979 3207 394982
rect 579797 393002 579863 393005
rect 583520 393002 584960 393092
rect 579797 393000 584960 393002
rect 579797 392944 579802 393000
rect 579858 392944 584960 393000
rect 579797 392942 584960 392944
rect 579797 392939 579863 392942
rect 583520 392852 584960 392942
rect 583520 381156 584960 381396
rect -960 380626 480 380716
rect 3417 380626 3483 380629
rect -960 380624 3483 380626
rect -960 380568 3422 380624
rect 3478 380568 3483 380624
rect -960 380566 3483 380568
rect -960 380476 480 380566
rect 3417 380563 3483 380566
rect 580165 369610 580231 369613
rect 583520 369610 584960 369700
rect 580165 369608 584960 369610
rect 580165 369552 580170 369608
rect 580226 369552 584960 369608
rect 580165 369550 584960 369552
rect 580165 369547 580231 369550
rect 583520 369460 584960 369550
rect -960 366210 480 366300
rect 2957 366210 3023 366213
rect -960 366208 3023 366210
rect -960 366152 2962 366208
rect 3018 366152 3023 366208
rect -960 366150 3023 366152
rect -960 366060 480 366150
rect 2957 366147 3023 366150
rect 580073 357914 580139 357917
rect 583520 357914 584960 358004
rect 580073 357912 584960 357914
rect 580073 357856 580078 357912
rect 580134 357856 584960 357912
rect 580073 357854 584960 357856
rect 580073 357851 580139 357854
rect 583520 357764 584960 357854
rect -960 351780 480 352020
rect 579797 346082 579863 346085
rect 583520 346082 584960 346172
rect 579797 346080 584960 346082
rect 579797 346024 579802 346080
rect 579858 346024 584960 346080
rect 579797 346022 584960 346024
rect 579797 346019 579863 346022
rect 583520 345932 584960 346022
rect 282637 338058 282703 338061
rect 288065 338058 288131 338061
rect 282637 338056 288131 338058
rect 282637 338000 282642 338056
rect 282698 338000 288070 338056
rect 288126 338000 288131 338056
rect 282637 337998 288131 338000
rect 282637 337995 282703 337998
rect 288065 337995 288131 337998
rect 280797 337922 280863 337925
rect 289537 337922 289603 337925
rect 280797 337920 289603 337922
rect 280797 337864 280802 337920
rect 280858 337864 289542 337920
rect 289598 337864 289603 337920
rect 280797 337862 289603 337864
rect 280797 337859 280863 337862
rect 289537 337859 289603 337862
rect 289813 337922 289879 337925
rect 291101 337922 291167 337925
rect 289813 337920 291167 337922
rect 289813 337864 289818 337920
rect 289874 337864 291106 337920
rect 291162 337864 291167 337920
rect 289813 337862 291167 337864
rect 289813 337859 289879 337862
rect 291101 337859 291167 337862
rect 281901 337786 281967 337789
rect 287697 337786 287763 337789
rect 281901 337784 287763 337786
rect 281901 337728 281906 337784
rect 281962 337728 287702 337784
rect 287758 337728 287763 337784
rect 281901 337726 287763 337728
rect 281901 337723 281967 337726
rect 287697 337723 287763 337726
rect -960 337514 480 337604
rect 3417 337514 3483 337517
rect -960 337512 3483 337514
rect -960 337456 3422 337512
rect 3478 337456 3483 337512
rect -960 337454 3483 337456
rect -960 337364 480 337454
rect 3417 337451 3483 337454
rect 263685 337106 263751 337109
rect 267733 337106 267799 337109
rect 263685 337104 267799 337106
rect 263685 337048 263690 337104
rect 263746 337048 267738 337104
rect 267794 337048 267799 337104
rect 263685 337046 267799 337048
rect 263685 337043 263751 337046
rect 267733 337043 267799 337046
rect 273621 336970 273687 336973
rect 285213 336970 285279 336973
rect 285581 336970 285647 336973
rect 273621 336968 273730 336970
rect 273621 336912 273626 336968
rect 273682 336912 273730 336968
rect 273621 336907 273730 336912
rect 285213 336968 285647 336970
rect 285213 336912 285218 336968
rect 285274 336912 285586 336968
rect 285642 336912 285647 336968
rect 285213 336910 285647 336912
rect 285213 336907 285279 336910
rect 285581 336907 285647 336910
rect 273670 336834 273730 336907
rect 273805 336834 273871 336837
rect 273670 336832 273871 336834
rect 273670 336776 273810 336832
rect 273866 336776 273871 336832
rect 273670 336774 273871 336776
rect 273805 336771 273871 336774
rect 277025 335610 277091 335613
rect 277025 335608 277226 335610
rect 277025 335552 277030 335608
rect 277086 335552 277226 335608
rect 277025 335550 277226 335552
rect 277025 335547 277091 335550
rect 277166 335372 277226 335550
rect 277301 335372 277367 335375
rect 277166 335370 277367 335372
rect 277166 335314 277306 335370
rect 277362 335314 277367 335370
rect 277166 335312 277367 335314
rect 277301 335309 277367 335312
rect 583520 334236 584960 334476
rect 307753 333808 307819 333811
rect 307710 333806 307819 333808
rect 307710 333750 307758 333806
rect 307814 333750 307819 333806
rect 307710 333745 307819 333750
rect 307710 333573 307770 333745
rect 307710 333568 307819 333573
rect 307710 333512 307758 333568
rect 307814 333512 307819 333568
rect 307710 333510 307819 333512
rect 307753 333507 307819 333510
rect 260373 324322 260439 324325
rect 260649 324322 260715 324325
rect 260373 324320 260715 324322
rect 260373 324264 260378 324320
rect 260434 324264 260654 324320
rect 260710 324264 260715 324320
rect 260373 324262 260715 324264
rect 260373 324259 260439 324262
rect 260649 324259 260715 324262
rect 262397 324322 262463 324325
rect 262673 324322 262739 324325
rect 262397 324320 262739 324322
rect 262397 324264 262402 324320
rect 262458 324264 262678 324320
rect 262734 324264 262739 324320
rect 262397 324262 262739 324264
rect 262397 324259 262463 324262
rect 262673 324259 262739 324262
rect 277025 324322 277091 324325
rect 277393 324322 277459 324325
rect 277025 324320 277459 324322
rect 277025 324264 277030 324320
rect 277086 324264 277398 324320
rect 277454 324264 277459 324320
rect 277025 324262 277459 324264
rect 277025 324259 277091 324262
rect 277393 324259 277459 324262
rect -960 323098 480 323188
rect 3969 323098 4035 323101
rect -960 323096 4035 323098
rect -960 323040 3974 323096
rect 4030 323040 4035 323096
rect -960 323038 4035 323040
rect -960 322948 480 323038
rect 3969 323035 4035 323038
rect 580165 322690 580231 322693
rect 583520 322690 584960 322780
rect 580165 322688 584960 322690
rect 580165 322632 580170 322688
rect 580226 322632 584960 322688
rect 580165 322630 584960 322632
rect 580165 322627 580231 322630
rect 583520 322540 584960 322630
rect 254710 314604 254716 314668
rect 254780 314666 254786 314668
rect 254853 314666 254919 314669
rect 254780 314664 254919 314666
rect 254780 314608 254858 314664
rect 254914 314608 254919 314664
rect 254780 314606 254919 314608
rect 254780 314604 254786 314606
rect 254853 314603 254919 314606
rect 256417 314666 256483 314669
rect 256601 314666 256667 314669
rect 256417 314664 256667 314666
rect 256417 314608 256422 314664
rect 256478 314608 256606 314664
rect 256662 314608 256667 314664
rect 256417 314606 256667 314608
rect 256417 314603 256483 314606
rect 256601 314603 256667 314606
rect 580165 310858 580231 310861
rect 583520 310858 584960 310948
rect 580165 310856 584960 310858
rect 580165 310800 580170 310856
rect 580226 310800 584960 310856
rect 580165 310798 584960 310800
rect 580165 310795 580231 310798
rect 583520 310708 584960 310798
rect -960 308818 480 308908
rect 3417 308818 3483 308821
rect -960 308816 3483 308818
rect -960 308760 3422 308816
rect 3478 308760 3483 308816
rect -960 308758 3483 308760
rect -960 308668 480 308758
rect 3417 308755 3483 308758
rect 264237 306370 264303 306373
rect 264421 306370 264487 306373
rect 264237 306368 264487 306370
rect 264237 306312 264242 306368
rect 264298 306312 264426 306368
rect 264482 306312 264487 306368
rect 264237 306310 264487 306312
rect 264237 306307 264303 306310
rect 264421 306307 264487 306310
rect 254761 305012 254827 305013
rect 254710 304948 254716 305012
rect 254780 305010 254827 305012
rect 256417 305010 256483 305013
rect 256601 305010 256667 305013
rect 254780 305008 254872 305010
rect 254822 304952 254872 305008
rect 254780 304950 254872 304952
rect 256417 305008 256667 305010
rect 256417 304952 256422 305008
rect 256478 304952 256606 305008
rect 256662 304952 256667 305008
rect 256417 304950 256667 304952
rect 254780 304948 254827 304950
rect 254761 304947 254827 304948
rect 256417 304947 256483 304950
rect 256601 304947 256667 304950
rect 579797 299162 579863 299165
rect 583520 299162 584960 299252
rect 579797 299160 584960 299162
rect 579797 299104 579802 299160
rect 579858 299104 584960 299160
rect 579797 299102 584960 299104
rect 579797 299099 579863 299102
rect 583520 299012 584960 299102
rect 254853 295354 254919 295357
rect 255037 295354 255103 295357
rect 254853 295352 255103 295354
rect 254853 295296 254858 295352
rect 254914 295296 255042 295352
rect 255098 295296 255103 295352
rect 254853 295294 255103 295296
rect 254853 295291 254919 295294
rect 255037 295291 255103 295294
rect 271597 295354 271663 295357
rect 271781 295354 271847 295357
rect 271597 295352 271847 295354
rect 271597 295296 271602 295352
rect 271658 295296 271786 295352
rect 271842 295296 271847 295352
rect 271597 295294 271847 295296
rect 271597 295291 271663 295294
rect 271781 295291 271847 295294
rect -960 294402 480 294492
rect 3049 294402 3115 294405
rect -960 294400 3115 294402
rect -960 294344 3054 294400
rect 3110 294344 3115 294400
rect -960 294342 3115 294344
rect -960 294252 480 294342
rect 3049 294339 3115 294342
rect 255630 289036 255636 289100
rect 255700 289098 255706 289100
rect 255773 289098 255839 289101
rect 255700 289096 255839 289098
rect 255700 289040 255778 289096
rect 255834 289040 255839 289096
rect 255700 289038 255839 289040
rect 255700 289036 255706 289038
rect 255773 289035 255839 289038
rect 583520 287316 584960 287556
rect 256417 285698 256483 285701
rect 256601 285698 256667 285701
rect 256417 285696 256667 285698
rect 256417 285640 256422 285696
rect 256478 285640 256606 285696
rect 256662 285640 256667 285696
rect 256417 285638 256667 285640
rect 256417 285635 256483 285638
rect 256601 285635 256667 285638
rect -960 280122 480 280212
rect 3785 280122 3851 280125
rect -960 280120 3851 280122
rect -960 280064 3790 280120
rect 3846 280064 3851 280120
rect -960 280062 3851 280064
rect -960 279972 480 280062
rect 3785 280059 3851 280062
rect 250253 280122 250319 280125
rect 250437 280122 250503 280125
rect 250253 280120 250503 280122
rect 250253 280064 250258 280120
rect 250314 280064 250442 280120
rect 250498 280064 250503 280120
rect 250253 280062 250503 280064
rect 250253 280059 250319 280062
rect 250437 280059 250503 280062
rect 255630 275980 255636 276044
rect 255700 276042 255706 276044
rect 255773 276042 255839 276045
rect 255700 276040 255839 276042
rect 255700 275984 255778 276040
rect 255834 275984 255839 276040
rect 255700 275982 255839 275984
rect 255700 275980 255706 275982
rect 255773 275979 255839 275982
rect 276841 276042 276907 276045
rect 277025 276042 277091 276045
rect 276841 276040 277091 276042
rect 276841 275984 276846 276040
rect 276902 275984 277030 276040
rect 277086 275984 277091 276040
rect 276841 275982 277091 275984
rect 276841 275979 276907 275982
rect 277025 275979 277091 275982
rect 580165 275770 580231 275773
rect 583520 275770 584960 275860
rect 580165 275768 584960 275770
rect 580165 275712 580170 275768
rect 580226 275712 584960 275768
rect 580165 275710 584960 275712
rect 580165 275707 580231 275710
rect 583520 275620 584960 275710
rect 260649 266522 260715 266525
rect 260606 266520 260715 266522
rect 260606 266464 260654 266520
rect 260710 266464 260715 266520
rect 260606 266459 260715 266464
rect 260606 266389 260666 266459
rect 260606 266384 260715 266389
rect 260606 266328 260654 266384
rect 260710 266328 260715 266384
rect 260606 266326 260715 266328
rect 260649 266323 260715 266326
rect -960 265706 480 265796
rect 2865 265706 2931 265709
rect -960 265704 2931 265706
rect -960 265648 2870 265704
rect 2926 265648 2931 265704
rect -960 265646 2931 265648
rect -960 265556 480 265646
rect 2865 265643 2931 265646
rect 580165 263938 580231 263941
rect 583520 263938 584960 264028
rect 580165 263936 584960 263938
rect 580165 263880 580170 263936
rect 580226 263880 584960 263936
rect 580165 263878 584960 263880
rect 580165 263875 580231 263878
rect 583520 263788 584960 263878
rect 250713 261082 250779 261085
rect 250302 261080 250779 261082
rect 250302 261024 250718 261080
rect 250774 261024 250779 261080
rect 250302 261022 250779 261024
rect 250302 260946 250362 261022
rect 250713 261019 250779 261022
rect 250437 260946 250503 260949
rect 250302 260944 250503 260946
rect 250302 260888 250442 260944
rect 250498 260888 250503 260944
rect 250302 260886 250503 260888
rect 250437 260883 250503 260886
rect 256969 259450 257035 259453
rect 257153 259450 257219 259453
rect 256969 259448 257219 259450
rect 256969 259392 256974 259448
rect 257030 259392 257158 259448
rect 257214 259392 257219 259448
rect 256969 259390 257219 259392
rect 256969 259387 257035 259390
rect 257153 259387 257219 259390
rect 579797 252242 579863 252245
rect 583520 252242 584960 252332
rect 579797 252240 584960 252242
rect 579797 252184 579802 252240
rect 579858 252184 584960 252240
rect 579797 252182 584960 252184
rect 579797 252179 579863 252182
rect 583520 252092 584960 252182
rect -960 251290 480 251380
rect 3417 251290 3483 251293
rect -960 251288 3483 251290
rect -960 251232 3422 251288
rect 3478 251232 3483 251288
rect -960 251230 3483 251232
rect -960 251140 480 251230
rect 3417 251227 3483 251230
rect 229553 241498 229619 241501
rect 229829 241498 229895 241501
rect 229553 241496 229895 241498
rect 229553 241440 229558 241496
rect 229614 241440 229834 241496
rect 229890 241440 229895 241496
rect 229553 241438 229895 241440
rect 229553 241435 229619 241438
rect 229829 241435 229895 241438
rect 234981 241498 235047 241501
rect 235165 241498 235231 241501
rect 234981 241496 235231 241498
rect 234981 241440 234986 241496
rect 235042 241440 235170 241496
rect 235226 241440 235231 241496
rect 234981 241438 235231 241440
rect 234981 241435 235047 241438
rect 235165 241435 235231 241438
rect 235533 241498 235599 241501
rect 235717 241498 235783 241501
rect 235533 241496 235783 241498
rect 235533 241440 235538 241496
rect 235594 241440 235722 241496
rect 235778 241440 235783 241496
rect 235533 241438 235783 241440
rect 235533 241435 235599 241438
rect 235717 241435 235783 241438
rect 583520 240396 584960 240636
rect 262489 237418 262555 237421
rect 262673 237418 262739 237421
rect 262489 237416 262739 237418
rect 262489 237360 262494 237416
rect 262550 237360 262678 237416
rect 262734 237360 262739 237416
rect 262489 237358 262739 237360
rect 262489 237355 262555 237358
rect 262673 237355 262739 237358
rect -960 237010 480 237100
rect 3601 237010 3667 237013
rect -960 237008 3667 237010
rect -960 236952 3606 237008
rect 3662 236952 3667 237008
rect -960 236950 3667 236952
rect -960 236860 480 236950
rect 3601 236947 3667 236950
rect 257245 229122 257311 229125
rect 257110 229120 257311 229122
rect 257110 229064 257250 229120
rect 257306 229064 257311 229120
rect 257110 229062 257311 229064
rect 257110 228986 257170 229062
rect 257245 229059 257311 229062
rect 257245 228986 257311 228989
rect 257110 228984 257311 228986
rect 257110 228928 257250 228984
rect 257306 228928 257311 228984
rect 257110 228926 257311 228928
rect 257245 228923 257311 228926
rect 583520 228850 584960 228940
rect 583342 228790 584960 228850
rect 248413 228034 248479 228037
rect 266261 228034 266327 228037
rect 328453 228034 328519 228037
rect 248413 228032 266327 228034
rect 248413 227976 248418 228032
rect 248474 227976 266266 228032
rect 266322 227976 266327 228032
rect 248413 227974 266327 227976
rect 248413 227971 248479 227974
rect 266261 227971 266327 227974
rect 328318 228032 328519 228034
rect 328318 227976 328458 228032
rect 328514 227976 328519 228032
rect 328318 227974 328519 227976
rect 237230 227836 237236 227900
rect 237300 227898 237306 227900
rect 248413 227898 248479 227901
rect 302141 227898 302207 227901
rect 237300 227896 248479 227898
rect 237300 227840 248418 227896
rect 248474 227840 248479 227896
rect 237300 227838 248479 227840
rect 237300 227836 237306 227838
rect 248413 227835 248479 227838
rect 292622 227896 302207 227898
rect 292622 227840 302146 227896
rect 302202 227840 302207 227896
rect 292622 227838 302207 227840
rect 255773 227762 255839 227765
rect 256049 227762 256115 227765
rect 255773 227760 256115 227762
rect 255773 227704 255778 227760
rect 255834 227704 256054 227760
rect 256110 227704 256115 227760
rect 255773 227702 256115 227704
rect 255773 227699 255839 227702
rect 256049 227699 256115 227702
rect 260557 227762 260623 227765
rect 260741 227762 260807 227765
rect 260557 227760 260807 227762
rect 260557 227704 260562 227760
rect 260618 227704 260746 227760
rect 260802 227704 260807 227760
rect 260557 227702 260807 227704
rect 260557 227699 260623 227702
rect 260741 227699 260807 227702
rect 266261 227762 266327 227765
rect 278681 227762 278747 227765
rect 266261 227760 278747 227762
rect 266261 227704 266266 227760
rect 266322 227704 278686 227760
rect 278742 227704 278747 227760
rect 266261 227702 278747 227704
rect 266261 227699 266327 227702
rect 278681 227699 278747 227702
rect 289721 227762 289787 227765
rect 292622 227762 292682 227838
rect 302141 227835 302207 227838
rect 312629 227898 312695 227901
rect 318742 227898 318748 227900
rect 312629 227896 318748 227898
rect 312629 227840 312634 227896
rect 312690 227840 318748 227896
rect 312629 227838 318748 227840
rect 312629 227835 312695 227838
rect 318742 227836 318748 227838
rect 318812 227836 318818 227900
rect 323577 227898 323643 227901
rect 328318 227898 328378 227974
rect 328453 227971 328519 227974
rect 338062 227972 338068 228036
rect 338132 228034 338138 228036
rect 418061 228034 418127 228037
rect 338132 227974 354690 228034
rect 338132 227972 338138 227974
rect 323577 227896 328378 227898
rect 323577 227840 323582 227896
rect 323638 227840 328378 227896
rect 323577 227838 328378 227840
rect 354630 227898 354690 227974
rect 364382 227974 374010 228034
rect 354630 227838 364258 227898
rect 323577 227835 323643 227838
rect 309133 227762 309199 227765
rect 338062 227762 338068 227764
rect 289721 227760 292682 227762
rect 289721 227704 289726 227760
rect 289782 227704 292682 227760
rect 289721 227702 292682 227704
rect 308998 227760 309199 227762
rect 308998 227704 309138 227760
rect 309194 227704 309199 227760
rect 308998 227702 309199 227704
rect 289721 227699 289787 227702
rect 302141 227490 302207 227493
rect 308998 227490 309058 227702
rect 309133 227699 309199 227702
rect 331446 227702 338068 227762
rect 318742 227564 318748 227628
rect 318812 227626 318818 227628
rect 323577 227626 323643 227629
rect 318812 227624 323643 227626
rect 318812 227568 323582 227624
rect 323638 227568 323643 227624
rect 318812 227566 323643 227568
rect 318812 227564 318818 227566
rect 323577 227563 323643 227566
rect 328545 227626 328611 227629
rect 331446 227626 331506 227702
rect 338062 227700 338068 227702
rect 338132 227700 338138 227764
rect 364198 227762 364258 227838
rect 364382 227762 364442 227974
rect 373950 227898 374010 227974
rect 383702 227974 408234 228034
rect 373950 227838 383578 227898
rect 364198 227702 364442 227762
rect 383518 227762 383578 227838
rect 383702 227762 383762 227974
rect 408174 227898 408234 227974
rect 415350 228032 418127 228034
rect 415350 227976 418066 228032
rect 418122 227976 418127 228032
rect 415350 227974 418127 227976
rect 415350 227898 415410 227974
rect 418061 227971 418127 227974
rect 424961 228034 425027 228037
rect 424961 228032 427738 228034
rect 424961 227976 424966 228032
rect 425022 227976 427738 228032
rect 424961 227974 427738 227976
rect 424961 227971 425027 227974
rect 408174 227838 415410 227898
rect 383518 227702 383762 227762
rect 427678 227762 427738 227974
rect 437381 227898 437447 227901
rect 456701 227898 456767 227901
rect 427862 227896 437447 227898
rect 427862 227840 437386 227896
rect 437442 227840 437447 227896
rect 427862 227838 437447 227840
rect 427862 227762 427922 227838
rect 437381 227835 437447 227838
rect 447182 227896 456767 227898
rect 447182 227840 456706 227896
rect 456762 227840 456767 227896
rect 447182 227838 456767 227840
rect 427678 227702 427922 227762
rect 444281 227762 444347 227765
rect 447182 227762 447242 227838
rect 456701 227835 456767 227838
rect 456885 227898 456951 227901
rect 476021 227898 476087 227901
rect 495341 227898 495407 227901
rect 456885 227896 466378 227898
rect 456885 227840 456890 227896
rect 456946 227840 466378 227896
rect 456885 227838 466378 227840
rect 456885 227835 456951 227838
rect 444281 227760 447242 227762
rect 444281 227704 444286 227760
rect 444342 227704 447242 227760
rect 444281 227702 447242 227704
rect 466318 227762 466378 227838
rect 466502 227896 476087 227898
rect 466502 227840 476026 227896
rect 476082 227840 476087 227896
rect 466502 227838 476087 227840
rect 466502 227762 466562 227838
rect 476021 227835 476087 227838
rect 485822 227896 495407 227898
rect 485822 227840 495346 227896
rect 495402 227840 495407 227896
rect 485822 227838 495407 227840
rect 466318 227702 466562 227762
rect 482921 227762 482987 227765
rect 485822 227762 485882 227838
rect 495341 227835 495407 227838
rect 496997 227898 497063 227901
rect 514661 227898 514727 227901
rect 533981 227898 534047 227901
rect 553301 227898 553367 227901
rect 496997 227896 505018 227898
rect 496997 227840 497002 227896
rect 497058 227840 505018 227896
rect 496997 227838 505018 227840
rect 496997 227835 497063 227838
rect 482921 227760 485882 227762
rect 482921 227704 482926 227760
rect 482982 227704 485882 227760
rect 482921 227702 485882 227704
rect 504958 227762 505018 227838
rect 505142 227896 514727 227898
rect 505142 227840 514666 227896
rect 514722 227840 514727 227896
rect 505142 227838 514727 227840
rect 505142 227762 505202 227838
rect 514661 227835 514727 227838
rect 524462 227896 534047 227898
rect 524462 227840 533986 227896
rect 534042 227840 534047 227896
rect 524462 227838 534047 227840
rect 504958 227702 505202 227762
rect 521561 227762 521627 227765
rect 524462 227762 524522 227838
rect 533981 227835 534047 227838
rect 543782 227896 553367 227898
rect 543782 227840 553306 227896
rect 553362 227840 553367 227896
rect 543782 227838 553367 227840
rect 521561 227760 524522 227762
rect 521561 227704 521566 227760
rect 521622 227704 524522 227760
rect 521561 227702 524522 227704
rect 540881 227762 540947 227765
rect 543782 227762 543842 227838
rect 553301 227835 553367 227838
rect 554589 227898 554655 227901
rect 583342 227898 583402 228790
rect 583520 228700 584960 228790
rect 554589 227896 562978 227898
rect 554589 227840 554594 227896
rect 554650 227840 562978 227896
rect 554589 227838 562978 227840
rect 554589 227835 554655 227838
rect 540881 227760 543842 227762
rect 540881 227704 540886 227760
rect 540942 227704 543842 227760
rect 540881 227702 543842 227704
rect 562918 227762 562978 227838
rect 576902 227838 583402 227898
rect 576902 227762 576962 227838
rect 562918 227702 576962 227762
rect 444281 227699 444347 227702
rect 482921 227699 482987 227702
rect 521561 227699 521627 227702
rect 540881 227699 540947 227702
rect 328545 227624 331506 227626
rect 328545 227568 328550 227624
rect 328606 227568 331506 227624
rect 328545 227566 331506 227568
rect 328545 227563 328611 227566
rect 302141 227488 309058 227490
rect 302141 227432 302146 227488
rect 302202 227432 309058 227488
rect 302141 227430 309058 227432
rect 302141 227427 302207 227430
rect -960 222594 480 222684
rect 3141 222594 3207 222597
rect -960 222592 3207 222594
rect -960 222536 3146 222592
rect 3202 222536 3207 222592
rect -960 222534 3207 222536
rect -960 222444 480 222534
rect 3141 222531 3207 222534
rect 229553 222186 229619 222189
rect 229829 222186 229895 222189
rect 229553 222184 229895 222186
rect 229553 222128 229558 222184
rect 229614 222128 229834 222184
rect 229890 222128 229895 222184
rect 229553 222126 229895 222128
rect 229553 222123 229619 222126
rect 229829 222123 229895 222126
rect 245009 222186 245075 222189
rect 245193 222186 245259 222189
rect 245009 222184 245259 222186
rect 245009 222128 245014 222184
rect 245070 222128 245198 222184
rect 245254 222128 245259 222184
rect 245009 222126 245259 222128
rect 245009 222123 245075 222126
rect 245193 222123 245259 222126
rect 234981 220826 235047 220829
rect 235165 220826 235231 220829
rect 234981 220824 235231 220826
rect 234981 220768 234986 220824
rect 235042 220768 235170 220824
rect 235226 220768 235231 220824
rect 234981 220766 235231 220768
rect 234981 220763 235047 220766
rect 235165 220763 235231 220766
rect 235533 220826 235599 220829
rect 235717 220826 235783 220829
rect 235533 220824 235783 220826
rect 235533 220768 235538 220824
rect 235594 220768 235722 220824
rect 235778 220768 235783 220824
rect 235533 220766 235783 220768
rect 235533 220763 235599 220766
rect 235717 220763 235783 220766
rect 580165 217018 580231 217021
rect 583520 217018 584960 217108
rect 580165 217016 584960 217018
rect 580165 216960 580170 217016
rect 580226 216960 584960 217016
rect 580165 216958 584960 216960
rect 580165 216955 580231 216958
rect 583520 216868 584960 216958
rect 277577 212530 277643 212533
rect 277761 212530 277827 212533
rect 277577 212528 277827 212530
rect 277577 212472 277582 212528
rect 277638 212472 277766 212528
rect 277822 212472 277827 212528
rect 277577 212470 277827 212472
rect 277577 212467 277643 212470
rect 277761 212467 277827 212470
rect 234981 211170 235047 211173
rect 235165 211170 235231 211173
rect 234981 211168 235231 211170
rect 234981 211112 234986 211168
rect 235042 211112 235170 211168
rect 235226 211112 235231 211168
rect 234981 211110 235231 211112
rect 234981 211107 235047 211110
rect 235165 211107 235231 211110
rect 235533 211170 235599 211173
rect 235717 211170 235783 211173
rect 235533 211168 235783 211170
rect 235533 211112 235538 211168
rect 235594 211112 235722 211168
rect 235778 211112 235783 211168
rect 235533 211110 235783 211112
rect 235533 211107 235599 211110
rect 235717 211107 235783 211110
rect 260925 208450 260991 208453
rect 260790 208448 260991 208450
rect 260790 208392 260930 208448
rect 260986 208392 260991 208448
rect 260790 208390 260991 208392
rect 260790 208317 260850 208390
rect 260925 208387 260991 208390
rect 260741 208312 260850 208317
rect -960 208178 480 208268
rect 260741 208256 260746 208312
rect 260802 208256 260850 208312
rect 260741 208254 260850 208256
rect 260741 208251 260807 208254
rect 3417 208178 3483 208181
rect -960 208176 3483 208178
rect -960 208120 3422 208176
rect 3478 208120 3483 208176
rect -960 208118 3483 208120
rect -960 208028 480 208118
rect 3417 208115 3483 208118
rect 579797 205322 579863 205325
rect 583520 205322 584960 205412
rect 579797 205320 584960 205322
rect 579797 205264 579802 205320
rect 579858 205264 584960 205320
rect 579797 205262 584960 205264
rect 579797 205259 579863 205262
rect 583520 205172 584960 205262
rect 229553 202874 229619 202877
rect 229829 202874 229895 202877
rect 229553 202872 229895 202874
rect 229553 202816 229558 202872
rect 229614 202816 229834 202872
rect 229890 202816 229895 202872
rect 229553 202814 229895 202816
rect 229553 202811 229619 202814
rect 229829 202811 229895 202814
rect 245009 202874 245075 202877
rect 245193 202874 245259 202877
rect 245009 202872 245259 202874
rect 245009 202816 245014 202872
rect 245070 202816 245198 202872
rect 245254 202816 245259 202872
rect 245009 202814 245259 202816
rect 245009 202811 245075 202814
rect 245193 202811 245259 202814
rect 3325 194578 3391 194581
rect 282862 194578 282868 194580
rect 3325 194576 282868 194578
rect 3325 194520 3330 194576
rect 3386 194520 282868 194576
rect 3325 194518 282868 194520
rect 3325 194515 3391 194518
rect 282862 194516 282868 194518
rect 282932 194516 282938 194580
rect -960 193898 480 193988
rect 3325 193898 3391 193901
rect -960 193896 3391 193898
rect -960 193840 3330 193896
rect 3386 193840 3391 193896
rect -960 193838 3391 193840
rect -960 193748 480 193838
rect 3325 193835 3391 193838
rect 583520 193476 584960 193716
rect 256417 193218 256483 193221
rect 256601 193218 256667 193221
rect 256417 193216 256667 193218
rect 256417 193160 256422 193216
rect 256478 193160 256606 193216
rect 256662 193160 256667 193216
rect 256417 193158 256667 193160
rect 256417 193155 256483 193158
rect 256601 193155 256667 193158
rect 268837 190498 268903 190501
rect 269021 190498 269087 190501
rect 268837 190496 269087 190498
rect 268837 190440 268842 190496
rect 268898 190440 269026 190496
rect 269082 190440 269087 190496
rect 268837 190438 269087 190440
rect 268837 190435 268903 190438
rect 269021 190435 269087 190438
rect 259913 189138 259979 189141
rect 259732 189136 259979 189138
rect 259732 189080 259918 189136
rect 259974 189080 259979 189136
rect 259732 189078 259979 189080
rect 259732 189005 259792 189078
rect 259913 189075 259979 189078
rect 259729 189000 259795 189005
rect 259729 188944 259734 189000
rect 259790 188944 259795 189000
rect 259729 188939 259795 188944
rect 229553 183562 229619 183565
rect 229829 183562 229895 183565
rect 229553 183560 229895 183562
rect 229553 183504 229558 183560
rect 229614 183504 229834 183560
rect 229890 183504 229895 183560
rect 229553 183502 229895 183504
rect 229553 183499 229619 183502
rect 229829 183499 229895 183502
rect 234981 183562 235047 183565
rect 235165 183562 235231 183565
rect 234981 183560 235231 183562
rect 234981 183504 234986 183560
rect 235042 183504 235170 183560
rect 235226 183504 235231 183560
rect 234981 183502 235231 183504
rect 234981 183499 235047 183502
rect 235165 183499 235231 183502
rect 245009 183562 245075 183565
rect 245193 183562 245259 183565
rect 245009 183560 245259 183562
rect 245009 183504 245014 183560
rect 245070 183504 245198 183560
rect 245254 183504 245259 183560
rect 245009 183502 245259 183504
rect 245009 183499 245075 183502
rect 245193 183499 245259 183502
rect 580165 181930 580231 181933
rect 583520 181930 584960 182020
rect 580165 181928 584960 181930
rect 580165 181872 580170 181928
rect 580226 181872 584960 181928
rect 580165 181870 584960 181872
rect 580165 181867 580231 181870
rect 583520 181780 584960 181870
rect -960 179482 480 179572
rect 3233 179482 3299 179485
rect -960 179480 3299 179482
rect -960 179424 3238 179480
rect 3294 179424 3299 179480
rect -960 179422 3299 179424
rect -960 179332 480 179422
rect 3233 179419 3299 179422
rect 260649 177986 260715 177989
rect 260833 177986 260899 177989
rect 260649 177984 260899 177986
rect 260649 177928 260654 177984
rect 260710 177928 260838 177984
rect 260894 177928 260899 177984
rect 260649 177926 260899 177928
rect 260649 177923 260715 177926
rect 260833 177923 260899 177926
rect 580165 170098 580231 170101
rect 583520 170098 584960 170188
rect 580165 170096 584960 170098
rect 580165 170040 580170 170096
rect 580226 170040 584960 170096
rect 580165 170038 584960 170040
rect 580165 170035 580231 170038
rect 583520 169948 584960 170038
rect 260649 168466 260715 168469
rect 260833 168466 260899 168469
rect 260649 168464 260899 168466
rect 260649 168408 260654 168464
rect 260710 168408 260838 168464
rect 260894 168408 260899 168464
rect 260649 168406 260899 168408
rect 260649 168403 260715 168406
rect 260833 168403 260899 168406
rect -960 165066 480 165156
rect 3509 165066 3575 165069
rect -960 165064 3575 165066
rect -960 165008 3514 165064
rect 3570 165008 3575 165064
rect -960 165006 3575 165008
rect -960 164916 480 165006
rect 3509 165003 3575 165006
rect 257245 164250 257311 164253
rect 257429 164250 257495 164253
rect 257245 164248 257495 164250
rect 257245 164192 257250 164248
rect 257306 164192 257434 164248
rect 257490 164192 257495 164248
rect 257245 164190 257495 164192
rect 257245 164187 257311 164190
rect 257429 164187 257495 164190
rect 234981 162890 235047 162893
rect 235165 162890 235231 162893
rect 234981 162888 235231 162890
rect 234981 162832 234986 162888
rect 235042 162832 235170 162888
rect 235226 162832 235231 162888
rect 234981 162830 235231 162832
rect 234981 162827 235047 162830
rect 235165 162827 235231 162830
rect 579797 158402 579863 158405
rect 583520 158402 584960 158492
rect 579797 158400 584960 158402
rect 579797 158344 579802 158400
rect 579858 158344 584960 158400
rect 579797 158342 584960 158344
rect 579797 158339 579863 158342
rect 583520 158252 584960 158342
rect 229645 154594 229711 154597
rect 229829 154594 229895 154597
rect 229645 154592 229895 154594
rect 229645 154536 229650 154592
rect 229706 154536 229834 154592
rect 229890 154536 229895 154592
rect 229645 154534 229895 154536
rect 229645 154531 229711 154534
rect 229829 154531 229895 154534
rect 238753 153234 238819 153237
rect 238937 153234 239003 153237
rect 238753 153232 239003 153234
rect 238753 153176 238758 153232
rect 238814 153176 238942 153232
rect 238998 153176 239003 153232
rect 238753 153174 239003 153176
rect 238753 153171 238819 153174
rect 238937 153171 239003 153174
rect -960 150786 480 150876
rect 3141 150786 3207 150789
rect -960 150784 3207 150786
rect -960 150728 3146 150784
rect 3202 150728 3207 150784
rect -960 150726 3207 150728
rect -960 150636 480 150726
rect 3141 150723 3207 150726
rect 583520 146556 584960 146796
rect 238937 145074 239003 145077
rect 238894 145072 239003 145074
rect 238894 145016 238942 145072
rect 238998 145016 239003 145072
rect 238894 145011 239003 145016
rect 233785 144938 233851 144941
rect 233969 144938 234035 144941
rect 233785 144936 234035 144938
rect 233785 144880 233790 144936
rect 233846 144880 233974 144936
rect 234030 144880 234035 144936
rect 233785 144878 234035 144880
rect 233785 144875 233851 144878
rect 233969 144875 234035 144878
rect 238753 144802 238819 144805
rect 238894 144802 238954 145011
rect 238753 144800 238954 144802
rect 238753 144744 238758 144800
rect 238814 144744 238954 144800
rect 238753 144742 238954 144744
rect 238753 144739 238819 144742
rect 245009 143578 245075 143581
rect 245193 143578 245259 143581
rect 245009 143576 245259 143578
rect 245009 143520 245014 143576
rect 245070 143520 245198 143576
rect 245254 143520 245259 143576
rect 245009 143518 245259 143520
rect 245009 143515 245075 143518
rect 245193 143515 245259 143518
rect 250713 142354 250779 142357
rect 250486 142352 250779 142354
rect 250486 142296 250718 142352
rect 250774 142296 250779 142352
rect 250486 142294 250779 142296
rect 250486 142218 250546 142294
rect 250713 142291 250779 142294
rect 250621 142218 250687 142221
rect 250486 142216 250687 142218
rect 250486 142160 250626 142216
rect 250682 142160 250687 142216
rect 250486 142158 250687 142160
rect 250621 142155 250687 142158
rect -960 136370 480 136460
rect 3233 136370 3299 136373
rect -960 136368 3299 136370
rect -960 136312 3238 136368
rect 3294 136312 3299 136368
rect -960 136310 3299 136312
rect -960 136220 480 136310
rect 3233 136307 3299 136310
rect 229461 135282 229527 135285
rect 229645 135282 229711 135285
rect 229461 135280 229711 135282
rect 229461 135224 229466 135280
rect 229522 135224 229650 135280
rect 229706 135224 229711 135280
rect 229461 135222 229711 135224
rect 229461 135219 229527 135222
rect 229645 135219 229711 135222
rect 238753 135282 238819 135285
rect 238937 135282 239003 135285
rect 238753 135280 239003 135282
rect 238753 135224 238758 135280
rect 238814 135224 238942 135280
rect 238998 135224 239003 135280
rect 238753 135222 239003 135224
rect 238753 135219 238819 135222
rect 238937 135219 239003 135222
rect 580165 134874 580231 134877
rect 583520 134874 584960 134964
rect 580165 134872 584960 134874
rect 580165 134816 580170 134872
rect 580226 134816 584960 134872
rect 580165 134814 584960 134816
rect 580165 134811 580231 134814
rect 583520 134724 584960 134814
rect 238937 125762 239003 125765
rect 238894 125760 239003 125762
rect 238894 125704 238942 125760
rect 238998 125704 239003 125760
rect 238894 125699 239003 125704
rect 238753 125354 238819 125357
rect 238894 125354 238954 125699
rect 255865 125626 255931 125629
rect 256049 125626 256115 125629
rect 255865 125624 256115 125626
rect 255865 125568 255870 125624
rect 255926 125568 256054 125624
rect 256110 125568 256115 125624
rect 255865 125566 256115 125568
rect 255865 125563 255931 125566
rect 256049 125563 256115 125566
rect 238753 125352 238954 125354
rect 238753 125296 238758 125352
rect 238814 125296 238954 125352
rect 238753 125294 238954 125296
rect 238753 125291 238819 125294
rect 580165 123178 580231 123181
rect 583520 123178 584960 123268
rect 580165 123176 584960 123178
rect 580165 123120 580170 123176
rect 580226 123120 584960 123176
rect 580165 123118 584960 123120
rect 580165 123115 580231 123118
rect 583520 123028 584960 123118
rect -960 122090 480 122180
rect 3417 122090 3483 122093
rect -960 122088 3483 122090
rect -960 122032 3422 122088
rect 3478 122032 3483 122088
rect -960 122030 3483 122032
rect -960 121940 480 122030
rect 3417 122027 3483 122030
rect 229461 115970 229527 115973
rect 229645 115970 229711 115973
rect 229461 115968 229711 115970
rect 229461 115912 229466 115968
rect 229522 115912 229650 115968
rect 229706 115912 229711 115968
rect 229461 115910 229711 115912
rect 229461 115907 229527 115910
rect 229645 115907 229711 115910
rect 238753 115970 238819 115973
rect 238937 115970 239003 115973
rect 238753 115968 239003 115970
rect 238753 115912 238758 115968
rect 238814 115912 238942 115968
rect 238998 115912 239003 115968
rect 238753 115910 239003 115912
rect 238753 115907 238819 115910
rect 238937 115907 239003 115910
rect 579797 111482 579863 111485
rect 583520 111482 584960 111572
rect 579797 111480 584960 111482
rect 579797 111424 579802 111480
rect 579858 111424 584960 111480
rect 579797 111422 584960 111424
rect 579797 111419 579863 111422
rect 583520 111332 584960 111422
rect 3417 109034 3483 109037
rect 285622 109034 285628 109036
rect 3417 109032 285628 109034
rect 3417 108976 3422 109032
rect 3478 108976 285628 109032
rect 3417 108974 285628 108976
rect 3417 108971 3483 108974
rect 285622 108972 285628 108974
rect 285692 108972 285698 109036
rect -960 107674 480 107764
rect 3417 107674 3483 107677
rect -960 107672 3483 107674
rect -960 107616 3422 107672
rect 3478 107616 3483 107672
rect -960 107614 3483 107616
rect -960 107524 480 107614
rect 3417 107611 3483 107614
rect 255865 106314 255931 106317
rect 256049 106314 256115 106317
rect 255865 106312 256115 106314
rect 255865 106256 255870 106312
rect 255926 106256 256054 106312
rect 256110 106256 256115 106312
rect 255865 106254 256115 106256
rect 255865 106251 255931 106254
rect 256049 106251 256115 106254
rect 260557 100738 260623 100741
rect 276933 100738 276999 100741
rect 277209 100738 277275 100741
rect 260557 100736 260666 100738
rect 260557 100680 260562 100736
rect 260618 100680 260666 100736
rect 260557 100675 260666 100680
rect 276933 100736 277275 100738
rect 276933 100680 276938 100736
rect 276994 100680 277214 100736
rect 277270 100680 277275 100736
rect 276933 100678 277275 100680
rect 276933 100675 276999 100678
rect 277209 100675 277275 100678
rect 260606 100605 260666 100675
rect 260606 100600 260715 100605
rect 260606 100544 260654 100600
rect 260710 100544 260715 100600
rect 260606 100542 260715 100544
rect 260649 100539 260715 100542
rect 583520 99636 584960 99876
rect 229461 96658 229527 96661
rect 229645 96658 229711 96661
rect 229461 96656 229711 96658
rect 229461 96600 229466 96656
rect 229522 96600 229650 96656
rect 229706 96600 229711 96656
rect 229461 96598 229711 96600
rect 229461 96595 229527 96598
rect 229645 96595 229711 96598
rect -960 93258 480 93348
rect 3417 93258 3483 93261
rect -960 93256 3483 93258
rect -960 93200 3422 93256
rect 3478 93200 3483 93256
rect -960 93198 3483 93200
rect -960 93108 480 93198
rect 3417 93195 3483 93198
rect 254761 91082 254827 91085
rect 255037 91082 255103 91085
rect 254761 91080 255103 91082
rect 254761 91024 254766 91080
rect 254822 91024 255042 91080
rect 255098 91024 255103 91080
rect 254761 91022 255103 91024
rect 254761 91019 254827 91022
rect 255037 91019 255103 91022
rect 273805 91082 273871 91085
rect 274081 91082 274147 91085
rect 273805 91080 274147 91082
rect 273805 91024 273810 91080
rect 273866 91024 274086 91080
rect 274142 91024 274147 91080
rect 273805 91022 274147 91024
rect 273805 91019 273871 91022
rect 274081 91019 274147 91022
rect 580165 87954 580231 87957
rect 583520 87954 584960 88044
rect 580165 87952 584960 87954
rect 580165 87896 580170 87952
rect 580226 87896 584960 87952
rect 580165 87894 584960 87896
rect 580165 87891 580231 87894
rect 583520 87804 584960 87894
rect 235533 87138 235599 87141
rect 235398 87136 235599 87138
rect 235398 87080 235538 87136
rect 235594 87080 235599 87136
rect 235398 87078 235599 87080
rect 235398 87005 235458 87078
rect 235533 87075 235599 87078
rect 233785 87002 233851 87005
rect 233969 87002 234035 87005
rect 233785 87000 234035 87002
rect 233785 86944 233790 87000
rect 233846 86944 233974 87000
rect 234030 86944 234035 87000
rect 233785 86942 234035 86944
rect 235398 87000 235507 87005
rect 235398 86944 235446 87000
rect 235502 86944 235507 87000
rect 235398 86942 235507 86944
rect 233785 86939 233851 86942
rect 233969 86939 234035 86942
rect 235441 86939 235507 86942
rect 254853 80066 254919 80069
rect 255037 80066 255103 80069
rect 254853 80064 255103 80066
rect 254853 80008 254858 80064
rect 254914 80008 255042 80064
rect 255098 80008 255103 80064
rect 254853 80006 255103 80008
rect 254853 80003 254919 80006
rect 255037 80003 255103 80006
rect -960 78978 480 79068
rect 3417 78978 3483 78981
rect -960 78976 3483 78978
rect -960 78920 3422 78976
rect 3478 78920 3483 78976
rect -960 78918 3483 78920
rect -960 78828 480 78918
rect 3417 78915 3483 78918
rect 521561 76530 521627 76533
rect 511950 76528 521627 76530
rect 511950 76472 521566 76528
rect 521622 76472 521627 76528
rect 511950 76470 521627 76472
rect 232998 76196 233004 76260
rect 233068 76258 233074 76260
rect 328453 76258 328519 76261
rect 233068 76198 234538 76258
rect 233068 76196 233074 76198
rect 234478 75986 234538 76198
rect 234662 76198 246314 76258
rect 234662 75986 234722 76198
rect 234478 75926 234722 75986
rect 246254 75986 246314 76198
rect 328318 76256 328519 76258
rect 328318 76200 328458 76256
rect 328514 76200 328519 76256
rect 328318 76198 328519 76200
rect 302141 76122 302207 76125
rect 292622 76120 302207 76122
rect 292622 76064 302146 76120
rect 302202 76064 302207 76120
rect 292622 76062 302207 76064
rect 292622 75986 292682 76062
rect 302141 76059 302207 76062
rect 313917 76122 313983 76125
rect 318742 76122 318748 76124
rect 313917 76120 318748 76122
rect 313917 76064 313922 76120
rect 313978 76064 318748 76120
rect 313917 76062 318748 76064
rect 313917 76059 313983 76062
rect 318742 76060 318748 76062
rect 318812 76060 318818 76124
rect 323577 76122 323643 76125
rect 328318 76122 328378 76198
rect 328453 76195 328519 76198
rect 338062 76196 338068 76260
rect 338132 76258 338138 76260
rect 510521 76258 510587 76261
rect 511950 76258 512010 76470
rect 521561 76467 521627 76470
rect 583520 76258 584960 76348
rect 338132 76198 354690 76258
rect 338132 76196 338138 76198
rect 323577 76120 328378 76122
rect 323577 76064 323582 76120
rect 323638 76064 328378 76120
rect 323577 76062 328378 76064
rect 354630 76122 354690 76198
rect 364382 76198 374010 76258
rect 354630 76062 364258 76122
rect 323577 76059 323643 76062
rect 309133 75986 309199 75989
rect 338062 75986 338068 75988
rect 246254 75926 292682 75986
rect 308998 75984 309199 75986
rect 308998 75928 309138 75984
rect 309194 75928 309199 75984
rect 308998 75926 309199 75928
rect 302141 75714 302207 75717
rect 308998 75714 309058 75926
rect 309133 75923 309199 75926
rect 331446 75926 338068 75986
rect 318742 75788 318748 75852
rect 318812 75850 318818 75852
rect 323577 75850 323643 75853
rect 318812 75848 323643 75850
rect 318812 75792 323582 75848
rect 323638 75792 323643 75848
rect 318812 75790 323643 75792
rect 318812 75788 318818 75790
rect 323577 75787 323643 75790
rect 328545 75850 328611 75853
rect 331446 75850 331506 75926
rect 338062 75924 338068 75926
rect 338132 75924 338138 75988
rect 364198 75986 364258 76062
rect 364382 75986 364442 76198
rect 373950 76122 374010 76198
rect 383702 76198 405842 76258
rect 373950 76062 383578 76122
rect 364198 75926 364442 75986
rect 383518 75986 383578 76062
rect 383702 75986 383762 76198
rect 405782 76122 405842 76198
rect 510521 76256 512010 76258
rect 510521 76200 510526 76256
rect 510582 76200 512010 76256
rect 510521 76198 512010 76200
rect 583342 76198 584960 76258
rect 510521 76195 510587 76198
rect 415301 76122 415367 76125
rect 437381 76122 437447 76125
rect 456701 76122 456767 76125
rect 405782 76120 415367 76122
rect 405782 76064 415306 76120
rect 415362 76064 415367 76120
rect 405782 76062 415367 76064
rect 415301 76059 415367 76062
rect 427862 76120 437447 76122
rect 427862 76064 437386 76120
rect 437442 76064 437447 76120
rect 427862 76062 437447 76064
rect 383518 75926 383762 75986
rect 415301 75986 415367 75989
rect 427862 75986 427922 76062
rect 437381 76059 437447 76062
rect 447182 76120 456767 76122
rect 447182 76064 456706 76120
rect 456762 76064 456767 76120
rect 447182 76062 456767 76064
rect 415301 75984 427922 75986
rect 415301 75928 415306 75984
rect 415362 75928 427922 75984
rect 415301 75926 427922 75928
rect 444281 75986 444347 75989
rect 447182 75986 447242 76062
rect 456701 76059 456767 76062
rect 456885 76122 456951 76125
rect 482921 76122 482987 76125
rect 492622 76122 492628 76124
rect 456885 76120 466378 76122
rect 456885 76064 456890 76120
rect 456946 76064 466378 76120
rect 456885 76062 466378 76064
rect 456885 76059 456951 76062
rect 444281 75984 447242 75986
rect 444281 75928 444286 75984
rect 444342 75928 447242 75984
rect 444281 75926 447242 75928
rect 466318 75986 466378 76062
rect 466502 76120 482987 76122
rect 466502 76064 482926 76120
rect 482982 76064 482987 76120
rect 466502 76062 482987 76064
rect 466502 75986 466562 76062
rect 482921 76059 482987 76062
rect 483062 76062 492628 76122
rect 466318 75926 466562 75986
rect 482921 75986 482987 75989
rect 483062 75986 483122 76062
rect 492622 76060 492628 76062
rect 492692 76060 492698 76124
rect 533981 76122 534047 76125
rect 553301 76122 553367 76125
rect 524462 76120 534047 76122
rect 524462 76064 533986 76120
rect 534042 76064 534047 76120
rect 524462 76062 534047 76064
rect 482921 75984 483122 75986
rect 482921 75928 482926 75984
rect 482982 75928 483122 75984
rect 482921 75926 483122 75928
rect 521561 75986 521627 75989
rect 524462 75986 524522 76062
rect 533981 76059 534047 76062
rect 543782 76120 553367 76122
rect 543782 76064 553306 76120
rect 553362 76064 553367 76120
rect 543782 76062 553367 76064
rect 521561 75984 524522 75986
rect 521561 75928 521566 75984
rect 521622 75928 524522 75984
rect 521561 75926 524522 75928
rect 540881 75986 540947 75989
rect 543782 75986 543842 76062
rect 553301 76059 553367 76062
rect 554589 76122 554655 76125
rect 583342 76122 583402 76198
rect 554589 76120 562978 76122
rect 554589 76064 554594 76120
rect 554650 76064 562978 76120
rect 554589 76062 562978 76064
rect 554589 76059 554655 76062
rect 540881 75984 543842 75986
rect 540881 75928 540886 75984
rect 540942 75928 543842 75984
rect 540881 75926 543842 75928
rect 562918 75986 562978 76062
rect 576902 76062 583402 76122
rect 583520 76108 584960 76198
rect 576902 75986 576962 76062
rect 562918 75926 576962 75986
rect 415301 75923 415367 75926
rect 444281 75923 444347 75926
rect 482921 75923 482987 75926
rect 521561 75923 521627 75926
rect 540881 75923 540947 75926
rect 328545 75848 331506 75850
rect 328545 75792 328550 75848
rect 328606 75792 331506 75848
rect 328545 75790 331506 75792
rect 328545 75787 328611 75790
rect 492622 75788 492628 75852
rect 492692 75850 492698 75852
rect 502241 75850 502307 75853
rect 492692 75848 502307 75850
rect 492692 75792 502246 75848
rect 502302 75792 502307 75848
rect 492692 75790 502307 75792
rect 492692 75788 492698 75790
rect 502241 75787 502307 75790
rect 302141 75712 309058 75714
rect 302141 75656 302146 75712
rect 302202 75656 309058 75712
rect 302141 75654 309058 75656
rect 302141 75651 302207 75654
rect 259729 71770 259795 71773
rect 260097 71770 260163 71773
rect 259729 71768 260163 71770
rect 259729 71712 259734 71768
rect 259790 71712 260102 71768
rect 260158 71712 260163 71768
rect 259729 71710 260163 71712
rect 259729 71707 259795 71710
rect 260097 71707 260163 71710
rect 254853 70410 254919 70413
rect 255037 70410 255103 70413
rect 254853 70408 255103 70410
rect 254853 70352 254858 70408
rect 254914 70352 255042 70408
rect 255098 70352 255103 70408
rect 254853 70350 255103 70352
rect 254853 70347 254919 70350
rect 255037 70347 255103 70350
rect -960 64562 480 64652
rect 3325 64562 3391 64565
rect -960 64560 3391 64562
rect -960 64504 3330 64560
rect 3386 64504 3391 64560
rect -960 64502 3391 64504
rect -960 64412 480 64502
rect 3325 64499 3391 64502
rect 579797 64562 579863 64565
rect 583520 64562 584960 64652
rect 579797 64560 584960 64562
rect 579797 64504 579802 64560
rect 579858 64504 584960 64560
rect 579797 64502 584960 64504
rect 579797 64499 579863 64502
rect 583520 64412 584960 64502
rect 256969 62114 257035 62117
rect 257153 62114 257219 62117
rect 256969 62112 257219 62114
rect 256969 62056 256974 62112
rect 257030 62056 257158 62112
rect 257214 62056 257219 62112
rect 256969 62054 257219 62056
rect 256969 62051 257035 62054
rect 257153 62051 257219 62054
rect 583520 52716 584960 52956
rect -960 50146 480 50236
rect 3417 50146 3483 50149
rect -960 50144 3483 50146
rect -960 50088 3422 50144
rect 3478 50088 3483 50144
rect -960 50086 3483 50088
rect -960 49996 480 50086
rect 3417 50083 3483 50086
rect 250437 44162 250503 44165
rect 250713 44162 250779 44165
rect 250437 44160 250779 44162
rect 250437 44104 250442 44160
rect 250498 44104 250718 44160
rect 250774 44104 250779 44160
rect 250437 44102 250779 44104
rect 250437 44099 250503 44102
rect 250713 44099 250779 44102
rect 580165 41034 580231 41037
rect 583520 41034 584960 41124
rect 580165 41032 584960 41034
rect 580165 40976 580170 41032
rect 580226 40976 584960 41032
rect 580165 40974 584960 40976
rect 580165 40971 580231 40974
rect 583520 40884 584960 40974
rect -960 35866 480 35956
rect 3417 35866 3483 35869
rect -960 35864 3483 35866
rect -960 35808 3422 35864
rect 3478 35808 3483 35864
rect -960 35806 3483 35808
rect -960 35716 480 35806
rect 3417 35803 3483 35806
rect 236318 29414 251098 29474
rect 231710 29004 231716 29068
rect 231780 29066 231786 29068
rect 236318 29066 236378 29414
rect 231780 29006 236378 29066
rect 251038 29066 251098 29414
rect 405641 29338 405707 29341
rect 424961 29338 425027 29341
rect 444281 29338 444347 29341
rect 463601 29338 463667 29341
rect 482921 29338 482987 29341
rect 502241 29338 502307 29341
rect 521561 29338 521627 29341
rect 540881 29338 540947 29341
rect 560201 29338 560267 29341
rect 583520 29338 584960 29428
rect 302190 29278 321570 29338
rect 280245 29066 280311 29069
rect 251038 29064 280311 29066
rect 251038 29008 280250 29064
rect 280306 29008 280311 29064
rect 251038 29006 280311 29008
rect 231780 29004 231786 29006
rect 280245 29003 280311 29006
rect 289721 29066 289787 29069
rect 302190 29066 302250 29278
rect 321510 29202 321570 29278
rect 335310 29278 344938 29338
rect 321510 29142 331138 29202
rect 289721 29064 302250 29066
rect 289721 29008 289726 29064
rect 289782 29008 302250 29064
rect 289721 29006 302250 29008
rect 331078 29066 331138 29142
rect 335310 29066 335370 29278
rect 331078 29006 335370 29066
rect 344878 29066 344938 29278
rect 345062 29278 354690 29338
rect 345062 29066 345122 29278
rect 354630 29202 354690 29278
rect 364382 29278 374010 29338
rect 354630 29142 364258 29202
rect 344878 29006 345122 29066
rect 364198 29066 364258 29142
rect 364382 29066 364442 29278
rect 373950 29202 374010 29278
rect 383702 29278 389282 29338
rect 373950 29142 383578 29202
rect 364198 29006 364442 29066
rect 383518 29066 383578 29142
rect 383702 29066 383762 29278
rect 389222 29202 389282 29278
rect 405641 29336 408602 29338
rect 405641 29280 405646 29336
rect 405702 29280 408602 29336
rect 405641 29278 408602 29280
rect 405641 29275 405707 29278
rect 398097 29202 398163 29205
rect 389222 29200 398163 29202
rect 389222 29144 398102 29200
rect 398158 29144 398163 29200
rect 389222 29142 398163 29144
rect 408542 29202 408602 29278
rect 424961 29336 427922 29338
rect 424961 29280 424966 29336
rect 425022 29280 427922 29336
rect 424961 29278 427922 29280
rect 424961 29275 425027 29278
rect 417325 29202 417391 29205
rect 408542 29200 417391 29202
rect 408542 29144 417330 29200
rect 417386 29144 417391 29200
rect 408542 29142 417391 29144
rect 427862 29202 427922 29278
rect 444281 29336 447242 29338
rect 444281 29280 444286 29336
rect 444342 29280 447242 29336
rect 444281 29278 447242 29280
rect 444281 29275 444347 29278
rect 436737 29202 436803 29205
rect 427862 29200 436803 29202
rect 427862 29144 436742 29200
rect 436798 29144 436803 29200
rect 427862 29142 436803 29144
rect 447182 29202 447242 29278
rect 463601 29336 466562 29338
rect 463601 29280 463606 29336
rect 463662 29280 466562 29336
rect 463601 29278 466562 29280
rect 463601 29275 463667 29278
rect 456701 29202 456767 29205
rect 447182 29200 456767 29202
rect 447182 29144 456706 29200
rect 456762 29144 456767 29200
rect 447182 29142 456767 29144
rect 466502 29202 466562 29278
rect 482921 29336 485882 29338
rect 482921 29280 482926 29336
rect 482982 29280 485882 29336
rect 482921 29278 485882 29280
rect 482921 29275 482987 29278
rect 475285 29202 475351 29205
rect 466502 29200 475351 29202
rect 466502 29144 475290 29200
rect 475346 29144 475351 29200
rect 466502 29142 475351 29144
rect 485822 29202 485882 29278
rect 502241 29336 505202 29338
rect 502241 29280 502246 29336
rect 502302 29280 505202 29336
rect 502241 29278 505202 29280
rect 502241 29275 502307 29278
rect 495157 29202 495223 29205
rect 485822 29200 495223 29202
rect 485822 29144 495162 29200
rect 495218 29144 495223 29200
rect 485822 29142 495223 29144
rect 505142 29202 505202 29278
rect 521561 29336 524522 29338
rect 521561 29280 521566 29336
rect 521622 29280 524522 29336
rect 521561 29278 524522 29280
rect 521561 29275 521627 29278
rect 513557 29202 513623 29205
rect 505142 29200 513623 29202
rect 505142 29144 513562 29200
rect 513618 29144 513623 29200
rect 505142 29142 513623 29144
rect 524462 29202 524522 29278
rect 540881 29336 543842 29338
rect 540881 29280 540886 29336
rect 540942 29280 543842 29336
rect 540881 29278 543842 29280
rect 540881 29275 540947 29278
rect 533797 29202 533863 29205
rect 524462 29200 533863 29202
rect 524462 29144 533802 29200
rect 533858 29144 533863 29200
rect 524462 29142 533863 29144
rect 543782 29202 543842 29278
rect 560201 29336 572730 29338
rect 560201 29280 560206 29336
rect 560262 29280 572730 29336
rect 560201 29278 572730 29280
rect 560201 29275 560267 29278
rect 552473 29202 552539 29205
rect 543782 29200 552539 29202
rect 543782 29144 552478 29200
rect 552534 29144 552539 29200
rect 543782 29142 552539 29144
rect 398097 29139 398163 29142
rect 417325 29139 417391 29142
rect 436737 29139 436803 29142
rect 456701 29139 456767 29142
rect 475285 29139 475351 29142
rect 495157 29139 495223 29142
rect 513557 29139 513623 29142
rect 533797 29139 533863 29142
rect 552473 29139 552539 29142
rect 383518 29006 383762 29066
rect 572670 29066 572730 29278
rect 583342 29278 584960 29338
rect 583342 29066 583402 29278
rect 583520 29188 584960 29278
rect 572670 29006 583402 29066
rect 289721 29003 289787 29006
rect -960 21450 480 21540
rect 3141 21450 3207 21453
rect -960 21448 3207 21450
rect -960 21392 3146 21448
rect 3202 21392 3207 21448
rect -960 21390 3207 21392
rect -960 21300 480 21390
rect 3141 21387 3207 21390
rect 579797 17642 579863 17645
rect 583520 17642 584960 17732
rect 579797 17640 584960 17642
rect 579797 17584 579802 17640
rect 579858 17584 584960 17640
rect 579797 17582 584960 17584
rect 579797 17579 579863 17582
rect 583520 17492 584960 17582
rect -960 7170 480 7260
rect 3417 7170 3483 7173
rect -960 7168 3483 7170
rect -960 7112 3422 7168
rect 3478 7112 3483 7168
rect -960 7110 3483 7112
rect -960 7020 480 7110
rect 3417 7107 3483 7110
rect 583520 5796 584960 6036
rect 32673 4042 32739 4045
rect 233601 4042 233667 4045
rect 32673 4040 233667 4042
rect 32673 3984 32678 4040
rect 32734 3984 233606 4040
rect 233662 3984 233667 4040
rect 32673 3982 233667 3984
rect 32673 3979 32739 3982
rect 233601 3979 233667 3982
rect 278129 4042 278195 4045
rect 464429 4042 464495 4045
rect 278129 4040 464495 4042
rect 278129 3984 278134 4040
rect 278190 3984 464434 4040
rect 464490 3984 464495 4040
rect 278129 3982 464495 3984
rect 278129 3979 278195 3982
rect 464429 3979 464495 3982
rect 25497 3906 25563 3909
rect 232957 3906 233023 3909
rect 25497 3904 233023 3906
rect 25497 3848 25502 3904
rect 25558 3848 232962 3904
rect 233018 3848 233023 3904
rect 25497 3846 233023 3848
rect 25497 3843 25563 3846
rect 232957 3843 233023 3846
rect 278037 3906 278103 3909
rect 467925 3906 467991 3909
rect 278037 3904 467991 3906
rect 278037 3848 278042 3904
rect 278098 3848 467930 3904
rect 467986 3848 467991 3904
rect 278037 3846 467991 3848
rect 278037 3843 278103 3846
rect 467925 3843 467991 3846
rect 24301 3770 24367 3773
rect 232773 3770 232839 3773
rect 24301 3768 232839 3770
rect 24301 3712 24306 3768
rect 24362 3712 232778 3768
rect 232834 3712 232839 3768
rect 24301 3710 232839 3712
rect 24301 3707 24367 3710
rect 232773 3707 232839 3710
rect 277853 3770 277919 3773
rect 471513 3770 471579 3773
rect 277853 3768 471579 3770
rect 277853 3712 277858 3768
rect 277914 3712 471518 3768
rect 471574 3712 471579 3768
rect 277853 3710 471579 3712
rect 277853 3707 277919 3710
rect 471513 3707 471579 3710
rect 16021 3634 16087 3637
rect 231577 3634 231643 3637
rect 16021 3632 231643 3634
rect 16021 3576 16026 3632
rect 16082 3576 231582 3632
rect 231638 3576 231643 3632
rect 16021 3574 231643 3576
rect 16021 3571 16087 3574
rect 231577 3571 231643 3574
rect 279969 3634 280035 3637
rect 475101 3634 475167 3637
rect 279969 3632 475167 3634
rect 279969 3576 279974 3632
rect 280030 3576 475106 3632
rect 475162 3576 475167 3632
rect 279969 3574 475167 3576
rect 279969 3571 280035 3574
rect 475101 3571 475167 3574
rect 14825 3498 14891 3501
rect 231393 3498 231459 3501
rect 14825 3496 231459 3498
rect 14825 3440 14830 3496
rect 14886 3440 231398 3496
rect 231454 3440 231459 3496
rect 14825 3438 231459 3440
rect 14825 3435 14891 3438
rect 231393 3435 231459 3438
rect 279877 3498 279943 3501
rect 478689 3498 478755 3501
rect 279877 3496 478755 3498
rect 279877 3440 279882 3496
rect 279938 3440 478694 3496
rect 478750 3440 478755 3496
rect 279877 3438 478755 3440
rect 279877 3435 279943 3438
rect 478689 3435 478755 3438
rect 6453 3362 6519 3365
rect 231117 3362 231183 3365
rect 6453 3360 231183 3362
rect 6453 3304 6458 3360
rect 6514 3304 231122 3360
rect 231178 3304 231183 3360
rect 6453 3302 231183 3304
rect 6453 3299 6519 3302
rect 231117 3299 231183 3302
rect 279785 3362 279851 3365
rect 482277 3362 482343 3365
rect 279785 3360 482343 3362
rect 279785 3304 279790 3360
rect 279846 3304 482282 3360
rect 482338 3304 482343 3360
rect 279785 3302 482343 3304
rect 279785 3299 279851 3302
rect 482277 3299 482343 3302
rect 224953 3226 225019 3229
rect 229829 3226 229895 3229
rect 224953 3224 229895 3226
rect 224953 3168 224958 3224
rect 225014 3168 229834 3224
rect 229890 3168 229895 3224
rect 224953 3166 229895 3168
rect 224953 3163 225019 3166
rect 229829 3163 229895 3166
<< via3 >>
rect 231716 399332 231780 399396
rect 233004 399392 233068 399396
rect 233004 399336 233018 399392
rect 233018 399336 233068 399392
rect 233004 399332 233068 399336
rect 237236 399392 237300 399396
rect 237236 399336 237250 399392
rect 237250 399336 237300 399392
rect 237236 399332 237300 399336
rect 238156 399332 238220 399396
rect 242756 399332 242820 399396
rect 276796 399392 276860 399396
rect 276796 399336 276846 399392
rect 276846 399336 276860 399392
rect 276796 399332 276860 399336
rect 282868 399332 282932 399396
rect 284340 399332 284404 399396
rect 285628 399332 285692 399396
rect 287284 399392 287348 399396
rect 287284 399336 287334 399392
rect 287334 399336 287348 399392
rect 287284 399332 287348 399336
rect 287836 399392 287900 399396
rect 287836 399336 287886 399392
rect 287886 399336 287900 399392
rect 287836 399332 287900 399336
rect 276796 398652 276860 398716
rect 238156 398516 238220 398580
rect 242756 398380 242820 398444
rect 287284 398244 287348 398308
rect 287836 398108 287900 398172
rect 284340 397972 284404 398036
rect 254716 314604 254780 314668
rect 254716 305008 254780 305012
rect 254716 304952 254766 305008
rect 254766 304952 254780 305008
rect 254716 304948 254780 304952
rect 255636 289036 255700 289100
rect 255636 275980 255700 276044
rect 237236 227836 237300 227900
rect 318748 227836 318812 227900
rect 338068 227972 338132 228036
rect 318748 227564 318812 227628
rect 338068 227700 338132 227764
rect 282868 194516 282932 194580
rect 285628 108972 285692 109036
rect 233004 76196 233068 76260
rect 318748 76060 318812 76124
rect 338068 76196 338132 76260
rect 318748 75788 318812 75852
rect 338068 75924 338132 75988
rect 492628 76060 492692 76124
rect 492628 75788 492692 75852
rect 231716 29004 231780 29068
<< metal4 >>
rect -8436 711278 -7836 711300
rect -8436 711042 -8254 711278
rect -8018 711042 -7836 711278
rect -8436 710958 -7836 711042
rect -8436 710722 -8254 710958
rect -8018 710722 -7836 710958
rect -8436 679254 -7836 710722
rect -8436 679018 -8254 679254
rect -8018 679018 -7836 679254
rect -8436 678934 -7836 679018
rect -8436 678698 -8254 678934
rect -8018 678698 -7836 678934
rect -8436 643254 -7836 678698
rect -8436 643018 -8254 643254
rect -8018 643018 -7836 643254
rect -8436 642934 -7836 643018
rect -8436 642698 -8254 642934
rect -8018 642698 -7836 642934
rect -8436 607254 -7836 642698
rect -8436 607018 -8254 607254
rect -8018 607018 -7836 607254
rect -8436 606934 -7836 607018
rect -8436 606698 -8254 606934
rect -8018 606698 -7836 606934
rect -8436 571254 -7836 606698
rect -8436 571018 -8254 571254
rect -8018 571018 -7836 571254
rect -8436 570934 -7836 571018
rect -8436 570698 -8254 570934
rect -8018 570698 -7836 570934
rect -8436 535254 -7836 570698
rect -8436 535018 -8254 535254
rect -8018 535018 -7836 535254
rect -8436 534934 -7836 535018
rect -8436 534698 -8254 534934
rect -8018 534698 -7836 534934
rect -8436 499254 -7836 534698
rect -8436 499018 -8254 499254
rect -8018 499018 -7836 499254
rect -8436 498934 -7836 499018
rect -8436 498698 -8254 498934
rect -8018 498698 -7836 498934
rect -8436 463254 -7836 498698
rect -8436 463018 -8254 463254
rect -8018 463018 -7836 463254
rect -8436 462934 -7836 463018
rect -8436 462698 -8254 462934
rect -8018 462698 -7836 462934
rect -8436 427254 -7836 462698
rect -8436 427018 -8254 427254
rect -8018 427018 -7836 427254
rect -8436 426934 -7836 427018
rect -8436 426698 -8254 426934
rect -8018 426698 -7836 426934
rect -8436 391254 -7836 426698
rect -8436 391018 -8254 391254
rect -8018 391018 -7836 391254
rect -8436 390934 -7836 391018
rect -8436 390698 -8254 390934
rect -8018 390698 -7836 390934
rect -8436 355254 -7836 390698
rect -8436 355018 -8254 355254
rect -8018 355018 -7836 355254
rect -8436 354934 -7836 355018
rect -8436 354698 -8254 354934
rect -8018 354698 -7836 354934
rect -8436 319254 -7836 354698
rect -8436 319018 -8254 319254
rect -8018 319018 -7836 319254
rect -8436 318934 -7836 319018
rect -8436 318698 -8254 318934
rect -8018 318698 -7836 318934
rect -8436 283254 -7836 318698
rect -8436 283018 -8254 283254
rect -8018 283018 -7836 283254
rect -8436 282934 -7836 283018
rect -8436 282698 -8254 282934
rect -8018 282698 -7836 282934
rect -8436 247254 -7836 282698
rect -8436 247018 -8254 247254
rect -8018 247018 -7836 247254
rect -8436 246934 -7836 247018
rect -8436 246698 -8254 246934
rect -8018 246698 -7836 246934
rect -8436 211254 -7836 246698
rect -8436 211018 -8254 211254
rect -8018 211018 -7836 211254
rect -8436 210934 -7836 211018
rect -8436 210698 -8254 210934
rect -8018 210698 -7836 210934
rect -8436 175254 -7836 210698
rect -8436 175018 -8254 175254
rect -8018 175018 -7836 175254
rect -8436 174934 -7836 175018
rect -8436 174698 -8254 174934
rect -8018 174698 -7836 174934
rect -8436 139254 -7836 174698
rect -8436 139018 -8254 139254
rect -8018 139018 -7836 139254
rect -8436 138934 -7836 139018
rect -8436 138698 -8254 138934
rect -8018 138698 -7836 138934
rect -8436 103254 -7836 138698
rect -8436 103018 -8254 103254
rect -8018 103018 -7836 103254
rect -8436 102934 -7836 103018
rect -8436 102698 -8254 102934
rect -8018 102698 -7836 102934
rect -8436 67254 -7836 102698
rect -8436 67018 -8254 67254
rect -8018 67018 -7836 67254
rect -8436 66934 -7836 67018
rect -8436 66698 -8254 66934
rect -8018 66698 -7836 66934
rect -8436 31254 -7836 66698
rect -8436 31018 -8254 31254
rect -8018 31018 -7836 31254
rect -8436 30934 -7836 31018
rect -8436 30698 -8254 30934
rect -8018 30698 -7836 30934
rect -8436 -6786 -7836 30698
rect -7516 710358 -6916 710380
rect -7516 710122 -7334 710358
rect -7098 710122 -6916 710358
rect -7516 710038 -6916 710122
rect -7516 709802 -7334 710038
rect -7098 709802 -6916 710038
rect -7516 697254 -6916 709802
rect 11604 710358 12204 711300
rect 11604 710122 11786 710358
rect 12022 710122 12204 710358
rect 11604 710038 12204 710122
rect 11604 709802 11786 710038
rect 12022 709802 12204 710038
rect -7516 697018 -7334 697254
rect -7098 697018 -6916 697254
rect -7516 696934 -6916 697018
rect -7516 696698 -7334 696934
rect -7098 696698 -6916 696934
rect -7516 661254 -6916 696698
rect -7516 661018 -7334 661254
rect -7098 661018 -6916 661254
rect -7516 660934 -6916 661018
rect -7516 660698 -7334 660934
rect -7098 660698 -6916 660934
rect -7516 625254 -6916 660698
rect -7516 625018 -7334 625254
rect -7098 625018 -6916 625254
rect -7516 624934 -6916 625018
rect -7516 624698 -7334 624934
rect -7098 624698 -6916 624934
rect -7516 589254 -6916 624698
rect -7516 589018 -7334 589254
rect -7098 589018 -6916 589254
rect -7516 588934 -6916 589018
rect -7516 588698 -7334 588934
rect -7098 588698 -6916 588934
rect -7516 553254 -6916 588698
rect -7516 553018 -7334 553254
rect -7098 553018 -6916 553254
rect -7516 552934 -6916 553018
rect -7516 552698 -7334 552934
rect -7098 552698 -6916 552934
rect -7516 517254 -6916 552698
rect -7516 517018 -7334 517254
rect -7098 517018 -6916 517254
rect -7516 516934 -6916 517018
rect -7516 516698 -7334 516934
rect -7098 516698 -6916 516934
rect -7516 481254 -6916 516698
rect -7516 481018 -7334 481254
rect -7098 481018 -6916 481254
rect -7516 480934 -6916 481018
rect -7516 480698 -7334 480934
rect -7098 480698 -6916 480934
rect -7516 445254 -6916 480698
rect -7516 445018 -7334 445254
rect -7098 445018 -6916 445254
rect -7516 444934 -6916 445018
rect -7516 444698 -7334 444934
rect -7098 444698 -6916 444934
rect -7516 409254 -6916 444698
rect -7516 409018 -7334 409254
rect -7098 409018 -6916 409254
rect -7516 408934 -6916 409018
rect -7516 408698 -7334 408934
rect -7098 408698 -6916 408934
rect -7516 373254 -6916 408698
rect -7516 373018 -7334 373254
rect -7098 373018 -6916 373254
rect -7516 372934 -6916 373018
rect -7516 372698 -7334 372934
rect -7098 372698 -6916 372934
rect -7516 337254 -6916 372698
rect -7516 337018 -7334 337254
rect -7098 337018 -6916 337254
rect -7516 336934 -6916 337018
rect -7516 336698 -7334 336934
rect -7098 336698 -6916 336934
rect -7516 301254 -6916 336698
rect -7516 301018 -7334 301254
rect -7098 301018 -6916 301254
rect -7516 300934 -6916 301018
rect -7516 300698 -7334 300934
rect -7098 300698 -6916 300934
rect -7516 265254 -6916 300698
rect -7516 265018 -7334 265254
rect -7098 265018 -6916 265254
rect -7516 264934 -6916 265018
rect -7516 264698 -7334 264934
rect -7098 264698 -6916 264934
rect -7516 229254 -6916 264698
rect -7516 229018 -7334 229254
rect -7098 229018 -6916 229254
rect -7516 228934 -6916 229018
rect -7516 228698 -7334 228934
rect -7098 228698 -6916 228934
rect -7516 193254 -6916 228698
rect -7516 193018 -7334 193254
rect -7098 193018 -6916 193254
rect -7516 192934 -6916 193018
rect -7516 192698 -7334 192934
rect -7098 192698 -6916 192934
rect -7516 157254 -6916 192698
rect -7516 157018 -7334 157254
rect -7098 157018 -6916 157254
rect -7516 156934 -6916 157018
rect -7516 156698 -7334 156934
rect -7098 156698 -6916 156934
rect -7516 121254 -6916 156698
rect -7516 121018 -7334 121254
rect -7098 121018 -6916 121254
rect -7516 120934 -6916 121018
rect -7516 120698 -7334 120934
rect -7098 120698 -6916 120934
rect -7516 85254 -6916 120698
rect -7516 85018 -7334 85254
rect -7098 85018 -6916 85254
rect -7516 84934 -6916 85018
rect -7516 84698 -7334 84934
rect -7098 84698 -6916 84934
rect -7516 49254 -6916 84698
rect -7516 49018 -7334 49254
rect -7098 49018 -6916 49254
rect -7516 48934 -6916 49018
rect -7516 48698 -7334 48934
rect -7098 48698 -6916 48934
rect -7516 13254 -6916 48698
rect -7516 13018 -7334 13254
rect -7098 13018 -6916 13254
rect -7516 12934 -6916 13018
rect -7516 12698 -7334 12934
rect -7098 12698 -6916 12934
rect -7516 -5866 -6916 12698
rect -6596 709438 -5996 709460
rect -6596 709202 -6414 709438
rect -6178 709202 -5996 709438
rect -6596 709118 -5996 709202
rect -6596 708882 -6414 709118
rect -6178 708882 -5996 709118
rect -6596 675654 -5996 708882
rect -6596 675418 -6414 675654
rect -6178 675418 -5996 675654
rect -6596 675334 -5996 675418
rect -6596 675098 -6414 675334
rect -6178 675098 -5996 675334
rect -6596 639654 -5996 675098
rect -6596 639418 -6414 639654
rect -6178 639418 -5996 639654
rect -6596 639334 -5996 639418
rect -6596 639098 -6414 639334
rect -6178 639098 -5996 639334
rect -6596 603654 -5996 639098
rect -6596 603418 -6414 603654
rect -6178 603418 -5996 603654
rect -6596 603334 -5996 603418
rect -6596 603098 -6414 603334
rect -6178 603098 -5996 603334
rect -6596 567654 -5996 603098
rect -6596 567418 -6414 567654
rect -6178 567418 -5996 567654
rect -6596 567334 -5996 567418
rect -6596 567098 -6414 567334
rect -6178 567098 -5996 567334
rect -6596 531654 -5996 567098
rect -6596 531418 -6414 531654
rect -6178 531418 -5996 531654
rect -6596 531334 -5996 531418
rect -6596 531098 -6414 531334
rect -6178 531098 -5996 531334
rect -6596 495654 -5996 531098
rect -6596 495418 -6414 495654
rect -6178 495418 -5996 495654
rect -6596 495334 -5996 495418
rect -6596 495098 -6414 495334
rect -6178 495098 -5996 495334
rect -6596 459654 -5996 495098
rect -6596 459418 -6414 459654
rect -6178 459418 -5996 459654
rect -6596 459334 -5996 459418
rect -6596 459098 -6414 459334
rect -6178 459098 -5996 459334
rect -6596 423654 -5996 459098
rect -6596 423418 -6414 423654
rect -6178 423418 -5996 423654
rect -6596 423334 -5996 423418
rect -6596 423098 -6414 423334
rect -6178 423098 -5996 423334
rect -6596 387654 -5996 423098
rect -6596 387418 -6414 387654
rect -6178 387418 -5996 387654
rect -6596 387334 -5996 387418
rect -6596 387098 -6414 387334
rect -6178 387098 -5996 387334
rect -6596 351654 -5996 387098
rect -6596 351418 -6414 351654
rect -6178 351418 -5996 351654
rect -6596 351334 -5996 351418
rect -6596 351098 -6414 351334
rect -6178 351098 -5996 351334
rect -6596 315654 -5996 351098
rect -6596 315418 -6414 315654
rect -6178 315418 -5996 315654
rect -6596 315334 -5996 315418
rect -6596 315098 -6414 315334
rect -6178 315098 -5996 315334
rect -6596 279654 -5996 315098
rect -6596 279418 -6414 279654
rect -6178 279418 -5996 279654
rect -6596 279334 -5996 279418
rect -6596 279098 -6414 279334
rect -6178 279098 -5996 279334
rect -6596 243654 -5996 279098
rect -6596 243418 -6414 243654
rect -6178 243418 -5996 243654
rect -6596 243334 -5996 243418
rect -6596 243098 -6414 243334
rect -6178 243098 -5996 243334
rect -6596 207654 -5996 243098
rect -6596 207418 -6414 207654
rect -6178 207418 -5996 207654
rect -6596 207334 -5996 207418
rect -6596 207098 -6414 207334
rect -6178 207098 -5996 207334
rect -6596 171654 -5996 207098
rect -6596 171418 -6414 171654
rect -6178 171418 -5996 171654
rect -6596 171334 -5996 171418
rect -6596 171098 -6414 171334
rect -6178 171098 -5996 171334
rect -6596 135654 -5996 171098
rect -6596 135418 -6414 135654
rect -6178 135418 -5996 135654
rect -6596 135334 -5996 135418
rect -6596 135098 -6414 135334
rect -6178 135098 -5996 135334
rect -6596 99654 -5996 135098
rect -6596 99418 -6414 99654
rect -6178 99418 -5996 99654
rect -6596 99334 -5996 99418
rect -6596 99098 -6414 99334
rect -6178 99098 -5996 99334
rect -6596 63654 -5996 99098
rect -6596 63418 -6414 63654
rect -6178 63418 -5996 63654
rect -6596 63334 -5996 63418
rect -6596 63098 -6414 63334
rect -6178 63098 -5996 63334
rect -6596 27654 -5996 63098
rect -6596 27418 -6414 27654
rect -6178 27418 -5996 27654
rect -6596 27334 -5996 27418
rect -6596 27098 -6414 27334
rect -6178 27098 -5996 27334
rect -6596 -4946 -5996 27098
rect -5676 708518 -5076 708540
rect -5676 708282 -5494 708518
rect -5258 708282 -5076 708518
rect -5676 708198 -5076 708282
rect -5676 707962 -5494 708198
rect -5258 707962 -5076 708198
rect -5676 693654 -5076 707962
rect 8004 708518 8604 709460
rect 8004 708282 8186 708518
rect 8422 708282 8604 708518
rect 8004 708198 8604 708282
rect 8004 707962 8186 708198
rect 8422 707962 8604 708198
rect -5676 693418 -5494 693654
rect -5258 693418 -5076 693654
rect -5676 693334 -5076 693418
rect -5676 693098 -5494 693334
rect -5258 693098 -5076 693334
rect -5676 657654 -5076 693098
rect -5676 657418 -5494 657654
rect -5258 657418 -5076 657654
rect -5676 657334 -5076 657418
rect -5676 657098 -5494 657334
rect -5258 657098 -5076 657334
rect -5676 621654 -5076 657098
rect -5676 621418 -5494 621654
rect -5258 621418 -5076 621654
rect -5676 621334 -5076 621418
rect -5676 621098 -5494 621334
rect -5258 621098 -5076 621334
rect -5676 585654 -5076 621098
rect -5676 585418 -5494 585654
rect -5258 585418 -5076 585654
rect -5676 585334 -5076 585418
rect -5676 585098 -5494 585334
rect -5258 585098 -5076 585334
rect -5676 549654 -5076 585098
rect -5676 549418 -5494 549654
rect -5258 549418 -5076 549654
rect -5676 549334 -5076 549418
rect -5676 549098 -5494 549334
rect -5258 549098 -5076 549334
rect -5676 513654 -5076 549098
rect -5676 513418 -5494 513654
rect -5258 513418 -5076 513654
rect -5676 513334 -5076 513418
rect -5676 513098 -5494 513334
rect -5258 513098 -5076 513334
rect -5676 477654 -5076 513098
rect -5676 477418 -5494 477654
rect -5258 477418 -5076 477654
rect -5676 477334 -5076 477418
rect -5676 477098 -5494 477334
rect -5258 477098 -5076 477334
rect -5676 441654 -5076 477098
rect -5676 441418 -5494 441654
rect -5258 441418 -5076 441654
rect -5676 441334 -5076 441418
rect -5676 441098 -5494 441334
rect -5258 441098 -5076 441334
rect -5676 405654 -5076 441098
rect -5676 405418 -5494 405654
rect -5258 405418 -5076 405654
rect -5676 405334 -5076 405418
rect -5676 405098 -5494 405334
rect -5258 405098 -5076 405334
rect -5676 369654 -5076 405098
rect -5676 369418 -5494 369654
rect -5258 369418 -5076 369654
rect -5676 369334 -5076 369418
rect -5676 369098 -5494 369334
rect -5258 369098 -5076 369334
rect -5676 333654 -5076 369098
rect -5676 333418 -5494 333654
rect -5258 333418 -5076 333654
rect -5676 333334 -5076 333418
rect -5676 333098 -5494 333334
rect -5258 333098 -5076 333334
rect -5676 297654 -5076 333098
rect -5676 297418 -5494 297654
rect -5258 297418 -5076 297654
rect -5676 297334 -5076 297418
rect -5676 297098 -5494 297334
rect -5258 297098 -5076 297334
rect -5676 261654 -5076 297098
rect -5676 261418 -5494 261654
rect -5258 261418 -5076 261654
rect -5676 261334 -5076 261418
rect -5676 261098 -5494 261334
rect -5258 261098 -5076 261334
rect -5676 225654 -5076 261098
rect -5676 225418 -5494 225654
rect -5258 225418 -5076 225654
rect -5676 225334 -5076 225418
rect -5676 225098 -5494 225334
rect -5258 225098 -5076 225334
rect -5676 189654 -5076 225098
rect -5676 189418 -5494 189654
rect -5258 189418 -5076 189654
rect -5676 189334 -5076 189418
rect -5676 189098 -5494 189334
rect -5258 189098 -5076 189334
rect -5676 153654 -5076 189098
rect -5676 153418 -5494 153654
rect -5258 153418 -5076 153654
rect -5676 153334 -5076 153418
rect -5676 153098 -5494 153334
rect -5258 153098 -5076 153334
rect -5676 117654 -5076 153098
rect -5676 117418 -5494 117654
rect -5258 117418 -5076 117654
rect -5676 117334 -5076 117418
rect -5676 117098 -5494 117334
rect -5258 117098 -5076 117334
rect -5676 81654 -5076 117098
rect -5676 81418 -5494 81654
rect -5258 81418 -5076 81654
rect -5676 81334 -5076 81418
rect -5676 81098 -5494 81334
rect -5258 81098 -5076 81334
rect -5676 45654 -5076 81098
rect -5676 45418 -5494 45654
rect -5258 45418 -5076 45654
rect -5676 45334 -5076 45418
rect -5676 45098 -5494 45334
rect -5258 45098 -5076 45334
rect -5676 9654 -5076 45098
rect -5676 9418 -5494 9654
rect -5258 9418 -5076 9654
rect -5676 9334 -5076 9418
rect -5676 9098 -5494 9334
rect -5258 9098 -5076 9334
rect -5676 -4026 -5076 9098
rect -4756 707598 -4156 707620
rect -4756 707362 -4574 707598
rect -4338 707362 -4156 707598
rect -4756 707278 -4156 707362
rect -4756 707042 -4574 707278
rect -4338 707042 -4156 707278
rect -4756 672054 -4156 707042
rect -4756 671818 -4574 672054
rect -4338 671818 -4156 672054
rect -4756 671734 -4156 671818
rect -4756 671498 -4574 671734
rect -4338 671498 -4156 671734
rect -4756 636054 -4156 671498
rect -4756 635818 -4574 636054
rect -4338 635818 -4156 636054
rect -4756 635734 -4156 635818
rect -4756 635498 -4574 635734
rect -4338 635498 -4156 635734
rect -4756 600054 -4156 635498
rect -4756 599818 -4574 600054
rect -4338 599818 -4156 600054
rect -4756 599734 -4156 599818
rect -4756 599498 -4574 599734
rect -4338 599498 -4156 599734
rect -4756 564054 -4156 599498
rect -4756 563818 -4574 564054
rect -4338 563818 -4156 564054
rect -4756 563734 -4156 563818
rect -4756 563498 -4574 563734
rect -4338 563498 -4156 563734
rect -4756 528054 -4156 563498
rect -4756 527818 -4574 528054
rect -4338 527818 -4156 528054
rect -4756 527734 -4156 527818
rect -4756 527498 -4574 527734
rect -4338 527498 -4156 527734
rect -4756 492054 -4156 527498
rect -4756 491818 -4574 492054
rect -4338 491818 -4156 492054
rect -4756 491734 -4156 491818
rect -4756 491498 -4574 491734
rect -4338 491498 -4156 491734
rect -4756 456054 -4156 491498
rect -4756 455818 -4574 456054
rect -4338 455818 -4156 456054
rect -4756 455734 -4156 455818
rect -4756 455498 -4574 455734
rect -4338 455498 -4156 455734
rect -4756 420054 -4156 455498
rect -4756 419818 -4574 420054
rect -4338 419818 -4156 420054
rect -4756 419734 -4156 419818
rect -4756 419498 -4574 419734
rect -4338 419498 -4156 419734
rect -4756 384054 -4156 419498
rect -4756 383818 -4574 384054
rect -4338 383818 -4156 384054
rect -4756 383734 -4156 383818
rect -4756 383498 -4574 383734
rect -4338 383498 -4156 383734
rect -4756 348054 -4156 383498
rect -4756 347818 -4574 348054
rect -4338 347818 -4156 348054
rect -4756 347734 -4156 347818
rect -4756 347498 -4574 347734
rect -4338 347498 -4156 347734
rect -4756 312054 -4156 347498
rect -4756 311818 -4574 312054
rect -4338 311818 -4156 312054
rect -4756 311734 -4156 311818
rect -4756 311498 -4574 311734
rect -4338 311498 -4156 311734
rect -4756 276054 -4156 311498
rect -4756 275818 -4574 276054
rect -4338 275818 -4156 276054
rect -4756 275734 -4156 275818
rect -4756 275498 -4574 275734
rect -4338 275498 -4156 275734
rect -4756 240054 -4156 275498
rect -4756 239818 -4574 240054
rect -4338 239818 -4156 240054
rect -4756 239734 -4156 239818
rect -4756 239498 -4574 239734
rect -4338 239498 -4156 239734
rect -4756 204054 -4156 239498
rect -4756 203818 -4574 204054
rect -4338 203818 -4156 204054
rect -4756 203734 -4156 203818
rect -4756 203498 -4574 203734
rect -4338 203498 -4156 203734
rect -4756 168054 -4156 203498
rect -4756 167818 -4574 168054
rect -4338 167818 -4156 168054
rect -4756 167734 -4156 167818
rect -4756 167498 -4574 167734
rect -4338 167498 -4156 167734
rect -4756 132054 -4156 167498
rect -4756 131818 -4574 132054
rect -4338 131818 -4156 132054
rect -4756 131734 -4156 131818
rect -4756 131498 -4574 131734
rect -4338 131498 -4156 131734
rect -4756 96054 -4156 131498
rect -4756 95818 -4574 96054
rect -4338 95818 -4156 96054
rect -4756 95734 -4156 95818
rect -4756 95498 -4574 95734
rect -4338 95498 -4156 95734
rect -4756 60054 -4156 95498
rect -4756 59818 -4574 60054
rect -4338 59818 -4156 60054
rect -4756 59734 -4156 59818
rect -4756 59498 -4574 59734
rect -4338 59498 -4156 59734
rect -4756 24054 -4156 59498
rect -4756 23818 -4574 24054
rect -4338 23818 -4156 24054
rect -4756 23734 -4156 23818
rect -4756 23498 -4574 23734
rect -4338 23498 -4156 23734
rect -4756 -3106 -4156 23498
rect -3836 706678 -3236 706700
rect -3836 706442 -3654 706678
rect -3418 706442 -3236 706678
rect -3836 706358 -3236 706442
rect -3836 706122 -3654 706358
rect -3418 706122 -3236 706358
rect -3836 690054 -3236 706122
rect 4404 706678 5004 707620
rect 4404 706442 4586 706678
rect 4822 706442 5004 706678
rect 4404 706358 5004 706442
rect 4404 706122 4586 706358
rect 4822 706122 5004 706358
rect -3836 689818 -3654 690054
rect -3418 689818 -3236 690054
rect -3836 689734 -3236 689818
rect -3836 689498 -3654 689734
rect -3418 689498 -3236 689734
rect -3836 654054 -3236 689498
rect -3836 653818 -3654 654054
rect -3418 653818 -3236 654054
rect -3836 653734 -3236 653818
rect -3836 653498 -3654 653734
rect -3418 653498 -3236 653734
rect -3836 618054 -3236 653498
rect -3836 617818 -3654 618054
rect -3418 617818 -3236 618054
rect -3836 617734 -3236 617818
rect -3836 617498 -3654 617734
rect -3418 617498 -3236 617734
rect -3836 582054 -3236 617498
rect -3836 581818 -3654 582054
rect -3418 581818 -3236 582054
rect -3836 581734 -3236 581818
rect -3836 581498 -3654 581734
rect -3418 581498 -3236 581734
rect -3836 546054 -3236 581498
rect -3836 545818 -3654 546054
rect -3418 545818 -3236 546054
rect -3836 545734 -3236 545818
rect -3836 545498 -3654 545734
rect -3418 545498 -3236 545734
rect -3836 510054 -3236 545498
rect -3836 509818 -3654 510054
rect -3418 509818 -3236 510054
rect -3836 509734 -3236 509818
rect -3836 509498 -3654 509734
rect -3418 509498 -3236 509734
rect -3836 474054 -3236 509498
rect -3836 473818 -3654 474054
rect -3418 473818 -3236 474054
rect -3836 473734 -3236 473818
rect -3836 473498 -3654 473734
rect -3418 473498 -3236 473734
rect -3836 438054 -3236 473498
rect -3836 437818 -3654 438054
rect -3418 437818 -3236 438054
rect -3836 437734 -3236 437818
rect -3836 437498 -3654 437734
rect -3418 437498 -3236 437734
rect -3836 402054 -3236 437498
rect -3836 401818 -3654 402054
rect -3418 401818 -3236 402054
rect -3836 401734 -3236 401818
rect -3836 401498 -3654 401734
rect -3418 401498 -3236 401734
rect -3836 366054 -3236 401498
rect -3836 365818 -3654 366054
rect -3418 365818 -3236 366054
rect -3836 365734 -3236 365818
rect -3836 365498 -3654 365734
rect -3418 365498 -3236 365734
rect -3836 330054 -3236 365498
rect -3836 329818 -3654 330054
rect -3418 329818 -3236 330054
rect -3836 329734 -3236 329818
rect -3836 329498 -3654 329734
rect -3418 329498 -3236 329734
rect -3836 294054 -3236 329498
rect -3836 293818 -3654 294054
rect -3418 293818 -3236 294054
rect -3836 293734 -3236 293818
rect -3836 293498 -3654 293734
rect -3418 293498 -3236 293734
rect -3836 258054 -3236 293498
rect -3836 257818 -3654 258054
rect -3418 257818 -3236 258054
rect -3836 257734 -3236 257818
rect -3836 257498 -3654 257734
rect -3418 257498 -3236 257734
rect -3836 222054 -3236 257498
rect -3836 221818 -3654 222054
rect -3418 221818 -3236 222054
rect -3836 221734 -3236 221818
rect -3836 221498 -3654 221734
rect -3418 221498 -3236 221734
rect -3836 186054 -3236 221498
rect -3836 185818 -3654 186054
rect -3418 185818 -3236 186054
rect -3836 185734 -3236 185818
rect -3836 185498 -3654 185734
rect -3418 185498 -3236 185734
rect -3836 150054 -3236 185498
rect -3836 149818 -3654 150054
rect -3418 149818 -3236 150054
rect -3836 149734 -3236 149818
rect -3836 149498 -3654 149734
rect -3418 149498 -3236 149734
rect -3836 114054 -3236 149498
rect -3836 113818 -3654 114054
rect -3418 113818 -3236 114054
rect -3836 113734 -3236 113818
rect -3836 113498 -3654 113734
rect -3418 113498 -3236 113734
rect -3836 78054 -3236 113498
rect -3836 77818 -3654 78054
rect -3418 77818 -3236 78054
rect -3836 77734 -3236 77818
rect -3836 77498 -3654 77734
rect -3418 77498 -3236 77734
rect -3836 42054 -3236 77498
rect -3836 41818 -3654 42054
rect -3418 41818 -3236 42054
rect -3836 41734 -3236 41818
rect -3836 41498 -3654 41734
rect -3418 41498 -3236 41734
rect -3836 6054 -3236 41498
rect -3836 5818 -3654 6054
rect -3418 5818 -3236 6054
rect -3836 5734 -3236 5818
rect -3836 5498 -3654 5734
rect -3418 5498 -3236 5734
rect -3836 -2186 -3236 5498
rect -2916 705758 -2316 705780
rect -2916 705522 -2734 705758
rect -2498 705522 -2316 705758
rect -2916 705438 -2316 705522
rect -2916 705202 -2734 705438
rect -2498 705202 -2316 705438
rect -2916 668454 -2316 705202
rect -2916 668218 -2734 668454
rect -2498 668218 -2316 668454
rect -2916 668134 -2316 668218
rect -2916 667898 -2734 668134
rect -2498 667898 -2316 668134
rect -2916 632454 -2316 667898
rect -2916 632218 -2734 632454
rect -2498 632218 -2316 632454
rect -2916 632134 -2316 632218
rect -2916 631898 -2734 632134
rect -2498 631898 -2316 632134
rect -2916 596454 -2316 631898
rect -2916 596218 -2734 596454
rect -2498 596218 -2316 596454
rect -2916 596134 -2316 596218
rect -2916 595898 -2734 596134
rect -2498 595898 -2316 596134
rect -2916 560454 -2316 595898
rect -2916 560218 -2734 560454
rect -2498 560218 -2316 560454
rect -2916 560134 -2316 560218
rect -2916 559898 -2734 560134
rect -2498 559898 -2316 560134
rect -2916 524454 -2316 559898
rect -2916 524218 -2734 524454
rect -2498 524218 -2316 524454
rect -2916 524134 -2316 524218
rect -2916 523898 -2734 524134
rect -2498 523898 -2316 524134
rect -2916 488454 -2316 523898
rect -2916 488218 -2734 488454
rect -2498 488218 -2316 488454
rect -2916 488134 -2316 488218
rect -2916 487898 -2734 488134
rect -2498 487898 -2316 488134
rect -2916 452454 -2316 487898
rect -2916 452218 -2734 452454
rect -2498 452218 -2316 452454
rect -2916 452134 -2316 452218
rect -2916 451898 -2734 452134
rect -2498 451898 -2316 452134
rect -2916 416454 -2316 451898
rect -2916 416218 -2734 416454
rect -2498 416218 -2316 416454
rect -2916 416134 -2316 416218
rect -2916 415898 -2734 416134
rect -2498 415898 -2316 416134
rect -2916 380454 -2316 415898
rect -2916 380218 -2734 380454
rect -2498 380218 -2316 380454
rect -2916 380134 -2316 380218
rect -2916 379898 -2734 380134
rect -2498 379898 -2316 380134
rect -2916 344454 -2316 379898
rect -2916 344218 -2734 344454
rect -2498 344218 -2316 344454
rect -2916 344134 -2316 344218
rect -2916 343898 -2734 344134
rect -2498 343898 -2316 344134
rect -2916 308454 -2316 343898
rect -2916 308218 -2734 308454
rect -2498 308218 -2316 308454
rect -2916 308134 -2316 308218
rect -2916 307898 -2734 308134
rect -2498 307898 -2316 308134
rect -2916 272454 -2316 307898
rect -2916 272218 -2734 272454
rect -2498 272218 -2316 272454
rect -2916 272134 -2316 272218
rect -2916 271898 -2734 272134
rect -2498 271898 -2316 272134
rect -2916 236454 -2316 271898
rect -2916 236218 -2734 236454
rect -2498 236218 -2316 236454
rect -2916 236134 -2316 236218
rect -2916 235898 -2734 236134
rect -2498 235898 -2316 236134
rect -2916 200454 -2316 235898
rect -2916 200218 -2734 200454
rect -2498 200218 -2316 200454
rect -2916 200134 -2316 200218
rect -2916 199898 -2734 200134
rect -2498 199898 -2316 200134
rect -2916 164454 -2316 199898
rect -2916 164218 -2734 164454
rect -2498 164218 -2316 164454
rect -2916 164134 -2316 164218
rect -2916 163898 -2734 164134
rect -2498 163898 -2316 164134
rect -2916 128454 -2316 163898
rect -2916 128218 -2734 128454
rect -2498 128218 -2316 128454
rect -2916 128134 -2316 128218
rect -2916 127898 -2734 128134
rect -2498 127898 -2316 128134
rect -2916 92454 -2316 127898
rect -2916 92218 -2734 92454
rect -2498 92218 -2316 92454
rect -2916 92134 -2316 92218
rect -2916 91898 -2734 92134
rect -2498 91898 -2316 92134
rect -2916 56454 -2316 91898
rect -2916 56218 -2734 56454
rect -2498 56218 -2316 56454
rect -2916 56134 -2316 56218
rect -2916 55898 -2734 56134
rect -2498 55898 -2316 56134
rect -2916 20454 -2316 55898
rect -2916 20218 -2734 20454
rect -2498 20218 -2316 20454
rect -2916 20134 -2316 20218
rect -2916 19898 -2734 20134
rect -2498 19898 -2316 20134
rect -2916 -1266 -2316 19898
rect -1996 704838 -1396 704860
rect -1996 704602 -1814 704838
rect -1578 704602 -1396 704838
rect -1996 704518 -1396 704602
rect -1996 704282 -1814 704518
rect -1578 704282 -1396 704518
rect -1996 686454 -1396 704282
rect -1996 686218 -1814 686454
rect -1578 686218 -1396 686454
rect -1996 686134 -1396 686218
rect -1996 685898 -1814 686134
rect -1578 685898 -1396 686134
rect -1996 650454 -1396 685898
rect -1996 650218 -1814 650454
rect -1578 650218 -1396 650454
rect -1996 650134 -1396 650218
rect -1996 649898 -1814 650134
rect -1578 649898 -1396 650134
rect -1996 614454 -1396 649898
rect -1996 614218 -1814 614454
rect -1578 614218 -1396 614454
rect -1996 614134 -1396 614218
rect -1996 613898 -1814 614134
rect -1578 613898 -1396 614134
rect -1996 578454 -1396 613898
rect -1996 578218 -1814 578454
rect -1578 578218 -1396 578454
rect -1996 578134 -1396 578218
rect -1996 577898 -1814 578134
rect -1578 577898 -1396 578134
rect -1996 542454 -1396 577898
rect -1996 542218 -1814 542454
rect -1578 542218 -1396 542454
rect -1996 542134 -1396 542218
rect -1996 541898 -1814 542134
rect -1578 541898 -1396 542134
rect -1996 506454 -1396 541898
rect -1996 506218 -1814 506454
rect -1578 506218 -1396 506454
rect -1996 506134 -1396 506218
rect -1996 505898 -1814 506134
rect -1578 505898 -1396 506134
rect -1996 470454 -1396 505898
rect -1996 470218 -1814 470454
rect -1578 470218 -1396 470454
rect -1996 470134 -1396 470218
rect -1996 469898 -1814 470134
rect -1578 469898 -1396 470134
rect -1996 434454 -1396 469898
rect -1996 434218 -1814 434454
rect -1578 434218 -1396 434454
rect -1996 434134 -1396 434218
rect -1996 433898 -1814 434134
rect -1578 433898 -1396 434134
rect -1996 398454 -1396 433898
rect -1996 398218 -1814 398454
rect -1578 398218 -1396 398454
rect -1996 398134 -1396 398218
rect -1996 397898 -1814 398134
rect -1578 397898 -1396 398134
rect -1996 362454 -1396 397898
rect -1996 362218 -1814 362454
rect -1578 362218 -1396 362454
rect -1996 362134 -1396 362218
rect -1996 361898 -1814 362134
rect -1578 361898 -1396 362134
rect -1996 326454 -1396 361898
rect -1996 326218 -1814 326454
rect -1578 326218 -1396 326454
rect -1996 326134 -1396 326218
rect -1996 325898 -1814 326134
rect -1578 325898 -1396 326134
rect -1996 290454 -1396 325898
rect -1996 290218 -1814 290454
rect -1578 290218 -1396 290454
rect -1996 290134 -1396 290218
rect -1996 289898 -1814 290134
rect -1578 289898 -1396 290134
rect -1996 254454 -1396 289898
rect -1996 254218 -1814 254454
rect -1578 254218 -1396 254454
rect -1996 254134 -1396 254218
rect -1996 253898 -1814 254134
rect -1578 253898 -1396 254134
rect -1996 218454 -1396 253898
rect -1996 218218 -1814 218454
rect -1578 218218 -1396 218454
rect -1996 218134 -1396 218218
rect -1996 217898 -1814 218134
rect -1578 217898 -1396 218134
rect -1996 182454 -1396 217898
rect -1996 182218 -1814 182454
rect -1578 182218 -1396 182454
rect -1996 182134 -1396 182218
rect -1996 181898 -1814 182134
rect -1578 181898 -1396 182134
rect -1996 146454 -1396 181898
rect -1996 146218 -1814 146454
rect -1578 146218 -1396 146454
rect -1996 146134 -1396 146218
rect -1996 145898 -1814 146134
rect -1578 145898 -1396 146134
rect -1996 110454 -1396 145898
rect -1996 110218 -1814 110454
rect -1578 110218 -1396 110454
rect -1996 110134 -1396 110218
rect -1996 109898 -1814 110134
rect -1578 109898 -1396 110134
rect -1996 74454 -1396 109898
rect -1996 74218 -1814 74454
rect -1578 74218 -1396 74454
rect -1996 74134 -1396 74218
rect -1996 73898 -1814 74134
rect -1578 73898 -1396 74134
rect -1996 38454 -1396 73898
rect -1996 38218 -1814 38454
rect -1578 38218 -1396 38454
rect -1996 38134 -1396 38218
rect -1996 37898 -1814 38134
rect -1578 37898 -1396 38134
rect -1996 2454 -1396 37898
rect -1996 2218 -1814 2454
rect -1578 2218 -1396 2454
rect -1996 2134 -1396 2218
rect -1996 1898 -1814 2134
rect -1578 1898 -1396 2134
rect -1996 -346 -1396 1898
rect -1996 -582 -1814 -346
rect -1578 -582 -1396 -346
rect -1996 -666 -1396 -582
rect -1996 -902 -1814 -666
rect -1578 -902 -1396 -666
rect -1996 -924 -1396 -902
rect 804 704838 1404 705780
rect 804 704602 986 704838
rect 1222 704602 1404 704838
rect 804 704518 1404 704602
rect 804 704282 986 704518
rect 1222 704282 1404 704518
rect 804 686454 1404 704282
rect 804 686218 986 686454
rect 1222 686218 1404 686454
rect 804 686134 1404 686218
rect 804 685898 986 686134
rect 1222 685898 1404 686134
rect 804 650454 1404 685898
rect 804 650218 986 650454
rect 1222 650218 1404 650454
rect 804 650134 1404 650218
rect 804 649898 986 650134
rect 1222 649898 1404 650134
rect 804 614454 1404 649898
rect 804 614218 986 614454
rect 1222 614218 1404 614454
rect 804 614134 1404 614218
rect 804 613898 986 614134
rect 1222 613898 1404 614134
rect 804 578454 1404 613898
rect 804 578218 986 578454
rect 1222 578218 1404 578454
rect 804 578134 1404 578218
rect 804 577898 986 578134
rect 1222 577898 1404 578134
rect 804 542454 1404 577898
rect 804 542218 986 542454
rect 1222 542218 1404 542454
rect 804 542134 1404 542218
rect 804 541898 986 542134
rect 1222 541898 1404 542134
rect 804 506454 1404 541898
rect 804 506218 986 506454
rect 1222 506218 1404 506454
rect 804 506134 1404 506218
rect 804 505898 986 506134
rect 1222 505898 1404 506134
rect 804 470454 1404 505898
rect 804 470218 986 470454
rect 1222 470218 1404 470454
rect 804 470134 1404 470218
rect 804 469898 986 470134
rect 1222 469898 1404 470134
rect 804 434454 1404 469898
rect 804 434218 986 434454
rect 1222 434218 1404 434454
rect 804 434134 1404 434218
rect 804 433898 986 434134
rect 1222 433898 1404 434134
rect 804 398454 1404 433898
rect 804 398218 986 398454
rect 1222 398218 1404 398454
rect 804 398134 1404 398218
rect 804 397898 986 398134
rect 1222 397898 1404 398134
rect 804 362454 1404 397898
rect 804 362218 986 362454
rect 1222 362218 1404 362454
rect 804 362134 1404 362218
rect 804 361898 986 362134
rect 1222 361898 1404 362134
rect 804 326454 1404 361898
rect 804 326218 986 326454
rect 1222 326218 1404 326454
rect 804 326134 1404 326218
rect 804 325898 986 326134
rect 1222 325898 1404 326134
rect 804 290454 1404 325898
rect 804 290218 986 290454
rect 1222 290218 1404 290454
rect 804 290134 1404 290218
rect 804 289898 986 290134
rect 1222 289898 1404 290134
rect 804 254454 1404 289898
rect 804 254218 986 254454
rect 1222 254218 1404 254454
rect 804 254134 1404 254218
rect 804 253898 986 254134
rect 1222 253898 1404 254134
rect 804 218454 1404 253898
rect 804 218218 986 218454
rect 1222 218218 1404 218454
rect 804 218134 1404 218218
rect 804 217898 986 218134
rect 1222 217898 1404 218134
rect 804 182454 1404 217898
rect 804 182218 986 182454
rect 1222 182218 1404 182454
rect 804 182134 1404 182218
rect 804 181898 986 182134
rect 1222 181898 1404 182134
rect 804 146454 1404 181898
rect 804 146218 986 146454
rect 1222 146218 1404 146454
rect 804 146134 1404 146218
rect 804 145898 986 146134
rect 1222 145898 1404 146134
rect 804 110454 1404 145898
rect 804 110218 986 110454
rect 1222 110218 1404 110454
rect 804 110134 1404 110218
rect 804 109898 986 110134
rect 1222 109898 1404 110134
rect 804 74454 1404 109898
rect 804 74218 986 74454
rect 1222 74218 1404 74454
rect 804 74134 1404 74218
rect 804 73898 986 74134
rect 1222 73898 1404 74134
rect 804 38454 1404 73898
rect 804 38218 986 38454
rect 1222 38218 1404 38454
rect 804 38134 1404 38218
rect 804 37898 986 38134
rect 1222 37898 1404 38134
rect 804 2454 1404 37898
rect 804 2218 986 2454
rect 1222 2218 1404 2454
rect 804 2134 1404 2218
rect 804 1898 986 2134
rect 1222 1898 1404 2134
rect 804 -346 1404 1898
rect 804 -582 986 -346
rect 1222 -582 1404 -346
rect 804 -666 1404 -582
rect 804 -902 986 -666
rect 1222 -902 1404 -666
rect -2916 -1502 -2734 -1266
rect -2498 -1502 -2316 -1266
rect -2916 -1586 -2316 -1502
rect -2916 -1822 -2734 -1586
rect -2498 -1822 -2316 -1586
rect -2916 -1844 -2316 -1822
rect 804 -1844 1404 -902
rect 4404 690054 5004 706122
rect 4404 689818 4586 690054
rect 4822 689818 5004 690054
rect 4404 689734 5004 689818
rect 4404 689498 4586 689734
rect 4822 689498 5004 689734
rect 4404 654054 5004 689498
rect 4404 653818 4586 654054
rect 4822 653818 5004 654054
rect 4404 653734 5004 653818
rect 4404 653498 4586 653734
rect 4822 653498 5004 653734
rect 4404 618054 5004 653498
rect 4404 617818 4586 618054
rect 4822 617818 5004 618054
rect 4404 617734 5004 617818
rect 4404 617498 4586 617734
rect 4822 617498 5004 617734
rect 4404 582054 5004 617498
rect 4404 581818 4586 582054
rect 4822 581818 5004 582054
rect 4404 581734 5004 581818
rect 4404 581498 4586 581734
rect 4822 581498 5004 581734
rect 4404 546054 5004 581498
rect 4404 545818 4586 546054
rect 4822 545818 5004 546054
rect 4404 545734 5004 545818
rect 4404 545498 4586 545734
rect 4822 545498 5004 545734
rect 4404 510054 5004 545498
rect 4404 509818 4586 510054
rect 4822 509818 5004 510054
rect 4404 509734 5004 509818
rect 4404 509498 4586 509734
rect 4822 509498 5004 509734
rect 4404 474054 5004 509498
rect 4404 473818 4586 474054
rect 4822 473818 5004 474054
rect 4404 473734 5004 473818
rect 4404 473498 4586 473734
rect 4822 473498 5004 473734
rect 4404 438054 5004 473498
rect 4404 437818 4586 438054
rect 4822 437818 5004 438054
rect 4404 437734 5004 437818
rect 4404 437498 4586 437734
rect 4822 437498 5004 437734
rect 4404 402054 5004 437498
rect 4404 401818 4586 402054
rect 4822 401818 5004 402054
rect 4404 401734 5004 401818
rect 4404 401498 4586 401734
rect 4822 401498 5004 401734
rect 4404 366054 5004 401498
rect 4404 365818 4586 366054
rect 4822 365818 5004 366054
rect 4404 365734 5004 365818
rect 4404 365498 4586 365734
rect 4822 365498 5004 365734
rect 4404 330054 5004 365498
rect 4404 329818 4586 330054
rect 4822 329818 5004 330054
rect 4404 329734 5004 329818
rect 4404 329498 4586 329734
rect 4822 329498 5004 329734
rect 4404 294054 5004 329498
rect 4404 293818 4586 294054
rect 4822 293818 5004 294054
rect 4404 293734 5004 293818
rect 4404 293498 4586 293734
rect 4822 293498 5004 293734
rect 4404 258054 5004 293498
rect 4404 257818 4586 258054
rect 4822 257818 5004 258054
rect 4404 257734 5004 257818
rect 4404 257498 4586 257734
rect 4822 257498 5004 257734
rect 4404 222054 5004 257498
rect 4404 221818 4586 222054
rect 4822 221818 5004 222054
rect 4404 221734 5004 221818
rect 4404 221498 4586 221734
rect 4822 221498 5004 221734
rect 4404 186054 5004 221498
rect 4404 185818 4586 186054
rect 4822 185818 5004 186054
rect 4404 185734 5004 185818
rect 4404 185498 4586 185734
rect 4822 185498 5004 185734
rect 4404 150054 5004 185498
rect 4404 149818 4586 150054
rect 4822 149818 5004 150054
rect 4404 149734 5004 149818
rect 4404 149498 4586 149734
rect 4822 149498 5004 149734
rect 4404 114054 5004 149498
rect 4404 113818 4586 114054
rect 4822 113818 5004 114054
rect 4404 113734 5004 113818
rect 4404 113498 4586 113734
rect 4822 113498 5004 113734
rect 4404 78054 5004 113498
rect 4404 77818 4586 78054
rect 4822 77818 5004 78054
rect 4404 77734 5004 77818
rect 4404 77498 4586 77734
rect 4822 77498 5004 77734
rect 4404 42054 5004 77498
rect 4404 41818 4586 42054
rect 4822 41818 5004 42054
rect 4404 41734 5004 41818
rect 4404 41498 4586 41734
rect 4822 41498 5004 41734
rect 4404 6054 5004 41498
rect 4404 5818 4586 6054
rect 4822 5818 5004 6054
rect 4404 5734 5004 5818
rect 4404 5498 4586 5734
rect 4822 5498 5004 5734
rect -3836 -2422 -3654 -2186
rect -3418 -2422 -3236 -2186
rect -3836 -2506 -3236 -2422
rect -3836 -2742 -3654 -2506
rect -3418 -2742 -3236 -2506
rect -3836 -2764 -3236 -2742
rect 4404 -2186 5004 5498
rect 4404 -2422 4586 -2186
rect 4822 -2422 5004 -2186
rect 4404 -2506 5004 -2422
rect 4404 -2742 4586 -2506
rect 4822 -2742 5004 -2506
rect -4756 -3342 -4574 -3106
rect -4338 -3342 -4156 -3106
rect -4756 -3426 -4156 -3342
rect -4756 -3662 -4574 -3426
rect -4338 -3662 -4156 -3426
rect -4756 -3684 -4156 -3662
rect 4404 -3684 5004 -2742
rect 8004 693654 8604 707962
rect 8004 693418 8186 693654
rect 8422 693418 8604 693654
rect 8004 693334 8604 693418
rect 8004 693098 8186 693334
rect 8422 693098 8604 693334
rect 8004 657654 8604 693098
rect 8004 657418 8186 657654
rect 8422 657418 8604 657654
rect 8004 657334 8604 657418
rect 8004 657098 8186 657334
rect 8422 657098 8604 657334
rect 8004 621654 8604 657098
rect 8004 621418 8186 621654
rect 8422 621418 8604 621654
rect 8004 621334 8604 621418
rect 8004 621098 8186 621334
rect 8422 621098 8604 621334
rect 8004 585654 8604 621098
rect 8004 585418 8186 585654
rect 8422 585418 8604 585654
rect 8004 585334 8604 585418
rect 8004 585098 8186 585334
rect 8422 585098 8604 585334
rect 8004 549654 8604 585098
rect 8004 549418 8186 549654
rect 8422 549418 8604 549654
rect 8004 549334 8604 549418
rect 8004 549098 8186 549334
rect 8422 549098 8604 549334
rect 8004 513654 8604 549098
rect 8004 513418 8186 513654
rect 8422 513418 8604 513654
rect 8004 513334 8604 513418
rect 8004 513098 8186 513334
rect 8422 513098 8604 513334
rect 8004 477654 8604 513098
rect 8004 477418 8186 477654
rect 8422 477418 8604 477654
rect 8004 477334 8604 477418
rect 8004 477098 8186 477334
rect 8422 477098 8604 477334
rect 8004 441654 8604 477098
rect 8004 441418 8186 441654
rect 8422 441418 8604 441654
rect 8004 441334 8604 441418
rect 8004 441098 8186 441334
rect 8422 441098 8604 441334
rect 8004 405654 8604 441098
rect 8004 405418 8186 405654
rect 8422 405418 8604 405654
rect 8004 405334 8604 405418
rect 8004 405098 8186 405334
rect 8422 405098 8604 405334
rect 8004 369654 8604 405098
rect 8004 369418 8186 369654
rect 8422 369418 8604 369654
rect 8004 369334 8604 369418
rect 8004 369098 8186 369334
rect 8422 369098 8604 369334
rect 8004 333654 8604 369098
rect 8004 333418 8186 333654
rect 8422 333418 8604 333654
rect 8004 333334 8604 333418
rect 8004 333098 8186 333334
rect 8422 333098 8604 333334
rect 8004 297654 8604 333098
rect 8004 297418 8186 297654
rect 8422 297418 8604 297654
rect 8004 297334 8604 297418
rect 8004 297098 8186 297334
rect 8422 297098 8604 297334
rect 8004 261654 8604 297098
rect 8004 261418 8186 261654
rect 8422 261418 8604 261654
rect 8004 261334 8604 261418
rect 8004 261098 8186 261334
rect 8422 261098 8604 261334
rect 8004 225654 8604 261098
rect 8004 225418 8186 225654
rect 8422 225418 8604 225654
rect 8004 225334 8604 225418
rect 8004 225098 8186 225334
rect 8422 225098 8604 225334
rect 8004 189654 8604 225098
rect 8004 189418 8186 189654
rect 8422 189418 8604 189654
rect 8004 189334 8604 189418
rect 8004 189098 8186 189334
rect 8422 189098 8604 189334
rect 8004 153654 8604 189098
rect 8004 153418 8186 153654
rect 8422 153418 8604 153654
rect 8004 153334 8604 153418
rect 8004 153098 8186 153334
rect 8422 153098 8604 153334
rect 8004 117654 8604 153098
rect 8004 117418 8186 117654
rect 8422 117418 8604 117654
rect 8004 117334 8604 117418
rect 8004 117098 8186 117334
rect 8422 117098 8604 117334
rect 8004 81654 8604 117098
rect 8004 81418 8186 81654
rect 8422 81418 8604 81654
rect 8004 81334 8604 81418
rect 8004 81098 8186 81334
rect 8422 81098 8604 81334
rect 8004 45654 8604 81098
rect 8004 45418 8186 45654
rect 8422 45418 8604 45654
rect 8004 45334 8604 45418
rect 8004 45098 8186 45334
rect 8422 45098 8604 45334
rect 8004 9654 8604 45098
rect 8004 9418 8186 9654
rect 8422 9418 8604 9654
rect 8004 9334 8604 9418
rect 8004 9098 8186 9334
rect 8422 9098 8604 9334
rect -5676 -4262 -5494 -4026
rect -5258 -4262 -5076 -4026
rect -5676 -4346 -5076 -4262
rect -5676 -4582 -5494 -4346
rect -5258 -4582 -5076 -4346
rect -5676 -4604 -5076 -4582
rect 8004 -4026 8604 9098
rect 8004 -4262 8186 -4026
rect 8422 -4262 8604 -4026
rect 8004 -4346 8604 -4262
rect 8004 -4582 8186 -4346
rect 8422 -4582 8604 -4346
rect -6596 -5182 -6414 -4946
rect -6178 -5182 -5996 -4946
rect -6596 -5266 -5996 -5182
rect -6596 -5502 -6414 -5266
rect -6178 -5502 -5996 -5266
rect -6596 -5524 -5996 -5502
rect 8004 -5524 8604 -4582
rect 11604 697254 12204 709802
rect 29604 711278 30204 711300
rect 29604 711042 29786 711278
rect 30022 711042 30204 711278
rect 29604 710958 30204 711042
rect 29604 710722 29786 710958
rect 30022 710722 30204 710958
rect 26004 709438 26604 709460
rect 26004 709202 26186 709438
rect 26422 709202 26604 709438
rect 26004 709118 26604 709202
rect 26004 708882 26186 709118
rect 26422 708882 26604 709118
rect 22404 707598 23004 707620
rect 22404 707362 22586 707598
rect 22822 707362 23004 707598
rect 22404 707278 23004 707362
rect 22404 707042 22586 707278
rect 22822 707042 23004 707278
rect 11604 697018 11786 697254
rect 12022 697018 12204 697254
rect 11604 696934 12204 697018
rect 11604 696698 11786 696934
rect 12022 696698 12204 696934
rect 11604 661254 12204 696698
rect 11604 661018 11786 661254
rect 12022 661018 12204 661254
rect 11604 660934 12204 661018
rect 11604 660698 11786 660934
rect 12022 660698 12204 660934
rect 11604 625254 12204 660698
rect 11604 625018 11786 625254
rect 12022 625018 12204 625254
rect 11604 624934 12204 625018
rect 11604 624698 11786 624934
rect 12022 624698 12204 624934
rect 11604 589254 12204 624698
rect 11604 589018 11786 589254
rect 12022 589018 12204 589254
rect 11604 588934 12204 589018
rect 11604 588698 11786 588934
rect 12022 588698 12204 588934
rect 11604 553254 12204 588698
rect 11604 553018 11786 553254
rect 12022 553018 12204 553254
rect 11604 552934 12204 553018
rect 11604 552698 11786 552934
rect 12022 552698 12204 552934
rect 11604 517254 12204 552698
rect 11604 517018 11786 517254
rect 12022 517018 12204 517254
rect 11604 516934 12204 517018
rect 11604 516698 11786 516934
rect 12022 516698 12204 516934
rect 11604 481254 12204 516698
rect 11604 481018 11786 481254
rect 12022 481018 12204 481254
rect 11604 480934 12204 481018
rect 11604 480698 11786 480934
rect 12022 480698 12204 480934
rect 11604 445254 12204 480698
rect 11604 445018 11786 445254
rect 12022 445018 12204 445254
rect 11604 444934 12204 445018
rect 11604 444698 11786 444934
rect 12022 444698 12204 444934
rect 11604 409254 12204 444698
rect 11604 409018 11786 409254
rect 12022 409018 12204 409254
rect 11604 408934 12204 409018
rect 11604 408698 11786 408934
rect 12022 408698 12204 408934
rect 11604 373254 12204 408698
rect 11604 373018 11786 373254
rect 12022 373018 12204 373254
rect 11604 372934 12204 373018
rect 11604 372698 11786 372934
rect 12022 372698 12204 372934
rect 11604 337254 12204 372698
rect 11604 337018 11786 337254
rect 12022 337018 12204 337254
rect 11604 336934 12204 337018
rect 11604 336698 11786 336934
rect 12022 336698 12204 336934
rect 11604 301254 12204 336698
rect 11604 301018 11786 301254
rect 12022 301018 12204 301254
rect 11604 300934 12204 301018
rect 11604 300698 11786 300934
rect 12022 300698 12204 300934
rect 11604 265254 12204 300698
rect 11604 265018 11786 265254
rect 12022 265018 12204 265254
rect 11604 264934 12204 265018
rect 11604 264698 11786 264934
rect 12022 264698 12204 264934
rect 11604 229254 12204 264698
rect 11604 229018 11786 229254
rect 12022 229018 12204 229254
rect 11604 228934 12204 229018
rect 11604 228698 11786 228934
rect 12022 228698 12204 228934
rect 11604 193254 12204 228698
rect 11604 193018 11786 193254
rect 12022 193018 12204 193254
rect 11604 192934 12204 193018
rect 11604 192698 11786 192934
rect 12022 192698 12204 192934
rect 11604 157254 12204 192698
rect 11604 157018 11786 157254
rect 12022 157018 12204 157254
rect 11604 156934 12204 157018
rect 11604 156698 11786 156934
rect 12022 156698 12204 156934
rect 11604 121254 12204 156698
rect 11604 121018 11786 121254
rect 12022 121018 12204 121254
rect 11604 120934 12204 121018
rect 11604 120698 11786 120934
rect 12022 120698 12204 120934
rect 11604 85254 12204 120698
rect 11604 85018 11786 85254
rect 12022 85018 12204 85254
rect 11604 84934 12204 85018
rect 11604 84698 11786 84934
rect 12022 84698 12204 84934
rect 11604 49254 12204 84698
rect 11604 49018 11786 49254
rect 12022 49018 12204 49254
rect 11604 48934 12204 49018
rect 11604 48698 11786 48934
rect 12022 48698 12204 48934
rect 11604 13254 12204 48698
rect 11604 13018 11786 13254
rect 12022 13018 12204 13254
rect 11604 12934 12204 13018
rect 11604 12698 11786 12934
rect 12022 12698 12204 12934
rect -7516 -6102 -7334 -5866
rect -7098 -6102 -6916 -5866
rect -7516 -6186 -6916 -6102
rect -7516 -6422 -7334 -6186
rect -7098 -6422 -6916 -6186
rect -7516 -6444 -6916 -6422
rect 11604 -5866 12204 12698
rect 18804 705758 19404 705780
rect 18804 705522 18986 705758
rect 19222 705522 19404 705758
rect 18804 705438 19404 705522
rect 18804 705202 18986 705438
rect 19222 705202 19404 705438
rect 18804 668454 19404 705202
rect 18804 668218 18986 668454
rect 19222 668218 19404 668454
rect 18804 668134 19404 668218
rect 18804 667898 18986 668134
rect 19222 667898 19404 668134
rect 18804 632454 19404 667898
rect 18804 632218 18986 632454
rect 19222 632218 19404 632454
rect 18804 632134 19404 632218
rect 18804 631898 18986 632134
rect 19222 631898 19404 632134
rect 18804 596454 19404 631898
rect 18804 596218 18986 596454
rect 19222 596218 19404 596454
rect 18804 596134 19404 596218
rect 18804 595898 18986 596134
rect 19222 595898 19404 596134
rect 18804 560454 19404 595898
rect 18804 560218 18986 560454
rect 19222 560218 19404 560454
rect 18804 560134 19404 560218
rect 18804 559898 18986 560134
rect 19222 559898 19404 560134
rect 18804 524454 19404 559898
rect 18804 524218 18986 524454
rect 19222 524218 19404 524454
rect 18804 524134 19404 524218
rect 18804 523898 18986 524134
rect 19222 523898 19404 524134
rect 18804 488454 19404 523898
rect 18804 488218 18986 488454
rect 19222 488218 19404 488454
rect 18804 488134 19404 488218
rect 18804 487898 18986 488134
rect 19222 487898 19404 488134
rect 18804 452454 19404 487898
rect 18804 452218 18986 452454
rect 19222 452218 19404 452454
rect 18804 452134 19404 452218
rect 18804 451898 18986 452134
rect 19222 451898 19404 452134
rect 18804 416454 19404 451898
rect 18804 416218 18986 416454
rect 19222 416218 19404 416454
rect 18804 416134 19404 416218
rect 18804 415898 18986 416134
rect 19222 415898 19404 416134
rect 18804 380454 19404 415898
rect 18804 380218 18986 380454
rect 19222 380218 19404 380454
rect 18804 380134 19404 380218
rect 18804 379898 18986 380134
rect 19222 379898 19404 380134
rect 18804 344454 19404 379898
rect 18804 344218 18986 344454
rect 19222 344218 19404 344454
rect 18804 344134 19404 344218
rect 18804 343898 18986 344134
rect 19222 343898 19404 344134
rect 18804 308454 19404 343898
rect 18804 308218 18986 308454
rect 19222 308218 19404 308454
rect 18804 308134 19404 308218
rect 18804 307898 18986 308134
rect 19222 307898 19404 308134
rect 18804 272454 19404 307898
rect 18804 272218 18986 272454
rect 19222 272218 19404 272454
rect 18804 272134 19404 272218
rect 18804 271898 18986 272134
rect 19222 271898 19404 272134
rect 18804 236454 19404 271898
rect 18804 236218 18986 236454
rect 19222 236218 19404 236454
rect 18804 236134 19404 236218
rect 18804 235898 18986 236134
rect 19222 235898 19404 236134
rect 18804 200454 19404 235898
rect 18804 200218 18986 200454
rect 19222 200218 19404 200454
rect 18804 200134 19404 200218
rect 18804 199898 18986 200134
rect 19222 199898 19404 200134
rect 18804 164454 19404 199898
rect 18804 164218 18986 164454
rect 19222 164218 19404 164454
rect 18804 164134 19404 164218
rect 18804 163898 18986 164134
rect 19222 163898 19404 164134
rect 18804 128454 19404 163898
rect 18804 128218 18986 128454
rect 19222 128218 19404 128454
rect 18804 128134 19404 128218
rect 18804 127898 18986 128134
rect 19222 127898 19404 128134
rect 18804 92454 19404 127898
rect 18804 92218 18986 92454
rect 19222 92218 19404 92454
rect 18804 92134 19404 92218
rect 18804 91898 18986 92134
rect 19222 91898 19404 92134
rect 18804 56454 19404 91898
rect 18804 56218 18986 56454
rect 19222 56218 19404 56454
rect 18804 56134 19404 56218
rect 18804 55898 18986 56134
rect 19222 55898 19404 56134
rect 18804 20454 19404 55898
rect 18804 20218 18986 20454
rect 19222 20218 19404 20454
rect 18804 20134 19404 20218
rect 18804 19898 18986 20134
rect 19222 19898 19404 20134
rect 18804 -1266 19404 19898
rect 18804 -1502 18986 -1266
rect 19222 -1502 19404 -1266
rect 18804 -1586 19404 -1502
rect 18804 -1822 18986 -1586
rect 19222 -1822 19404 -1586
rect 18804 -1844 19404 -1822
rect 22404 672054 23004 707042
rect 22404 671818 22586 672054
rect 22822 671818 23004 672054
rect 22404 671734 23004 671818
rect 22404 671498 22586 671734
rect 22822 671498 23004 671734
rect 22404 636054 23004 671498
rect 22404 635818 22586 636054
rect 22822 635818 23004 636054
rect 22404 635734 23004 635818
rect 22404 635498 22586 635734
rect 22822 635498 23004 635734
rect 22404 600054 23004 635498
rect 22404 599818 22586 600054
rect 22822 599818 23004 600054
rect 22404 599734 23004 599818
rect 22404 599498 22586 599734
rect 22822 599498 23004 599734
rect 22404 564054 23004 599498
rect 22404 563818 22586 564054
rect 22822 563818 23004 564054
rect 22404 563734 23004 563818
rect 22404 563498 22586 563734
rect 22822 563498 23004 563734
rect 22404 528054 23004 563498
rect 22404 527818 22586 528054
rect 22822 527818 23004 528054
rect 22404 527734 23004 527818
rect 22404 527498 22586 527734
rect 22822 527498 23004 527734
rect 22404 492054 23004 527498
rect 22404 491818 22586 492054
rect 22822 491818 23004 492054
rect 22404 491734 23004 491818
rect 22404 491498 22586 491734
rect 22822 491498 23004 491734
rect 22404 456054 23004 491498
rect 22404 455818 22586 456054
rect 22822 455818 23004 456054
rect 22404 455734 23004 455818
rect 22404 455498 22586 455734
rect 22822 455498 23004 455734
rect 22404 420054 23004 455498
rect 22404 419818 22586 420054
rect 22822 419818 23004 420054
rect 22404 419734 23004 419818
rect 22404 419498 22586 419734
rect 22822 419498 23004 419734
rect 22404 384054 23004 419498
rect 22404 383818 22586 384054
rect 22822 383818 23004 384054
rect 22404 383734 23004 383818
rect 22404 383498 22586 383734
rect 22822 383498 23004 383734
rect 22404 348054 23004 383498
rect 22404 347818 22586 348054
rect 22822 347818 23004 348054
rect 22404 347734 23004 347818
rect 22404 347498 22586 347734
rect 22822 347498 23004 347734
rect 22404 312054 23004 347498
rect 22404 311818 22586 312054
rect 22822 311818 23004 312054
rect 22404 311734 23004 311818
rect 22404 311498 22586 311734
rect 22822 311498 23004 311734
rect 22404 276054 23004 311498
rect 22404 275818 22586 276054
rect 22822 275818 23004 276054
rect 22404 275734 23004 275818
rect 22404 275498 22586 275734
rect 22822 275498 23004 275734
rect 22404 240054 23004 275498
rect 22404 239818 22586 240054
rect 22822 239818 23004 240054
rect 22404 239734 23004 239818
rect 22404 239498 22586 239734
rect 22822 239498 23004 239734
rect 22404 204054 23004 239498
rect 22404 203818 22586 204054
rect 22822 203818 23004 204054
rect 22404 203734 23004 203818
rect 22404 203498 22586 203734
rect 22822 203498 23004 203734
rect 22404 168054 23004 203498
rect 22404 167818 22586 168054
rect 22822 167818 23004 168054
rect 22404 167734 23004 167818
rect 22404 167498 22586 167734
rect 22822 167498 23004 167734
rect 22404 132054 23004 167498
rect 22404 131818 22586 132054
rect 22822 131818 23004 132054
rect 22404 131734 23004 131818
rect 22404 131498 22586 131734
rect 22822 131498 23004 131734
rect 22404 96054 23004 131498
rect 22404 95818 22586 96054
rect 22822 95818 23004 96054
rect 22404 95734 23004 95818
rect 22404 95498 22586 95734
rect 22822 95498 23004 95734
rect 22404 60054 23004 95498
rect 22404 59818 22586 60054
rect 22822 59818 23004 60054
rect 22404 59734 23004 59818
rect 22404 59498 22586 59734
rect 22822 59498 23004 59734
rect 22404 24054 23004 59498
rect 22404 23818 22586 24054
rect 22822 23818 23004 24054
rect 22404 23734 23004 23818
rect 22404 23498 22586 23734
rect 22822 23498 23004 23734
rect 22404 -3106 23004 23498
rect 22404 -3342 22586 -3106
rect 22822 -3342 23004 -3106
rect 22404 -3426 23004 -3342
rect 22404 -3662 22586 -3426
rect 22822 -3662 23004 -3426
rect 22404 -3684 23004 -3662
rect 26004 675654 26604 708882
rect 26004 675418 26186 675654
rect 26422 675418 26604 675654
rect 26004 675334 26604 675418
rect 26004 675098 26186 675334
rect 26422 675098 26604 675334
rect 26004 639654 26604 675098
rect 26004 639418 26186 639654
rect 26422 639418 26604 639654
rect 26004 639334 26604 639418
rect 26004 639098 26186 639334
rect 26422 639098 26604 639334
rect 26004 603654 26604 639098
rect 26004 603418 26186 603654
rect 26422 603418 26604 603654
rect 26004 603334 26604 603418
rect 26004 603098 26186 603334
rect 26422 603098 26604 603334
rect 26004 567654 26604 603098
rect 26004 567418 26186 567654
rect 26422 567418 26604 567654
rect 26004 567334 26604 567418
rect 26004 567098 26186 567334
rect 26422 567098 26604 567334
rect 26004 531654 26604 567098
rect 26004 531418 26186 531654
rect 26422 531418 26604 531654
rect 26004 531334 26604 531418
rect 26004 531098 26186 531334
rect 26422 531098 26604 531334
rect 26004 495654 26604 531098
rect 26004 495418 26186 495654
rect 26422 495418 26604 495654
rect 26004 495334 26604 495418
rect 26004 495098 26186 495334
rect 26422 495098 26604 495334
rect 26004 459654 26604 495098
rect 26004 459418 26186 459654
rect 26422 459418 26604 459654
rect 26004 459334 26604 459418
rect 26004 459098 26186 459334
rect 26422 459098 26604 459334
rect 26004 423654 26604 459098
rect 26004 423418 26186 423654
rect 26422 423418 26604 423654
rect 26004 423334 26604 423418
rect 26004 423098 26186 423334
rect 26422 423098 26604 423334
rect 26004 387654 26604 423098
rect 26004 387418 26186 387654
rect 26422 387418 26604 387654
rect 26004 387334 26604 387418
rect 26004 387098 26186 387334
rect 26422 387098 26604 387334
rect 26004 351654 26604 387098
rect 26004 351418 26186 351654
rect 26422 351418 26604 351654
rect 26004 351334 26604 351418
rect 26004 351098 26186 351334
rect 26422 351098 26604 351334
rect 26004 315654 26604 351098
rect 26004 315418 26186 315654
rect 26422 315418 26604 315654
rect 26004 315334 26604 315418
rect 26004 315098 26186 315334
rect 26422 315098 26604 315334
rect 26004 279654 26604 315098
rect 26004 279418 26186 279654
rect 26422 279418 26604 279654
rect 26004 279334 26604 279418
rect 26004 279098 26186 279334
rect 26422 279098 26604 279334
rect 26004 243654 26604 279098
rect 26004 243418 26186 243654
rect 26422 243418 26604 243654
rect 26004 243334 26604 243418
rect 26004 243098 26186 243334
rect 26422 243098 26604 243334
rect 26004 207654 26604 243098
rect 26004 207418 26186 207654
rect 26422 207418 26604 207654
rect 26004 207334 26604 207418
rect 26004 207098 26186 207334
rect 26422 207098 26604 207334
rect 26004 171654 26604 207098
rect 26004 171418 26186 171654
rect 26422 171418 26604 171654
rect 26004 171334 26604 171418
rect 26004 171098 26186 171334
rect 26422 171098 26604 171334
rect 26004 135654 26604 171098
rect 26004 135418 26186 135654
rect 26422 135418 26604 135654
rect 26004 135334 26604 135418
rect 26004 135098 26186 135334
rect 26422 135098 26604 135334
rect 26004 99654 26604 135098
rect 26004 99418 26186 99654
rect 26422 99418 26604 99654
rect 26004 99334 26604 99418
rect 26004 99098 26186 99334
rect 26422 99098 26604 99334
rect 26004 63654 26604 99098
rect 26004 63418 26186 63654
rect 26422 63418 26604 63654
rect 26004 63334 26604 63418
rect 26004 63098 26186 63334
rect 26422 63098 26604 63334
rect 26004 27654 26604 63098
rect 26004 27418 26186 27654
rect 26422 27418 26604 27654
rect 26004 27334 26604 27418
rect 26004 27098 26186 27334
rect 26422 27098 26604 27334
rect 26004 -4946 26604 27098
rect 26004 -5182 26186 -4946
rect 26422 -5182 26604 -4946
rect 26004 -5266 26604 -5182
rect 26004 -5502 26186 -5266
rect 26422 -5502 26604 -5266
rect 26004 -5524 26604 -5502
rect 29604 679254 30204 710722
rect 47604 710358 48204 711300
rect 47604 710122 47786 710358
rect 48022 710122 48204 710358
rect 47604 710038 48204 710122
rect 47604 709802 47786 710038
rect 48022 709802 48204 710038
rect 44004 708518 44604 709460
rect 44004 708282 44186 708518
rect 44422 708282 44604 708518
rect 44004 708198 44604 708282
rect 44004 707962 44186 708198
rect 44422 707962 44604 708198
rect 40404 706678 41004 707620
rect 40404 706442 40586 706678
rect 40822 706442 41004 706678
rect 40404 706358 41004 706442
rect 40404 706122 40586 706358
rect 40822 706122 41004 706358
rect 29604 679018 29786 679254
rect 30022 679018 30204 679254
rect 29604 678934 30204 679018
rect 29604 678698 29786 678934
rect 30022 678698 30204 678934
rect 29604 643254 30204 678698
rect 29604 643018 29786 643254
rect 30022 643018 30204 643254
rect 29604 642934 30204 643018
rect 29604 642698 29786 642934
rect 30022 642698 30204 642934
rect 29604 607254 30204 642698
rect 29604 607018 29786 607254
rect 30022 607018 30204 607254
rect 29604 606934 30204 607018
rect 29604 606698 29786 606934
rect 30022 606698 30204 606934
rect 29604 571254 30204 606698
rect 29604 571018 29786 571254
rect 30022 571018 30204 571254
rect 29604 570934 30204 571018
rect 29604 570698 29786 570934
rect 30022 570698 30204 570934
rect 29604 535254 30204 570698
rect 29604 535018 29786 535254
rect 30022 535018 30204 535254
rect 29604 534934 30204 535018
rect 29604 534698 29786 534934
rect 30022 534698 30204 534934
rect 29604 499254 30204 534698
rect 29604 499018 29786 499254
rect 30022 499018 30204 499254
rect 29604 498934 30204 499018
rect 29604 498698 29786 498934
rect 30022 498698 30204 498934
rect 29604 463254 30204 498698
rect 29604 463018 29786 463254
rect 30022 463018 30204 463254
rect 29604 462934 30204 463018
rect 29604 462698 29786 462934
rect 30022 462698 30204 462934
rect 29604 427254 30204 462698
rect 29604 427018 29786 427254
rect 30022 427018 30204 427254
rect 29604 426934 30204 427018
rect 29604 426698 29786 426934
rect 30022 426698 30204 426934
rect 29604 391254 30204 426698
rect 29604 391018 29786 391254
rect 30022 391018 30204 391254
rect 29604 390934 30204 391018
rect 29604 390698 29786 390934
rect 30022 390698 30204 390934
rect 29604 355254 30204 390698
rect 29604 355018 29786 355254
rect 30022 355018 30204 355254
rect 29604 354934 30204 355018
rect 29604 354698 29786 354934
rect 30022 354698 30204 354934
rect 29604 319254 30204 354698
rect 29604 319018 29786 319254
rect 30022 319018 30204 319254
rect 29604 318934 30204 319018
rect 29604 318698 29786 318934
rect 30022 318698 30204 318934
rect 29604 283254 30204 318698
rect 29604 283018 29786 283254
rect 30022 283018 30204 283254
rect 29604 282934 30204 283018
rect 29604 282698 29786 282934
rect 30022 282698 30204 282934
rect 29604 247254 30204 282698
rect 29604 247018 29786 247254
rect 30022 247018 30204 247254
rect 29604 246934 30204 247018
rect 29604 246698 29786 246934
rect 30022 246698 30204 246934
rect 29604 211254 30204 246698
rect 29604 211018 29786 211254
rect 30022 211018 30204 211254
rect 29604 210934 30204 211018
rect 29604 210698 29786 210934
rect 30022 210698 30204 210934
rect 29604 175254 30204 210698
rect 29604 175018 29786 175254
rect 30022 175018 30204 175254
rect 29604 174934 30204 175018
rect 29604 174698 29786 174934
rect 30022 174698 30204 174934
rect 29604 139254 30204 174698
rect 29604 139018 29786 139254
rect 30022 139018 30204 139254
rect 29604 138934 30204 139018
rect 29604 138698 29786 138934
rect 30022 138698 30204 138934
rect 29604 103254 30204 138698
rect 29604 103018 29786 103254
rect 30022 103018 30204 103254
rect 29604 102934 30204 103018
rect 29604 102698 29786 102934
rect 30022 102698 30204 102934
rect 29604 67254 30204 102698
rect 29604 67018 29786 67254
rect 30022 67018 30204 67254
rect 29604 66934 30204 67018
rect 29604 66698 29786 66934
rect 30022 66698 30204 66934
rect 29604 31254 30204 66698
rect 29604 31018 29786 31254
rect 30022 31018 30204 31254
rect 29604 30934 30204 31018
rect 29604 30698 29786 30934
rect 30022 30698 30204 30934
rect 11604 -6102 11786 -5866
rect 12022 -6102 12204 -5866
rect 11604 -6186 12204 -6102
rect 11604 -6422 11786 -6186
rect 12022 -6422 12204 -6186
rect -8436 -7022 -8254 -6786
rect -8018 -7022 -7836 -6786
rect -8436 -7106 -7836 -7022
rect -8436 -7342 -8254 -7106
rect -8018 -7342 -7836 -7106
rect -8436 -7364 -7836 -7342
rect 11604 -7364 12204 -6422
rect 29604 -6786 30204 30698
rect 36804 704838 37404 705780
rect 36804 704602 36986 704838
rect 37222 704602 37404 704838
rect 36804 704518 37404 704602
rect 36804 704282 36986 704518
rect 37222 704282 37404 704518
rect 36804 686454 37404 704282
rect 36804 686218 36986 686454
rect 37222 686218 37404 686454
rect 36804 686134 37404 686218
rect 36804 685898 36986 686134
rect 37222 685898 37404 686134
rect 36804 650454 37404 685898
rect 36804 650218 36986 650454
rect 37222 650218 37404 650454
rect 36804 650134 37404 650218
rect 36804 649898 36986 650134
rect 37222 649898 37404 650134
rect 36804 614454 37404 649898
rect 36804 614218 36986 614454
rect 37222 614218 37404 614454
rect 36804 614134 37404 614218
rect 36804 613898 36986 614134
rect 37222 613898 37404 614134
rect 36804 578454 37404 613898
rect 36804 578218 36986 578454
rect 37222 578218 37404 578454
rect 36804 578134 37404 578218
rect 36804 577898 36986 578134
rect 37222 577898 37404 578134
rect 36804 542454 37404 577898
rect 36804 542218 36986 542454
rect 37222 542218 37404 542454
rect 36804 542134 37404 542218
rect 36804 541898 36986 542134
rect 37222 541898 37404 542134
rect 36804 506454 37404 541898
rect 36804 506218 36986 506454
rect 37222 506218 37404 506454
rect 36804 506134 37404 506218
rect 36804 505898 36986 506134
rect 37222 505898 37404 506134
rect 36804 470454 37404 505898
rect 36804 470218 36986 470454
rect 37222 470218 37404 470454
rect 36804 470134 37404 470218
rect 36804 469898 36986 470134
rect 37222 469898 37404 470134
rect 36804 434454 37404 469898
rect 36804 434218 36986 434454
rect 37222 434218 37404 434454
rect 36804 434134 37404 434218
rect 36804 433898 36986 434134
rect 37222 433898 37404 434134
rect 36804 398454 37404 433898
rect 36804 398218 36986 398454
rect 37222 398218 37404 398454
rect 36804 398134 37404 398218
rect 36804 397898 36986 398134
rect 37222 397898 37404 398134
rect 36804 362454 37404 397898
rect 36804 362218 36986 362454
rect 37222 362218 37404 362454
rect 36804 362134 37404 362218
rect 36804 361898 36986 362134
rect 37222 361898 37404 362134
rect 36804 326454 37404 361898
rect 36804 326218 36986 326454
rect 37222 326218 37404 326454
rect 36804 326134 37404 326218
rect 36804 325898 36986 326134
rect 37222 325898 37404 326134
rect 36804 290454 37404 325898
rect 36804 290218 36986 290454
rect 37222 290218 37404 290454
rect 36804 290134 37404 290218
rect 36804 289898 36986 290134
rect 37222 289898 37404 290134
rect 36804 254454 37404 289898
rect 36804 254218 36986 254454
rect 37222 254218 37404 254454
rect 36804 254134 37404 254218
rect 36804 253898 36986 254134
rect 37222 253898 37404 254134
rect 36804 218454 37404 253898
rect 36804 218218 36986 218454
rect 37222 218218 37404 218454
rect 36804 218134 37404 218218
rect 36804 217898 36986 218134
rect 37222 217898 37404 218134
rect 36804 182454 37404 217898
rect 36804 182218 36986 182454
rect 37222 182218 37404 182454
rect 36804 182134 37404 182218
rect 36804 181898 36986 182134
rect 37222 181898 37404 182134
rect 36804 146454 37404 181898
rect 36804 146218 36986 146454
rect 37222 146218 37404 146454
rect 36804 146134 37404 146218
rect 36804 145898 36986 146134
rect 37222 145898 37404 146134
rect 36804 110454 37404 145898
rect 36804 110218 36986 110454
rect 37222 110218 37404 110454
rect 36804 110134 37404 110218
rect 36804 109898 36986 110134
rect 37222 109898 37404 110134
rect 36804 74454 37404 109898
rect 36804 74218 36986 74454
rect 37222 74218 37404 74454
rect 36804 74134 37404 74218
rect 36804 73898 36986 74134
rect 37222 73898 37404 74134
rect 36804 38454 37404 73898
rect 36804 38218 36986 38454
rect 37222 38218 37404 38454
rect 36804 38134 37404 38218
rect 36804 37898 36986 38134
rect 37222 37898 37404 38134
rect 36804 2454 37404 37898
rect 36804 2218 36986 2454
rect 37222 2218 37404 2454
rect 36804 2134 37404 2218
rect 36804 1898 36986 2134
rect 37222 1898 37404 2134
rect 36804 -346 37404 1898
rect 36804 -582 36986 -346
rect 37222 -582 37404 -346
rect 36804 -666 37404 -582
rect 36804 -902 36986 -666
rect 37222 -902 37404 -666
rect 36804 -1844 37404 -902
rect 40404 690054 41004 706122
rect 40404 689818 40586 690054
rect 40822 689818 41004 690054
rect 40404 689734 41004 689818
rect 40404 689498 40586 689734
rect 40822 689498 41004 689734
rect 40404 654054 41004 689498
rect 40404 653818 40586 654054
rect 40822 653818 41004 654054
rect 40404 653734 41004 653818
rect 40404 653498 40586 653734
rect 40822 653498 41004 653734
rect 40404 618054 41004 653498
rect 40404 617818 40586 618054
rect 40822 617818 41004 618054
rect 40404 617734 41004 617818
rect 40404 617498 40586 617734
rect 40822 617498 41004 617734
rect 40404 582054 41004 617498
rect 40404 581818 40586 582054
rect 40822 581818 41004 582054
rect 40404 581734 41004 581818
rect 40404 581498 40586 581734
rect 40822 581498 41004 581734
rect 40404 546054 41004 581498
rect 40404 545818 40586 546054
rect 40822 545818 41004 546054
rect 40404 545734 41004 545818
rect 40404 545498 40586 545734
rect 40822 545498 41004 545734
rect 40404 510054 41004 545498
rect 40404 509818 40586 510054
rect 40822 509818 41004 510054
rect 40404 509734 41004 509818
rect 40404 509498 40586 509734
rect 40822 509498 41004 509734
rect 40404 474054 41004 509498
rect 40404 473818 40586 474054
rect 40822 473818 41004 474054
rect 40404 473734 41004 473818
rect 40404 473498 40586 473734
rect 40822 473498 41004 473734
rect 40404 438054 41004 473498
rect 40404 437818 40586 438054
rect 40822 437818 41004 438054
rect 40404 437734 41004 437818
rect 40404 437498 40586 437734
rect 40822 437498 41004 437734
rect 40404 402054 41004 437498
rect 40404 401818 40586 402054
rect 40822 401818 41004 402054
rect 40404 401734 41004 401818
rect 40404 401498 40586 401734
rect 40822 401498 41004 401734
rect 40404 366054 41004 401498
rect 40404 365818 40586 366054
rect 40822 365818 41004 366054
rect 40404 365734 41004 365818
rect 40404 365498 40586 365734
rect 40822 365498 41004 365734
rect 40404 330054 41004 365498
rect 40404 329818 40586 330054
rect 40822 329818 41004 330054
rect 40404 329734 41004 329818
rect 40404 329498 40586 329734
rect 40822 329498 41004 329734
rect 40404 294054 41004 329498
rect 40404 293818 40586 294054
rect 40822 293818 41004 294054
rect 40404 293734 41004 293818
rect 40404 293498 40586 293734
rect 40822 293498 41004 293734
rect 40404 258054 41004 293498
rect 40404 257818 40586 258054
rect 40822 257818 41004 258054
rect 40404 257734 41004 257818
rect 40404 257498 40586 257734
rect 40822 257498 41004 257734
rect 40404 222054 41004 257498
rect 40404 221818 40586 222054
rect 40822 221818 41004 222054
rect 40404 221734 41004 221818
rect 40404 221498 40586 221734
rect 40822 221498 41004 221734
rect 40404 186054 41004 221498
rect 40404 185818 40586 186054
rect 40822 185818 41004 186054
rect 40404 185734 41004 185818
rect 40404 185498 40586 185734
rect 40822 185498 41004 185734
rect 40404 150054 41004 185498
rect 40404 149818 40586 150054
rect 40822 149818 41004 150054
rect 40404 149734 41004 149818
rect 40404 149498 40586 149734
rect 40822 149498 41004 149734
rect 40404 114054 41004 149498
rect 40404 113818 40586 114054
rect 40822 113818 41004 114054
rect 40404 113734 41004 113818
rect 40404 113498 40586 113734
rect 40822 113498 41004 113734
rect 40404 78054 41004 113498
rect 40404 77818 40586 78054
rect 40822 77818 41004 78054
rect 40404 77734 41004 77818
rect 40404 77498 40586 77734
rect 40822 77498 41004 77734
rect 40404 42054 41004 77498
rect 40404 41818 40586 42054
rect 40822 41818 41004 42054
rect 40404 41734 41004 41818
rect 40404 41498 40586 41734
rect 40822 41498 41004 41734
rect 40404 6054 41004 41498
rect 40404 5818 40586 6054
rect 40822 5818 41004 6054
rect 40404 5734 41004 5818
rect 40404 5498 40586 5734
rect 40822 5498 41004 5734
rect 40404 -2186 41004 5498
rect 40404 -2422 40586 -2186
rect 40822 -2422 41004 -2186
rect 40404 -2506 41004 -2422
rect 40404 -2742 40586 -2506
rect 40822 -2742 41004 -2506
rect 40404 -3684 41004 -2742
rect 44004 693654 44604 707962
rect 44004 693418 44186 693654
rect 44422 693418 44604 693654
rect 44004 693334 44604 693418
rect 44004 693098 44186 693334
rect 44422 693098 44604 693334
rect 44004 657654 44604 693098
rect 44004 657418 44186 657654
rect 44422 657418 44604 657654
rect 44004 657334 44604 657418
rect 44004 657098 44186 657334
rect 44422 657098 44604 657334
rect 44004 621654 44604 657098
rect 44004 621418 44186 621654
rect 44422 621418 44604 621654
rect 44004 621334 44604 621418
rect 44004 621098 44186 621334
rect 44422 621098 44604 621334
rect 44004 585654 44604 621098
rect 44004 585418 44186 585654
rect 44422 585418 44604 585654
rect 44004 585334 44604 585418
rect 44004 585098 44186 585334
rect 44422 585098 44604 585334
rect 44004 549654 44604 585098
rect 44004 549418 44186 549654
rect 44422 549418 44604 549654
rect 44004 549334 44604 549418
rect 44004 549098 44186 549334
rect 44422 549098 44604 549334
rect 44004 513654 44604 549098
rect 44004 513418 44186 513654
rect 44422 513418 44604 513654
rect 44004 513334 44604 513418
rect 44004 513098 44186 513334
rect 44422 513098 44604 513334
rect 44004 477654 44604 513098
rect 44004 477418 44186 477654
rect 44422 477418 44604 477654
rect 44004 477334 44604 477418
rect 44004 477098 44186 477334
rect 44422 477098 44604 477334
rect 44004 441654 44604 477098
rect 44004 441418 44186 441654
rect 44422 441418 44604 441654
rect 44004 441334 44604 441418
rect 44004 441098 44186 441334
rect 44422 441098 44604 441334
rect 44004 405654 44604 441098
rect 44004 405418 44186 405654
rect 44422 405418 44604 405654
rect 44004 405334 44604 405418
rect 44004 405098 44186 405334
rect 44422 405098 44604 405334
rect 44004 369654 44604 405098
rect 44004 369418 44186 369654
rect 44422 369418 44604 369654
rect 44004 369334 44604 369418
rect 44004 369098 44186 369334
rect 44422 369098 44604 369334
rect 44004 333654 44604 369098
rect 44004 333418 44186 333654
rect 44422 333418 44604 333654
rect 44004 333334 44604 333418
rect 44004 333098 44186 333334
rect 44422 333098 44604 333334
rect 44004 297654 44604 333098
rect 44004 297418 44186 297654
rect 44422 297418 44604 297654
rect 44004 297334 44604 297418
rect 44004 297098 44186 297334
rect 44422 297098 44604 297334
rect 44004 261654 44604 297098
rect 44004 261418 44186 261654
rect 44422 261418 44604 261654
rect 44004 261334 44604 261418
rect 44004 261098 44186 261334
rect 44422 261098 44604 261334
rect 44004 225654 44604 261098
rect 44004 225418 44186 225654
rect 44422 225418 44604 225654
rect 44004 225334 44604 225418
rect 44004 225098 44186 225334
rect 44422 225098 44604 225334
rect 44004 189654 44604 225098
rect 44004 189418 44186 189654
rect 44422 189418 44604 189654
rect 44004 189334 44604 189418
rect 44004 189098 44186 189334
rect 44422 189098 44604 189334
rect 44004 153654 44604 189098
rect 44004 153418 44186 153654
rect 44422 153418 44604 153654
rect 44004 153334 44604 153418
rect 44004 153098 44186 153334
rect 44422 153098 44604 153334
rect 44004 117654 44604 153098
rect 44004 117418 44186 117654
rect 44422 117418 44604 117654
rect 44004 117334 44604 117418
rect 44004 117098 44186 117334
rect 44422 117098 44604 117334
rect 44004 81654 44604 117098
rect 44004 81418 44186 81654
rect 44422 81418 44604 81654
rect 44004 81334 44604 81418
rect 44004 81098 44186 81334
rect 44422 81098 44604 81334
rect 44004 45654 44604 81098
rect 44004 45418 44186 45654
rect 44422 45418 44604 45654
rect 44004 45334 44604 45418
rect 44004 45098 44186 45334
rect 44422 45098 44604 45334
rect 44004 9654 44604 45098
rect 44004 9418 44186 9654
rect 44422 9418 44604 9654
rect 44004 9334 44604 9418
rect 44004 9098 44186 9334
rect 44422 9098 44604 9334
rect 44004 -4026 44604 9098
rect 44004 -4262 44186 -4026
rect 44422 -4262 44604 -4026
rect 44004 -4346 44604 -4262
rect 44004 -4582 44186 -4346
rect 44422 -4582 44604 -4346
rect 44004 -5524 44604 -4582
rect 47604 697254 48204 709802
rect 65604 711278 66204 711300
rect 65604 711042 65786 711278
rect 66022 711042 66204 711278
rect 65604 710958 66204 711042
rect 65604 710722 65786 710958
rect 66022 710722 66204 710958
rect 62004 709438 62604 709460
rect 62004 709202 62186 709438
rect 62422 709202 62604 709438
rect 62004 709118 62604 709202
rect 62004 708882 62186 709118
rect 62422 708882 62604 709118
rect 58404 707598 59004 707620
rect 58404 707362 58586 707598
rect 58822 707362 59004 707598
rect 58404 707278 59004 707362
rect 58404 707042 58586 707278
rect 58822 707042 59004 707278
rect 47604 697018 47786 697254
rect 48022 697018 48204 697254
rect 47604 696934 48204 697018
rect 47604 696698 47786 696934
rect 48022 696698 48204 696934
rect 47604 661254 48204 696698
rect 47604 661018 47786 661254
rect 48022 661018 48204 661254
rect 47604 660934 48204 661018
rect 47604 660698 47786 660934
rect 48022 660698 48204 660934
rect 47604 625254 48204 660698
rect 47604 625018 47786 625254
rect 48022 625018 48204 625254
rect 47604 624934 48204 625018
rect 47604 624698 47786 624934
rect 48022 624698 48204 624934
rect 47604 589254 48204 624698
rect 47604 589018 47786 589254
rect 48022 589018 48204 589254
rect 47604 588934 48204 589018
rect 47604 588698 47786 588934
rect 48022 588698 48204 588934
rect 47604 553254 48204 588698
rect 47604 553018 47786 553254
rect 48022 553018 48204 553254
rect 47604 552934 48204 553018
rect 47604 552698 47786 552934
rect 48022 552698 48204 552934
rect 47604 517254 48204 552698
rect 47604 517018 47786 517254
rect 48022 517018 48204 517254
rect 47604 516934 48204 517018
rect 47604 516698 47786 516934
rect 48022 516698 48204 516934
rect 47604 481254 48204 516698
rect 47604 481018 47786 481254
rect 48022 481018 48204 481254
rect 47604 480934 48204 481018
rect 47604 480698 47786 480934
rect 48022 480698 48204 480934
rect 47604 445254 48204 480698
rect 47604 445018 47786 445254
rect 48022 445018 48204 445254
rect 47604 444934 48204 445018
rect 47604 444698 47786 444934
rect 48022 444698 48204 444934
rect 47604 409254 48204 444698
rect 47604 409018 47786 409254
rect 48022 409018 48204 409254
rect 47604 408934 48204 409018
rect 47604 408698 47786 408934
rect 48022 408698 48204 408934
rect 47604 373254 48204 408698
rect 47604 373018 47786 373254
rect 48022 373018 48204 373254
rect 47604 372934 48204 373018
rect 47604 372698 47786 372934
rect 48022 372698 48204 372934
rect 47604 337254 48204 372698
rect 47604 337018 47786 337254
rect 48022 337018 48204 337254
rect 47604 336934 48204 337018
rect 47604 336698 47786 336934
rect 48022 336698 48204 336934
rect 47604 301254 48204 336698
rect 47604 301018 47786 301254
rect 48022 301018 48204 301254
rect 47604 300934 48204 301018
rect 47604 300698 47786 300934
rect 48022 300698 48204 300934
rect 47604 265254 48204 300698
rect 47604 265018 47786 265254
rect 48022 265018 48204 265254
rect 47604 264934 48204 265018
rect 47604 264698 47786 264934
rect 48022 264698 48204 264934
rect 47604 229254 48204 264698
rect 47604 229018 47786 229254
rect 48022 229018 48204 229254
rect 47604 228934 48204 229018
rect 47604 228698 47786 228934
rect 48022 228698 48204 228934
rect 47604 193254 48204 228698
rect 47604 193018 47786 193254
rect 48022 193018 48204 193254
rect 47604 192934 48204 193018
rect 47604 192698 47786 192934
rect 48022 192698 48204 192934
rect 47604 157254 48204 192698
rect 47604 157018 47786 157254
rect 48022 157018 48204 157254
rect 47604 156934 48204 157018
rect 47604 156698 47786 156934
rect 48022 156698 48204 156934
rect 47604 121254 48204 156698
rect 47604 121018 47786 121254
rect 48022 121018 48204 121254
rect 47604 120934 48204 121018
rect 47604 120698 47786 120934
rect 48022 120698 48204 120934
rect 47604 85254 48204 120698
rect 47604 85018 47786 85254
rect 48022 85018 48204 85254
rect 47604 84934 48204 85018
rect 47604 84698 47786 84934
rect 48022 84698 48204 84934
rect 47604 49254 48204 84698
rect 47604 49018 47786 49254
rect 48022 49018 48204 49254
rect 47604 48934 48204 49018
rect 47604 48698 47786 48934
rect 48022 48698 48204 48934
rect 47604 13254 48204 48698
rect 47604 13018 47786 13254
rect 48022 13018 48204 13254
rect 47604 12934 48204 13018
rect 47604 12698 47786 12934
rect 48022 12698 48204 12934
rect 29604 -7022 29786 -6786
rect 30022 -7022 30204 -6786
rect 29604 -7106 30204 -7022
rect 29604 -7342 29786 -7106
rect 30022 -7342 30204 -7106
rect 29604 -7364 30204 -7342
rect 47604 -5866 48204 12698
rect 54804 705758 55404 705780
rect 54804 705522 54986 705758
rect 55222 705522 55404 705758
rect 54804 705438 55404 705522
rect 54804 705202 54986 705438
rect 55222 705202 55404 705438
rect 54804 668454 55404 705202
rect 54804 668218 54986 668454
rect 55222 668218 55404 668454
rect 54804 668134 55404 668218
rect 54804 667898 54986 668134
rect 55222 667898 55404 668134
rect 54804 632454 55404 667898
rect 54804 632218 54986 632454
rect 55222 632218 55404 632454
rect 54804 632134 55404 632218
rect 54804 631898 54986 632134
rect 55222 631898 55404 632134
rect 54804 596454 55404 631898
rect 54804 596218 54986 596454
rect 55222 596218 55404 596454
rect 54804 596134 55404 596218
rect 54804 595898 54986 596134
rect 55222 595898 55404 596134
rect 54804 560454 55404 595898
rect 54804 560218 54986 560454
rect 55222 560218 55404 560454
rect 54804 560134 55404 560218
rect 54804 559898 54986 560134
rect 55222 559898 55404 560134
rect 54804 524454 55404 559898
rect 54804 524218 54986 524454
rect 55222 524218 55404 524454
rect 54804 524134 55404 524218
rect 54804 523898 54986 524134
rect 55222 523898 55404 524134
rect 54804 488454 55404 523898
rect 54804 488218 54986 488454
rect 55222 488218 55404 488454
rect 54804 488134 55404 488218
rect 54804 487898 54986 488134
rect 55222 487898 55404 488134
rect 54804 452454 55404 487898
rect 54804 452218 54986 452454
rect 55222 452218 55404 452454
rect 54804 452134 55404 452218
rect 54804 451898 54986 452134
rect 55222 451898 55404 452134
rect 54804 416454 55404 451898
rect 54804 416218 54986 416454
rect 55222 416218 55404 416454
rect 54804 416134 55404 416218
rect 54804 415898 54986 416134
rect 55222 415898 55404 416134
rect 54804 380454 55404 415898
rect 54804 380218 54986 380454
rect 55222 380218 55404 380454
rect 54804 380134 55404 380218
rect 54804 379898 54986 380134
rect 55222 379898 55404 380134
rect 54804 344454 55404 379898
rect 54804 344218 54986 344454
rect 55222 344218 55404 344454
rect 54804 344134 55404 344218
rect 54804 343898 54986 344134
rect 55222 343898 55404 344134
rect 54804 308454 55404 343898
rect 54804 308218 54986 308454
rect 55222 308218 55404 308454
rect 54804 308134 55404 308218
rect 54804 307898 54986 308134
rect 55222 307898 55404 308134
rect 54804 272454 55404 307898
rect 54804 272218 54986 272454
rect 55222 272218 55404 272454
rect 54804 272134 55404 272218
rect 54804 271898 54986 272134
rect 55222 271898 55404 272134
rect 54804 236454 55404 271898
rect 54804 236218 54986 236454
rect 55222 236218 55404 236454
rect 54804 236134 55404 236218
rect 54804 235898 54986 236134
rect 55222 235898 55404 236134
rect 54804 200454 55404 235898
rect 54804 200218 54986 200454
rect 55222 200218 55404 200454
rect 54804 200134 55404 200218
rect 54804 199898 54986 200134
rect 55222 199898 55404 200134
rect 54804 164454 55404 199898
rect 54804 164218 54986 164454
rect 55222 164218 55404 164454
rect 54804 164134 55404 164218
rect 54804 163898 54986 164134
rect 55222 163898 55404 164134
rect 54804 128454 55404 163898
rect 54804 128218 54986 128454
rect 55222 128218 55404 128454
rect 54804 128134 55404 128218
rect 54804 127898 54986 128134
rect 55222 127898 55404 128134
rect 54804 92454 55404 127898
rect 54804 92218 54986 92454
rect 55222 92218 55404 92454
rect 54804 92134 55404 92218
rect 54804 91898 54986 92134
rect 55222 91898 55404 92134
rect 54804 56454 55404 91898
rect 54804 56218 54986 56454
rect 55222 56218 55404 56454
rect 54804 56134 55404 56218
rect 54804 55898 54986 56134
rect 55222 55898 55404 56134
rect 54804 20454 55404 55898
rect 54804 20218 54986 20454
rect 55222 20218 55404 20454
rect 54804 20134 55404 20218
rect 54804 19898 54986 20134
rect 55222 19898 55404 20134
rect 54804 -1266 55404 19898
rect 54804 -1502 54986 -1266
rect 55222 -1502 55404 -1266
rect 54804 -1586 55404 -1502
rect 54804 -1822 54986 -1586
rect 55222 -1822 55404 -1586
rect 54804 -1844 55404 -1822
rect 58404 672054 59004 707042
rect 58404 671818 58586 672054
rect 58822 671818 59004 672054
rect 58404 671734 59004 671818
rect 58404 671498 58586 671734
rect 58822 671498 59004 671734
rect 58404 636054 59004 671498
rect 58404 635818 58586 636054
rect 58822 635818 59004 636054
rect 58404 635734 59004 635818
rect 58404 635498 58586 635734
rect 58822 635498 59004 635734
rect 58404 600054 59004 635498
rect 58404 599818 58586 600054
rect 58822 599818 59004 600054
rect 58404 599734 59004 599818
rect 58404 599498 58586 599734
rect 58822 599498 59004 599734
rect 58404 564054 59004 599498
rect 58404 563818 58586 564054
rect 58822 563818 59004 564054
rect 58404 563734 59004 563818
rect 58404 563498 58586 563734
rect 58822 563498 59004 563734
rect 58404 528054 59004 563498
rect 58404 527818 58586 528054
rect 58822 527818 59004 528054
rect 58404 527734 59004 527818
rect 58404 527498 58586 527734
rect 58822 527498 59004 527734
rect 58404 492054 59004 527498
rect 58404 491818 58586 492054
rect 58822 491818 59004 492054
rect 58404 491734 59004 491818
rect 58404 491498 58586 491734
rect 58822 491498 59004 491734
rect 58404 456054 59004 491498
rect 58404 455818 58586 456054
rect 58822 455818 59004 456054
rect 58404 455734 59004 455818
rect 58404 455498 58586 455734
rect 58822 455498 59004 455734
rect 58404 420054 59004 455498
rect 58404 419818 58586 420054
rect 58822 419818 59004 420054
rect 58404 419734 59004 419818
rect 58404 419498 58586 419734
rect 58822 419498 59004 419734
rect 58404 384054 59004 419498
rect 58404 383818 58586 384054
rect 58822 383818 59004 384054
rect 58404 383734 59004 383818
rect 58404 383498 58586 383734
rect 58822 383498 59004 383734
rect 58404 348054 59004 383498
rect 58404 347818 58586 348054
rect 58822 347818 59004 348054
rect 58404 347734 59004 347818
rect 58404 347498 58586 347734
rect 58822 347498 59004 347734
rect 58404 312054 59004 347498
rect 58404 311818 58586 312054
rect 58822 311818 59004 312054
rect 58404 311734 59004 311818
rect 58404 311498 58586 311734
rect 58822 311498 59004 311734
rect 58404 276054 59004 311498
rect 58404 275818 58586 276054
rect 58822 275818 59004 276054
rect 58404 275734 59004 275818
rect 58404 275498 58586 275734
rect 58822 275498 59004 275734
rect 58404 240054 59004 275498
rect 58404 239818 58586 240054
rect 58822 239818 59004 240054
rect 58404 239734 59004 239818
rect 58404 239498 58586 239734
rect 58822 239498 59004 239734
rect 58404 204054 59004 239498
rect 58404 203818 58586 204054
rect 58822 203818 59004 204054
rect 58404 203734 59004 203818
rect 58404 203498 58586 203734
rect 58822 203498 59004 203734
rect 58404 168054 59004 203498
rect 58404 167818 58586 168054
rect 58822 167818 59004 168054
rect 58404 167734 59004 167818
rect 58404 167498 58586 167734
rect 58822 167498 59004 167734
rect 58404 132054 59004 167498
rect 58404 131818 58586 132054
rect 58822 131818 59004 132054
rect 58404 131734 59004 131818
rect 58404 131498 58586 131734
rect 58822 131498 59004 131734
rect 58404 96054 59004 131498
rect 58404 95818 58586 96054
rect 58822 95818 59004 96054
rect 58404 95734 59004 95818
rect 58404 95498 58586 95734
rect 58822 95498 59004 95734
rect 58404 60054 59004 95498
rect 58404 59818 58586 60054
rect 58822 59818 59004 60054
rect 58404 59734 59004 59818
rect 58404 59498 58586 59734
rect 58822 59498 59004 59734
rect 58404 24054 59004 59498
rect 58404 23818 58586 24054
rect 58822 23818 59004 24054
rect 58404 23734 59004 23818
rect 58404 23498 58586 23734
rect 58822 23498 59004 23734
rect 58404 -3106 59004 23498
rect 58404 -3342 58586 -3106
rect 58822 -3342 59004 -3106
rect 58404 -3426 59004 -3342
rect 58404 -3662 58586 -3426
rect 58822 -3662 59004 -3426
rect 58404 -3684 59004 -3662
rect 62004 675654 62604 708882
rect 62004 675418 62186 675654
rect 62422 675418 62604 675654
rect 62004 675334 62604 675418
rect 62004 675098 62186 675334
rect 62422 675098 62604 675334
rect 62004 639654 62604 675098
rect 62004 639418 62186 639654
rect 62422 639418 62604 639654
rect 62004 639334 62604 639418
rect 62004 639098 62186 639334
rect 62422 639098 62604 639334
rect 62004 603654 62604 639098
rect 62004 603418 62186 603654
rect 62422 603418 62604 603654
rect 62004 603334 62604 603418
rect 62004 603098 62186 603334
rect 62422 603098 62604 603334
rect 62004 567654 62604 603098
rect 62004 567418 62186 567654
rect 62422 567418 62604 567654
rect 62004 567334 62604 567418
rect 62004 567098 62186 567334
rect 62422 567098 62604 567334
rect 62004 531654 62604 567098
rect 62004 531418 62186 531654
rect 62422 531418 62604 531654
rect 62004 531334 62604 531418
rect 62004 531098 62186 531334
rect 62422 531098 62604 531334
rect 62004 495654 62604 531098
rect 62004 495418 62186 495654
rect 62422 495418 62604 495654
rect 62004 495334 62604 495418
rect 62004 495098 62186 495334
rect 62422 495098 62604 495334
rect 62004 459654 62604 495098
rect 62004 459418 62186 459654
rect 62422 459418 62604 459654
rect 62004 459334 62604 459418
rect 62004 459098 62186 459334
rect 62422 459098 62604 459334
rect 62004 423654 62604 459098
rect 62004 423418 62186 423654
rect 62422 423418 62604 423654
rect 62004 423334 62604 423418
rect 62004 423098 62186 423334
rect 62422 423098 62604 423334
rect 62004 387654 62604 423098
rect 62004 387418 62186 387654
rect 62422 387418 62604 387654
rect 62004 387334 62604 387418
rect 62004 387098 62186 387334
rect 62422 387098 62604 387334
rect 62004 351654 62604 387098
rect 62004 351418 62186 351654
rect 62422 351418 62604 351654
rect 62004 351334 62604 351418
rect 62004 351098 62186 351334
rect 62422 351098 62604 351334
rect 62004 315654 62604 351098
rect 62004 315418 62186 315654
rect 62422 315418 62604 315654
rect 62004 315334 62604 315418
rect 62004 315098 62186 315334
rect 62422 315098 62604 315334
rect 62004 279654 62604 315098
rect 62004 279418 62186 279654
rect 62422 279418 62604 279654
rect 62004 279334 62604 279418
rect 62004 279098 62186 279334
rect 62422 279098 62604 279334
rect 62004 243654 62604 279098
rect 62004 243418 62186 243654
rect 62422 243418 62604 243654
rect 62004 243334 62604 243418
rect 62004 243098 62186 243334
rect 62422 243098 62604 243334
rect 62004 207654 62604 243098
rect 62004 207418 62186 207654
rect 62422 207418 62604 207654
rect 62004 207334 62604 207418
rect 62004 207098 62186 207334
rect 62422 207098 62604 207334
rect 62004 171654 62604 207098
rect 62004 171418 62186 171654
rect 62422 171418 62604 171654
rect 62004 171334 62604 171418
rect 62004 171098 62186 171334
rect 62422 171098 62604 171334
rect 62004 135654 62604 171098
rect 62004 135418 62186 135654
rect 62422 135418 62604 135654
rect 62004 135334 62604 135418
rect 62004 135098 62186 135334
rect 62422 135098 62604 135334
rect 62004 99654 62604 135098
rect 62004 99418 62186 99654
rect 62422 99418 62604 99654
rect 62004 99334 62604 99418
rect 62004 99098 62186 99334
rect 62422 99098 62604 99334
rect 62004 63654 62604 99098
rect 62004 63418 62186 63654
rect 62422 63418 62604 63654
rect 62004 63334 62604 63418
rect 62004 63098 62186 63334
rect 62422 63098 62604 63334
rect 62004 27654 62604 63098
rect 62004 27418 62186 27654
rect 62422 27418 62604 27654
rect 62004 27334 62604 27418
rect 62004 27098 62186 27334
rect 62422 27098 62604 27334
rect 62004 -4946 62604 27098
rect 62004 -5182 62186 -4946
rect 62422 -5182 62604 -4946
rect 62004 -5266 62604 -5182
rect 62004 -5502 62186 -5266
rect 62422 -5502 62604 -5266
rect 62004 -5524 62604 -5502
rect 65604 679254 66204 710722
rect 83604 710358 84204 711300
rect 83604 710122 83786 710358
rect 84022 710122 84204 710358
rect 83604 710038 84204 710122
rect 83604 709802 83786 710038
rect 84022 709802 84204 710038
rect 80004 708518 80604 709460
rect 80004 708282 80186 708518
rect 80422 708282 80604 708518
rect 80004 708198 80604 708282
rect 80004 707962 80186 708198
rect 80422 707962 80604 708198
rect 76404 706678 77004 707620
rect 76404 706442 76586 706678
rect 76822 706442 77004 706678
rect 76404 706358 77004 706442
rect 76404 706122 76586 706358
rect 76822 706122 77004 706358
rect 65604 679018 65786 679254
rect 66022 679018 66204 679254
rect 65604 678934 66204 679018
rect 65604 678698 65786 678934
rect 66022 678698 66204 678934
rect 65604 643254 66204 678698
rect 65604 643018 65786 643254
rect 66022 643018 66204 643254
rect 65604 642934 66204 643018
rect 65604 642698 65786 642934
rect 66022 642698 66204 642934
rect 65604 607254 66204 642698
rect 65604 607018 65786 607254
rect 66022 607018 66204 607254
rect 65604 606934 66204 607018
rect 65604 606698 65786 606934
rect 66022 606698 66204 606934
rect 65604 571254 66204 606698
rect 65604 571018 65786 571254
rect 66022 571018 66204 571254
rect 65604 570934 66204 571018
rect 65604 570698 65786 570934
rect 66022 570698 66204 570934
rect 65604 535254 66204 570698
rect 65604 535018 65786 535254
rect 66022 535018 66204 535254
rect 65604 534934 66204 535018
rect 65604 534698 65786 534934
rect 66022 534698 66204 534934
rect 65604 499254 66204 534698
rect 65604 499018 65786 499254
rect 66022 499018 66204 499254
rect 65604 498934 66204 499018
rect 65604 498698 65786 498934
rect 66022 498698 66204 498934
rect 65604 463254 66204 498698
rect 65604 463018 65786 463254
rect 66022 463018 66204 463254
rect 65604 462934 66204 463018
rect 65604 462698 65786 462934
rect 66022 462698 66204 462934
rect 65604 427254 66204 462698
rect 65604 427018 65786 427254
rect 66022 427018 66204 427254
rect 65604 426934 66204 427018
rect 65604 426698 65786 426934
rect 66022 426698 66204 426934
rect 65604 391254 66204 426698
rect 65604 391018 65786 391254
rect 66022 391018 66204 391254
rect 65604 390934 66204 391018
rect 65604 390698 65786 390934
rect 66022 390698 66204 390934
rect 65604 355254 66204 390698
rect 65604 355018 65786 355254
rect 66022 355018 66204 355254
rect 65604 354934 66204 355018
rect 65604 354698 65786 354934
rect 66022 354698 66204 354934
rect 65604 319254 66204 354698
rect 65604 319018 65786 319254
rect 66022 319018 66204 319254
rect 65604 318934 66204 319018
rect 65604 318698 65786 318934
rect 66022 318698 66204 318934
rect 65604 283254 66204 318698
rect 65604 283018 65786 283254
rect 66022 283018 66204 283254
rect 65604 282934 66204 283018
rect 65604 282698 65786 282934
rect 66022 282698 66204 282934
rect 65604 247254 66204 282698
rect 65604 247018 65786 247254
rect 66022 247018 66204 247254
rect 65604 246934 66204 247018
rect 65604 246698 65786 246934
rect 66022 246698 66204 246934
rect 65604 211254 66204 246698
rect 65604 211018 65786 211254
rect 66022 211018 66204 211254
rect 65604 210934 66204 211018
rect 65604 210698 65786 210934
rect 66022 210698 66204 210934
rect 65604 175254 66204 210698
rect 65604 175018 65786 175254
rect 66022 175018 66204 175254
rect 65604 174934 66204 175018
rect 65604 174698 65786 174934
rect 66022 174698 66204 174934
rect 65604 139254 66204 174698
rect 65604 139018 65786 139254
rect 66022 139018 66204 139254
rect 65604 138934 66204 139018
rect 65604 138698 65786 138934
rect 66022 138698 66204 138934
rect 65604 103254 66204 138698
rect 65604 103018 65786 103254
rect 66022 103018 66204 103254
rect 65604 102934 66204 103018
rect 65604 102698 65786 102934
rect 66022 102698 66204 102934
rect 65604 67254 66204 102698
rect 65604 67018 65786 67254
rect 66022 67018 66204 67254
rect 65604 66934 66204 67018
rect 65604 66698 65786 66934
rect 66022 66698 66204 66934
rect 65604 31254 66204 66698
rect 65604 31018 65786 31254
rect 66022 31018 66204 31254
rect 65604 30934 66204 31018
rect 65604 30698 65786 30934
rect 66022 30698 66204 30934
rect 47604 -6102 47786 -5866
rect 48022 -6102 48204 -5866
rect 47604 -6186 48204 -6102
rect 47604 -6422 47786 -6186
rect 48022 -6422 48204 -6186
rect 47604 -7364 48204 -6422
rect 65604 -6786 66204 30698
rect 72804 704838 73404 705780
rect 72804 704602 72986 704838
rect 73222 704602 73404 704838
rect 72804 704518 73404 704602
rect 72804 704282 72986 704518
rect 73222 704282 73404 704518
rect 72804 686454 73404 704282
rect 72804 686218 72986 686454
rect 73222 686218 73404 686454
rect 72804 686134 73404 686218
rect 72804 685898 72986 686134
rect 73222 685898 73404 686134
rect 72804 650454 73404 685898
rect 72804 650218 72986 650454
rect 73222 650218 73404 650454
rect 72804 650134 73404 650218
rect 72804 649898 72986 650134
rect 73222 649898 73404 650134
rect 72804 614454 73404 649898
rect 72804 614218 72986 614454
rect 73222 614218 73404 614454
rect 72804 614134 73404 614218
rect 72804 613898 72986 614134
rect 73222 613898 73404 614134
rect 72804 578454 73404 613898
rect 72804 578218 72986 578454
rect 73222 578218 73404 578454
rect 72804 578134 73404 578218
rect 72804 577898 72986 578134
rect 73222 577898 73404 578134
rect 72804 542454 73404 577898
rect 72804 542218 72986 542454
rect 73222 542218 73404 542454
rect 72804 542134 73404 542218
rect 72804 541898 72986 542134
rect 73222 541898 73404 542134
rect 72804 506454 73404 541898
rect 72804 506218 72986 506454
rect 73222 506218 73404 506454
rect 72804 506134 73404 506218
rect 72804 505898 72986 506134
rect 73222 505898 73404 506134
rect 72804 470454 73404 505898
rect 72804 470218 72986 470454
rect 73222 470218 73404 470454
rect 72804 470134 73404 470218
rect 72804 469898 72986 470134
rect 73222 469898 73404 470134
rect 72804 434454 73404 469898
rect 72804 434218 72986 434454
rect 73222 434218 73404 434454
rect 72804 434134 73404 434218
rect 72804 433898 72986 434134
rect 73222 433898 73404 434134
rect 72804 398454 73404 433898
rect 72804 398218 72986 398454
rect 73222 398218 73404 398454
rect 72804 398134 73404 398218
rect 72804 397898 72986 398134
rect 73222 397898 73404 398134
rect 72804 362454 73404 397898
rect 72804 362218 72986 362454
rect 73222 362218 73404 362454
rect 72804 362134 73404 362218
rect 72804 361898 72986 362134
rect 73222 361898 73404 362134
rect 72804 326454 73404 361898
rect 72804 326218 72986 326454
rect 73222 326218 73404 326454
rect 72804 326134 73404 326218
rect 72804 325898 72986 326134
rect 73222 325898 73404 326134
rect 72804 290454 73404 325898
rect 72804 290218 72986 290454
rect 73222 290218 73404 290454
rect 72804 290134 73404 290218
rect 72804 289898 72986 290134
rect 73222 289898 73404 290134
rect 72804 254454 73404 289898
rect 72804 254218 72986 254454
rect 73222 254218 73404 254454
rect 72804 254134 73404 254218
rect 72804 253898 72986 254134
rect 73222 253898 73404 254134
rect 72804 218454 73404 253898
rect 72804 218218 72986 218454
rect 73222 218218 73404 218454
rect 72804 218134 73404 218218
rect 72804 217898 72986 218134
rect 73222 217898 73404 218134
rect 72804 182454 73404 217898
rect 72804 182218 72986 182454
rect 73222 182218 73404 182454
rect 72804 182134 73404 182218
rect 72804 181898 72986 182134
rect 73222 181898 73404 182134
rect 72804 146454 73404 181898
rect 72804 146218 72986 146454
rect 73222 146218 73404 146454
rect 72804 146134 73404 146218
rect 72804 145898 72986 146134
rect 73222 145898 73404 146134
rect 72804 110454 73404 145898
rect 72804 110218 72986 110454
rect 73222 110218 73404 110454
rect 72804 110134 73404 110218
rect 72804 109898 72986 110134
rect 73222 109898 73404 110134
rect 72804 74454 73404 109898
rect 72804 74218 72986 74454
rect 73222 74218 73404 74454
rect 72804 74134 73404 74218
rect 72804 73898 72986 74134
rect 73222 73898 73404 74134
rect 72804 38454 73404 73898
rect 72804 38218 72986 38454
rect 73222 38218 73404 38454
rect 72804 38134 73404 38218
rect 72804 37898 72986 38134
rect 73222 37898 73404 38134
rect 72804 2454 73404 37898
rect 72804 2218 72986 2454
rect 73222 2218 73404 2454
rect 72804 2134 73404 2218
rect 72804 1898 72986 2134
rect 73222 1898 73404 2134
rect 72804 -346 73404 1898
rect 72804 -582 72986 -346
rect 73222 -582 73404 -346
rect 72804 -666 73404 -582
rect 72804 -902 72986 -666
rect 73222 -902 73404 -666
rect 72804 -1844 73404 -902
rect 76404 690054 77004 706122
rect 76404 689818 76586 690054
rect 76822 689818 77004 690054
rect 76404 689734 77004 689818
rect 76404 689498 76586 689734
rect 76822 689498 77004 689734
rect 76404 654054 77004 689498
rect 76404 653818 76586 654054
rect 76822 653818 77004 654054
rect 76404 653734 77004 653818
rect 76404 653498 76586 653734
rect 76822 653498 77004 653734
rect 76404 618054 77004 653498
rect 76404 617818 76586 618054
rect 76822 617818 77004 618054
rect 76404 617734 77004 617818
rect 76404 617498 76586 617734
rect 76822 617498 77004 617734
rect 76404 582054 77004 617498
rect 76404 581818 76586 582054
rect 76822 581818 77004 582054
rect 76404 581734 77004 581818
rect 76404 581498 76586 581734
rect 76822 581498 77004 581734
rect 76404 546054 77004 581498
rect 76404 545818 76586 546054
rect 76822 545818 77004 546054
rect 76404 545734 77004 545818
rect 76404 545498 76586 545734
rect 76822 545498 77004 545734
rect 76404 510054 77004 545498
rect 76404 509818 76586 510054
rect 76822 509818 77004 510054
rect 76404 509734 77004 509818
rect 76404 509498 76586 509734
rect 76822 509498 77004 509734
rect 76404 474054 77004 509498
rect 76404 473818 76586 474054
rect 76822 473818 77004 474054
rect 76404 473734 77004 473818
rect 76404 473498 76586 473734
rect 76822 473498 77004 473734
rect 76404 438054 77004 473498
rect 76404 437818 76586 438054
rect 76822 437818 77004 438054
rect 76404 437734 77004 437818
rect 76404 437498 76586 437734
rect 76822 437498 77004 437734
rect 76404 402054 77004 437498
rect 76404 401818 76586 402054
rect 76822 401818 77004 402054
rect 76404 401734 77004 401818
rect 76404 401498 76586 401734
rect 76822 401498 77004 401734
rect 76404 366054 77004 401498
rect 76404 365818 76586 366054
rect 76822 365818 77004 366054
rect 76404 365734 77004 365818
rect 76404 365498 76586 365734
rect 76822 365498 77004 365734
rect 76404 330054 77004 365498
rect 76404 329818 76586 330054
rect 76822 329818 77004 330054
rect 76404 329734 77004 329818
rect 76404 329498 76586 329734
rect 76822 329498 77004 329734
rect 76404 294054 77004 329498
rect 76404 293818 76586 294054
rect 76822 293818 77004 294054
rect 76404 293734 77004 293818
rect 76404 293498 76586 293734
rect 76822 293498 77004 293734
rect 76404 258054 77004 293498
rect 76404 257818 76586 258054
rect 76822 257818 77004 258054
rect 76404 257734 77004 257818
rect 76404 257498 76586 257734
rect 76822 257498 77004 257734
rect 76404 222054 77004 257498
rect 76404 221818 76586 222054
rect 76822 221818 77004 222054
rect 76404 221734 77004 221818
rect 76404 221498 76586 221734
rect 76822 221498 77004 221734
rect 76404 186054 77004 221498
rect 76404 185818 76586 186054
rect 76822 185818 77004 186054
rect 76404 185734 77004 185818
rect 76404 185498 76586 185734
rect 76822 185498 77004 185734
rect 76404 150054 77004 185498
rect 76404 149818 76586 150054
rect 76822 149818 77004 150054
rect 76404 149734 77004 149818
rect 76404 149498 76586 149734
rect 76822 149498 77004 149734
rect 76404 114054 77004 149498
rect 76404 113818 76586 114054
rect 76822 113818 77004 114054
rect 76404 113734 77004 113818
rect 76404 113498 76586 113734
rect 76822 113498 77004 113734
rect 76404 78054 77004 113498
rect 76404 77818 76586 78054
rect 76822 77818 77004 78054
rect 76404 77734 77004 77818
rect 76404 77498 76586 77734
rect 76822 77498 77004 77734
rect 76404 42054 77004 77498
rect 76404 41818 76586 42054
rect 76822 41818 77004 42054
rect 76404 41734 77004 41818
rect 76404 41498 76586 41734
rect 76822 41498 77004 41734
rect 76404 6054 77004 41498
rect 76404 5818 76586 6054
rect 76822 5818 77004 6054
rect 76404 5734 77004 5818
rect 76404 5498 76586 5734
rect 76822 5498 77004 5734
rect 76404 -2186 77004 5498
rect 76404 -2422 76586 -2186
rect 76822 -2422 77004 -2186
rect 76404 -2506 77004 -2422
rect 76404 -2742 76586 -2506
rect 76822 -2742 77004 -2506
rect 76404 -3684 77004 -2742
rect 80004 693654 80604 707962
rect 80004 693418 80186 693654
rect 80422 693418 80604 693654
rect 80004 693334 80604 693418
rect 80004 693098 80186 693334
rect 80422 693098 80604 693334
rect 80004 657654 80604 693098
rect 80004 657418 80186 657654
rect 80422 657418 80604 657654
rect 80004 657334 80604 657418
rect 80004 657098 80186 657334
rect 80422 657098 80604 657334
rect 80004 621654 80604 657098
rect 80004 621418 80186 621654
rect 80422 621418 80604 621654
rect 80004 621334 80604 621418
rect 80004 621098 80186 621334
rect 80422 621098 80604 621334
rect 80004 585654 80604 621098
rect 80004 585418 80186 585654
rect 80422 585418 80604 585654
rect 80004 585334 80604 585418
rect 80004 585098 80186 585334
rect 80422 585098 80604 585334
rect 80004 549654 80604 585098
rect 80004 549418 80186 549654
rect 80422 549418 80604 549654
rect 80004 549334 80604 549418
rect 80004 549098 80186 549334
rect 80422 549098 80604 549334
rect 80004 513654 80604 549098
rect 80004 513418 80186 513654
rect 80422 513418 80604 513654
rect 80004 513334 80604 513418
rect 80004 513098 80186 513334
rect 80422 513098 80604 513334
rect 80004 477654 80604 513098
rect 80004 477418 80186 477654
rect 80422 477418 80604 477654
rect 80004 477334 80604 477418
rect 80004 477098 80186 477334
rect 80422 477098 80604 477334
rect 80004 441654 80604 477098
rect 80004 441418 80186 441654
rect 80422 441418 80604 441654
rect 80004 441334 80604 441418
rect 80004 441098 80186 441334
rect 80422 441098 80604 441334
rect 80004 405654 80604 441098
rect 80004 405418 80186 405654
rect 80422 405418 80604 405654
rect 80004 405334 80604 405418
rect 80004 405098 80186 405334
rect 80422 405098 80604 405334
rect 80004 369654 80604 405098
rect 80004 369418 80186 369654
rect 80422 369418 80604 369654
rect 80004 369334 80604 369418
rect 80004 369098 80186 369334
rect 80422 369098 80604 369334
rect 80004 333654 80604 369098
rect 80004 333418 80186 333654
rect 80422 333418 80604 333654
rect 80004 333334 80604 333418
rect 80004 333098 80186 333334
rect 80422 333098 80604 333334
rect 80004 297654 80604 333098
rect 80004 297418 80186 297654
rect 80422 297418 80604 297654
rect 80004 297334 80604 297418
rect 80004 297098 80186 297334
rect 80422 297098 80604 297334
rect 80004 261654 80604 297098
rect 80004 261418 80186 261654
rect 80422 261418 80604 261654
rect 80004 261334 80604 261418
rect 80004 261098 80186 261334
rect 80422 261098 80604 261334
rect 80004 225654 80604 261098
rect 80004 225418 80186 225654
rect 80422 225418 80604 225654
rect 80004 225334 80604 225418
rect 80004 225098 80186 225334
rect 80422 225098 80604 225334
rect 80004 189654 80604 225098
rect 80004 189418 80186 189654
rect 80422 189418 80604 189654
rect 80004 189334 80604 189418
rect 80004 189098 80186 189334
rect 80422 189098 80604 189334
rect 80004 153654 80604 189098
rect 80004 153418 80186 153654
rect 80422 153418 80604 153654
rect 80004 153334 80604 153418
rect 80004 153098 80186 153334
rect 80422 153098 80604 153334
rect 80004 117654 80604 153098
rect 80004 117418 80186 117654
rect 80422 117418 80604 117654
rect 80004 117334 80604 117418
rect 80004 117098 80186 117334
rect 80422 117098 80604 117334
rect 80004 81654 80604 117098
rect 80004 81418 80186 81654
rect 80422 81418 80604 81654
rect 80004 81334 80604 81418
rect 80004 81098 80186 81334
rect 80422 81098 80604 81334
rect 80004 45654 80604 81098
rect 80004 45418 80186 45654
rect 80422 45418 80604 45654
rect 80004 45334 80604 45418
rect 80004 45098 80186 45334
rect 80422 45098 80604 45334
rect 80004 9654 80604 45098
rect 80004 9418 80186 9654
rect 80422 9418 80604 9654
rect 80004 9334 80604 9418
rect 80004 9098 80186 9334
rect 80422 9098 80604 9334
rect 80004 -4026 80604 9098
rect 80004 -4262 80186 -4026
rect 80422 -4262 80604 -4026
rect 80004 -4346 80604 -4262
rect 80004 -4582 80186 -4346
rect 80422 -4582 80604 -4346
rect 80004 -5524 80604 -4582
rect 83604 697254 84204 709802
rect 101604 711278 102204 711300
rect 101604 711042 101786 711278
rect 102022 711042 102204 711278
rect 101604 710958 102204 711042
rect 101604 710722 101786 710958
rect 102022 710722 102204 710958
rect 98004 709438 98604 709460
rect 98004 709202 98186 709438
rect 98422 709202 98604 709438
rect 98004 709118 98604 709202
rect 98004 708882 98186 709118
rect 98422 708882 98604 709118
rect 94404 707598 95004 707620
rect 94404 707362 94586 707598
rect 94822 707362 95004 707598
rect 94404 707278 95004 707362
rect 94404 707042 94586 707278
rect 94822 707042 95004 707278
rect 83604 697018 83786 697254
rect 84022 697018 84204 697254
rect 83604 696934 84204 697018
rect 83604 696698 83786 696934
rect 84022 696698 84204 696934
rect 83604 661254 84204 696698
rect 83604 661018 83786 661254
rect 84022 661018 84204 661254
rect 83604 660934 84204 661018
rect 83604 660698 83786 660934
rect 84022 660698 84204 660934
rect 83604 625254 84204 660698
rect 83604 625018 83786 625254
rect 84022 625018 84204 625254
rect 83604 624934 84204 625018
rect 83604 624698 83786 624934
rect 84022 624698 84204 624934
rect 83604 589254 84204 624698
rect 83604 589018 83786 589254
rect 84022 589018 84204 589254
rect 83604 588934 84204 589018
rect 83604 588698 83786 588934
rect 84022 588698 84204 588934
rect 83604 553254 84204 588698
rect 83604 553018 83786 553254
rect 84022 553018 84204 553254
rect 83604 552934 84204 553018
rect 83604 552698 83786 552934
rect 84022 552698 84204 552934
rect 83604 517254 84204 552698
rect 83604 517018 83786 517254
rect 84022 517018 84204 517254
rect 83604 516934 84204 517018
rect 83604 516698 83786 516934
rect 84022 516698 84204 516934
rect 83604 481254 84204 516698
rect 83604 481018 83786 481254
rect 84022 481018 84204 481254
rect 83604 480934 84204 481018
rect 83604 480698 83786 480934
rect 84022 480698 84204 480934
rect 83604 445254 84204 480698
rect 83604 445018 83786 445254
rect 84022 445018 84204 445254
rect 83604 444934 84204 445018
rect 83604 444698 83786 444934
rect 84022 444698 84204 444934
rect 83604 409254 84204 444698
rect 83604 409018 83786 409254
rect 84022 409018 84204 409254
rect 83604 408934 84204 409018
rect 83604 408698 83786 408934
rect 84022 408698 84204 408934
rect 83604 373254 84204 408698
rect 83604 373018 83786 373254
rect 84022 373018 84204 373254
rect 83604 372934 84204 373018
rect 83604 372698 83786 372934
rect 84022 372698 84204 372934
rect 83604 337254 84204 372698
rect 83604 337018 83786 337254
rect 84022 337018 84204 337254
rect 83604 336934 84204 337018
rect 83604 336698 83786 336934
rect 84022 336698 84204 336934
rect 83604 301254 84204 336698
rect 83604 301018 83786 301254
rect 84022 301018 84204 301254
rect 83604 300934 84204 301018
rect 83604 300698 83786 300934
rect 84022 300698 84204 300934
rect 83604 265254 84204 300698
rect 83604 265018 83786 265254
rect 84022 265018 84204 265254
rect 83604 264934 84204 265018
rect 83604 264698 83786 264934
rect 84022 264698 84204 264934
rect 83604 229254 84204 264698
rect 83604 229018 83786 229254
rect 84022 229018 84204 229254
rect 83604 228934 84204 229018
rect 83604 228698 83786 228934
rect 84022 228698 84204 228934
rect 83604 193254 84204 228698
rect 83604 193018 83786 193254
rect 84022 193018 84204 193254
rect 83604 192934 84204 193018
rect 83604 192698 83786 192934
rect 84022 192698 84204 192934
rect 83604 157254 84204 192698
rect 83604 157018 83786 157254
rect 84022 157018 84204 157254
rect 83604 156934 84204 157018
rect 83604 156698 83786 156934
rect 84022 156698 84204 156934
rect 83604 121254 84204 156698
rect 83604 121018 83786 121254
rect 84022 121018 84204 121254
rect 83604 120934 84204 121018
rect 83604 120698 83786 120934
rect 84022 120698 84204 120934
rect 83604 85254 84204 120698
rect 83604 85018 83786 85254
rect 84022 85018 84204 85254
rect 83604 84934 84204 85018
rect 83604 84698 83786 84934
rect 84022 84698 84204 84934
rect 83604 49254 84204 84698
rect 83604 49018 83786 49254
rect 84022 49018 84204 49254
rect 83604 48934 84204 49018
rect 83604 48698 83786 48934
rect 84022 48698 84204 48934
rect 83604 13254 84204 48698
rect 83604 13018 83786 13254
rect 84022 13018 84204 13254
rect 83604 12934 84204 13018
rect 83604 12698 83786 12934
rect 84022 12698 84204 12934
rect 65604 -7022 65786 -6786
rect 66022 -7022 66204 -6786
rect 65604 -7106 66204 -7022
rect 65604 -7342 65786 -7106
rect 66022 -7342 66204 -7106
rect 65604 -7364 66204 -7342
rect 83604 -5866 84204 12698
rect 90804 705758 91404 705780
rect 90804 705522 90986 705758
rect 91222 705522 91404 705758
rect 90804 705438 91404 705522
rect 90804 705202 90986 705438
rect 91222 705202 91404 705438
rect 90804 668454 91404 705202
rect 90804 668218 90986 668454
rect 91222 668218 91404 668454
rect 90804 668134 91404 668218
rect 90804 667898 90986 668134
rect 91222 667898 91404 668134
rect 90804 632454 91404 667898
rect 90804 632218 90986 632454
rect 91222 632218 91404 632454
rect 90804 632134 91404 632218
rect 90804 631898 90986 632134
rect 91222 631898 91404 632134
rect 90804 596454 91404 631898
rect 90804 596218 90986 596454
rect 91222 596218 91404 596454
rect 90804 596134 91404 596218
rect 90804 595898 90986 596134
rect 91222 595898 91404 596134
rect 90804 560454 91404 595898
rect 90804 560218 90986 560454
rect 91222 560218 91404 560454
rect 90804 560134 91404 560218
rect 90804 559898 90986 560134
rect 91222 559898 91404 560134
rect 90804 524454 91404 559898
rect 90804 524218 90986 524454
rect 91222 524218 91404 524454
rect 90804 524134 91404 524218
rect 90804 523898 90986 524134
rect 91222 523898 91404 524134
rect 90804 488454 91404 523898
rect 90804 488218 90986 488454
rect 91222 488218 91404 488454
rect 90804 488134 91404 488218
rect 90804 487898 90986 488134
rect 91222 487898 91404 488134
rect 90804 452454 91404 487898
rect 90804 452218 90986 452454
rect 91222 452218 91404 452454
rect 90804 452134 91404 452218
rect 90804 451898 90986 452134
rect 91222 451898 91404 452134
rect 90804 416454 91404 451898
rect 90804 416218 90986 416454
rect 91222 416218 91404 416454
rect 90804 416134 91404 416218
rect 90804 415898 90986 416134
rect 91222 415898 91404 416134
rect 90804 380454 91404 415898
rect 90804 380218 90986 380454
rect 91222 380218 91404 380454
rect 90804 380134 91404 380218
rect 90804 379898 90986 380134
rect 91222 379898 91404 380134
rect 90804 344454 91404 379898
rect 90804 344218 90986 344454
rect 91222 344218 91404 344454
rect 90804 344134 91404 344218
rect 90804 343898 90986 344134
rect 91222 343898 91404 344134
rect 90804 308454 91404 343898
rect 90804 308218 90986 308454
rect 91222 308218 91404 308454
rect 90804 308134 91404 308218
rect 90804 307898 90986 308134
rect 91222 307898 91404 308134
rect 90804 272454 91404 307898
rect 90804 272218 90986 272454
rect 91222 272218 91404 272454
rect 90804 272134 91404 272218
rect 90804 271898 90986 272134
rect 91222 271898 91404 272134
rect 90804 236454 91404 271898
rect 90804 236218 90986 236454
rect 91222 236218 91404 236454
rect 90804 236134 91404 236218
rect 90804 235898 90986 236134
rect 91222 235898 91404 236134
rect 90804 200454 91404 235898
rect 90804 200218 90986 200454
rect 91222 200218 91404 200454
rect 90804 200134 91404 200218
rect 90804 199898 90986 200134
rect 91222 199898 91404 200134
rect 90804 164454 91404 199898
rect 90804 164218 90986 164454
rect 91222 164218 91404 164454
rect 90804 164134 91404 164218
rect 90804 163898 90986 164134
rect 91222 163898 91404 164134
rect 90804 128454 91404 163898
rect 90804 128218 90986 128454
rect 91222 128218 91404 128454
rect 90804 128134 91404 128218
rect 90804 127898 90986 128134
rect 91222 127898 91404 128134
rect 90804 92454 91404 127898
rect 90804 92218 90986 92454
rect 91222 92218 91404 92454
rect 90804 92134 91404 92218
rect 90804 91898 90986 92134
rect 91222 91898 91404 92134
rect 90804 56454 91404 91898
rect 90804 56218 90986 56454
rect 91222 56218 91404 56454
rect 90804 56134 91404 56218
rect 90804 55898 90986 56134
rect 91222 55898 91404 56134
rect 90804 20454 91404 55898
rect 90804 20218 90986 20454
rect 91222 20218 91404 20454
rect 90804 20134 91404 20218
rect 90804 19898 90986 20134
rect 91222 19898 91404 20134
rect 90804 -1266 91404 19898
rect 90804 -1502 90986 -1266
rect 91222 -1502 91404 -1266
rect 90804 -1586 91404 -1502
rect 90804 -1822 90986 -1586
rect 91222 -1822 91404 -1586
rect 90804 -1844 91404 -1822
rect 94404 672054 95004 707042
rect 94404 671818 94586 672054
rect 94822 671818 95004 672054
rect 94404 671734 95004 671818
rect 94404 671498 94586 671734
rect 94822 671498 95004 671734
rect 94404 636054 95004 671498
rect 94404 635818 94586 636054
rect 94822 635818 95004 636054
rect 94404 635734 95004 635818
rect 94404 635498 94586 635734
rect 94822 635498 95004 635734
rect 94404 600054 95004 635498
rect 94404 599818 94586 600054
rect 94822 599818 95004 600054
rect 94404 599734 95004 599818
rect 94404 599498 94586 599734
rect 94822 599498 95004 599734
rect 94404 564054 95004 599498
rect 94404 563818 94586 564054
rect 94822 563818 95004 564054
rect 94404 563734 95004 563818
rect 94404 563498 94586 563734
rect 94822 563498 95004 563734
rect 94404 528054 95004 563498
rect 94404 527818 94586 528054
rect 94822 527818 95004 528054
rect 94404 527734 95004 527818
rect 94404 527498 94586 527734
rect 94822 527498 95004 527734
rect 94404 492054 95004 527498
rect 94404 491818 94586 492054
rect 94822 491818 95004 492054
rect 94404 491734 95004 491818
rect 94404 491498 94586 491734
rect 94822 491498 95004 491734
rect 94404 456054 95004 491498
rect 94404 455818 94586 456054
rect 94822 455818 95004 456054
rect 94404 455734 95004 455818
rect 94404 455498 94586 455734
rect 94822 455498 95004 455734
rect 94404 420054 95004 455498
rect 94404 419818 94586 420054
rect 94822 419818 95004 420054
rect 94404 419734 95004 419818
rect 94404 419498 94586 419734
rect 94822 419498 95004 419734
rect 94404 384054 95004 419498
rect 94404 383818 94586 384054
rect 94822 383818 95004 384054
rect 94404 383734 95004 383818
rect 94404 383498 94586 383734
rect 94822 383498 95004 383734
rect 94404 348054 95004 383498
rect 94404 347818 94586 348054
rect 94822 347818 95004 348054
rect 94404 347734 95004 347818
rect 94404 347498 94586 347734
rect 94822 347498 95004 347734
rect 94404 312054 95004 347498
rect 94404 311818 94586 312054
rect 94822 311818 95004 312054
rect 94404 311734 95004 311818
rect 94404 311498 94586 311734
rect 94822 311498 95004 311734
rect 94404 276054 95004 311498
rect 94404 275818 94586 276054
rect 94822 275818 95004 276054
rect 94404 275734 95004 275818
rect 94404 275498 94586 275734
rect 94822 275498 95004 275734
rect 94404 240054 95004 275498
rect 94404 239818 94586 240054
rect 94822 239818 95004 240054
rect 94404 239734 95004 239818
rect 94404 239498 94586 239734
rect 94822 239498 95004 239734
rect 94404 204054 95004 239498
rect 94404 203818 94586 204054
rect 94822 203818 95004 204054
rect 94404 203734 95004 203818
rect 94404 203498 94586 203734
rect 94822 203498 95004 203734
rect 94404 168054 95004 203498
rect 94404 167818 94586 168054
rect 94822 167818 95004 168054
rect 94404 167734 95004 167818
rect 94404 167498 94586 167734
rect 94822 167498 95004 167734
rect 94404 132054 95004 167498
rect 94404 131818 94586 132054
rect 94822 131818 95004 132054
rect 94404 131734 95004 131818
rect 94404 131498 94586 131734
rect 94822 131498 95004 131734
rect 94404 96054 95004 131498
rect 94404 95818 94586 96054
rect 94822 95818 95004 96054
rect 94404 95734 95004 95818
rect 94404 95498 94586 95734
rect 94822 95498 95004 95734
rect 94404 60054 95004 95498
rect 94404 59818 94586 60054
rect 94822 59818 95004 60054
rect 94404 59734 95004 59818
rect 94404 59498 94586 59734
rect 94822 59498 95004 59734
rect 94404 24054 95004 59498
rect 94404 23818 94586 24054
rect 94822 23818 95004 24054
rect 94404 23734 95004 23818
rect 94404 23498 94586 23734
rect 94822 23498 95004 23734
rect 94404 -3106 95004 23498
rect 94404 -3342 94586 -3106
rect 94822 -3342 95004 -3106
rect 94404 -3426 95004 -3342
rect 94404 -3662 94586 -3426
rect 94822 -3662 95004 -3426
rect 94404 -3684 95004 -3662
rect 98004 675654 98604 708882
rect 98004 675418 98186 675654
rect 98422 675418 98604 675654
rect 98004 675334 98604 675418
rect 98004 675098 98186 675334
rect 98422 675098 98604 675334
rect 98004 639654 98604 675098
rect 98004 639418 98186 639654
rect 98422 639418 98604 639654
rect 98004 639334 98604 639418
rect 98004 639098 98186 639334
rect 98422 639098 98604 639334
rect 98004 603654 98604 639098
rect 98004 603418 98186 603654
rect 98422 603418 98604 603654
rect 98004 603334 98604 603418
rect 98004 603098 98186 603334
rect 98422 603098 98604 603334
rect 98004 567654 98604 603098
rect 98004 567418 98186 567654
rect 98422 567418 98604 567654
rect 98004 567334 98604 567418
rect 98004 567098 98186 567334
rect 98422 567098 98604 567334
rect 98004 531654 98604 567098
rect 98004 531418 98186 531654
rect 98422 531418 98604 531654
rect 98004 531334 98604 531418
rect 98004 531098 98186 531334
rect 98422 531098 98604 531334
rect 98004 495654 98604 531098
rect 98004 495418 98186 495654
rect 98422 495418 98604 495654
rect 98004 495334 98604 495418
rect 98004 495098 98186 495334
rect 98422 495098 98604 495334
rect 98004 459654 98604 495098
rect 98004 459418 98186 459654
rect 98422 459418 98604 459654
rect 98004 459334 98604 459418
rect 98004 459098 98186 459334
rect 98422 459098 98604 459334
rect 98004 423654 98604 459098
rect 98004 423418 98186 423654
rect 98422 423418 98604 423654
rect 98004 423334 98604 423418
rect 98004 423098 98186 423334
rect 98422 423098 98604 423334
rect 98004 387654 98604 423098
rect 98004 387418 98186 387654
rect 98422 387418 98604 387654
rect 98004 387334 98604 387418
rect 98004 387098 98186 387334
rect 98422 387098 98604 387334
rect 98004 351654 98604 387098
rect 98004 351418 98186 351654
rect 98422 351418 98604 351654
rect 98004 351334 98604 351418
rect 98004 351098 98186 351334
rect 98422 351098 98604 351334
rect 98004 315654 98604 351098
rect 98004 315418 98186 315654
rect 98422 315418 98604 315654
rect 98004 315334 98604 315418
rect 98004 315098 98186 315334
rect 98422 315098 98604 315334
rect 98004 279654 98604 315098
rect 98004 279418 98186 279654
rect 98422 279418 98604 279654
rect 98004 279334 98604 279418
rect 98004 279098 98186 279334
rect 98422 279098 98604 279334
rect 98004 243654 98604 279098
rect 98004 243418 98186 243654
rect 98422 243418 98604 243654
rect 98004 243334 98604 243418
rect 98004 243098 98186 243334
rect 98422 243098 98604 243334
rect 98004 207654 98604 243098
rect 98004 207418 98186 207654
rect 98422 207418 98604 207654
rect 98004 207334 98604 207418
rect 98004 207098 98186 207334
rect 98422 207098 98604 207334
rect 98004 171654 98604 207098
rect 98004 171418 98186 171654
rect 98422 171418 98604 171654
rect 98004 171334 98604 171418
rect 98004 171098 98186 171334
rect 98422 171098 98604 171334
rect 98004 135654 98604 171098
rect 98004 135418 98186 135654
rect 98422 135418 98604 135654
rect 98004 135334 98604 135418
rect 98004 135098 98186 135334
rect 98422 135098 98604 135334
rect 98004 99654 98604 135098
rect 98004 99418 98186 99654
rect 98422 99418 98604 99654
rect 98004 99334 98604 99418
rect 98004 99098 98186 99334
rect 98422 99098 98604 99334
rect 98004 63654 98604 99098
rect 98004 63418 98186 63654
rect 98422 63418 98604 63654
rect 98004 63334 98604 63418
rect 98004 63098 98186 63334
rect 98422 63098 98604 63334
rect 98004 27654 98604 63098
rect 98004 27418 98186 27654
rect 98422 27418 98604 27654
rect 98004 27334 98604 27418
rect 98004 27098 98186 27334
rect 98422 27098 98604 27334
rect 98004 -4946 98604 27098
rect 98004 -5182 98186 -4946
rect 98422 -5182 98604 -4946
rect 98004 -5266 98604 -5182
rect 98004 -5502 98186 -5266
rect 98422 -5502 98604 -5266
rect 98004 -5524 98604 -5502
rect 101604 679254 102204 710722
rect 119604 710358 120204 711300
rect 119604 710122 119786 710358
rect 120022 710122 120204 710358
rect 119604 710038 120204 710122
rect 119604 709802 119786 710038
rect 120022 709802 120204 710038
rect 116004 708518 116604 709460
rect 116004 708282 116186 708518
rect 116422 708282 116604 708518
rect 116004 708198 116604 708282
rect 116004 707962 116186 708198
rect 116422 707962 116604 708198
rect 112404 706678 113004 707620
rect 112404 706442 112586 706678
rect 112822 706442 113004 706678
rect 112404 706358 113004 706442
rect 112404 706122 112586 706358
rect 112822 706122 113004 706358
rect 101604 679018 101786 679254
rect 102022 679018 102204 679254
rect 101604 678934 102204 679018
rect 101604 678698 101786 678934
rect 102022 678698 102204 678934
rect 101604 643254 102204 678698
rect 101604 643018 101786 643254
rect 102022 643018 102204 643254
rect 101604 642934 102204 643018
rect 101604 642698 101786 642934
rect 102022 642698 102204 642934
rect 101604 607254 102204 642698
rect 101604 607018 101786 607254
rect 102022 607018 102204 607254
rect 101604 606934 102204 607018
rect 101604 606698 101786 606934
rect 102022 606698 102204 606934
rect 101604 571254 102204 606698
rect 101604 571018 101786 571254
rect 102022 571018 102204 571254
rect 101604 570934 102204 571018
rect 101604 570698 101786 570934
rect 102022 570698 102204 570934
rect 101604 535254 102204 570698
rect 101604 535018 101786 535254
rect 102022 535018 102204 535254
rect 101604 534934 102204 535018
rect 101604 534698 101786 534934
rect 102022 534698 102204 534934
rect 101604 499254 102204 534698
rect 101604 499018 101786 499254
rect 102022 499018 102204 499254
rect 101604 498934 102204 499018
rect 101604 498698 101786 498934
rect 102022 498698 102204 498934
rect 101604 463254 102204 498698
rect 101604 463018 101786 463254
rect 102022 463018 102204 463254
rect 101604 462934 102204 463018
rect 101604 462698 101786 462934
rect 102022 462698 102204 462934
rect 101604 427254 102204 462698
rect 101604 427018 101786 427254
rect 102022 427018 102204 427254
rect 101604 426934 102204 427018
rect 101604 426698 101786 426934
rect 102022 426698 102204 426934
rect 101604 391254 102204 426698
rect 101604 391018 101786 391254
rect 102022 391018 102204 391254
rect 101604 390934 102204 391018
rect 101604 390698 101786 390934
rect 102022 390698 102204 390934
rect 101604 355254 102204 390698
rect 101604 355018 101786 355254
rect 102022 355018 102204 355254
rect 101604 354934 102204 355018
rect 101604 354698 101786 354934
rect 102022 354698 102204 354934
rect 101604 319254 102204 354698
rect 101604 319018 101786 319254
rect 102022 319018 102204 319254
rect 101604 318934 102204 319018
rect 101604 318698 101786 318934
rect 102022 318698 102204 318934
rect 101604 283254 102204 318698
rect 101604 283018 101786 283254
rect 102022 283018 102204 283254
rect 101604 282934 102204 283018
rect 101604 282698 101786 282934
rect 102022 282698 102204 282934
rect 101604 247254 102204 282698
rect 101604 247018 101786 247254
rect 102022 247018 102204 247254
rect 101604 246934 102204 247018
rect 101604 246698 101786 246934
rect 102022 246698 102204 246934
rect 101604 211254 102204 246698
rect 101604 211018 101786 211254
rect 102022 211018 102204 211254
rect 101604 210934 102204 211018
rect 101604 210698 101786 210934
rect 102022 210698 102204 210934
rect 101604 175254 102204 210698
rect 101604 175018 101786 175254
rect 102022 175018 102204 175254
rect 101604 174934 102204 175018
rect 101604 174698 101786 174934
rect 102022 174698 102204 174934
rect 101604 139254 102204 174698
rect 101604 139018 101786 139254
rect 102022 139018 102204 139254
rect 101604 138934 102204 139018
rect 101604 138698 101786 138934
rect 102022 138698 102204 138934
rect 101604 103254 102204 138698
rect 101604 103018 101786 103254
rect 102022 103018 102204 103254
rect 101604 102934 102204 103018
rect 101604 102698 101786 102934
rect 102022 102698 102204 102934
rect 101604 67254 102204 102698
rect 101604 67018 101786 67254
rect 102022 67018 102204 67254
rect 101604 66934 102204 67018
rect 101604 66698 101786 66934
rect 102022 66698 102204 66934
rect 101604 31254 102204 66698
rect 101604 31018 101786 31254
rect 102022 31018 102204 31254
rect 101604 30934 102204 31018
rect 101604 30698 101786 30934
rect 102022 30698 102204 30934
rect 83604 -6102 83786 -5866
rect 84022 -6102 84204 -5866
rect 83604 -6186 84204 -6102
rect 83604 -6422 83786 -6186
rect 84022 -6422 84204 -6186
rect 83604 -7364 84204 -6422
rect 101604 -6786 102204 30698
rect 108804 704838 109404 705780
rect 108804 704602 108986 704838
rect 109222 704602 109404 704838
rect 108804 704518 109404 704602
rect 108804 704282 108986 704518
rect 109222 704282 109404 704518
rect 108804 686454 109404 704282
rect 108804 686218 108986 686454
rect 109222 686218 109404 686454
rect 108804 686134 109404 686218
rect 108804 685898 108986 686134
rect 109222 685898 109404 686134
rect 108804 650454 109404 685898
rect 108804 650218 108986 650454
rect 109222 650218 109404 650454
rect 108804 650134 109404 650218
rect 108804 649898 108986 650134
rect 109222 649898 109404 650134
rect 108804 614454 109404 649898
rect 108804 614218 108986 614454
rect 109222 614218 109404 614454
rect 108804 614134 109404 614218
rect 108804 613898 108986 614134
rect 109222 613898 109404 614134
rect 108804 578454 109404 613898
rect 108804 578218 108986 578454
rect 109222 578218 109404 578454
rect 108804 578134 109404 578218
rect 108804 577898 108986 578134
rect 109222 577898 109404 578134
rect 108804 542454 109404 577898
rect 108804 542218 108986 542454
rect 109222 542218 109404 542454
rect 108804 542134 109404 542218
rect 108804 541898 108986 542134
rect 109222 541898 109404 542134
rect 108804 506454 109404 541898
rect 108804 506218 108986 506454
rect 109222 506218 109404 506454
rect 108804 506134 109404 506218
rect 108804 505898 108986 506134
rect 109222 505898 109404 506134
rect 108804 470454 109404 505898
rect 108804 470218 108986 470454
rect 109222 470218 109404 470454
rect 108804 470134 109404 470218
rect 108804 469898 108986 470134
rect 109222 469898 109404 470134
rect 108804 434454 109404 469898
rect 108804 434218 108986 434454
rect 109222 434218 109404 434454
rect 108804 434134 109404 434218
rect 108804 433898 108986 434134
rect 109222 433898 109404 434134
rect 108804 398454 109404 433898
rect 108804 398218 108986 398454
rect 109222 398218 109404 398454
rect 108804 398134 109404 398218
rect 108804 397898 108986 398134
rect 109222 397898 109404 398134
rect 108804 362454 109404 397898
rect 108804 362218 108986 362454
rect 109222 362218 109404 362454
rect 108804 362134 109404 362218
rect 108804 361898 108986 362134
rect 109222 361898 109404 362134
rect 108804 326454 109404 361898
rect 108804 326218 108986 326454
rect 109222 326218 109404 326454
rect 108804 326134 109404 326218
rect 108804 325898 108986 326134
rect 109222 325898 109404 326134
rect 108804 290454 109404 325898
rect 108804 290218 108986 290454
rect 109222 290218 109404 290454
rect 108804 290134 109404 290218
rect 108804 289898 108986 290134
rect 109222 289898 109404 290134
rect 108804 254454 109404 289898
rect 108804 254218 108986 254454
rect 109222 254218 109404 254454
rect 108804 254134 109404 254218
rect 108804 253898 108986 254134
rect 109222 253898 109404 254134
rect 108804 218454 109404 253898
rect 108804 218218 108986 218454
rect 109222 218218 109404 218454
rect 108804 218134 109404 218218
rect 108804 217898 108986 218134
rect 109222 217898 109404 218134
rect 108804 182454 109404 217898
rect 108804 182218 108986 182454
rect 109222 182218 109404 182454
rect 108804 182134 109404 182218
rect 108804 181898 108986 182134
rect 109222 181898 109404 182134
rect 108804 146454 109404 181898
rect 108804 146218 108986 146454
rect 109222 146218 109404 146454
rect 108804 146134 109404 146218
rect 108804 145898 108986 146134
rect 109222 145898 109404 146134
rect 108804 110454 109404 145898
rect 108804 110218 108986 110454
rect 109222 110218 109404 110454
rect 108804 110134 109404 110218
rect 108804 109898 108986 110134
rect 109222 109898 109404 110134
rect 108804 74454 109404 109898
rect 108804 74218 108986 74454
rect 109222 74218 109404 74454
rect 108804 74134 109404 74218
rect 108804 73898 108986 74134
rect 109222 73898 109404 74134
rect 108804 38454 109404 73898
rect 108804 38218 108986 38454
rect 109222 38218 109404 38454
rect 108804 38134 109404 38218
rect 108804 37898 108986 38134
rect 109222 37898 109404 38134
rect 108804 2454 109404 37898
rect 108804 2218 108986 2454
rect 109222 2218 109404 2454
rect 108804 2134 109404 2218
rect 108804 1898 108986 2134
rect 109222 1898 109404 2134
rect 108804 -346 109404 1898
rect 108804 -582 108986 -346
rect 109222 -582 109404 -346
rect 108804 -666 109404 -582
rect 108804 -902 108986 -666
rect 109222 -902 109404 -666
rect 108804 -1844 109404 -902
rect 112404 690054 113004 706122
rect 112404 689818 112586 690054
rect 112822 689818 113004 690054
rect 112404 689734 113004 689818
rect 112404 689498 112586 689734
rect 112822 689498 113004 689734
rect 112404 654054 113004 689498
rect 112404 653818 112586 654054
rect 112822 653818 113004 654054
rect 112404 653734 113004 653818
rect 112404 653498 112586 653734
rect 112822 653498 113004 653734
rect 112404 618054 113004 653498
rect 112404 617818 112586 618054
rect 112822 617818 113004 618054
rect 112404 617734 113004 617818
rect 112404 617498 112586 617734
rect 112822 617498 113004 617734
rect 112404 582054 113004 617498
rect 112404 581818 112586 582054
rect 112822 581818 113004 582054
rect 112404 581734 113004 581818
rect 112404 581498 112586 581734
rect 112822 581498 113004 581734
rect 112404 546054 113004 581498
rect 112404 545818 112586 546054
rect 112822 545818 113004 546054
rect 112404 545734 113004 545818
rect 112404 545498 112586 545734
rect 112822 545498 113004 545734
rect 112404 510054 113004 545498
rect 112404 509818 112586 510054
rect 112822 509818 113004 510054
rect 112404 509734 113004 509818
rect 112404 509498 112586 509734
rect 112822 509498 113004 509734
rect 112404 474054 113004 509498
rect 112404 473818 112586 474054
rect 112822 473818 113004 474054
rect 112404 473734 113004 473818
rect 112404 473498 112586 473734
rect 112822 473498 113004 473734
rect 112404 438054 113004 473498
rect 112404 437818 112586 438054
rect 112822 437818 113004 438054
rect 112404 437734 113004 437818
rect 112404 437498 112586 437734
rect 112822 437498 113004 437734
rect 112404 402054 113004 437498
rect 112404 401818 112586 402054
rect 112822 401818 113004 402054
rect 112404 401734 113004 401818
rect 112404 401498 112586 401734
rect 112822 401498 113004 401734
rect 112404 366054 113004 401498
rect 112404 365818 112586 366054
rect 112822 365818 113004 366054
rect 112404 365734 113004 365818
rect 112404 365498 112586 365734
rect 112822 365498 113004 365734
rect 112404 330054 113004 365498
rect 112404 329818 112586 330054
rect 112822 329818 113004 330054
rect 112404 329734 113004 329818
rect 112404 329498 112586 329734
rect 112822 329498 113004 329734
rect 112404 294054 113004 329498
rect 112404 293818 112586 294054
rect 112822 293818 113004 294054
rect 112404 293734 113004 293818
rect 112404 293498 112586 293734
rect 112822 293498 113004 293734
rect 112404 258054 113004 293498
rect 112404 257818 112586 258054
rect 112822 257818 113004 258054
rect 112404 257734 113004 257818
rect 112404 257498 112586 257734
rect 112822 257498 113004 257734
rect 112404 222054 113004 257498
rect 112404 221818 112586 222054
rect 112822 221818 113004 222054
rect 112404 221734 113004 221818
rect 112404 221498 112586 221734
rect 112822 221498 113004 221734
rect 112404 186054 113004 221498
rect 112404 185818 112586 186054
rect 112822 185818 113004 186054
rect 112404 185734 113004 185818
rect 112404 185498 112586 185734
rect 112822 185498 113004 185734
rect 112404 150054 113004 185498
rect 112404 149818 112586 150054
rect 112822 149818 113004 150054
rect 112404 149734 113004 149818
rect 112404 149498 112586 149734
rect 112822 149498 113004 149734
rect 112404 114054 113004 149498
rect 112404 113818 112586 114054
rect 112822 113818 113004 114054
rect 112404 113734 113004 113818
rect 112404 113498 112586 113734
rect 112822 113498 113004 113734
rect 112404 78054 113004 113498
rect 112404 77818 112586 78054
rect 112822 77818 113004 78054
rect 112404 77734 113004 77818
rect 112404 77498 112586 77734
rect 112822 77498 113004 77734
rect 112404 42054 113004 77498
rect 112404 41818 112586 42054
rect 112822 41818 113004 42054
rect 112404 41734 113004 41818
rect 112404 41498 112586 41734
rect 112822 41498 113004 41734
rect 112404 6054 113004 41498
rect 112404 5818 112586 6054
rect 112822 5818 113004 6054
rect 112404 5734 113004 5818
rect 112404 5498 112586 5734
rect 112822 5498 113004 5734
rect 112404 -2186 113004 5498
rect 112404 -2422 112586 -2186
rect 112822 -2422 113004 -2186
rect 112404 -2506 113004 -2422
rect 112404 -2742 112586 -2506
rect 112822 -2742 113004 -2506
rect 112404 -3684 113004 -2742
rect 116004 693654 116604 707962
rect 116004 693418 116186 693654
rect 116422 693418 116604 693654
rect 116004 693334 116604 693418
rect 116004 693098 116186 693334
rect 116422 693098 116604 693334
rect 116004 657654 116604 693098
rect 116004 657418 116186 657654
rect 116422 657418 116604 657654
rect 116004 657334 116604 657418
rect 116004 657098 116186 657334
rect 116422 657098 116604 657334
rect 116004 621654 116604 657098
rect 116004 621418 116186 621654
rect 116422 621418 116604 621654
rect 116004 621334 116604 621418
rect 116004 621098 116186 621334
rect 116422 621098 116604 621334
rect 116004 585654 116604 621098
rect 116004 585418 116186 585654
rect 116422 585418 116604 585654
rect 116004 585334 116604 585418
rect 116004 585098 116186 585334
rect 116422 585098 116604 585334
rect 116004 549654 116604 585098
rect 116004 549418 116186 549654
rect 116422 549418 116604 549654
rect 116004 549334 116604 549418
rect 116004 549098 116186 549334
rect 116422 549098 116604 549334
rect 116004 513654 116604 549098
rect 116004 513418 116186 513654
rect 116422 513418 116604 513654
rect 116004 513334 116604 513418
rect 116004 513098 116186 513334
rect 116422 513098 116604 513334
rect 116004 477654 116604 513098
rect 116004 477418 116186 477654
rect 116422 477418 116604 477654
rect 116004 477334 116604 477418
rect 116004 477098 116186 477334
rect 116422 477098 116604 477334
rect 116004 441654 116604 477098
rect 116004 441418 116186 441654
rect 116422 441418 116604 441654
rect 116004 441334 116604 441418
rect 116004 441098 116186 441334
rect 116422 441098 116604 441334
rect 116004 405654 116604 441098
rect 116004 405418 116186 405654
rect 116422 405418 116604 405654
rect 116004 405334 116604 405418
rect 116004 405098 116186 405334
rect 116422 405098 116604 405334
rect 116004 369654 116604 405098
rect 116004 369418 116186 369654
rect 116422 369418 116604 369654
rect 116004 369334 116604 369418
rect 116004 369098 116186 369334
rect 116422 369098 116604 369334
rect 116004 333654 116604 369098
rect 116004 333418 116186 333654
rect 116422 333418 116604 333654
rect 116004 333334 116604 333418
rect 116004 333098 116186 333334
rect 116422 333098 116604 333334
rect 116004 297654 116604 333098
rect 116004 297418 116186 297654
rect 116422 297418 116604 297654
rect 116004 297334 116604 297418
rect 116004 297098 116186 297334
rect 116422 297098 116604 297334
rect 116004 261654 116604 297098
rect 116004 261418 116186 261654
rect 116422 261418 116604 261654
rect 116004 261334 116604 261418
rect 116004 261098 116186 261334
rect 116422 261098 116604 261334
rect 116004 225654 116604 261098
rect 116004 225418 116186 225654
rect 116422 225418 116604 225654
rect 116004 225334 116604 225418
rect 116004 225098 116186 225334
rect 116422 225098 116604 225334
rect 116004 189654 116604 225098
rect 116004 189418 116186 189654
rect 116422 189418 116604 189654
rect 116004 189334 116604 189418
rect 116004 189098 116186 189334
rect 116422 189098 116604 189334
rect 116004 153654 116604 189098
rect 116004 153418 116186 153654
rect 116422 153418 116604 153654
rect 116004 153334 116604 153418
rect 116004 153098 116186 153334
rect 116422 153098 116604 153334
rect 116004 117654 116604 153098
rect 116004 117418 116186 117654
rect 116422 117418 116604 117654
rect 116004 117334 116604 117418
rect 116004 117098 116186 117334
rect 116422 117098 116604 117334
rect 116004 81654 116604 117098
rect 116004 81418 116186 81654
rect 116422 81418 116604 81654
rect 116004 81334 116604 81418
rect 116004 81098 116186 81334
rect 116422 81098 116604 81334
rect 116004 45654 116604 81098
rect 116004 45418 116186 45654
rect 116422 45418 116604 45654
rect 116004 45334 116604 45418
rect 116004 45098 116186 45334
rect 116422 45098 116604 45334
rect 116004 9654 116604 45098
rect 116004 9418 116186 9654
rect 116422 9418 116604 9654
rect 116004 9334 116604 9418
rect 116004 9098 116186 9334
rect 116422 9098 116604 9334
rect 116004 -4026 116604 9098
rect 116004 -4262 116186 -4026
rect 116422 -4262 116604 -4026
rect 116004 -4346 116604 -4262
rect 116004 -4582 116186 -4346
rect 116422 -4582 116604 -4346
rect 116004 -5524 116604 -4582
rect 119604 697254 120204 709802
rect 137604 711278 138204 711300
rect 137604 711042 137786 711278
rect 138022 711042 138204 711278
rect 137604 710958 138204 711042
rect 137604 710722 137786 710958
rect 138022 710722 138204 710958
rect 134004 709438 134604 709460
rect 134004 709202 134186 709438
rect 134422 709202 134604 709438
rect 134004 709118 134604 709202
rect 134004 708882 134186 709118
rect 134422 708882 134604 709118
rect 130404 707598 131004 707620
rect 130404 707362 130586 707598
rect 130822 707362 131004 707598
rect 130404 707278 131004 707362
rect 130404 707042 130586 707278
rect 130822 707042 131004 707278
rect 119604 697018 119786 697254
rect 120022 697018 120204 697254
rect 119604 696934 120204 697018
rect 119604 696698 119786 696934
rect 120022 696698 120204 696934
rect 119604 661254 120204 696698
rect 119604 661018 119786 661254
rect 120022 661018 120204 661254
rect 119604 660934 120204 661018
rect 119604 660698 119786 660934
rect 120022 660698 120204 660934
rect 119604 625254 120204 660698
rect 119604 625018 119786 625254
rect 120022 625018 120204 625254
rect 119604 624934 120204 625018
rect 119604 624698 119786 624934
rect 120022 624698 120204 624934
rect 119604 589254 120204 624698
rect 119604 589018 119786 589254
rect 120022 589018 120204 589254
rect 119604 588934 120204 589018
rect 119604 588698 119786 588934
rect 120022 588698 120204 588934
rect 119604 553254 120204 588698
rect 119604 553018 119786 553254
rect 120022 553018 120204 553254
rect 119604 552934 120204 553018
rect 119604 552698 119786 552934
rect 120022 552698 120204 552934
rect 119604 517254 120204 552698
rect 119604 517018 119786 517254
rect 120022 517018 120204 517254
rect 119604 516934 120204 517018
rect 119604 516698 119786 516934
rect 120022 516698 120204 516934
rect 119604 481254 120204 516698
rect 119604 481018 119786 481254
rect 120022 481018 120204 481254
rect 119604 480934 120204 481018
rect 119604 480698 119786 480934
rect 120022 480698 120204 480934
rect 119604 445254 120204 480698
rect 119604 445018 119786 445254
rect 120022 445018 120204 445254
rect 119604 444934 120204 445018
rect 119604 444698 119786 444934
rect 120022 444698 120204 444934
rect 119604 409254 120204 444698
rect 119604 409018 119786 409254
rect 120022 409018 120204 409254
rect 119604 408934 120204 409018
rect 119604 408698 119786 408934
rect 120022 408698 120204 408934
rect 119604 373254 120204 408698
rect 119604 373018 119786 373254
rect 120022 373018 120204 373254
rect 119604 372934 120204 373018
rect 119604 372698 119786 372934
rect 120022 372698 120204 372934
rect 119604 337254 120204 372698
rect 119604 337018 119786 337254
rect 120022 337018 120204 337254
rect 119604 336934 120204 337018
rect 119604 336698 119786 336934
rect 120022 336698 120204 336934
rect 119604 301254 120204 336698
rect 119604 301018 119786 301254
rect 120022 301018 120204 301254
rect 119604 300934 120204 301018
rect 119604 300698 119786 300934
rect 120022 300698 120204 300934
rect 119604 265254 120204 300698
rect 119604 265018 119786 265254
rect 120022 265018 120204 265254
rect 119604 264934 120204 265018
rect 119604 264698 119786 264934
rect 120022 264698 120204 264934
rect 119604 229254 120204 264698
rect 119604 229018 119786 229254
rect 120022 229018 120204 229254
rect 119604 228934 120204 229018
rect 119604 228698 119786 228934
rect 120022 228698 120204 228934
rect 119604 193254 120204 228698
rect 119604 193018 119786 193254
rect 120022 193018 120204 193254
rect 119604 192934 120204 193018
rect 119604 192698 119786 192934
rect 120022 192698 120204 192934
rect 119604 157254 120204 192698
rect 119604 157018 119786 157254
rect 120022 157018 120204 157254
rect 119604 156934 120204 157018
rect 119604 156698 119786 156934
rect 120022 156698 120204 156934
rect 119604 121254 120204 156698
rect 119604 121018 119786 121254
rect 120022 121018 120204 121254
rect 119604 120934 120204 121018
rect 119604 120698 119786 120934
rect 120022 120698 120204 120934
rect 119604 85254 120204 120698
rect 119604 85018 119786 85254
rect 120022 85018 120204 85254
rect 119604 84934 120204 85018
rect 119604 84698 119786 84934
rect 120022 84698 120204 84934
rect 119604 49254 120204 84698
rect 119604 49018 119786 49254
rect 120022 49018 120204 49254
rect 119604 48934 120204 49018
rect 119604 48698 119786 48934
rect 120022 48698 120204 48934
rect 119604 13254 120204 48698
rect 119604 13018 119786 13254
rect 120022 13018 120204 13254
rect 119604 12934 120204 13018
rect 119604 12698 119786 12934
rect 120022 12698 120204 12934
rect 101604 -7022 101786 -6786
rect 102022 -7022 102204 -6786
rect 101604 -7106 102204 -7022
rect 101604 -7342 101786 -7106
rect 102022 -7342 102204 -7106
rect 101604 -7364 102204 -7342
rect 119604 -5866 120204 12698
rect 126804 705758 127404 705780
rect 126804 705522 126986 705758
rect 127222 705522 127404 705758
rect 126804 705438 127404 705522
rect 126804 705202 126986 705438
rect 127222 705202 127404 705438
rect 126804 668454 127404 705202
rect 126804 668218 126986 668454
rect 127222 668218 127404 668454
rect 126804 668134 127404 668218
rect 126804 667898 126986 668134
rect 127222 667898 127404 668134
rect 126804 632454 127404 667898
rect 126804 632218 126986 632454
rect 127222 632218 127404 632454
rect 126804 632134 127404 632218
rect 126804 631898 126986 632134
rect 127222 631898 127404 632134
rect 126804 596454 127404 631898
rect 126804 596218 126986 596454
rect 127222 596218 127404 596454
rect 126804 596134 127404 596218
rect 126804 595898 126986 596134
rect 127222 595898 127404 596134
rect 126804 560454 127404 595898
rect 126804 560218 126986 560454
rect 127222 560218 127404 560454
rect 126804 560134 127404 560218
rect 126804 559898 126986 560134
rect 127222 559898 127404 560134
rect 126804 524454 127404 559898
rect 126804 524218 126986 524454
rect 127222 524218 127404 524454
rect 126804 524134 127404 524218
rect 126804 523898 126986 524134
rect 127222 523898 127404 524134
rect 126804 488454 127404 523898
rect 126804 488218 126986 488454
rect 127222 488218 127404 488454
rect 126804 488134 127404 488218
rect 126804 487898 126986 488134
rect 127222 487898 127404 488134
rect 126804 452454 127404 487898
rect 126804 452218 126986 452454
rect 127222 452218 127404 452454
rect 126804 452134 127404 452218
rect 126804 451898 126986 452134
rect 127222 451898 127404 452134
rect 126804 416454 127404 451898
rect 126804 416218 126986 416454
rect 127222 416218 127404 416454
rect 126804 416134 127404 416218
rect 126804 415898 126986 416134
rect 127222 415898 127404 416134
rect 126804 380454 127404 415898
rect 126804 380218 126986 380454
rect 127222 380218 127404 380454
rect 126804 380134 127404 380218
rect 126804 379898 126986 380134
rect 127222 379898 127404 380134
rect 126804 344454 127404 379898
rect 126804 344218 126986 344454
rect 127222 344218 127404 344454
rect 126804 344134 127404 344218
rect 126804 343898 126986 344134
rect 127222 343898 127404 344134
rect 126804 308454 127404 343898
rect 126804 308218 126986 308454
rect 127222 308218 127404 308454
rect 126804 308134 127404 308218
rect 126804 307898 126986 308134
rect 127222 307898 127404 308134
rect 126804 272454 127404 307898
rect 126804 272218 126986 272454
rect 127222 272218 127404 272454
rect 126804 272134 127404 272218
rect 126804 271898 126986 272134
rect 127222 271898 127404 272134
rect 126804 236454 127404 271898
rect 126804 236218 126986 236454
rect 127222 236218 127404 236454
rect 126804 236134 127404 236218
rect 126804 235898 126986 236134
rect 127222 235898 127404 236134
rect 126804 200454 127404 235898
rect 126804 200218 126986 200454
rect 127222 200218 127404 200454
rect 126804 200134 127404 200218
rect 126804 199898 126986 200134
rect 127222 199898 127404 200134
rect 126804 164454 127404 199898
rect 126804 164218 126986 164454
rect 127222 164218 127404 164454
rect 126804 164134 127404 164218
rect 126804 163898 126986 164134
rect 127222 163898 127404 164134
rect 126804 128454 127404 163898
rect 126804 128218 126986 128454
rect 127222 128218 127404 128454
rect 126804 128134 127404 128218
rect 126804 127898 126986 128134
rect 127222 127898 127404 128134
rect 126804 92454 127404 127898
rect 126804 92218 126986 92454
rect 127222 92218 127404 92454
rect 126804 92134 127404 92218
rect 126804 91898 126986 92134
rect 127222 91898 127404 92134
rect 126804 56454 127404 91898
rect 126804 56218 126986 56454
rect 127222 56218 127404 56454
rect 126804 56134 127404 56218
rect 126804 55898 126986 56134
rect 127222 55898 127404 56134
rect 126804 20454 127404 55898
rect 126804 20218 126986 20454
rect 127222 20218 127404 20454
rect 126804 20134 127404 20218
rect 126804 19898 126986 20134
rect 127222 19898 127404 20134
rect 126804 -1266 127404 19898
rect 126804 -1502 126986 -1266
rect 127222 -1502 127404 -1266
rect 126804 -1586 127404 -1502
rect 126804 -1822 126986 -1586
rect 127222 -1822 127404 -1586
rect 126804 -1844 127404 -1822
rect 130404 672054 131004 707042
rect 130404 671818 130586 672054
rect 130822 671818 131004 672054
rect 130404 671734 131004 671818
rect 130404 671498 130586 671734
rect 130822 671498 131004 671734
rect 130404 636054 131004 671498
rect 130404 635818 130586 636054
rect 130822 635818 131004 636054
rect 130404 635734 131004 635818
rect 130404 635498 130586 635734
rect 130822 635498 131004 635734
rect 130404 600054 131004 635498
rect 130404 599818 130586 600054
rect 130822 599818 131004 600054
rect 130404 599734 131004 599818
rect 130404 599498 130586 599734
rect 130822 599498 131004 599734
rect 130404 564054 131004 599498
rect 130404 563818 130586 564054
rect 130822 563818 131004 564054
rect 130404 563734 131004 563818
rect 130404 563498 130586 563734
rect 130822 563498 131004 563734
rect 130404 528054 131004 563498
rect 130404 527818 130586 528054
rect 130822 527818 131004 528054
rect 130404 527734 131004 527818
rect 130404 527498 130586 527734
rect 130822 527498 131004 527734
rect 130404 492054 131004 527498
rect 130404 491818 130586 492054
rect 130822 491818 131004 492054
rect 130404 491734 131004 491818
rect 130404 491498 130586 491734
rect 130822 491498 131004 491734
rect 130404 456054 131004 491498
rect 130404 455818 130586 456054
rect 130822 455818 131004 456054
rect 130404 455734 131004 455818
rect 130404 455498 130586 455734
rect 130822 455498 131004 455734
rect 130404 420054 131004 455498
rect 130404 419818 130586 420054
rect 130822 419818 131004 420054
rect 130404 419734 131004 419818
rect 130404 419498 130586 419734
rect 130822 419498 131004 419734
rect 130404 384054 131004 419498
rect 130404 383818 130586 384054
rect 130822 383818 131004 384054
rect 130404 383734 131004 383818
rect 130404 383498 130586 383734
rect 130822 383498 131004 383734
rect 130404 348054 131004 383498
rect 130404 347818 130586 348054
rect 130822 347818 131004 348054
rect 130404 347734 131004 347818
rect 130404 347498 130586 347734
rect 130822 347498 131004 347734
rect 130404 312054 131004 347498
rect 130404 311818 130586 312054
rect 130822 311818 131004 312054
rect 130404 311734 131004 311818
rect 130404 311498 130586 311734
rect 130822 311498 131004 311734
rect 130404 276054 131004 311498
rect 130404 275818 130586 276054
rect 130822 275818 131004 276054
rect 130404 275734 131004 275818
rect 130404 275498 130586 275734
rect 130822 275498 131004 275734
rect 130404 240054 131004 275498
rect 130404 239818 130586 240054
rect 130822 239818 131004 240054
rect 130404 239734 131004 239818
rect 130404 239498 130586 239734
rect 130822 239498 131004 239734
rect 130404 204054 131004 239498
rect 130404 203818 130586 204054
rect 130822 203818 131004 204054
rect 130404 203734 131004 203818
rect 130404 203498 130586 203734
rect 130822 203498 131004 203734
rect 130404 168054 131004 203498
rect 130404 167818 130586 168054
rect 130822 167818 131004 168054
rect 130404 167734 131004 167818
rect 130404 167498 130586 167734
rect 130822 167498 131004 167734
rect 130404 132054 131004 167498
rect 130404 131818 130586 132054
rect 130822 131818 131004 132054
rect 130404 131734 131004 131818
rect 130404 131498 130586 131734
rect 130822 131498 131004 131734
rect 130404 96054 131004 131498
rect 130404 95818 130586 96054
rect 130822 95818 131004 96054
rect 130404 95734 131004 95818
rect 130404 95498 130586 95734
rect 130822 95498 131004 95734
rect 130404 60054 131004 95498
rect 130404 59818 130586 60054
rect 130822 59818 131004 60054
rect 130404 59734 131004 59818
rect 130404 59498 130586 59734
rect 130822 59498 131004 59734
rect 130404 24054 131004 59498
rect 130404 23818 130586 24054
rect 130822 23818 131004 24054
rect 130404 23734 131004 23818
rect 130404 23498 130586 23734
rect 130822 23498 131004 23734
rect 130404 -3106 131004 23498
rect 130404 -3342 130586 -3106
rect 130822 -3342 131004 -3106
rect 130404 -3426 131004 -3342
rect 130404 -3662 130586 -3426
rect 130822 -3662 131004 -3426
rect 130404 -3684 131004 -3662
rect 134004 675654 134604 708882
rect 134004 675418 134186 675654
rect 134422 675418 134604 675654
rect 134004 675334 134604 675418
rect 134004 675098 134186 675334
rect 134422 675098 134604 675334
rect 134004 639654 134604 675098
rect 134004 639418 134186 639654
rect 134422 639418 134604 639654
rect 134004 639334 134604 639418
rect 134004 639098 134186 639334
rect 134422 639098 134604 639334
rect 134004 603654 134604 639098
rect 134004 603418 134186 603654
rect 134422 603418 134604 603654
rect 134004 603334 134604 603418
rect 134004 603098 134186 603334
rect 134422 603098 134604 603334
rect 134004 567654 134604 603098
rect 134004 567418 134186 567654
rect 134422 567418 134604 567654
rect 134004 567334 134604 567418
rect 134004 567098 134186 567334
rect 134422 567098 134604 567334
rect 134004 531654 134604 567098
rect 134004 531418 134186 531654
rect 134422 531418 134604 531654
rect 134004 531334 134604 531418
rect 134004 531098 134186 531334
rect 134422 531098 134604 531334
rect 134004 495654 134604 531098
rect 134004 495418 134186 495654
rect 134422 495418 134604 495654
rect 134004 495334 134604 495418
rect 134004 495098 134186 495334
rect 134422 495098 134604 495334
rect 134004 459654 134604 495098
rect 134004 459418 134186 459654
rect 134422 459418 134604 459654
rect 134004 459334 134604 459418
rect 134004 459098 134186 459334
rect 134422 459098 134604 459334
rect 134004 423654 134604 459098
rect 134004 423418 134186 423654
rect 134422 423418 134604 423654
rect 134004 423334 134604 423418
rect 134004 423098 134186 423334
rect 134422 423098 134604 423334
rect 134004 387654 134604 423098
rect 134004 387418 134186 387654
rect 134422 387418 134604 387654
rect 134004 387334 134604 387418
rect 134004 387098 134186 387334
rect 134422 387098 134604 387334
rect 134004 351654 134604 387098
rect 134004 351418 134186 351654
rect 134422 351418 134604 351654
rect 134004 351334 134604 351418
rect 134004 351098 134186 351334
rect 134422 351098 134604 351334
rect 134004 315654 134604 351098
rect 134004 315418 134186 315654
rect 134422 315418 134604 315654
rect 134004 315334 134604 315418
rect 134004 315098 134186 315334
rect 134422 315098 134604 315334
rect 134004 279654 134604 315098
rect 134004 279418 134186 279654
rect 134422 279418 134604 279654
rect 134004 279334 134604 279418
rect 134004 279098 134186 279334
rect 134422 279098 134604 279334
rect 134004 243654 134604 279098
rect 134004 243418 134186 243654
rect 134422 243418 134604 243654
rect 134004 243334 134604 243418
rect 134004 243098 134186 243334
rect 134422 243098 134604 243334
rect 134004 207654 134604 243098
rect 134004 207418 134186 207654
rect 134422 207418 134604 207654
rect 134004 207334 134604 207418
rect 134004 207098 134186 207334
rect 134422 207098 134604 207334
rect 134004 171654 134604 207098
rect 134004 171418 134186 171654
rect 134422 171418 134604 171654
rect 134004 171334 134604 171418
rect 134004 171098 134186 171334
rect 134422 171098 134604 171334
rect 134004 135654 134604 171098
rect 134004 135418 134186 135654
rect 134422 135418 134604 135654
rect 134004 135334 134604 135418
rect 134004 135098 134186 135334
rect 134422 135098 134604 135334
rect 134004 99654 134604 135098
rect 134004 99418 134186 99654
rect 134422 99418 134604 99654
rect 134004 99334 134604 99418
rect 134004 99098 134186 99334
rect 134422 99098 134604 99334
rect 134004 63654 134604 99098
rect 134004 63418 134186 63654
rect 134422 63418 134604 63654
rect 134004 63334 134604 63418
rect 134004 63098 134186 63334
rect 134422 63098 134604 63334
rect 134004 27654 134604 63098
rect 134004 27418 134186 27654
rect 134422 27418 134604 27654
rect 134004 27334 134604 27418
rect 134004 27098 134186 27334
rect 134422 27098 134604 27334
rect 134004 -4946 134604 27098
rect 134004 -5182 134186 -4946
rect 134422 -5182 134604 -4946
rect 134004 -5266 134604 -5182
rect 134004 -5502 134186 -5266
rect 134422 -5502 134604 -5266
rect 134004 -5524 134604 -5502
rect 137604 679254 138204 710722
rect 155604 710358 156204 711300
rect 155604 710122 155786 710358
rect 156022 710122 156204 710358
rect 155604 710038 156204 710122
rect 155604 709802 155786 710038
rect 156022 709802 156204 710038
rect 152004 708518 152604 709460
rect 152004 708282 152186 708518
rect 152422 708282 152604 708518
rect 152004 708198 152604 708282
rect 152004 707962 152186 708198
rect 152422 707962 152604 708198
rect 148404 706678 149004 707620
rect 148404 706442 148586 706678
rect 148822 706442 149004 706678
rect 148404 706358 149004 706442
rect 148404 706122 148586 706358
rect 148822 706122 149004 706358
rect 137604 679018 137786 679254
rect 138022 679018 138204 679254
rect 137604 678934 138204 679018
rect 137604 678698 137786 678934
rect 138022 678698 138204 678934
rect 137604 643254 138204 678698
rect 137604 643018 137786 643254
rect 138022 643018 138204 643254
rect 137604 642934 138204 643018
rect 137604 642698 137786 642934
rect 138022 642698 138204 642934
rect 137604 607254 138204 642698
rect 137604 607018 137786 607254
rect 138022 607018 138204 607254
rect 137604 606934 138204 607018
rect 137604 606698 137786 606934
rect 138022 606698 138204 606934
rect 137604 571254 138204 606698
rect 137604 571018 137786 571254
rect 138022 571018 138204 571254
rect 137604 570934 138204 571018
rect 137604 570698 137786 570934
rect 138022 570698 138204 570934
rect 137604 535254 138204 570698
rect 137604 535018 137786 535254
rect 138022 535018 138204 535254
rect 137604 534934 138204 535018
rect 137604 534698 137786 534934
rect 138022 534698 138204 534934
rect 137604 499254 138204 534698
rect 137604 499018 137786 499254
rect 138022 499018 138204 499254
rect 137604 498934 138204 499018
rect 137604 498698 137786 498934
rect 138022 498698 138204 498934
rect 137604 463254 138204 498698
rect 137604 463018 137786 463254
rect 138022 463018 138204 463254
rect 137604 462934 138204 463018
rect 137604 462698 137786 462934
rect 138022 462698 138204 462934
rect 137604 427254 138204 462698
rect 137604 427018 137786 427254
rect 138022 427018 138204 427254
rect 137604 426934 138204 427018
rect 137604 426698 137786 426934
rect 138022 426698 138204 426934
rect 137604 391254 138204 426698
rect 137604 391018 137786 391254
rect 138022 391018 138204 391254
rect 137604 390934 138204 391018
rect 137604 390698 137786 390934
rect 138022 390698 138204 390934
rect 137604 355254 138204 390698
rect 137604 355018 137786 355254
rect 138022 355018 138204 355254
rect 137604 354934 138204 355018
rect 137604 354698 137786 354934
rect 138022 354698 138204 354934
rect 137604 319254 138204 354698
rect 137604 319018 137786 319254
rect 138022 319018 138204 319254
rect 137604 318934 138204 319018
rect 137604 318698 137786 318934
rect 138022 318698 138204 318934
rect 137604 283254 138204 318698
rect 137604 283018 137786 283254
rect 138022 283018 138204 283254
rect 137604 282934 138204 283018
rect 137604 282698 137786 282934
rect 138022 282698 138204 282934
rect 137604 247254 138204 282698
rect 137604 247018 137786 247254
rect 138022 247018 138204 247254
rect 137604 246934 138204 247018
rect 137604 246698 137786 246934
rect 138022 246698 138204 246934
rect 137604 211254 138204 246698
rect 137604 211018 137786 211254
rect 138022 211018 138204 211254
rect 137604 210934 138204 211018
rect 137604 210698 137786 210934
rect 138022 210698 138204 210934
rect 137604 175254 138204 210698
rect 137604 175018 137786 175254
rect 138022 175018 138204 175254
rect 137604 174934 138204 175018
rect 137604 174698 137786 174934
rect 138022 174698 138204 174934
rect 137604 139254 138204 174698
rect 137604 139018 137786 139254
rect 138022 139018 138204 139254
rect 137604 138934 138204 139018
rect 137604 138698 137786 138934
rect 138022 138698 138204 138934
rect 137604 103254 138204 138698
rect 137604 103018 137786 103254
rect 138022 103018 138204 103254
rect 137604 102934 138204 103018
rect 137604 102698 137786 102934
rect 138022 102698 138204 102934
rect 137604 67254 138204 102698
rect 137604 67018 137786 67254
rect 138022 67018 138204 67254
rect 137604 66934 138204 67018
rect 137604 66698 137786 66934
rect 138022 66698 138204 66934
rect 137604 31254 138204 66698
rect 137604 31018 137786 31254
rect 138022 31018 138204 31254
rect 137604 30934 138204 31018
rect 137604 30698 137786 30934
rect 138022 30698 138204 30934
rect 119604 -6102 119786 -5866
rect 120022 -6102 120204 -5866
rect 119604 -6186 120204 -6102
rect 119604 -6422 119786 -6186
rect 120022 -6422 120204 -6186
rect 119604 -7364 120204 -6422
rect 137604 -6786 138204 30698
rect 144804 704838 145404 705780
rect 144804 704602 144986 704838
rect 145222 704602 145404 704838
rect 144804 704518 145404 704602
rect 144804 704282 144986 704518
rect 145222 704282 145404 704518
rect 144804 686454 145404 704282
rect 144804 686218 144986 686454
rect 145222 686218 145404 686454
rect 144804 686134 145404 686218
rect 144804 685898 144986 686134
rect 145222 685898 145404 686134
rect 144804 650454 145404 685898
rect 144804 650218 144986 650454
rect 145222 650218 145404 650454
rect 144804 650134 145404 650218
rect 144804 649898 144986 650134
rect 145222 649898 145404 650134
rect 144804 614454 145404 649898
rect 144804 614218 144986 614454
rect 145222 614218 145404 614454
rect 144804 614134 145404 614218
rect 144804 613898 144986 614134
rect 145222 613898 145404 614134
rect 144804 578454 145404 613898
rect 144804 578218 144986 578454
rect 145222 578218 145404 578454
rect 144804 578134 145404 578218
rect 144804 577898 144986 578134
rect 145222 577898 145404 578134
rect 144804 542454 145404 577898
rect 144804 542218 144986 542454
rect 145222 542218 145404 542454
rect 144804 542134 145404 542218
rect 144804 541898 144986 542134
rect 145222 541898 145404 542134
rect 144804 506454 145404 541898
rect 144804 506218 144986 506454
rect 145222 506218 145404 506454
rect 144804 506134 145404 506218
rect 144804 505898 144986 506134
rect 145222 505898 145404 506134
rect 144804 470454 145404 505898
rect 144804 470218 144986 470454
rect 145222 470218 145404 470454
rect 144804 470134 145404 470218
rect 144804 469898 144986 470134
rect 145222 469898 145404 470134
rect 144804 434454 145404 469898
rect 144804 434218 144986 434454
rect 145222 434218 145404 434454
rect 144804 434134 145404 434218
rect 144804 433898 144986 434134
rect 145222 433898 145404 434134
rect 144804 398454 145404 433898
rect 144804 398218 144986 398454
rect 145222 398218 145404 398454
rect 144804 398134 145404 398218
rect 144804 397898 144986 398134
rect 145222 397898 145404 398134
rect 144804 362454 145404 397898
rect 144804 362218 144986 362454
rect 145222 362218 145404 362454
rect 144804 362134 145404 362218
rect 144804 361898 144986 362134
rect 145222 361898 145404 362134
rect 144804 326454 145404 361898
rect 144804 326218 144986 326454
rect 145222 326218 145404 326454
rect 144804 326134 145404 326218
rect 144804 325898 144986 326134
rect 145222 325898 145404 326134
rect 144804 290454 145404 325898
rect 144804 290218 144986 290454
rect 145222 290218 145404 290454
rect 144804 290134 145404 290218
rect 144804 289898 144986 290134
rect 145222 289898 145404 290134
rect 144804 254454 145404 289898
rect 144804 254218 144986 254454
rect 145222 254218 145404 254454
rect 144804 254134 145404 254218
rect 144804 253898 144986 254134
rect 145222 253898 145404 254134
rect 144804 218454 145404 253898
rect 144804 218218 144986 218454
rect 145222 218218 145404 218454
rect 144804 218134 145404 218218
rect 144804 217898 144986 218134
rect 145222 217898 145404 218134
rect 144804 182454 145404 217898
rect 144804 182218 144986 182454
rect 145222 182218 145404 182454
rect 144804 182134 145404 182218
rect 144804 181898 144986 182134
rect 145222 181898 145404 182134
rect 144804 146454 145404 181898
rect 144804 146218 144986 146454
rect 145222 146218 145404 146454
rect 144804 146134 145404 146218
rect 144804 145898 144986 146134
rect 145222 145898 145404 146134
rect 144804 110454 145404 145898
rect 144804 110218 144986 110454
rect 145222 110218 145404 110454
rect 144804 110134 145404 110218
rect 144804 109898 144986 110134
rect 145222 109898 145404 110134
rect 144804 74454 145404 109898
rect 144804 74218 144986 74454
rect 145222 74218 145404 74454
rect 144804 74134 145404 74218
rect 144804 73898 144986 74134
rect 145222 73898 145404 74134
rect 144804 38454 145404 73898
rect 144804 38218 144986 38454
rect 145222 38218 145404 38454
rect 144804 38134 145404 38218
rect 144804 37898 144986 38134
rect 145222 37898 145404 38134
rect 144804 2454 145404 37898
rect 144804 2218 144986 2454
rect 145222 2218 145404 2454
rect 144804 2134 145404 2218
rect 144804 1898 144986 2134
rect 145222 1898 145404 2134
rect 144804 -346 145404 1898
rect 144804 -582 144986 -346
rect 145222 -582 145404 -346
rect 144804 -666 145404 -582
rect 144804 -902 144986 -666
rect 145222 -902 145404 -666
rect 144804 -1844 145404 -902
rect 148404 690054 149004 706122
rect 148404 689818 148586 690054
rect 148822 689818 149004 690054
rect 148404 689734 149004 689818
rect 148404 689498 148586 689734
rect 148822 689498 149004 689734
rect 148404 654054 149004 689498
rect 148404 653818 148586 654054
rect 148822 653818 149004 654054
rect 148404 653734 149004 653818
rect 148404 653498 148586 653734
rect 148822 653498 149004 653734
rect 148404 618054 149004 653498
rect 148404 617818 148586 618054
rect 148822 617818 149004 618054
rect 148404 617734 149004 617818
rect 148404 617498 148586 617734
rect 148822 617498 149004 617734
rect 148404 582054 149004 617498
rect 148404 581818 148586 582054
rect 148822 581818 149004 582054
rect 148404 581734 149004 581818
rect 148404 581498 148586 581734
rect 148822 581498 149004 581734
rect 148404 546054 149004 581498
rect 148404 545818 148586 546054
rect 148822 545818 149004 546054
rect 148404 545734 149004 545818
rect 148404 545498 148586 545734
rect 148822 545498 149004 545734
rect 148404 510054 149004 545498
rect 148404 509818 148586 510054
rect 148822 509818 149004 510054
rect 148404 509734 149004 509818
rect 148404 509498 148586 509734
rect 148822 509498 149004 509734
rect 148404 474054 149004 509498
rect 148404 473818 148586 474054
rect 148822 473818 149004 474054
rect 148404 473734 149004 473818
rect 148404 473498 148586 473734
rect 148822 473498 149004 473734
rect 148404 438054 149004 473498
rect 148404 437818 148586 438054
rect 148822 437818 149004 438054
rect 148404 437734 149004 437818
rect 148404 437498 148586 437734
rect 148822 437498 149004 437734
rect 148404 402054 149004 437498
rect 148404 401818 148586 402054
rect 148822 401818 149004 402054
rect 148404 401734 149004 401818
rect 148404 401498 148586 401734
rect 148822 401498 149004 401734
rect 148404 366054 149004 401498
rect 148404 365818 148586 366054
rect 148822 365818 149004 366054
rect 148404 365734 149004 365818
rect 148404 365498 148586 365734
rect 148822 365498 149004 365734
rect 148404 330054 149004 365498
rect 148404 329818 148586 330054
rect 148822 329818 149004 330054
rect 148404 329734 149004 329818
rect 148404 329498 148586 329734
rect 148822 329498 149004 329734
rect 148404 294054 149004 329498
rect 148404 293818 148586 294054
rect 148822 293818 149004 294054
rect 148404 293734 149004 293818
rect 148404 293498 148586 293734
rect 148822 293498 149004 293734
rect 148404 258054 149004 293498
rect 148404 257818 148586 258054
rect 148822 257818 149004 258054
rect 148404 257734 149004 257818
rect 148404 257498 148586 257734
rect 148822 257498 149004 257734
rect 148404 222054 149004 257498
rect 148404 221818 148586 222054
rect 148822 221818 149004 222054
rect 148404 221734 149004 221818
rect 148404 221498 148586 221734
rect 148822 221498 149004 221734
rect 148404 186054 149004 221498
rect 148404 185818 148586 186054
rect 148822 185818 149004 186054
rect 148404 185734 149004 185818
rect 148404 185498 148586 185734
rect 148822 185498 149004 185734
rect 148404 150054 149004 185498
rect 148404 149818 148586 150054
rect 148822 149818 149004 150054
rect 148404 149734 149004 149818
rect 148404 149498 148586 149734
rect 148822 149498 149004 149734
rect 148404 114054 149004 149498
rect 148404 113818 148586 114054
rect 148822 113818 149004 114054
rect 148404 113734 149004 113818
rect 148404 113498 148586 113734
rect 148822 113498 149004 113734
rect 148404 78054 149004 113498
rect 148404 77818 148586 78054
rect 148822 77818 149004 78054
rect 148404 77734 149004 77818
rect 148404 77498 148586 77734
rect 148822 77498 149004 77734
rect 148404 42054 149004 77498
rect 148404 41818 148586 42054
rect 148822 41818 149004 42054
rect 148404 41734 149004 41818
rect 148404 41498 148586 41734
rect 148822 41498 149004 41734
rect 148404 6054 149004 41498
rect 148404 5818 148586 6054
rect 148822 5818 149004 6054
rect 148404 5734 149004 5818
rect 148404 5498 148586 5734
rect 148822 5498 149004 5734
rect 148404 -2186 149004 5498
rect 148404 -2422 148586 -2186
rect 148822 -2422 149004 -2186
rect 148404 -2506 149004 -2422
rect 148404 -2742 148586 -2506
rect 148822 -2742 149004 -2506
rect 148404 -3684 149004 -2742
rect 152004 693654 152604 707962
rect 152004 693418 152186 693654
rect 152422 693418 152604 693654
rect 152004 693334 152604 693418
rect 152004 693098 152186 693334
rect 152422 693098 152604 693334
rect 152004 657654 152604 693098
rect 152004 657418 152186 657654
rect 152422 657418 152604 657654
rect 152004 657334 152604 657418
rect 152004 657098 152186 657334
rect 152422 657098 152604 657334
rect 152004 621654 152604 657098
rect 152004 621418 152186 621654
rect 152422 621418 152604 621654
rect 152004 621334 152604 621418
rect 152004 621098 152186 621334
rect 152422 621098 152604 621334
rect 152004 585654 152604 621098
rect 152004 585418 152186 585654
rect 152422 585418 152604 585654
rect 152004 585334 152604 585418
rect 152004 585098 152186 585334
rect 152422 585098 152604 585334
rect 152004 549654 152604 585098
rect 152004 549418 152186 549654
rect 152422 549418 152604 549654
rect 152004 549334 152604 549418
rect 152004 549098 152186 549334
rect 152422 549098 152604 549334
rect 152004 513654 152604 549098
rect 152004 513418 152186 513654
rect 152422 513418 152604 513654
rect 152004 513334 152604 513418
rect 152004 513098 152186 513334
rect 152422 513098 152604 513334
rect 152004 477654 152604 513098
rect 152004 477418 152186 477654
rect 152422 477418 152604 477654
rect 152004 477334 152604 477418
rect 152004 477098 152186 477334
rect 152422 477098 152604 477334
rect 152004 441654 152604 477098
rect 152004 441418 152186 441654
rect 152422 441418 152604 441654
rect 152004 441334 152604 441418
rect 152004 441098 152186 441334
rect 152422 441098 152604 441334
rect 152004 405654 152604 441098
rect 152004 405418 152186 405654
rect 152422 405418 152604 405654
rect 152004 405334 152604 405418
rect 152004 405098 152186 405334
rect 152422 405098 152604 405334
rect 152004 369654 152604 405098
rect 152004 369418 152186 369654
rect 152422 369418 152604 369654
rect 152004 369334 152604 369418
rect 152004 369098 152186 369334
rect 152422 369098 152604 369334
rect 152004 333654 152604 369098
rect 152004 333418 152186 333654
rect 152422 333418 152604 333654
rect 152004 333334 152604 333418
rect 152004 333098 152186 333334
rect 152422 333098 152604 333334
rect 152004 297654 152604 333098
rect 152004 297418 152186 297654
rect 152422 297418 152604 297654
rect 152004 297334 152604 297418
rect 152004 297098 152186 297334
rect 152422 297098 152604 297334
rect 152004 261654 152604 297098
rect 152004 261418 152186 261654
rect 152422 261418 152604 261654
rect 152004 261334 152604 261418
rect 152004 261098 152186 261334
rect 152422 261098 152604 261334
rect 152004 225654 152604 261098
rect 152004 225418 152186 225654
rect 152422 225418 152604 225654
rect 152004 225334 152604 225418
rect 152004 225098 152186 225334
rect 152422 225098 152604 225334
rect 152004 189654 152604 225098
rect 152004 189418 152186 189654
rect 152422 189418 152604 189654
rect 152004 189334 152604 189418
rect 152004 189098 152186 189334
rect 152422 189098 152604 189334
rect 152004 153654 152604 189098
rect 152004 153418 152186 153654
rect 152422 153418 152604 153654
rect 152004 153334 152604 153418
rect 152004 153098 152186 153334
rect 152422 153098 152604 153334
rect 152004 117654 152604 153098
rect 152004 117418 152186 117654
rect 152422 117418 152604 117654
rect 152004 117334 152604 117418
rect 152004 117098 152186 117334
rect 152422 117098 152604 117334
rect 152004 81654 152604 117098
rect 152004 81418 152186 81654
rect 152422 81418 152604 81654
rect 152004 81334 152604 81418
rect 152004 81098 152186 81334
rect 152422 81098 152604 81334
rect 152004 45654 152604 81098
rect 152004 45418 152186 45654
rect 152422 45418 152604 45654
rect 152004 45334 152604 45418
rect 152004 45098 152186 45334
rect 152422 45098 152604 45334
rect 152004 9654 152604 45098
rect 152004 9418 152186 9654
rect 152422 9418 152604 9654
rect 152004 9334 152604 9418
rect 152004 9098 152186 9334
rect 152422 9098 152604 9334
rect 152004 -4026 152604 9098
rect 152004 -4262 152186 -4026
rect 152422 -4262 152604 -4026
rect 152004 -4346 152604 -4262
rect 152004 -4582 152186 -4346
rect 152422 -4582 152604 -4346
rect 152004 -5524 152604 -4582
rect 155604 697254 156204 709802
rect 173604 711278 174204 711300
rect 173604 711042 173786 711278
rect 174022 711042 174204 711278
rect 173604 710958 174204 711042
rect 173604 710722 173786 710958
rect 174022 710722 174204 710958
rect 170004 709438 170604 709460
rect 170004 709202 170186 709438
rect 170422 709202 170604 709438
rect 170004 709118 170604 709202
rect 170004 708882 170186 709118
rect 170422 708882 170604 709118
rect 166404 707598 167004 707620
rect 166404 707362 166586 707598
rect 166822 707362 167004 707598
rect 166404 707278 167004 707362
rect 166404 707042 166586 707278
rect 166822 707042 167004 707278
rect 155604 697018 155786 697254
rect 156022 697018 156204 697254
rect 155604 696934 156204 697018
rect 155604 696698 155786 696934
rect 156022 696698 156204 696934
rect 155604 661254 156204 696698
rect 155604 661018 155786 661254
rect 156022 661018 156204 661254
rect 155604 660934 156204 661018
rect 155604 660698 155786 660934
rect 156022 660698 156204 660934
rect 155604 625254 156204 660698
rect 155604 625018 155786 625254
rect 156022 625018 156204 625254
rect 155604 624934 156204 625018
rect 155604 624698 155786 624934
rect 156022 624698 156204 624934
rect 155604 589254 156204 624698
rect 155604 589018 155786 589254
rect 156022 589018 156204 589254
rect 155604 588934 156204 589018
rect 155604 588698 155786 588934
rect 156022 588698 156204 588934
rect 155604 553254 156204 588698
rect 155604 553018 155786 553254
rect 156022 553018 156204 553254
rect 155604 552934 156204 553018
rect 155604 552698 155786 552934
rect 156022 552698 156204 552934
rect 155604 517254 156204 552698
rect 155604 517018 155786 517254
rect 156022 517018 156204 517254
rect 155604 516934 156204 517018
rect 155604 516698 155786 516934
rect 156022 516698 156204 516934
rect 155604 481254 156204 516698
rect 155604 481018 155786 481254
rect 156022 481018 156204 481254
rect 155604 480934 156204 481018
rect 155604 480698 155786 480934
rect 156022 480698 156204 480934
rect 155604 445254 156204 480698
rect 155604 445018 155786 445254
rect 156022 445018 156204 445254
rect 155604 444934 156204 445018
rect 155604 444698 155786 444934
rect 156022 444698 156204 444934
rect 155604 409254 156204 444698
rect 155604 409018 155786 409254
rect 156022 409018 156204 409254
rect 155604 408934 156204 409018
rect 155604 408698 155786 408934
rect 156022 408698 156204 408934
rect 155604 373254 156204 408698
rect 155604 373018 155786 373254
rect 156022 373018 156204 373254
rect 155604 372934 156204 373018
rect 155604 372698 155786 372934
rect 156022 372698 156204 372934
rect 155604 337254 156204 372698
rect 155604 337018 155786 337254
rect 156022 337018 156204 337254
rect 155604 336934 156204 337018
rect 155604 336698 155786 336934
rect 156022 336698 156204 336934
rect 155604 301254 156204 336698
rect 155604 301018 155786 301254
rect 156022 301018 156204 301254
rect 155604 300934 156204 301018
rect 155604 300698 155786 300934
rect 156022 300698 156204 300934
rect 155604 265254 156204 300698
rect 155604 265018 155786 265254
rect 156022 265018 156204 265254
rect 155604 264934 156204 265018
rect 155604 264698 155786 264934
rect 156022 264698 156204 264934
rect 155604 229254 156204 264698
rect 155604 229018 155786 229254
rect 156022 229018 156204 229254
rect 155604 228934 156204 229018
rect 155604 228698 155786 228934
rect 156022 228698 156204 228934
rect 155604 193254 156204 228698
rect 155604 193018 155786 193254
rect 156022 193018 156204 193254
rect 155604 192934 156204 193018
rect 155604 192698 155786 192934
rect 156022 192698 156204 192934
rect 155604 157254 156204 192698
rect 155604 157018 155786 157254
rect 156022 157018 156204 157254
rect 155604 156934 156204 157018
rect 155604 156698 155786 156934
rect 156022 156698 156204 156934
rect 155604 121254 156204 156698
rect 155604 121018 155786 121254
rect 156022 121018 156204 121254
rect 155604 120934 156204 121018
rect 155604 120698 155786 120934
rect 156022 120698 156204 120934
rect 155604 85254 156204 120698
rect 155604 85018 155786 85254
rect 156022 85018 156204 85254
rect 155604 84934 156204 85018
rect 155604 84698 155786 84934
rect 156022 84698 156204 84934
rect 155604 49254 156204 84698
rect 155604 49018 155786 49254
rect 156022 49018 156204 49254
rect 155604 48934 156204 49018
rect 155604 48698 155786 48934
rect 156022 48698 156204 48934
rect 155604 13254 156204 48698
rect 155604 13018 155786 13254
rect 156022 13018 156204 13254
rect 155604 12934 156204 13018
rect 155604 12698 155786 12934
rect 156022 12698 156204 12934
rect 137604 -7022 137786 -6786
rect 138022 -7022 138204 -6786
rect 137604 -7106 138204 -7022
rect 137604 -7342 137786 -7106
rect 138022 -7342 138204 -7106
rect 137604 -7364 138204 -7342
rect 155604 -5866 156204 12698
rect 162804 705758 163404 705780
rect 162804 705522 162986 705758
rect 163222 705522 163404 705758
rect 162804 705438 163404 705522
rect 162804 705202 162986 705438
rect 163222 705202 163404 705438
rect 162804 668454 163404 705202
rect 162804 668218 162986 668454
rect 163222 668218 163404 668454
rect 162804 668134 163404 668218
rect 162804 667898 162986 668134
rect 163222 667898 163404 668134
rect 162804 632454 163404 667898
rect 162804 632218 162986 632454
rect 163222 632218 163404 632454
rect 162804 632134 163404 632218
rect 162804 631898 162986 632134
rect 163222 631898 163404 632134
rect 162804 596454 163404 631898
rect 162804 596218 162986 596454
rect 163222 596218 163404 596454
rect 162804 596134 163404 596218
rect 162804 595898 162986 596134
rect 163222 595898 163404 596134
rect 162804 560454 163404 595898
rect 162804 560218 162986 560454
rect 163222 560218 163404 560454
rect 162804 560134 163404 560218
rect 162804 559898 162986 560134
rect 163222 559898 163404 560134
rect 162804 524454 163404 559898
rect 162804 524218 162986 524454
rect 163222 524218 163404 524454
rect 162804 524134 163404 524218
rect 162804 523898 162986 524134
rect 163222 523898 163404 524134
rect 162804 488454 163404 523898
rect 162804 488218 162986 488454
rect 163222 488218 163404 488454
rect 162804 488134 163404 488218
rect 162804 487898 162986 488134
rect 163222 487898 163404 488134
rect 162804 452454 163404 487898
rect 162804 452218 162986 452454
rect 163222 452218 163404 452454
rect 162804 452134 163404 452218
rect 162804 451898 162986 452134
rect 163222 451898 163404 452134
rect 162804 416454 163404 451898
rect 162804 416218 162986 416454
rect 163222 416218 163404 416454
rect 162804 416134 163404 416218
rect 162804 415898 162986 416134
rect 163222 415898 163404 416134
rect 162804 380454 163404 415898
rect 162804 380218 162986 380454
rect 163222 380218 163404 380454
rect 162804 380134 163404 380218
rect 162804 379898 162986 380134
rect 163222 379898 163404 380134
rect 162804 344454 163404 379898
rect 162804 344218 162986 344454
rect 163222 344218 163404 344454
rect 162804 344134 163404 344218
rect 162804 343898 162986 344134
rect 163222 343898 163404 344134
rect 162804 308454 163404 343898
rect 162804 308218 162986 308454
rect 163222 308218 163404 308454
rect 162804 308134 163404 308218
rect 162804 307898 162986 308134
rect 163222 307898 163404 308134
rect 162804 272454 163404 307898
rect 162804 272218 162986 272454
rect 163222 272218 163404 272454
rect 162804 272134 163404 272218
rect 162804 271898 162986 272134
rect 163222 271898 163404 272134
rect 162804 236454 163404 271898
rect 162804 236218 162986 236454
rect 163222 236218 163404 236454
rect 162804 236134 163404 236218
rect 162804 235898 162986 236134
rect 163222 235898 163404 236134
rect 162804 200454 163404 235898
rect 162804 200218 162986 200454
rect 163222 200218 163404 200454
rect 162804 200134 163404 200218
rect 162804 199898 162986 200134
rect 163222 199898 163404 200134
rect 162804 164454 163404 199898
rect 162804 164218 162986 164454
rect 163222 164218 163404 164454
rect 162804 164134 163404 164218
rect 162804 163898 162986 164134
rect 163222 163898 163404 164134
rect 162804 128454 163404 163898
rect 162804 128218 162986 128454
rect 163222 128218 163404 128454
rect 162804 128134 163404 128218
rect 162804 127898 162986 128134
rect 163222 127898 163404 128134
rect 162804 92454 163404 127898
rect 162804 92218 162986 92454
rect 163222 92218 163404 92454
rect 162804 92134 163404 92218
rect 162804 91898 162986 92134
rect 163222 91898 163404 92134
rect 162804 56454 163404 91898
rect 162804 56218 162986 56454
rect 163222 56218 163404 56454
rect 162804 56134 163404 56218
rect 162804 55898 162986 56134
rect 163222 55898 163404 56134
rect 162804 20454 163404 55898
rect 162804 20218 162986 20454
rect 163222 20218 163404 20454
rect 162804 20134 163404 20218
rect 162804 19898 162986 20134
rect 163222 19898 163404 20134
rect 162804 -1266 163404 19898
rect 162804 -1502 162986 -1266
rect 163222 -1502 163404 -1266
rect 162804 -1586 163404 -1502
rect 162804 -1822 162986 -1586
rect 163222 -1822 163404 -1586
rect 162804 -1844 163404 -1822
rect 166404 672054 167004 707042
rect 166404 671818 166586 672054
rect 166822 671818 167004 672054
rect 166404 671734 167004 671818
rect 166404 671498 166586 671734
rect 166822 671498 167004 671734
rect 166404 636054 167004 671498
rect 166404 635818 166586 636054
rect 166822 635818 167004 636054
rect 166404 635734 167004 635818
rect 166404 635498 166586 635734
rect 166822 635498 167004 635734
rect 166404 600054 167004 635498
rect 166404 599818 166586 600054
rect 166822 599818 167004 600054
rect 166404 599734 167004 599818
rect 166404 599498 166586 599734
rect 166822 599498 167004 599734
rect 166404 564054 167004 599498
rect 166404 563818 166586 564054
rect 166822 563818 167004 564054
rect 166404 563734 167004 563818
rect 166404 563498 166586 563734
rect 166822 563498 167004 563734
rect 166404 528054 167004 563498
rect 166404 527818 166586 528054
rect 166822 527818 167004 528054
rect 166404 527734 167004 527818
rect 166404 527498 166586 527734
rect 166822 527498 167004 527734
rect 166404 492054 167004 527498
rect 166404 491818 166586 492054
rect 166822 491818 167004 492054
rect 166404 491734 167004 491818
rect 166404 491498 166586 491734
rect 166822 491498 167004 491734
rect 166404 456054 167004 491498
rect 166404 455818 166586 456054
rect 166822 455818 167004 456054
rect 166404 455734 167004 455818
rect 166404 455498 166586 455734
rect 166822 455498 167004 455734
rect 166404 420054 167004 455498
rect 166404 419818 166586 420054
rect 166822 419818 167004 420054
rect 166404 419734 167004 419818
rect 166404 419498 166586 419734
rect 166822 419498 167004 419734
rect 166404 384054 167004 419498
rect 166404 383818 166586 384054
rect 166822 383818 167004 384054
rect 166404 383734 167004 383818
rect 166404 383498 166586 383734
rect 166822 383498 167004 383734
rect 166404 348054 167004 383498
rect 166404 347818 166586 348054
rect 166822 347818 167004 348054
rect 166404 347734 167004 347818
rect 166404 347498 166586 347734
rect 166822 347498 167004 347734
rect 166404 312054 167004 347498
rect 166404 311818 166586 312054
rect 166822 311818 167004 312054
rect 166404 311734 167004 311818
rect 166404 311498 166586 311734
rect 166822 311498 167004 311734
rect 166404 276054 167004 311498
rect 166404 275818 166586 276054
rect 166822 275818 167004 276054
rect 166404 275734 167004 275818
rect 166404 275498 166586 275734
rect 166822 275498 167004 275734
rect 166404 240054 167004 275498
rect 166404 239818 166586 240054
rect 166822 239818 167004 240054
rect 166404 239734 167004 239818
rect 166404 239498 166586 239734
rect 166822 239498 167004 239734
rect 166404 204054 167004 239498
rect 166404 203818 166586 204054
rect 166822 203818 167004 204054
rect 166404 203734 167004 203818
rect 166404 203498 166586 203734
rect 166822 203498 167004 203734
rect 166404 168054 167004 203498
rect 166404 167818 166586 168054
rect 166822 167818 167004 168054
rect 166404 167734 167004 167818
rect 166404 167498 166586 167734
rect 166822 167498 167004 167734
rect 166404 132054 167004 167498
rect 166404 131818 166586 132054
rect 166822 131818 167004 132054
rect 166404 131734 167004 131818
rect 166404 131498 166586 131734
rect 166822 131498 167004 131734
rect 166404 96054 167004 131498
rect 166404 95818 166586 96054
rect 166822 95818 167004 96054
rect 166404 95734 167004 95818
rect 166404 95498 166586 95734
rect 166822 95498 167004 95734
rect 166404 60054 167004 95498
rect 166404 59818 166586 60054
rect 166822 59818 167004 60054
rect 166404 59734 167004 59818
rect 166404 59498 166586 59734
rect 166822 59498 167004 59734
rect 166404 24054 167004 59498
rect 166404 23818 166586 24054
rect 166822 23818 167004 24054
rect 166404 23734 167004 23818
rect 166404 23498 166586 23734
rect 166822 23498 167004 23734
rect 166404 -3106 167004 23498
rect 166404 -3342 166586 -3106
rect 166822 -3342 167004 -3106
rect 166404 -3426 167004 -3342
rect 166404 -3662 166586 -3426
rect 166822 -3662 167004 -3426
rect 166404 -3684 167004 -3662
rect 170004 675654 170604 708882
rect 170004 675418 170186 675654
rect 170422 675418 170604 675654
rect 170004 675334 170604 675418
rect 170004 675098 170186 675334
rect 170422 675098 170604 675334
rect 170004 639654 170604 675098
rect 170004 639418 170186 639654
rect 170422 639418 170604 639654
rect 170004 639334 170604 639418
rect 170004 639098 170186 639334
rect 170422 639098 170604 639334
rect 170004 603654 170604 639098
rect 170004 603418 170186 603654
rect 170422 603418 170604 603654
rect 170004 603334 170604 603418
rect 170004 603098 170186 603334
rect 170422 603098 170604 603334
rect 170004 567654 170604 603098
rect 170004 567418 170186 567654
rect 170422 567418 170604 567654
rect 170004 567334 170604 567418
rect 170004 567098 170186 567334
rect 170422 567098 170604 567334
rect 170004 531654 170604 567098
rect 170004 531418 170186 531654
rect 170422 531418 170604 531654
rect 170004 531334 170604 531418
rect 170004 531098 170186 531334
rect 170422 531098 170604 531334
rect 170004 495654 170604 531098
rect 170004 495418 170186 495654
rect 170422 495418 170604 495654
rect 170004 495334 170604 495418
rect 170004 495098 170186 495334
rect 170422 495098 170604 495334
rect 170004 459654 170604 495098
rect 170004 459418 170186 459654
rect 170422 459418 170604 459654
rect 170004 459334 170604 459418
rect 170004 459098 170186 459334
rect 170422 459098 170604 459334
rect 170004 423654 170604 459098
rect 170004 423418 170186 423654
rect 170422 423418 170604 423654
rect 170004 423334 170604 423418
rect 170004 423098 170186 423334
rect 170422 423098 170604 423334
rect 170004 387654 170604 423098
rect 170004 387418 170186 387654
rect 170422 387418 170604 387654
rect 170004 387334 170604 387418
rect 170004 387098 170186 387334
rect 170422 387098 170604 387334
rect 170004 351654 170604 387098
rect 170004 351418 170186 351654
rect 170422 351418 170604 351654
rect 170004 351334 170604 351418
rect 170004 351098 170186 351334
rect 170422 351098 170604 351334
rect 170004 315654 170604 351098
rect 170004 315418 170186 315654
rect 170422 315418 170604 315654
rect 170004 315334 170604 315418
rect 170004 315098 170186 315334
rect 170422 315098 170604 315334
rect 170004 279654 170604 315098
rect 170004 279418 170186 279654
rect 170422 279418 170604 279654
rect 170004 279334 170604 279418
rect 170004 279098 170186 279334
rect 170422 279098 170604 279334
rect 170004 243654 170604 279098
rect 170004 243418 170186 243654
rect 170422 243418 170604 243654
rect 170004 243334 170604 243418
rect 170004 243098 170186 243334
rect 170422 243098 170604 243334
rect 170004 207654 170604 243098
rect 170004 207418 170186 207654
rect 170422 207418 170604 207654
rect 170004 207334 170604 207418
rect 170004 207098 170186 207334
rect 170422 207098 170604 207334
rect 170004 171654 170604 207098
rect 170004 171418 170186 171654
rect 170422 171418 170604 171654
rect 170004 171334 170604 171418
rect 170004 171098 170186 171334
rect 170422 171098 170604 171334
rect 170004 135654 170604 171098
rect 170004 135418 170186 135654
rect 170422 135418 170604 135654
rect 170004 135334 170604 135418
rect 170004 135098 170186 135334
rect 170422 135098 170604 135334
rect 170004 99654 170604 135098
rect 170004 99418 170186 99654
rect 170422 99418 170604 99654
rect 170004 99334 170604 99418
rect 170004 99098 170186 99334
rect 170422 99098 170604 99334
rect 170004 63654 170604 99098
rect 170004 63418 170186 63654
rect 170422 63418 170604 63654
rect 170004 63334 170604 63418
rect 170004 63098 170186 63334
rect 170422 63098 170604 63334
rect 170004 27654 170604 63098
rect 170004 27418 170186 27654
rect 170422 27418 170604 27654
rect 170004 27334 170604 27418
rect 170004 27098 170186 27334
rect 170422 27098 170604 27334
rect 170004 -4946 170604 27098
rect 170004 -5182 170186 -4946
rect 170422 -5182 170604 -4946
rect 170004 -5266 170604 -5182
rect 170004 -5502 170186 -5266
rect 170422 -5502 170604 -5266
rect 170004 -5524 170604 -5502
rect 173604 679254 174204 710722
rect 191604 710358 192204 711300
rect 191604 710122 191786 710358
rect 192022 710122 192204 710358
rect 191604 710038 192204 710122
rect 191604 709802 191786 710038
rect 192022 709802 192204 710038
rect 188004 708518 188604 709460
rect 188004 708282 188186 708518
rect 188422 708282 188604 708518
rect 188004 708198 188604 708282
rect 188004 707962 188186 708198
rect 188422 707962 188604 708198
rect 184404 706678 185004 707620
rect 184404 706442 184586 706678
rect 184822 706442 185004 706678
rect 184404 706358 185004 706442
rect 184404 706122 184586 706358
rect 184822 706122 185004 706358
rect 173604 679018 173786 679254
rect 174022 679018 174204 679254
rect 173604 678934 174204 679018
rect 173604 678698 173786 678934
rect 174022 678698 174204 678934
rect 173604 643254 174204 678698
rect 173604 643018 173786 643254
rect 174022 643018 174204 643254
rect 173604 642934 174204 643018
rect 173604 642698 173786 642934
rect 174022 642698 174204 642934
rect 173604 607254 174204 642698
rect 173604 607018 173786 607254
rect 174022 607018 174204 607254
rect 173604 606934 174204 607018
rect 173604 606698 173786 606934
rect 174022 606698 174204 606934
rect 173604 571254 174204 606698
rect 173604 571018 173786 571254
rect 174022 571018 174204 571254
rect 173604 570934 174204 571018
rect 173604 570698 173786 570934
rect 174022 570698 174204 570934
rect 173604 535254 174204 570698
rect 173604 535018 173786 535254
rect 174022 535018 174204 535254
rect 173604 534934 174204 535018
rect 173604 534698 173786 534934
rect 174022 534698 174204 534934
rect 173604 499254 174204 534698
rect 173604 499018 173786 499254
rect 174022 499018 174204 499254
rect 173604 498934 174204 499018
rect 173604 498698 173786 498934
rect 174022 498698 174204 498934
rect 173604 463254 174204 498698
rect 173604 463018 173786 463254
rect 174022 463018 174204 463254
rect 173604 462934 174204 463018
rect 173604 462698 173786 462934
rect 174022 462698 174204 462934
rect 173604 427254 174204 462698
rect 173604 427018 173786 427254
rect 174022 427018 174204 427254
rect 173604 426934 174204 427018
rect 173604 426698 173786 426934
rect 174022 426698 174204 426934
rect 173604 391254 174204 426698
rect 173604 391018 173786 391254
rect 174022 391018 174204 391254
rect 173604 390934 174204 391018
rect 173604 390698 173786 390934
rect 174022 390698 174204 390934
rect 173604 355254 174204 390698
rect 173604 355018 173786 355254
rect 174022 355018 174204 355254
rect 173604 354934 174204 355018
rect 173604 354698 173786 354934
rect 174022 354698 174204 354934
rect 173604 319254 174204 354698
rect 173604 319018 173786 319254
rect 174022 319018 174204 319254
rect 173604 318934 174204 319018
rect 173604 318698 173786 318934
rect 174022 318698 174204 318934
rect 173604 283254 174204 318698
rect 173604 283018 173786 283254
rect 174022 283018 174204 283254
rect 173604 282934 174204 283018
rect 173604 282698 173786 282934
rect 174022 282698 174204 282934
rect 173604 247254 174204 282698
rect 173604 247018 173786 247254
rect 174022 247018 174204 247254
rect 173604 246934 174204 247018
rect 173604 246698 173786 246934
rect 174022 246698 174204 246934
rect 173604 211254 174204 246698
rect 173604 211018 173786 211254
rect 174022 211018 174204 211254
rect 173604 210934 174204 211018
rect 173604 210698 173786 210934
rect 174022 210698 174204 210934
rect 173604 175254 174204 210698
rect 173604 175018 173786 175254
rect 174022 175018 174204 175254
rect 173604 174934 174204 175018
rect 173604 174698 173786 174934
rect 174022 174698 174204 174934
rect 173604 139254 174204 174698
rect 173604 139018 173786 139254
rect 174022 139018 174204 139254
rect 173604 138934 174204 139018
rect 173604 138698 173786 138934
rect 174022 138698 174204 138934
rect 173604 103254 174204 138698
rect 173604 103018 173786 103254
rect 174022 103018 174204 103254
rect 173604 102934 174204 103018
rect 173604 102698 173786 102934
rect 174022 102698 174204 102934
rect 173604 67254 174204 102698
rect 173604 67018 173786 67254
rect 174022 67018 174204 67254
rect 173604 66934 174204 67018
rect 173604 66698 173786 66934
rect 174022 66698 174204 66934
rect 173604 31254 174204 66698
rect 173604 31018 173786 31254
rect 174022 31018 174204 31254
rect 173604 30934 174204 31018
rect 173604 30698 173786 30934
rect 174022 30698 174204 30934
rect 155604 -6102 155786 -5866
rect 156022 -6102 156204 -5866
rect 155604 -6186 156204 -6102
rect 155604 -6422 155786 -6186
rect 156022 -6422 156204 -6186
rect 155604 -7364 156204 -6422
rect 173604 -6786 174204 30698
rect 180804 704838 181404 705780
rect 180804 704602 180986 704838
rect 181222 704602 181404 704838
rect 180804 704518 181404 704602
rect 180804 704282 180986 704518
rect 181222 704282 181404 704518
rect 180804 686454 181404 704282
rect 180804 686218 180986 686454
rect 181222 686218 181404 686454
rect 180804 686134 181404 686218
rect 180804 685898 180986 686134
rect 181222 685898 181404 686134
rect 180804 650454 181404 685898
rect 180804 650218 180986 650454
rect 181222 650218 181404 650454
rect 180804 650134 181404 650218
rect 180804 649898 180986 650134
rect 181222 649898 181404 650134
rect 180804 614454 181404 649898
rect 180804 614218 180986 614454
rect 181222 614218 181404 614454
rect 180804 614134 181404 614218
rect 180804 613898 180986 614134
rect 181222 613898 181404 614134
rect 180804 578454 181404 613898
rect 180804 578218 180986 578454
rect 181222 578218 181404 578454
rect 180804 578134 181404 578218
rect 180804 577898 180986 578134
rect 181222 577898 181404 578134
rect 180804 542454 181404 577898
rect 180804 542218 180986 542454
rect 181222 542218 181404 542454
rect 180804 542134 181404 542218
rect 180804 541898 180986 542134
rect 181222 541898 181404 542134
rect 180804 506454 181404 541898
rect 180804 506218 180986 506454
rect 181222 506218 181404 506454
rect 180804 506134 181404 506218
rect 180804 505898 180986 506134
rect 181222 505898 181404 506134
rect 180804 470454 181404 505898
rect 180804 470218 180986 470454
rect 181222 470218 181404 470454
rect 180804 470134 181404 470218
rect 180804 469898 180986 470134
rect 181222 469898 181404 470134
rect 180804 434454 181404 469898
rect 180804 434218 180986 434454
rect 181222 434218 181404 434454
rect 180804 434134 181404 434218
rect 180804 433898 180986 434134
rect 181222 433898 181404 434134
rect 180804 398454 181404 433898
rect 180804 398218 180986 398454
rect 181222 398218 181404 398454
rect 180804 398134 181404 398218
rect 180804 397898 180986 398134
rect 181222 397898 181404 398134
rect 180804 362454 181404 397898
rect 180804 362218 180986 362454
rect 181222 362218 181404 362454
rect 180804 362134 181404 362218
rect 180804 361898 180986 362134
rect 181222 361898 181404 362134
rect 180804 326454 181404 361898
rect 180804 326218 180986 326454
rect 181222 326218 181404 326454
rect 180804 326134 181404 326218
rect 180804 325898 180986 326134
rect 181222 325898 181404 326134
rect 180804 290454 181404 325898
rect 180804 290218 180986 290454
rect 181222 290218 181404 290454
rect 180804 290134 181404 290218
rect 180804 289898 180986 290134
rect 181222 289898 181404 290134
rect 180804 254454 181404 289898
rect 180804 254218 180986 254454
rect 181222 254218 181404 254454
rect 180804 254134 181404 254218
rect 180804 253898 180986 254134
rect 181222 253898 181404 254134
rect 180804 218454 181404 253898
rect 180804 218218 180986 218454
rect 181222 218218 181404 218454
rect 180804 218134 181404 218218
rect 180804 217898 180986 218134
rect 181222 217898 181404 218134
rect 180804 182454 181404 217898
rect 180804 182218 180986 182454
rect 181222 182218 181404 182454
rect 180804 182134 181404 182218
rect 180804 181898 180986 182134
rect 181222 181898 181404 182134
rect 180804 146454 181404 181898
rect 180804 146218 180986 146454
rect 181222 146218 181404 146454
rect 180804 146134 181404 146218
rect 180804 145898 180986 146134
rect 181222 145898 181404 146134
rect 180804 110454 181404 145898
rect 180804 110218 180986 110454
rect 181222 110218 181404 110454
rect 180804 110134 181404 110218
rect 180804 109898 180986 110134
rect 181222 109898 181404 110134
rect 180804 74454 181404 109898
rect 180804 74218 180986 74454
rect 181222 74218 181404 74454
rect 180804 74134 181404 74218
rect 180804 73898 180986 74134
rect 181222 73898 181404 74134
rect 180804 38454 181404 73898
rect 180804 38218 180986 38454
rect 181222 38218 181404 38454
rect 180804 38134 181404 38218
rect 180804 37898 180986 38134
rect 181222 37898 181404 38134
rect 180804 2454 181404 37898
rect 180804 2218 180986 2454
rect 181222 2218 181404 2454
rect 180804 2134 181404 2218
rect 180804 1898 180986 2134
rect 181222 1898 181404 2134
rect 180804 -346 181404 1898
rect 180804 -582 180986 -346
rect 181222 -582 181404 -346
rect 180804 -666 181404 -582
rect 180804 -902 180986 -666
rect 181222 -902 181404 -666
rect 180804 -1844 181404 -902
rect 184404 690054 185004 706122
rect 184404 689818 184586 690054
rect 184822 689818 185004 690054
rect 184404 689734 185004 689818
rect 184404 689498 184586 689734
rect 184822 689498 185004 689734
rect 184404 654054 185004 689498
rect 184404 653818 184586 654054
rect 184822 653818 185004 654054
rect 184404 653734 185004 653818
rect 184404 653498 184586 653734
rect 184822 653498 185004 653734
rect 184404 618054 185004 653498
rect 184404 617818 184586 618054
rect 184822 617818 185004 618054
rect 184404 617734 185004 617818
rect 184404 617498 184586 617734
rect 184822 617498 185004 617734
rect 184404 582054 185004 617498
rect 184404 581818 184586 582054
rect 184822 581818 185004 582054
rect 184404 581734 185004 581818
rect 184404 581498 184586 581734
rect 184822 581498 185004 581734
rect 184404 546054 185004 581498
rect 184404 545818 184586 546054
rect 184822 545818 185004 546054
rect 184404 545734 185004 545818
rect 184404 545498 184586 545734
rect 184822 545498 185004 545734
rect 184404 510054 185004 545498
rect 184404 509818 184586 510054
rect 184822 509818 185004 510054
rect 184404 509734 185004 509818
rect 184404 509498 184586 509734
rect 184822 509498 185004 509734
rect 184404 474054 185004 509498
rect 184404 473818 184586 474054
rect 184822 473818 185004 474054
rect 184404 473734 185004 473818
rect 184404 473498 184586 473734
rect 184822 473498 185004 473734
rect 184404 438054 185004 473498
rect 184404 437818 184586 438054
rect 184822 437818 185004 438054
rect 184404 437734 185004 437818
rect 184404 437498 184586 437734
rect 184822 437498 185004 437734
rect 184404 402054 185004 437498
rect 184404 401818 184586 402054
rect 184822 401818 185004 402054
rect 184404 401734 185004 401818
rect 184404 401498 184586 401734
rect 184822 401498 185004 401734
rect 184404 366054 185004 401498
rect 184404 365818 184586 366054
rect 184822 365818 185004 366054
rect 184404 365734 185004 365818
rect 184404 365498 184586 365734
rect 184822 365498 185004 365734
rect 184404 330054 185004 365498
rect 184404 329818 184586 330054
rect 184822 329818 185004 330054
rect 184404 329734 185004 329818
rect 184404 329498 184586 329734
rect 184822 329498 185004 329734
rect 184404 294054 185004 329498
rect 184404 293818 184586 294054
rect 184822 293818 185004 294054
rect 184404 293734 185004 293818
rect 184404 293498 184586 293734
rect 184822 293498 185004 293734
rect 184404 258054 185004 293498
rect 184404 257818 184586 258054
rect 184822 257818 185004 258054
rect 184404 257734 185004 257818
rect 184404 257498 184586 257734
rect 184822 257498 185004 257734
rect 184404 222054 185004 257498
rect 184404 221818 184586 222054
rect 184822 221818 185004 222054
rect 184404 221734 185004 221818
rect 184404 221498 184586 221734
rect 184822 221498 185004 221734
rect 184404 186054 185004 221498
rect 184404 185818 184586 186054
rect 184822 185818 185004 186054
rect 184404 185734 185004 185818
rect 184404 185498 184586 185734
rect 184822 185498 185004 185734
rect 184404 150054 185004 185498
rect 184404 149818 184586 150054
rect 184822 149818 185004 150054
rect 184404 149734 185004 149818
rect 184404 149498 184586 149734
rect 184822 149498 185004 149734
rect 184404 114054 185004 149498
rect 184404 113818 184586 114054
rect 184822 113818 185004 114054
rect 184404 113734 185004 113818
rect 184404 113498 184586 113734
rect 184822 113498 185004 113734
rect 184404 78054 185004 113498
rect 184404 77818 184586 78054
rect 184822 77818 185004 78054
rect 184404 77734 185004 77818
rect 184404 77498 184586 77734
rect 184822 77498 185004 77734
rect 184404 42054 185004 77498
rect 184404 41818 184586 42054
rect 184822 41818 185004 42054
rect 184404 41734 185004 41818
rect 184404 41498 184586 41734
rect 184822 41498 185004 41734
rect 184404 6054 185004 41498
rect 184404 5818 184586 6054
rect 184822 5818 185004 6054
rect 184404 5734 185004 5818
rect 184404 5498 184586 5734
rect 184822 5498 185004 5734
rect 184404 -2186 185004 5498
rect 184404 -2422 184586 -2186
rect 184822 -2422 185004 -2186
rect 184404 -2506 185004 -2422
rect 184404 -2742 184586 -2506
rect 184822 -2742 185004 -2506
rect 184404 -3684 185004 -2742
rect 188004 693654 188604 707962
rect 188004 693418 188186 693654
rect 188422 693418 188604 693654
rect 188004 693334 188604 693418
rect 188004 693098 188186 693334
rect 188422 693098 188604 693334
rect 188004 657654 188604 693098
rect 188004 657418 188186 657654
rect 188422 657418 188604 657654
rect 188004 657334 188604 657418
rect 188004 657098 188186 657334
rect 188422 657098 188604 657334
rect 188004 621654 188604 657098
rect 188004 621418 188186 621654
rect 188422 621418 188604 621654
rect 188004 621334 188604 621418
rect 188004 621098 188186 621334
rect 188422 621098 188604 621334
rect 188004 585654 188604 621098
rect 188004 585418 188186 585654
rect 188422 585418 188604 585654
rect 188004 585334 188604 585418
rect 188004 585098 188186 585334
rect 188422 585098 188604 585334
rect 188004 549654 188604 585098
rect 188004 549418 188186 549654
rect 188422 549418 188604 549654
rect 188004 549334 188604 549418
rect 188004 549098 188186 549334
rect 188422 549098 188604 549334
rect 188004 513654 188604 549098
rect 188004 513418 188186 513654
rect 188422 513418 188604 513654
rect 188004 513334 188604 513418
rect 188004 513098 188186 513334
rect 188422 513098 188604 513334
rect 188004 477654 188604 513098
rect 188004 477418 188186 477654
rect 188422 477418 188604 477654
rect 188004 477334 188604 477418
rect 188004 477098 188186 477334
rect 188422 477098 188604 477334
rect 188004 441654 188604 477098
rect 188004 441418 188186 441654
rect 188422 441418 188604 441654
rect 188004 441334 188604 441418
rect 188004 441098 188186 441334
rect 188422 441098 188604 441334
rect 188004 405654 188604 441098
rect 188004 405418 188186 405654
rect 188422 405418 188604 405654
rect 188004 405334 188604 405418
rect 188004 405098 188186 405334
rect 188422 405098 188604 405334
rect 188004 369654 188604 405098
rect 188004 369418 188186 369654
rect 188422 369418 188604 369654
rect 188004 369334 188604 369418
rect 188004 369098 188186 369334
rect 188422 369098 188604 369334
rect 188004 333654 188604 369098
rect 188004 333418 188186 333654
rect 188422 333418 188604 333654
rect 188004 333334 188604 333418
rect 188004 333098 188186 333334
rect 188422 333098 188604 333334
rect 188004 297654 188604 333098
rect 188004 297418 188186 297654
rect 188422 297418 188604 297654
rect 188004 297334 188604 297418
rect 188004 297098 188186 297334
rect 188422 297098 188604 297334
rect 188004 261654 188604 297098
rect 188004 261418 188186 261654
rect 188422 261418 188604 261654
rect 188004 261334 188604 261418
rect 188004 261098 188186 261334
rect 188422 261098 188604 261334
rect 188004 225654 188604 261098
rect 188004 225418 188186 225654
rect 188422 225418 188604 225654
rect 188004 225334 188604 225418
rect 188004 225098 188186 225334
rect 188422 225098 188604 225334
rect 188004 189654 188604 225098
rect 188004 189418 188186 189654
rect 188422 189418 188604 189654
rect 188004 189334 188604 189418
rect 188004 189098 188186 189334
rect 188422 189098 188604 189334
rect 188004 153654 188604 189098
rect 188004 153418 188186 153654
rect 188422 153418 188604 153654
rect 188004 153334 188604 153418
rect 188004 153098 188186 153334
rect 188422 153098 188604 153334
rect 188004 117654 188604 153098
rect 188004 117418 188186 117654
rect 188422 117418 188604 117654
rect 188004 117334 188604 117418
rect 188004 117098 188186 117334
rect 188422 117098 188604 117334
rect 188004 81654 188604 117098
rect 188004 81418 188186 81654
rect 188422 81418 188604 81654
rect 188004 81334 188604 81418
rect 188004 81098 188186 81334
rect 188422 81098 188604 81334
rect 188004 45654 188604 81098
rect 188004 45418 188186 45654
rect 188422 45418 188604 45654
rect 188004 45334 188604 45418
rect 188004 45098 188186 45334
rect 188422 45098 188604 45334
rect 188004 9654 188604 45098
rect 188004 9418 188186 9654
rect 188422 9418 188604 9654
rect 188004 9334 188604 9418
rect 188004 9098 188186 9334
rect 188422 9098 188604 9334
rect 188004 -4026 188604 9098
rect 188004 -4262 188186 -4026
rect 188422 -4262 188604 -4026
rect 188004 -4346 188604 -4262
rect 188004 -4582 188186 -4346
rect 188422 -4582 188604 -4346
rect 188004 -5524 188604 -4582
rect 191604 697254 192204 709802
rect 209604 711278 210204 711300
rect 209604 711042 209786 711278
rect 210022 711042 210204 711278
rect 209604 710958 210204 711042
rect 209604 710722 209786 710958
rect 210022 710722 210204 710958
rect 206004 709438 206604 709460
rect 206004 709202 206186 709438
rect 206422 709202 206604 709438
rect 206004 709118 206604 709202
rect 206004 708882 206186 709118
rect 206422 708882 206604 709118
rect 202404 707598 203004 707620
rect 202404 707362 202586 707598
rect 202822 707362 203004 707598
rect 202404 707278 203004 707362
rect 202404 707042 202586 707278
rect 202822 707042 203004 707278
rect 191604 697018 191786 697254
rect 192022 697018 192204 697254
rect 191604 696934 192204 697018
rect 191604 696698 191786 696934
rect 192022 696698 192204 696934
rect 191604 661254 192204 696698
rect 191604 661018 191786 661254
rect 192022 661018 192204 661254
rect 191604 660934 192204 661018
rect 191604 660698 191786 660934
rect 192022 660698 192204 660934
rect 191604 625254 192204 660698
rect 191604 625018 191786 625254
rect 192022 625018 192204 625254
rect 191604 624934 192204 625018
rect 191604 624698 191786 624934
rect 192022 624698 192204 624934
rect 191604 589254 192204 624698
rect 191604 589018 191786 589254
rect 192022 589018 192204 589254
rect 191604 588934 192204 589018
rect 191604 588698 191786 588934
rect 192022 588698 192204 588934
rect 191604 553254 192204 588698
rect 191604 553018 191786 553254
rect 192022 553018 192204 553254
rect 191604 552934 192204 553018
rect 191604 552698 191786 552934
rect 192022 552698 192204 552934
rect 191604 517254 192204 552698
rect 191604 517018 191786 517254
rect 192022 517018 192204 517254
rect 191604 516934 192204 517018
rect 191604 516698 191786 516934
rect 192022 516698 192204 516934
rect 191604 481254 192204 516698
rect 191604 481018 191786 481254
rect 192022 481018 192204 481254
rect 191604 480934 192204 481018
rect 191604 480698 191786 480934
rect 192022 480698 192204 480934
rect 191604 445254 192204 480698
rect 191604 445018 191786 445254
rect 192022 445018 192204 445254
rect 191604 444934 192204 445018
rect 191604 444698 191786 444934
rect 192022 444698 192204 444934
rect 191604 409254 192204 444698
rect 191604 409018 191786 409254
rect 192022 409018 192204 409254
rect 191604 408934 192204 409018
rect 191604 408698 191786 408934
rect 192022 408698 192204 408934
rect 191604 373254 192204 408698
rect 191604 373018 191786 373254
rect 192022 373018 192204 373254
rect 191604 372934 192204 373018
rect 191604 372698 191786 372934
rect 192022 372698 192204 372934
rect 191604 337254 192204 372698
rect 191604 337018 191786 337254
rect 192022 337018 192204 337254
rect 191604 336934 192204 337018
rect 191604 336698 191786 336934
rect 192022 336698 192204 336934
rect 191604 301254 192204 336698
rect 191604 301018 191786 301254
rect 192022 301018 192204 301254
rect 191604 300934 192204 301018
rect 191604 300698 191786 300934
rect 192022 300698 192204 300934
rect 191604 265254 192204 300698
rect 191604 265018 191786 265254
rect 192022 265018 192204 265254
rect 191604 264934 192204 265018
rect 191604 264698 191786 264934
rect 192022 264698 192204 264934
rect 191604 229254 192204 264698
rect 191604 229018 191786 229254
rect 192022 229018 192204 229254
rect 191604 228934 192204 229018
rect 191604 228698 191786 228934
rect 192022 228698 192204 228934
rect 191604 193254 192204 228698
rect 191604 193018 191786 193254
rect 192022 193018 192204 193254
rect 191604 192934 192204 193018
rect 191604 192698 191786 192934
rect 192022 192698 192204 192934
rect 191604 157254 192204 192698
rect 191604 157018 191786 157254
rect 192022 157018 192204 157254
rect 191604 156934 192204 157018
rect 191604 156698 191786 156934
rect 192022 156698 192204 156934
rect 191604 121254 192204 156698
rect 191604 121018 191786 121254
rect 192022 121018 192204 121254
rect 191604 120934 192204 121018
rect 191604 120698 191786 120934
rect 192022 120698 192204 120934
rect 191604 85254 192204 120698
rect 191604 85018 191786 85254
rect 192022 85018 192204 85254
rect 191604 84934 192204 85018
rect 191604 84698 191786 84934
rect 192022 84698 192204 84934
rect 191604 49254 192204 84698
rect 191604 49018 191786 49254
rect 192022 49018 192204 49254
rect 191604 48934 192204 49018
rect 191604 48698 191786 48934
rect 192022 48698 192204 48934
rect 191604 13254 192204 48698
rect 191604 13018 191786 13254
rect 192022 13018 192204 13254
rect 191604 12934 192204 13018
rect 191604 12698 191786 12934
rect 192022 12698 192204 12934
rect 173604 -7022 173786 -6786
rect 174022 -7022 174204 -6786
rect 173604 -7106 174204 -7022
rect 173604 -7342 173786 -7106
rect 174022 -7342 174204 -7106
rect 173604 -7364 174204 -7342
rect 191604 -5866 192204 12698
rect 198804 705758 199404 705780
rect 198804 705522 198986 705758
rect 199222 705522 199404 705758
rect 198804 705438 199404 705522
rect 198804 705202 198986 705438
rect 199222 705202 199404 705438
rect 198804 668454 199404 705202
rect 198804 668218 198986 668454
rect 199222 668218 199404 668454
rect 198804 668134 199404 668218
rect 198804 667898 198986 668134
rect 199222 667898 199404 668134
rect 198804 632454 199404 667898
rect 198804 632218 198986 632454
rect 199222 632218 199404 632454
rect 198804 632134 199404 632218
rect 198804 631898 198986 632134
rect 199222 631898 199404 632134
rect 198804 596454 199404 631898
rect 198804 596218 198986 596454
rect 199222 596218 199404 596454
rect 198804 596134 199404 596218
rect 198804 595898 198986 596134
rect 199222 595898 199404 596134
rect 198804 560454 199404 595898
rect 198804 560218 198986 560454
rect 199222 560218 199404 560454
rect 198804 560134 199404 560218
rect 198804 559898 198986 560134
rect 199222 559898 199404 560134
rect 198804 524454 199404 559898
rect 198804 524218 198986 524454
rect 199222 524218 199404 524454
rect 198804 524134 199404 524218
rect 198804 523898 198986 524134
rect 199222 523898 199404 524134
rect 198804 488454 199404 523898
rect 198804 488218 198986 488454
rect 199222 488218 199404 488454
rect 198804 488134 199404 488218
rect 198804 487898 198986 488134
rect 199222 487898 199404 488134
rect 198804 452454 199404 487898
rect 198804 452218 198986 452454
rect 199222 452218 199404 452454
rect 198804 452134 199404 452218
rect 198804 451898 198986 452134
rect 199222 451898 199404 452134
rect 198804 416454 199404 451898
rect 198804 416218 198986 416454
rect 199222 416218 199404 416454
rect 198804 416134 199404 416218
rect 198804 415898 198986 416134
rect 199222 415898 199404 416134
rect 198804 380454 199404 415898
rect 198804 380218 198986 380454
rect 199222 380218 199404 380454
rect 198804 380134 199404 380218
rect 198804 379898 198986 380134
rect 199222 379898 199404 380134
rect 198804 344454 199404 379898
rect 198804 344218 198986 344454
rect 199222 344218 199404 344454
rect 198804 344134 199404 344218
rect 198804 343898 198986 344134
rect 199222 343898 199404 344134
rect 198804 308454 199404 343898
rect 198804 308218 198986 308454
rect 199222 308218 199404 308454
rect 198804 308134 199404 308218
rect 198804 307898 198986 308134
rect 199222 307898 199404 308134
rect 198804 272454 199404 307898
rect 198804 272218 198986 272454
rect 199222 272218 199404 272454
rect 198804 272134 199404 272218
rect 198804 271898 198986 272134
rect 199222 271898 199404 272134
rect 198804 236454 199404 271898
rect 198804 236218 198986 236454
rect 199222 236218 199404 236454
rect 198804 236134 199404 236218
rect 198804 235898 198986 236134
rect 199222 235898 199404 236134
rect 198804 200454 199404 235898
rect 198804 200218 198986 200454
rect 199222 200218 199404 200454
rect 198804 200134 199404 200218
rect 198804 199898 198986 200134
rect 199222 199898 199404 200134
rect 198804 164454 199404 199898
rect 198804 164218 198986 164454
rect 199222 164218 199404 164454
rect 198804 164134 199404 164218
rect 198804 163898 198986 164134
rect 199222 163898 199404 164134
rect 198804 128454 199404 163898
rect 198804 128218 198986 128454
rect 199222 128218 199404 128454
rect 198804 128134 199404 128218
rect 198804 127898 198986 128134
rect 199222 127898 199404 128134
rect 198804 92454 199404 127898
rect 198804 92218 198986 92454
rect 199222 92218 199404 92454
rect 198804 92134 199404 92218
rect 198804 91898 198986 92134
rect 199222 91898 199404 92134
rect 198804 56454 199404 91898
rect 198804 56218 198986 56454
rect 199222 56218 199404 56454
rect 198804 56134 199404 56218
rect 198804 55898 198986 56134
rect 199222 55898 199404 56134
rect 198804 20454 199404 55898
rect 198804 20218 198986 20454
rect 199222 20218 199404 20454
rect 198804 20134 199404 20218
rect 198804 19898 198986 20134
rect 199222 19898 199404 20134
rect 198804 -1266 199404 19898
rect 198804 -1502 198986 -1266
rect 199222 -1502 199404 -1266
rect 198804 -1586 199404 -1502
rect 198804 -1822 198986 -1586
rect 199222 -1822 199404 -1586
rect 198804 -1844 199404 -1822
rect 202404 672054 203004 707042
rect 202404 671818 202586 672054
rect 202822 671818 203004 672054
rect 202404 671734 203004 671818
rect 202404 671498 202586 671734
rect 202822 671498 203004 671734
rect 202404 636054 203004 671498
rect 202404 635818 202586 636054
rect 202822 635818 203004 636054
rect 202404 635734 203004 635818
rect 202404 635498 202586 635734
rect 202822 635498 203004 635734
rect 202404 600054 203004 635498
rect 202404 599818 202586 600054
rect 202822 599818 203004 600054
rect 202404 599734 203004 599818
rect 202404 599498 202586 599734
rect 202822 599498 203004 599734
rect 202404 564054 203004 599498
rect 202404 563818 202586 564054
rect 202822 563818 203004 564054
rect 202404 563734 203004 563818
rect 202404 563498 202586 563734
rect 202822 563498 203004 563734
rect 202404 528054 203004 563498
rect 202404 527818 202586 528054
rect 202822 527818 203004 528054
rect 202404 527734 203004 527818
rect 202404 527498 202586 527734
rect 202822 527498 203004 527734
rect 202404 492054 203004 527498
rect 202404 491818 202586 492054
rect 202822 491818 203004 492054
rect 202404 491734 203004 491818
rect 202404 491498 202586 491734
rect 202822 491498 203004 491734
rect 202404 456054 203004 491498
rect 202404 455818 202586 456054
rect 202822 455818 203004 456054
rect 202404 455734 203004 455818
rect 202404 455498 202586 455734
rect 202822 455498 203004 455734
rect 202404 420054 203004 455498
rect 202404 419818 202586 420054
rect 202822 419818 203004 420054
rect 202404 419734 203004 419818
rect 202404 419498 202586 419734
rect 202822 419498 203004 419734
rect 202404 384054 203004 419498
rect 202404 383818 202586 384054
rect 202822 383818 203004 384054
rect 202404 383734 203004 383818
rect 202404 383498 202586 383734
rect 202822 383498 203004 383734
rect 202404 348054 203004 383498
rect 202404 347818 202586 348054
rect 202822 347818 203004 348054
rect 202404 347734 203004 347818
rect 202404 347498 202586 347734
rect 202822 347498 203004 347734
rect 202404 312054 203004 347498
rect 202404 311818 202586 312054
rect 202822 311818 203004 312054
rect 202404 311734 203004 311818
rect 202404 311498 202586 311734
rect 202822 311498 203004 311734
rect 202404 276054 203004 311498
rect 202404 275818 202586 276054
rect 202822 275818 203004 276054
rect 202404 275734 203004 275818
rect 202404 275498 202586 275734
rect 202822 275498 203004 275734
rect 202404 240054 203004 275498
rect 202404 239818 202586 240054
rect 202822 239818 203004 240054
rect 202404 239734 203004 239818
rect 202404 239498 202586 239734
rect 202822 239498 203004 239734
rect 202404 204054 203004 239498
rect 202404 203818 202586 204054
rect 202822 203818 203004 204054
rect 202404 203734 203004 203818
rect 202404 203498 202586 203734
rect 202822 203498 203004 203734
rect 202404 168054 203004 203498
rect 202404 167818 202586 168054
rect 202822 167818 203004 168054
rect 202404 167734 203004 167818
rect 202404 167498 202586 167734
rect 202822 167498 203004 167734
rect 202404 132054 203004 167498
rect 202404 131818 202586 132054
rect 202822 131818 203004 132054
rect 202404 131734 203004 131818
rect 202404 131498 202586 131734
rect 202822 131498 203004 131734
rect 202404 96054 203004 131498
rect 202404 95818 202586 96054
rect 202822 95818 203004 96054
rect 202404 95734 203004 95818
rect 202404 95498 202586 95734
rect 202822 95498 203004 95734
rect 202404 60054 203004 95498
rect 202404 59818 202586 60054
rect 202822 59818 203004 60054
rect 202404 59734 203004 59818
rect 202404 59498 202586 59734
rect 202822 59498 203004 59734
rect 202404 24054 203004 59498
rect 202404 23818 202586 24054
rect 202822 23818 203004 24054
rect 202404 23734 203004 23818
rect 202404 23498 202586 23734
rect 202822 23498 203004 23734
rect 202404 -3106 203004 23498
rect 202404 -3342 202586 -3106
rect 202822 -3342 203004 -3106
rect 202404 -3426 203004 -3342
rect 202404 -3662 202586 -3426
rect 202822 -3662 203004 -3426
rect 202404 -3684 203004 -3662
rect 206004 675654 206604 708882
rect 206004 675418 206186 675654
rect 206422 675418 206604 675654
rect 206004 675334 206604 675418
rect 206004 675098 206186 675334
rect 206422 675098 206604 675334
rect 206004 639654 206604 675098
rect 206004 639418 206186 639654
rect 206422 639418 206604 639654
rect 206004 639334 206604 639418
rect 206004 639098 206186 639334
rect 206422 639098 206604 639334
rect 206004 603654 206604 639098
rect 206004 603418 206186 603654
rect 206422 603418 206604 603654
rect 206004 603334 206604 603418
rect 206004 603098 206186 603334
rect 206422 603098 206604 603334
rect 206004 567654 206604 603098
rect 206004 567418 206186 567654
rect 206422 567418 206604 567654
rect 206004 567334 206604 567418
rect 206004 567098 206186 567334
rect 206422 567098 206604 567334
rect 206004 531654 206604 567098
rect 206004 531418 206186 531654
rect 206422 531418 206604 531654
rect 206004 531334 206604 531418
rect 206004 531098 206186 531334
rect 206422 531098 206604 531334
rect 206004 495654 206604 531098
rect 206004 495418 206186 495654
rect 206422 495418 206604 495654
rect 206004 495334 206604 495418
rect 206004 495098 206186 495334
rect 206422 495098 206604 495334
rect 206004 459654 206604 495098
rect 206004 459418 206186 459654
rect 206422 459418 206604 459654
rect 206004 459334 206604 459418
rect 206004 459098 206186 459334
rect 206422 459098 206604 459334
rect 206004 423654 206604 459098
rect 206004 423418 206186 423654
rect 206422 423418 206604 423654
rect 206004 423334 206604 423418
rect 206004 423098 206186 423334
rect 206422 423098 206604 423334
rect 206004 387654 206604 423098
rect 206004 387418 206186 387654
rect 206422 387418 206604 387654
rect 206004 387334 206604 387418
rect 206004 387098 206186 387334
rect 206422 387098 206604 387334
rect 206004 351654 206604 387098
rect 206004 351418 206186 351654
rect 206422 351418 206604 351654
rect 206004 351334 206604 351418
rect 206004 351098 206186 351334
rect 206422 351098 206604 351334
rect 206004 315654 206604 351098
rect 206004 315418 206186 315654
rect 206422 315418 206604 315654
rect 206004 315334 206604 315418
rect 206004 315098 206186 315334
rect 206422 315098 206604 315334
rect 206004 279654 206604 315098
rect 206004 279418 206186 279654
rect 206422 279418 206604 279654
rect 206004 279334 206604 279418
rect 206004 279098 206186 279334
rect 206422 279098 206604 279334
rect 206004 243654 206604 279098
rect 206004 243418 206186 243654
rect 206422 243418 206604 243654
rect 206004 243334 206604 243418
rect 206004 243098 206186 243334
rect 206422 243098 206604 243334
rect 206004 207654 206604 243098
rect 206004 207418 206186 207654
rect 206422 207418 206604 207654
rect 206004 207334 206604 207418
rect 206004 207098 206186 207334
rect 206422 207098 206604 207334
rect 206004 171654 206604 207098
rect 206004 171418 206186 171654
rect 206422 171418 206604 171654
rect 206004 171334 206604 171418
rect 206004 171098 206186 171334
rect 206422 171098 206604 171334
rect 206004 135654 206604 171098
rect 206004 135418 206186 135654
rect 206422 135418 206604 135654
rect 206004 135334 206604 135418
rect 206004 135098 206186 135334
rect 206422 135098 206604 135334
rect 206004 99654 206604 135098
rect 206004 99418 206186 99654
rect 206422 99418 206604 99654
rect 206004 99334 206604 99418
rect 206004 99098 206186 99334
rect 206422 99098 206604 99334
rect 206004 63654 206604 99098
rect 206004 63418 206186 63654
rect 206422 63418 206604 63654
rect 206004 63334 206604 63418
rect 206004 63098 206186 63334
rect 206422 63098 206604 63334
rect 206004 27654 206604 63098
rect 206004 27418 206186 27654
rect 206422 27418 206604 27654
rect 206004 27334 206604 27418
rect 206004 27098 206186 27334
rect 206422 27098 206604 27334
rect 206004 -4946 206604 27098
rect 206004 -5182 206186 -4946
rect 206422 -5182 206604 -4946
rect 206004 -5266 206604 -5182
rect 206004 -5502 206186 -5266
rect 206422 -5502 206604 -5266
rect 206004 -5524 206604 -5502
rect 209604 679254 210204 710722
rect 227604 710358 228204 711300
rect 227604 710122 227786 710358
rect 228022 710122 228204 710358
rect 227604 710038 228204 710122
rect 227604 709802 227786 710038
rect 228022 709802 228204 710038
rect 224004 708518 224604 709460
rect 224004 708282 224186 708518
rect 224422 708282 224604 708518
rect 224004 708198 224604 708282
rect 224004 707962 224186 708198
rect 224422 707962 224604 708198
rect 220404 706678 221004 707620
rect 220404 706442 220586 706678
rect 220822 706442 221004 706678
rect 220404 706358 221004 706442
rect 220404 706122 220586 706358
rect 220822 706122 221004 706358
rect 209604 679018 209786 679254
rect 210022 679018 210204 679254
rect 209604 678934 210204 679018
rect 209604 678698 209786 678934
rect 210022 678698 210204 678934
rect 209604 643254 210204 678698
rect 209604 643018 209786 643254
rect 210022 643018 210204 643254
rect 209604 642934 210204 643018
rect 209604 642698 209786 642934
rect 210022 642698 210204 642934
rect 209604 607254 210204 642698
rect 209604 607018 209786 607254
rect 210022 607018 210204 607254
rect 209604 606934 210204 607018
rect 209604 606698 209786 606934
rect 210022 606698 210204 606934
rect 209604 571254 210204 606698
rect 209604 571018 209786 571254
rect 210022 571018 210204 571254
rect 209604 570934 210204 571018
rect 209604 570698 209786 570934
rect 210022 570698 210204 570934
rect 209604 535254 210204 570698
rect 209604 535018 209786 535254
rect 210022 535018 210204 535254
rect 209604 534934 210204 535018
rect 209604 534698 209786 534934
rect 210022 534698 210204 534934
rect 209604 499254 210204 534698
rect 209604 499018 209786 499254
rect 210022 499018 210204 499254
rect 209604 498934 210204 499018
rect 209604 498698 209786 498934
rect 210022 498698 210204 498934
rect 209604 463254 210204 498698
rect 209604 463018 209786 463254
rect 210022 463018 210204 463254
rect 209604 462934 210204 463018
rect 209604 462698 209786 462934
rect 210022 462698 210204 462934
rect 209604 427254 210204 462698
rect 209604 427018 209786 427254
rect 210022 427018 210204 427254
rect 209604 426934 210204 427018
rect 209604 426698 209786 426934
rect 210022 426698 210204 426934
rect 209604 391254 210204 426698
rect 209604 391018 209786 391254
rect 210022 391018 210204 391254
rect 209604 390934 210204 391018
rect 209604 390698 209786 390934
rect 210022 390698 210204 390934
rect 209604 355254 210204 390698
rect 209604 355018 209786 355254
rect 210022 355018 210204 355254
rect 209604 354934 210204 355018
rect 209604 354698 209786 354934
rect 210022 354698 210204 354934
rect 209604 319254 210204 354698
rect 209604 319018 209786 319254
rect 210022 319018 210204 319254
rect 209604 318934 210204 319018
rect 209604 318698 209786 318934
rect 210022 318698 210204 318934
rect 209604 283254 210204 318698
rect 209604 283018 209786 283254
rect 210022 283018 210204 283254
rect 209604 282934 210204 283018
rect 209604 282698 209786 282934
rect 210022 282698 210204 282934
rect 209604 247254 210204 282698
rect 209604 247018 209786 247254
rect 210022 247018 210204 247254
rect 209604 246934 210204 247018
rect 209604 246698 209786 246934
rect 210022 246698 210204 246934
rect 209604 211254 210204 246698
rect 209604 211018 209786 211254
rect 210022 211018 210204 211254
rect 209604 210934 210204 211018
rect 209604 210698 209786 210934
rect 210022 210698 210204 210934
rect 209604 175254 210204 210698
rect 209604 175018 209786 175254
rect 210022 175018 210204 175254
rect 209604 174934 210204 175018
rect 209604 174698 209786 174934
rect 210022 174698 210204 174934
rect 209604 139254 210204 174698
rect 209604 139018 209786 139254
rect 210022 139018 210204 139254
rect 209604 138934 210204 139018
rect 209604 138698 209786 138934
rect 210022 138698 210204 138934
rect 209604 103254 210204 138698
rect 209604 103018 209786 103254
rect 210022 103018 210204 103254
rect 209604 102934 210204 103018
rect 209604 102698 209786 102934
rect 210022 102698 210204 102934
rect 209604 67254 210204 102698
rect 209604 67018 209786 67254
rect 210022 67018 210204 67254
rect 209604 66934 210204 67018
rect 209604 66698 209786 66934
rect 210022 66698 210204 66934
rect 209604 31254 210204 66698
rect 209604 31018 209786 31254
rect 210022 31018 210204 31254
rect 209604 30934 210204 31018
rect 209604 30698 209786 30934
rect 210022 30698 210204 30934
rect 191604 -6102 191786 -5866
rect 192022 -6102 192204 -5866
rect 191604 -6186 192204 -6102
rect 191604 -6422 191786 -6186
rect 192022 -6422 192204 -6186
rect 191604 -7364 192204 -6422
rect 209604 -6786 210204 30698
rect 216804 704838 217404 705780
rect 216804 704602 216986 704838
rect 217222 704602 217404 704838
rect 216804 704518 217404 704602
rect 216804 704282 216986 704518
rect 217222 704282 217404 704518
rect 216804 686454 217404 704282
rect 216804 686218 216986 686454
rect 217222 686218 217404 686454
rect 216804 686134 217404 686218
rect 216804 685898 216986 686134
rect 217222 685898 217404 686134
rect 216804 650454 217404 685898
rect 216804 650218 216986 650454
rect 217222 650218 217404 650454
rect 216804 650134 217404 650218
rect 216804 649898 216986 650134
rect 217222 649898 217404 650134
rect 216804 614454 217404 649898
rect 216804 614218 216986 614454
rect 217222 614218 217404 614454
rect 216804 614134 217404 614218
rect 216804 613898 216986 614134
rect 217222 613898 217404 614134
rect 216804 578454 217404 613898
rect 216804 578218 216986 578454
rect 217222 578218 217404 578454
rect 216804 578134 217404 578218
rect 216804 577898 216986 578134
rect 217222 577898 217404 578134
rect 216804 542454 217404 577898
rect 216804 542218 216986 542454
rect 217222 542218 217404 542454
rect 216804 542134 217404 542218
rect 216804 541898 216986 542134
rect 217222 541898 217404 542134
rect 216804 506454 217404 541898
rect 216804 506218 216986 506454
rect 217222 506218 217404 506454
rect 216804 506134 217404 506218
rect 216804 505898 216986 506134
rect 217222 505898 217404 506134
rect 216804 470454 217404 505898
rect 216804 470218 216986 470454
rect 217222 470218 217404 470454
rect 216804 470134 217404 470218
rect 216804 469898 216986 470134
rect 217222 469898 217404 470134
rect 216804 434454 217404 469898
rect 216804 434218 216986 434454
rect 217222 434218 217404 434454
rect 216804 434134 217404 434218
rect 216804 433898 216986 434134
rect 217222 433898 217404 434134
rect 216804 398454 217404 433898
rect 216804 398218 216986 398454
rect 217222 398218 217404 398454
rect 216804 398134 217404 398218
rect 216804 397898 216986 398134
rect 217222 397898 217404 398134
rect 216804 362454 217404 397898
rect 216804 362218 216986 362454
rect 217222 362218 217404 362454
rect 216804 362134 217404 362218
rect 216804 361898 216986 362134
rect 217222 361898 217404 362134
rect 216804 326454 217404 361898
rect 216804 326218 216986 326454
rect 217222 326218 217404 326454
rect 216804 326134 217404 326218
rect 216804 325898 216986 326134
rect 217222 325898 217404 326134
rect 216804 290454 217404 325898
rect 216804 290218 216986 290454
rect 217222 290218 217404 290454
rect 216804 290134 217404 290218
rect 216804 289898 216986 290134
rect 217222 289898 217404 290134
rect 216804 254454 217404 289898
rect 216804 254218 216986 254454
rect 217222 254218 217404 254454
rect 216804 254134 217404 254218
rect 216804 253898 216986 254134
rect 217222 253898 217404 254134
rect 216804 218454 217404 253898
rect 216804 218218 216986 218454
rect 217222 218218 217404 218454
rect 216804 218134 217404 218218
rect 216804 217898 216986 218134
rect 217222 217898 217404 218134
rect 216804 182454 217404 217898
rect 216804 182218 216986 182454
rect 217222 182218 217404 182454
rect 216804 182134 217404 182218
rect 216804 181898 216986 182134
rect 217222 181898 217404 182134
rect 216804 146454 217404 181898
rect 216804 146218 216986 146454
rect 217222 146218 217404 146454
rect 216804 146134 217404 146218
rect 216804 145898 216986 146134
rect 217222 145898 217404 146134
rect 216804 110454 217404 145898
rect 216804 110218 216986 110454
rect 217222 110218 217404 110454
rect 216804 110134 217404 110218
rect 216804 109898 216986 110134
rect 217222 109898 217404 110134
rect 216804 74454 217404 109898
rect 216804 74218 216986 74454
rect 217222 74218 217404 74454
rect 216804 74134 217404 74218
rect 216804 73898 216986 74134
rect 217222 73898 217404 74134
rect 216804 38454 217404 73898
rect 216804 38218 216986 38454
rect 217222 38218 217404 38454
rect 216804 38134 217404 38218
rect 216804 37898 216986 38134
rect 217222 37898 217404 38134
rect 216804 2454 217404 37898
rect 216804 2218 216986 2454
rect 217222 2218 217404 2454
rect 216804 2134 217404 2218
rect 216804 1898 216986 2134
rect 217222 1898 217404 2134
rect 216804 -346 217404 1898
rect 216804 -582 216986 -346
rect 217222 -582 217404 -346
rect 216804 -666 217404 -582
rect 216804 -902 216986 -666
rect 217222 -902 217404 -666
rect 216804 -1844 217404 -902
rect 220404 690054 221004 706122
rect 220404 689818 220586 690054
rect 220822 689818 221004 690054
rect 220404 689734 221004 689818
rect 220404 689498 220586 689734
rect 220822 689498 221004 689734
rect 220404 654054 221004 689498
rect 220404 653818 220586 654054
rect 220822 653818 221004 654054
rect 220404 653734 221004 653818
rect 220404 653498 220586 653734
rect 220822 653498 221004 653734
rect 220404 618054 221004 653498
rect 220404 617818 220586 618054
rect 220822 617818 221004 618054
rect 220404 617734 221004 617818
rect 220404 617498 220586 617734
rect 220822 617498 221004 617734
rect 220404 582054 221004 617498
rect 220404 581818 220586 582054
rect 220822 581818 221004 582054
rect 220404 581734 221004 581818
rect 220404 581498 220586 581734
rect 220822 581498 221004 581734
rect 220404 546054 221004 581498
rect 220404 545818 220586 546054
rect 220822 545818 221004 546054
rect 220404 545734 221004 545818
rect 220404 545498 220586 545734
rect 220822 545498 221004 545734
rect 220404 510054 221004 545498
rect 220404 509818 220586 510054
rect 220822 509818 221004 510054
rect 220404 509734 221004 509818
rect 220404 509498 220586 509734
rect 220822 509498 221004 509734
rect 220404 474054 221004 509498
rect 220404 473818 220586 474054
rect 220822 473818 221004 474054
rect 220404 473734 221004 473818
rect 220404 473498 220586 473734
rect 220822 473498 221004 473734
rect 220404 438054 221004 473498
rect 220404 437818 220586 438054
rect 220822 437818 221004 438054
rect 220404 437734 221004 437818
rect 220404 437498 220586 437734
rect 220822 437498 221004 437734
rect 220404 402054 221004 437498
rect 220404 401818 220586 402054
rect 220822 401818 221004 402054
rect 220404 401734 221004 401818
rect 220404 401498 220586 401734
rect 220822 401498 221004 401734
rect 220404 366054 221004 401498
rect 220404 365818 220586 366054
rect 220822 365818 221004 366054
rect 220404 365734 221004 365818
rect 220404 365498 220586 365734
rect 220822 365498 221004 365734
rect 220404 330054 221004 365498
rect 220404 329818 220586 330054
rect 220822 329818 221004 330054
rect 220404 329734 221004 329818
rect 220404 329498 220586 329734
rect 220822 329498 221004 329734
rect 220404 294054 221004 329498
rect 220404 293818 220586 294054
rect 220822 293818 221004 294054
rect 220404 293734 221004 293818
rect 220404 293498 220586 293734
rect 220822 293498 221004 293734
rect 220404 258054 221004 293498
rect 220404 257818 220586 258054
rect 220822 257818 221004 258054
rect 220404 257734 221004 257818
rect 220404 257498 220586 257734
rect 220822 257498 221004 257734
rect 220404 222054 221004 257498
rect 220404 221818 220586 222054
rect 220822 221818 221004 222054
rect 220404 221734 221004 221818
rect 220404 221498 220586 221734
rect 220822 221498 221004 221734
rect 220404 186054 221004 221498
rect 220404 185818 220586 186054
rect 220822 185818 221004 186054
rect 220404 185734 221004 185818
rect 220404 185498 220586 185734
rect 220822 185498 221004 185734
rect 220404 150054 221004 185498
rect 220404 149818 220586 150054
rect 220822 149818 221004 150054
rect 220404 149734 221004 149818
rect 220404 149498 220586 149734
rect 220822 149498 221004 149734
rect 220404 114054 221004 149498
rect 220404 113818 220586 114054
rect 220822 113818 221004 114054
rect 220404 113734 221004 113818
rect 220404 113498 220586 113734
rect 220822 113498 221004 113734
rect 220404 78054 221004 113498
rect 220404 77818 220586 78054
rect 220822 77818 221004 78054
rect 220404 77734 221004 77818
rect 220404 77498 220586 77734
rect 220822 77498 221004 77734
rect 220404 42054 221004 77498
rect 220404 41818 220586 42054
rect 220822 41818 221004 42054
rect 220404 41734 221004 41818
rect 220404 41498 220586 41734
rect 220822 41498 221004 41734
rect 220404 6054 221004 41498
rect 220404 5818 220586 6054
rect 220822 5818 221004 6054
rect 220404 5734 221004 5818
rect 220404 5498 220586 5734
rect 220822 5498 221004 5734
rect 220404 -2186 221004 5498
rect 220404 -2422 220586 -2186
rect 220822 -2422 221004 -2186
rect 220404 -2506 221004 -2422
rect 220404 -2742 220586 -2506
rect 220822 -2742 221004 -2506
rect 220404 -3684 221004 -2742
rect 224004 693654 224604 707962
rect 224004 693418 224186 693654
rect 224422 693418 224604 693654
rect 224004 693334 224604 693418
rect 224004 693098 224186 693334
rect 224422 693098 224604 693334
rect 224004 657654 224604 693098
rect 224004 657418 224186 657654
rect 224422 657418 224604 657654
rect 224004 657334 224604 657418
rect 224004 657098 224186 657334
rect 224422 657098 224604 657334
rect 224004 621654 224604 657098
rect 224004 621418 224186 621654
rect 224422 621418 224604 621654
rect 224004 621334 224604 621418
rect 224004 621098 224186 621334
rect 224422 621098 224604 621334
rect 224004 585654 224604 621098
rect 224004 585418 224186 585654
rect 224422 585418 224604 585654
rect 224004 585334 224604 585418
rect 224004 585098 224186 585334
rect 224422 585098 224604 585334
rect 224004 549654 224604 585098
rect 224004 549418 224186 549654
rect 224422 549418 224604 549654
rect 224004 549334 224604 549418
rect 224004 549098 224186 549334
rect 224422 549098 224604 549334
rect 224004 513654 224604 549098
rect 224004 513418 224186 513654
rect 224422 513418 224604 513654
rect 224004 513334 224604 513418
rect 224004 513098 224186 513334
rect 224422 513098 224604 513334
rect 224004 477654 224604 513098
rect 224004 477418 224186 477654
rect 224422 477418 224604 477654
rect 224004 477334 224604 477418
rect 224004 477098 224186 477334
rect 224422 477098 224604 477334
rect 224004 441654 224604 477098
rect 224004 441418 224186 441654
rect 224422 441418 224604 441654
rect 224004 441334 224604 441418
rect 224004 441098 224186 441334
rect 224422 441098 224604 441334
rect 224004 405654 224604 441098
rect 224004 405418 224186 405654
rect 224422 405418 224604 405654
rect 224004 405334 224604 405418
rect 224004 405098 224186 405334
rect 224422 405098 224604 405334
rect 224004 369654 224604 405098
rect 224004 369418 224186 369654
rect 224422 369418 224604 369654
rect 224004 369334 224604 369418
rect 224004 369098 224186 369334
rect 224422 369098 224604 369334
rect 224004 333654 224604 369098
rect 224004 333418 224186 333654
rect 224422 333418 224604 333654
rect 224004 333334 224604 333418
rect 224004 333098 224186 333334
rect 224422 333098 224604 333334
rect 224004 297654 224604 333098
rect 224004 297418 224186 297654
rect 224422 297418 224604 297654
rect 224004 297334 224604 297418
rect 224004 297098 224186 297334
rect 224422 297098 224604 297334
rect 224004 261654 224604 297098
rect 224004 261418 224186 261654
rect 224422 261418 224604 261654
rect 224004 261334 224604 261418
rect 224004 261098 224186 261334
rect 224422 261098 224604 261334
rect 224004 225654 224604 261098
rect 224004 225418 224186 225654
rect 224422 225418 224604 225654
rect 224004 225334 224604 225418
rect 224004 225098 224186 225334
rect 224422 225098 224604 225334
rect 224004 189654 224604 225098
rect 224004 189418 224186 189654
rect 224422 189418 224604 189654
rect 224004 189334 224604 189418
rect 224004 189098 224186 189334
rect 224422 189098 224604 189334
rect 224004 153654 224604 189098
rect 224004 153418 224186 153654
rect 224422 153418 224604 153654
rect 224004 153334 224604 153418
rect 224004 153098 224186 153334
rect 224422 153098 224604 153334
rect 224004 117654 224604 153098
rect 224004 117418 224186 117654
rect 224422 117418 224604 117654
rect 224004 117334 224604 117418
rect 224004 117098 224186 117334
rect 224422 117098 224604 117334
rect 224004 81654 224604 117098
rect 224004 81418 224186 81654
rect 224422 81418 224604 81654
rect 224004 81334 224604 81418
rect 224004 81098 224186 81334
rect 224422 81098 224604 81334
rect 224004 45654 224604 81098
rect 224004 45418 224186 45654
rect 224422 45418 224604 45654
rect 224004 45334 224604 45418
rect 224004 45098 224186 45334
rect 224422 45098 224604 45334
rect 224004 9654 224604 45098
rect 224004 9418 224186 9654
rect 224422 9418 224604 9654
rect 224004 9334 224604 9418
rect 224004 9098 224186 9334
rect 224422 9098 224604 9334
rect 224004 -4026 224604 9098
rect 224004 -4262 224186 -4026
rect 224422 -4262 224604 -4026
rect 224004 -4346 224604 -4262
rect 224004 -4582 224186 -4346
rect 224422 -4582 224604 -4346
rect 224004 -5524 224604 -4582
rect 227604 697254 228204 709802
rect 245604 711278 246204 711300
rect 245604 711042 245786 711278
rect 246022 711042 246204 711278
rect 245604 710958 246204 711042
rect 245604 710722 245786 710958
rect 246022 710722 246204 710958
rect 242004 709438 242604 709460
rect 242004 709202 242186 709438
rect 242422 709202 242604 709438
rect 242004 709118 242604 709202
rect 242004 708882 242186 709118
rect 242422 708882 242604 709118
rect 238404 707598 239004 707620
rect 238404 707362 238586 707598
rect 238822 707362 239004 707598
rect 238404 707278 239004 707362
rect 238404 707042 238586 707278
rect 238822 707042 239004 707278
rect 227604 697018 227786 697254
rect 228022 697018 228204 697254
rect 227604 696934 228204 697018
rect 227604 696698 227786 696934
rect 228022 696698 228204 696934
rect 227604 661254 228204 696698
rect 227604 661018 227786 661254
rect 228022 661018 228204 661254
rect 227604 660934 228204 661018
rect 227604 660698 227786 660934
rect 228022 660698 228204 660934
rect 227604 625254 228204 660698
rect 227604 625018 227786 625254
rect 228022 625018 228204 625254
rect 227604 624934 228204 625018
rect 227604 624698 227786 624934
rect 228022 624698 228204 624934
rect 227604 589254 228204 624698
rect 227604 589018 227786 589254
rect 228022 589018 228204 589254
rect 227604 588934 228204 589018
rect 227604 588698 227786 588934
rect 228022 588698 228204 588934
rect 227604 553254 228204 588698
rect 227604 553018 227786 553254
rect 228022 553018 228204 553254
rect 227604 552934 228204 553018
rect 227604 552698 227786 552934
rect 228022 552698 228204 552934
rect 227604 517254 228204 552698
rect 227604 517018 227786 517254
rect 228022 517018 228204 517254
rect 227604 516934 228204 517018
rect 227604 516698 227786 516934
rect 228022 516698 228204 516934
rect 227604 481254 228204 516698
rect 227604 481018 227786 481254
rect 228022 481018 228204 481254
rect 227604 480934 228204 481018
rect 227604 480698 227786 480934
rect 228022 480698 228204 480934
rect 227604 445254 228204 480698
rect 227604 445018 227786 445254
rect 228022 445018 228204 445254
rect 227604 444934 228204 445018
rect 227604 444698 227786 444934
rect 228022 444698 228204 444934
rect 227604 409254 228204 444698
rect 227604 409018 227786 409254
rect 228022 409018 228204 409254
rect 227604 408934 228204 409018
rect 227604 408698 227786 408934
rect 228022 408698 228204 408934
rect 227604 373254 228204 408698
rect 234804 705758 235404 705780
rect 234804 705522 234986 705758
rect 235222 705522 235404 705758
rect 234804 705438 235404 705522
rect 234804 705202 234986 705438
rect 235222 705202 235404 705438
rect 234804 668454 235404 705202
rect 234804 668218 234986 668454
rect 235222 668218 235404 668454
rect 234804 668134 235404 668218
rect 234804 667898 234986 668134
rect 235222 667898 235404 668134
rect 234804 632454 235404 667898
rect 234804 632218 234986 632454
rect 235222 632218 235404 632454
rect 234804 632134 235404 632218
rect 234804 631898 234986 632134
rect 235222 631898 235404 632134
rect 234804 596454 235404 631898
rect 234804 596218 234986 596454
rect 235222 596218 235404 596454
rect 234804 596134 235404 596218
rect 234804 595898 234986 596134
rect 235222 595898 235404 596134
rect 234804 560454 235404 595898
rect 234804 560218 234986 560454
rect 235222 560218 235404 560454
rect 234804 560134 235404 560218
rect 234804 559898 234986 560134
rect 235222 559898 235404 560134
rect 234804 524454 235404 559898
rect 234804 524218 234986 524454
rect 235222 524218 235404 524454
rect 234804 524134 235404 524218
rect 234804 523898 234986 524134
rect 235222 523898 235404 524134
rect 234804 488454 235404 523898
rect 234804 488218 234986 488454
rect 235222 488218 235404 488454
rect 234804 488134 235404 488218
rect 234804 487898 234986 488134
rect 235222 487898 235404 488134
rect 234804 452454 235404 487898
rect 234804 452218 234986 452454
rect 235222 452218 235404 452454
rect 234804 452134 235404 452218
rect 234804 451898 234986 452134
rect 235222 451898 235404 452134
rect 234804 416454 235404 451898
rect 234804 416218 234986 416454
rect 235222 416218 235404 416454
rect 234804 416134 235404 416218
rect 234804 415898 234986 416134
rect 235222 415898 235404 416134
rect 231715 399396 231781 399397
rect 231715 399332 231716 399396
rect 231780 399332 231781 399396
rect 231715 399331 231781 399332
rect 233003 399396 233069 399397
rect 233003 399332 233004 399396
rect 233068 399332 233069 399396
rect 233003 399331 233069 399332
rect 227604 373018 227786 373254
rect 228022 373018 228204 373254
rect 227604 372934 228204 373018
rect 227604 372698 227786 372934
rect 228022 372698 228204 372934
rect 227604 337254 228204 372698
rect 227604 337018 227786 337254
rect 228022 337018 228204 337254
rect 227604 336934 228204 337018
rect 227604 336698 227786 336934
rect 228022 336698 228204 336934
rect 227604 301254 228204 336698
rect 227604 301018 227786 301254
rect 228022 301018 228204 301254
rect 227604 300934 228204 301018
rect 227604 300698 227786 300934
rect 228022 300698 228204 300934
rect 227604 265254 228204 300698
rect 227604 265018 227786 265254
rect 228022 265018 228204 265254
rect 227604 264934 228204 265018
rect 227604 264698 227786 264934
rect 228022 264698 228204 264934
rect 227604 229254 228204 264698
rect 227604 229018 227786 229254
rect 228022 229018 228204 229254
rect 227604 228934 228204 229018
rect 227604 228698 227786 228934
rect 228022 228698 228204 228934
rect 227604 193254 228204 228698
rect 227604 193018 227786 193254
rect 228022 193018 228204 193254
rect 227604 192934 228204 193018
rect 227604 192698 227786 192934
rect 228022 192698 228204 192934
rect 227604 157254 228204 192698
rect 227604 157018 227786 157254
rect 228022 157018 228204 157254
rect 227604 156934 228204 157018
rect 227604 156698 227786 156934
rect 228022 156698 228204 156934
rect 227604 121254 228204 156698
rect 227604 121018 227786 121254
rect 228022 121018 228204 121254
rect 227604 120934 228204 121018
rect 227604 120698 227786 120934
rect 228022 120698 228204 120934
rect 227604 85254 228204 120698
rect 227604 85018 227786 85254
rect 228022 85018 228204 85254
rect 227604 84934 228204 85018
rect 227604 84698 227786 84934
rect 228022 84698 228204 84934
rect 227604 49254 228204 84698
rect 227604 49018 227786 49254
rect 228022 49018 228204 49254
rect 227604 48934 228204 49018
rect 227604 48698 227786 48934
rect 228022 48698 228204 48934
rect 227604 13254 228204 48698
rect 231718 29069 231778 399331
rect 233006 76261 233066 399331
rect 234804 380454 235404 415898
rect 238404 672054 239004 707042
rect 238404 671818 238586 672054
rect 238822 671818 239004 672054
rect 238404 671734 239004 671818
rect 238404 671498 238586 671734
rect 238822 671498 239004 671734
rect 238404 636054 239004 671498
rect 238404 635818 238586 636054
rect 238822 635818 239004 636054
rect 238404 635734 239004 635818
rect 238404 635498 238586 635734
rect 238822 635498 239004 635734
rect 238404 600054 239004 635498
rect 238404 599818 238586 600054
rect 238822 599818 239004 600054
rect 238404 599734 239004 599818
rect 238404 599498 238586 599734
rect 238822 599498 239004 599734
rect 238404 564054 239004 599498
rect 238404 563818 238586 564054
rect 238822 563818 239004 564054
rect 238404 563734 239004 563818
rect 238404 563498 238586 563734
rect 238822 563498 239004 563734
rect 238404 528054 239004 563498
rect 238404 527818 238586 528054
rect 238822 527818 239004 528054
rect 238404 527734 239004 527818
rect 238404 527498 238586 527734
rect 238822 527498 239004 527734
rect 238404 492054 239004 527498
rect 238404 491818 238586 492054
rect 238822 491818 239004 492054
rect 238404 491734 239004 491818
rect 238404 491498 238586 491734
rect 238822 491498 239004 491734
rect 238404 456054 239004 491498
rect 238404 455818 238586 456054
rect 238822 455818 239004 456054
rect 238404 455734 239004 455818
rect 238404 455498 238586 455734
rect 238822 455498 239004 455734
rect 238404 420054 239004 455498
rect 238404 419818 238586 420054
rect 238822 419818 239004 420054
rect 238404 419734 239004 419818
rect 238404 419498 238586 419734
rect 238822 419498 239004 419734
rect 237235 399396 237301 399397
rect 237235 399332 237236 399396
rect 237300 399332 237301 399396
rect 237235 399331 237301 399332
rect 238155 399396 238221 399397
rect 238155 399332 238156 399396
rect 238220 399332 238221 399396
rect 238155 399331 238221 399332
rect 234804 380218 234986 380454
rect 235222 380218 235404 380454
rect 234804 380134 235404 380218
rect 234804 379898 234986 380134
rect 235222 379898 235404 380134
rect 234804 344454 235404 379898
rect 234804 344218 234986 344454
rect 235222 344218 235404 344454
rect 234804 344134 235404 344218
rect 234804 343898 234986 344134
rect 235222 343898 235404 344134
rect 234804 308454 235404 343898
rect 234804 308218 234986 308454
rect 235222 308218 235404 308454
rect 234804 308134 235404 308218
rect 234804 307898 234986 308134
rect 235222 307898 235404 308134
rect 234804 272454 235404 307898
rect 234804 272218 234986 272454
rect 235222 272218 235404 272454
rect 234804 272134 235404 272218
rect 234804 271898 234986 272134
rect 235222 271898 235404 272134
rect 234804 236454 235404 271898
rect 234804 236218 234986 236454
rect 235222 236218 235404 236454
rect 234804 236134 235404 236218
rect 234804 235898 234986 236134
rect 235222 235898 235404 236134
rect 234804 200454 235404 235898
rect 237238 227901 237298 399331
rect 238158 398581 238218 399331
rect 238155 398580 238221 398581
rect 238155 398516 238156 398580
rect 238220 398516 238221 398580
rect 238155 398515 238221 398516
rect 238404 384054 239004 419498
rect 238404 383818 238586 384054
rect 238822 383818 239004 384054
rect 238404 383734 239004 383818
rect 238404 383498 238586 383734
rect 238822 383498 239004 383734
rect 238404 348054 239004 383498
rect 238404 347818 238586 348054
rect 238822 347818 239004 348054
rect 238404 347734 239004 347818
rect 238404 347498 238586 347734
rect 238822 347498 239004 347734
rect 238404 312054 239004 347498
rect 238404 311818 238586 312054
rect 238822 311818 239004 312054
rect 238404 311734 239004 311818
rect 238404 311498 238586 311734
rect 238822 311498 239004 311734
rect 238404 276054 239004 311498
rect 238404 275818 238586 276054
rect 238822 275818 239004 276054
rect 238404 275734 239004 275818
rect 238404 275498 238586 275734
rect 238822 275498 239004 275734
rect 238404 240054 239004 275498
rect 238404 239818 238586 240054
rect 238822 239818 239004 240054
rect 238404 239734 239004 239818
rect 238404 239498 238586 239734
rect 238822 239498 239004 239734
rect 237235 227900 237301 227901
rect 237235 227836 237236 227900
rect 237300 227836 237301 227900
rect 237235 227835 237301 227836
rect 234804 200218 234986 200454
rect 235222 200218 235404 200454
rect 234804 200134 235404 200218
rect 234804 199898 234986 200134
rect 235222 199898 235404 200134
rect 234804 164454 235404 199898
rect 234804 164218 234986 164454
rect 235222 164218 235404 164454
rect 234804 164134 235404 164218
rect 234804 163898 234986 164134
rect 235222 163898 235404 164134
rect 234804 128454 235404 163898
rect 234804 128218 234986 128454
rect 235222 128218 235404 128454
rect 234804 128134 235404 128218
rect 234804 127898 234986 128134
rect 235222 127898 235404 128134
rect 234804 92454 235404 127898
rect 234804 92218 234986 92454
rect 235222 92218 235404 92454
rect 234804 92134 235404 92218
rect 234804 91898 234986 92134
rect 235222 91898 235404 92134
rect 233003 76260 233069 76261
rect 233003 76196 233004 76260
rect 233068 76196 233069 76260
rect 233003 76195 233069 76196
rect 234804 56454 235404 91898
rect 234804 56218 234986 56454
rect 235222 56218 235404 56454
rect 234804 56134 235404 56218
rect 234804 55898 234986 56134
rect 235222 55898 235404 56134
rect 231715 29068 231781 29069
rect 231715 29004 231716 29068
rect 231780 29004 231781 29068
rect 231715 29003 231781 29004
rect 227604 13018 227786 13254
rect 228022 13018 228204 13254
rect 227604 12934 228204 13018
rect 227604 12698 227786 12934
rect 228022 12698 228204 12934
rect 209604 -7022 209786 -6786
rect 210022 -7022 210204 -6786
rect 209604 -7106 210204 -7022
rect 209604 -7342 209786 -7106
rect 210022 -7342 210204 -7106
rect 209604 -7364 210204 -7342
rect 227604 -5866 228204 12698
rect 234804 20454 235404 55898
rect 234804 20218 234986 20454
rect 235222 20218 235404 20454
rect 234804 20134 235404 20218
rect 234804 19898 234986 20134
rect 235222 19898 235404 20134
rect 234804 -1266 235404 19898
rect 234804 -1502 234986 -1266
rect 235222 -1502 235404 -1266
rect 234804 -1586 235404 -1502
rect 234804 -1822 234986 -1586
rect 235222 -1822 235404 -1586
rect 234804 -1844 235404 -1822
rect 238404 204054 239004 239498
rect 238404 203818 238586 204054
rect 238822 203818 239004 204054
rect 238404 203734 239004 203818
rect 238404 203498 238586 203734
rect 238822 203498 239004 203734
rect 238404 168054 239004 203498
rect 238404 167818 238586 168054
rect 238822 167818 239004 168054
rect 238404 167734 239004 167818
rect 238404 167498 238586 167734
rect 238822 167498 239004 167734
rect 238404 132054 239004 167498
rect 238404 131818 238586 132054
rect 238822 131818 239004 132054
rect 238404 131734 239004 131818
rect 238404 131498 238586 131734
rect 238822 131498 239004 131734
rect 238404 96054 239004 131498
rect 238404 95818 238586 96054
rect 238822 95818 239004 96054
rect 238404 95734 239004 95818
rect 238404 95498 238586 95734
rect 238822 95498 239004 95734
rect 238404 60054 239004 95498
rect 238404 59818 238586 60054
rect 238822 59818 239004 60054
rect 238404 59734 239004 59818
rect 238404 59498 238586 59734
rect 238822 59498 239004 59734
rect 238404 24054 239004 59498
rect 238404 23818 238586 24054
rect 238822 23818 239004 24054
rect 238404 23734 239004 23818
rect 238404 23498 238586 23734
rect 238822 23498 239004 23734
rect 238404 -3106 239004 23498
rect 238404 -3342 238586 -3106
rect 238822 -3342 239004 -3106
rect 238404 -3426 239004 -3342
rect 238404 -3662 238586 -3426
rect 238822 -3662 239004 -3426
rect 238404 -3684 239004 -3662
rect 242004 675654 242604 708882
rect 242004 675418 242186 675654
rect 242422 675418 242604 675654
rect 242004 675334 242604 675418
rect 242004 675098 242186 675334
rect 242422 675098 242604 675334
rect 242004 639654 242604 675098
rect 242004 639418 242186 639654
rect 242422 639418 242604 639654
rect 242004 639334 242604 639418
rect 242004 639098 242186 639334
rect 242422 639098 242604 639334
rect 242004 603654 242604 639098
rect 242004 603418 242186 603654
rect 242422 603418 242604 603654
rect 242004 603334 242604 603418
rect 242004 603098 242186 603334
rect 242422 603098 242604 603334
rect 242004 567654 242604 603098
rect 242004 567418 242186 567654
rect 242422 567418 242604 567654
rect 242004 567334 242604 567418
rect 242004 567098 242186 567334
rect 242422 567098 242604 567334
rect 242004 531654 242604 567098
rect 242004 531418 242186 531654
rect 242422 531418 242604 531654
rect 242004 531334 242604 531418
rect 242004 531098 242186 531334
rect 242422 531098 242604 531334
rect 242004 495654 242604 531098
rect 242004 495418 242186 495654
rect 242422 495418 242604 495654
rect 242004 495334 242604 495418
rect 242004 495098 242186 495334
rect 242422 495098 242604 495334
rect 242004 459654 242604 495098
rect 242004 459418 242186 459654
rect 242422 459418 242604 459654
rect 242004 459334 242604 459418
rect 242004 459098 242186 459334
rect 242422 459098 242604 459334
rect 242004 423654 242604 459098
rect 242004 423418 242186 423654
rect 242422 423418 242604 423654
rect 242004 423334 242604 423418
rect 242004 423098 242186 423334
rect 242422 423098 242604 423334
rect 242004 387654 242604 423098
rect 245604 679254 246204 710722
rect 263604 710358 264204 711300
rect 263604 710122 263786 710358
rect 264022 710122 264204 710358
rect 263604 710038 264204 710122
rect 263604 709802 263786 710038
rect 264022 709802 264204 710038
rect 260004 708518 260604 709460
rect 260004 708282 260186 708518
rect 260422 708282 260604 708518
rect 260004 708198 260604 708282
rect 260004 707962 260186 708198
rect 260422 707962 260604 708198
rect 256404 706678 257004 707620
rect 256404 706442 256586 706678
rect 256822 706442 257004 706678
rect 256404 706358 257004 706442
rect 256404 706122 256586 706358
rect 256822 706122 257004 706358
rect 245604 679018 245786 679254
rect 246022 679018 246204 679254
rect 245604 678934 246204 679018
rect 245604 678698 245786 678934
rect 246022 678698 246204 678934
rect 245604 643254 246204 678698
rect 245604 643018 245786 643254
rect 246022 643018 246204 643254
rect 245604 642934 246204 643018
rect 245604 642698 245786 642934
rect 246022 642698 246204 642934
rect 245604 607254 246204 642698
rect 245604 607018 245786 607254
rect 246022 607018 246204 607254
rect 245604 606934 246204 607018
rect 245604 606698 245786 606934
rect 246022 606698 246204 606934
rect 245604 571254 246204 606698
rect 245604 571018 245786 571254
rect 246022 571018 246204 571254
rect 245604 570934 246204 571018
rect 245604 570698 245786 570934
rect 246022 570698 246204 570934
rect 245604 535254 246204 570698
rect 245604 535018 245786 535254
rect 246022 535018 246204 535254
rect 245604 534934 246204 535018
rect 245604 534698 245786 534934
rect 246022 534698 246204 534934
rect 245604 499254 246204 534698
rect 245604 499018 245786 499254
rect 246022 499018 246204 499254
rect 245604 498934 246204 499018
rect 245604 498698 245786 498934
rect 246022 498698 246204 498934
rect 245604 463254 246204 498698
rect 245604 463018 245786 463254
rect 246022 463018 246204 463254
rect 245604 462934 246204 463018
rect 245604 462698 245786 462934
rect 246022 462698 246204 462934
rect 245604 427254 246204 462698
rect 245604 427018 245786 427254
rect 246022 427018 246204 427254
rect 245604 426934 246204 427018
rect 245604 426698 245786 426934
rect 246022 426698 246204 426934
rect 242755 399396 242821 399397
rect 242755 399332 242756 399396
rect 242820 399332 242821 399396
rect 242755 399331 242821 399332
rect 242758 398445 242818 399331
rect 242755 398444 242821 398445
rect 242755 398380 242756 398444
rect 242820 398380 242821 398444
rect 242755 398379 242821 398380
rect 242004 387418 242186 387654
rect 242422 387418 242604 387654
rect 242004 387334 242604 387418
rect 242004 387098 242186 387334
rect 242422 387098 242604 387334
rect 242004 351654 242604 387098
rect 242004 351418 242186 351654
rect 242422 351418 242604 351654
rect 242004 351334 242604 351418
rect 242004 351098 242186 351334
rect 242422 351098 242604 351334
rect 242004 315654 242604 351098
rect 242004 315418 242186 315654
rect 242422 315418 242604 315654
rect 242004 315334 242604 315418
rect 242004 315098 242186 315334
rect 242422 315098 242604 315334
rect 242004 279654 242604 315098
rect 242004 279418 242186 279654
rect 242422 279418 242604 279654
rect 242004 279334 242604 279418
rect 242004 279098 242186 279334
rect 242422 279098 242604 279334
rect 242004 243654 242604 279098
rect 242004 243418 242186 243654
rect 242422 243418 242604 243654
rect 242004 243334 242604 243418
rect 242004 243098 242186 243334
rect 242422 243098 242604 243334
rect 242004 207654 242604 243098
rect 242004 207418 242186 207654
rect 242422 207418 242604 207654
rect 242004 207334 242604 207418
rect 242004 207098 242186 207334
rect 242422 207098 242604 207334
rect 242004 171654 242604 207098
rect 242004 171418 242186 171654
rect 242422 171418 242604 171654
rect 242004 171334 242604 171418
rect 242004 171098 242186 171334
rect 242422 171098 242604 171334
rect 242004 135654 242604 171098
rect 242004 135418 242186 135654
rect 242422 135418 242604 135654
rect 242004 135334 242604 135418
rect 242004 135098 242186 135334
rect 242422 135098 242604 135334
rect 242004 99654 242604 135098
rect 242004 99418 242186 99654
rect 242422 99418 242604 99654
rect 242004 99334 242604 99418
rect 242004 99098 242186 99334
rect 242422 99098 242604 99334
rect 242004 63654 242604 99098
rect 242004 63418 242186 63654
rect 242422 63418 242604 63654
rect 242004 63334 242604 63418
rect 242004 63098 242186 63334
rect 242422 63098 242604 63334
rect 242004 27654 242604 63098
rect 242004 27418 242186 27654
rect 242422 27418 242604 27654
rect 242004 27334 242604 27418
rect 242004 27098 242186 27334
rect 242422 27098 242604 27334
rect 242004 -4946 242604 27098
rect 242004 -5182 242186 -4946
rect 242422 -5182 242604 -4946
rect 242004 -5266 242604 -5182
rect 242004 -5502 242186 -5266
rect 242422 -5502 242604 -5266
rect 242004 -5524 242604 -5502
rect 245604 391254 246204 426698
rect 245604 391018 245786 391254
rect 246022 391018 246204 391254
rect 245604 390934 246204 391018
rect 245604 390698 245786 390934
rect 246022 390698 246204 390934
rect 245604 355254 246204 390698
rect 245604 355018 245786 355254
rect 246022 355018 246204 355254
rect 245604 354934 246204 355018
rect 245604 354698 245786 354934
rect 246022 354698 246204 354934
rect 245604 319254 246204 354698
rect 245604 319018 245786 319254
rect 246022 319018 246204 319254
rect 245604 318934 246204 319018
rect 245604 318698 245786 318934
rect 246022 318698 246204 318934
rect 245604 283254 246204 318698
rect 245604 283018 245786 283254
rect 246022 283018 246204 283254
rect 245604 282934 246204 283018
rect 245604 282698 245786 282934
rect 246022 282698 246204 282934
rect 245604 247254 246204 282698
rect 245604 247018 245786 247254
rect 246022 247018 246204 247254
rect 245604 246934 246204 247018
rect 245604 246698 245786 246934
rect 246022 246698 246204 246934
rect 245604 211254 246204 246698
rect 245604 211018 245786 211254
rect 246022 211018 246204 211254
rect 245604 210934 246204 211018
rect 245604 210698 245786 210934
rect 246022 210698 246204 210934
rect 245604 175254 246204 210698
rect 245604 175018 245786 175254
rect 246022 175018 246204 175254
rect 245604 174934 246204 175018
rect 245604 174698 245786 174934
rect 246022 174698 246204 174934
rect 245604 139254 246204 174698
rect 245604 139018 245786 139254
rect 246022 139018 246204 139254
rect 245604 138934 246204 139018
rect 245604 138698 245786 138934
rect 246022 138698 246204 138934
rect 245604 103254 246204 138698
rect 245604 103018 245786 103254
rect 246022 103018 246204 103254
rect 245604 102934 246204 103018
rect 245604 102698 245786 102934
rect 246022 102698 246204 102934
rect 245604 67254 246204 102698
rect 245604 67018 245786 67254
rect 246022 67018 246204 67254
rect 245604 66934 246204 67018
rect 245604 66698 245786 66934
rect 246022 66698 246204 66934
rect 245604 31254 246204 66698
rect 245604 31018 245786 31254
rect 246022 31018 246204 31254
rect 245604 30934 246204 31018
rect 245604 30698 245786 30934
rect 246022 30698 246204 30934
rect 227604 -6102 227786 -5866
rect 228022 -6102 228204 -5866
rect 227604 -6186 228204 -6102
rect 227604 -6422 227786 -6186
rect 228022 -6422 228204 -6186
rect 227604 -7364 228204 -6422
rect 245604 -6786 246204 30698
rect 252804 704838 253404 705780
rect 252804 704602 252986 704838
rect 253222 704602 253404 704838
rect 252804 704518 253404 704602
rect 252804 704282 252986 704518
rect 253222 704282 253404 704518
rect 252804 686454 253404 704282
rect 252804 686218 252986 686454
rect 253222 686218 253404 686454
rect 252804 686134 253404 686218
rect 252804 685898 252986 686134
rect 253222 685898 253404 686134
rect 252804 650454 253404 685898
rect 252804 650218 252986 650454
rect 253222 650218 253404 650454
rect 252804 650134 253404 650218
rect 252804 649898 252986 650134
rect 253222 649898 253404 650134
rect 252804 614454 253404 649898
rect 252804 614218 252986 614454
rect 253222 614218 253404 614454
rect 252804 614134 253404 614218
rect 252804 613898 252986 614134
rect 253222 613898 253404 614134
rect 252804 578454 253404 613898
rect 252804 578218 252986 578454
rect 253222 578218 253404 578454
rect 252804 578134 253404 578218
rect 252804 577898 252986 578134
rect 253222 577898 253404 578134
rect 252804 542454 253404 577898
rect 252804 542218 252986 542454
rect 253222 542218 253404 542454
rect 252804 542134 253404 542218
rect 252804 541898 252986 542134
rect 253222 541898 253404 542134
rect 252804 506454 253404 541898
rect 252804 506218 252986 506454
rect 253222 506218 253404 506454
rect 252804 506134 253404 506218
rect 252804 505898 252986 506134
rect 253222 505898 253404 506134
rect 252804 470454 253404 505898
rect 252804 470218 252986 470454
rect 253222 470218 253404 470454
rect 252804 470134 253404 470218
rect 252804 469898 252986 470134
rect 253222 469898 253404 470134
rect 252804 434454 253404 469898
rect 252804 434218 252986 434454
rect 253222 434218 253404 434454
rect 252804 434134 253404 434218
rect 252804 433898 252986 434134
rect 253222 433898 253404 434134
rect 252804 398454 253404 433898
rect 252804 398218 252986 398454
rect 253222 398218 253404 398454
rect 252804 398134 253404 398218
rect 252804 397898 252986 398134
rect 253222 397898 253404 398134
rect 252804 362454 253404 397898
rect 252804 362218 252986 362454
rect 253222 362218 253404 362454
rect 252804 362134 253404 362218
rect 252804 361898 252986 362134
rect 253222 361898 253404 362134
rect 252804 326454 253404 361898
rect 252804 326218 252986 326454
rect 253222 326218 253404 326454
rect 252804 326134 253404 326218
rect 252804 325898 252986 326134
rect 253222 325898 253404 326134
rect 252804 290454 253404 325898
rect 256404 690054 257004 706122
rect 256404 689818 256586 690054
rect 256822 689818 257004 690054
rect 256404 689734 257004 689818
rect 256404 689498 256586 689734
rect 256822 689498 257004 689734
rect 256404 654054 257004 689498
rect 256404 653818 256586 654054
rect 256822 653818 257004 654054
rect 256404 653734 257004 653818
rect 256404 653498 256586 653734
rect 256822 653498 257004 653734
rect 256404 618054 257004 653498
rect 256404 617818 256586 618054
rect 256822 617818 257004 618054
rect 256404 617734 257004 617818
rect 256404 617498 256586 617734
rect 256822 617498 257004 617734
rect 256404 582054 257004 617498
rect 256404 581818 256586 582054
rect 256822 581818 257004 582054
rect 256404 581734 257004 581818
rect 256404 581498 256586 581734
rect 256822 581498 257004 581734
rect 256404 546054 257004 581498
rect 256404 545818 256586 546054
rect 256822 545818 257004 546054
rect 256404 545734 257004 545818
rect 256404 545498 256586 545734
rect 256822 545498 257004 545734
rect 256404 510054 257004 545498
rect 256404 509818 256586 510054
rect 256822 509818 257004 510054
rect 256404 509734 257004 509818
rect 256404 509498 256586 509734
rect 256822 509498 257004 509734
rect 256404 474054 257004 509498
rect 256404 473818 256586 474054
rect 256822 473818 257004 474054
rect 256404 473734 257004 473818
rect 256404 473498 256586 473734
rect 256822 473498 257004 473734
rect 256404 438054 257004 473498
rect 256404 437818 256586 438054
rect 256822 437818 257004 438054
rect 256404 437734 257004 437818
rect 256404 437498 256586 437734
rect 256822 437498 257004 437734
rect 256404 402054 257004 437498
rect 256404 401818 256586 402054
rect 256822 401818 257004 402054
rect 256404 401734 257004 401818
rect 256404 401498 256586 401734
rect 256822 401498 257004 401734
rect 256404 366054 257004 401498
rect 256404 365818 256586 366054
rect 256822 365818 257004 366054
rect 256404 365734 257004 365818
rect 256404 365498 256586 365734
rect 256822 365498 257004 365734
rect 256404 330054 257004 365498
rect 256404 329818 256586 330054
rect 256822 329818 257004 330054
rect 256404 329734 257004 329818
rect 256404 329498 256586 329734
rect 256822 329498 257004 329734
rect 254715 314668 254781 314669
rect 254715 314604 254716 314668
rect 254780 314604 254781 314668
rect 254715 314603 254781 314604
rect 254718 305013 254778 314603
rect 254715 305012 254781 305013
rect 254715 304948 254716 305012
rect 254780 304948 254781 305012
rect 254715 304947 254781 304948
rect 252804 290218 252986 290454
rect 253222 290218 253404 290454
rect 252804 290134 253404 290218
rect 252804 289898 252986 290134
rect 253222 289898 253404 290134
rect 252804 254454 253404 289898
rect 256404 294054 257004 329498
rect 256404 293818 256586 294054
rect 256822 293818 257004 294054
rect 256404 293734 257004 293818
rect 256404 293498 256586 293734
rect 256822 293498 257004 293734
rect 255635 289100 255701 289101
rect 255635 289036 255636 289100
rect 255700 289036 255701 289100
rect 255635 289035 255701 289036
rect 255638 276045 255698 289035
rect 255635 276044 255701 276045
rect 255635 275980 255636 276044
rect 255700 275980 255701 276044
rect 255635 275979 255701 275980
rect 252804 254218 252986 254454
rect 253222 254218 253404 254454
rect 252804 254134 253404 254218
rect 252804 253898 252986 254134
rect 253222 253898 253404 254134
rect 252804 218454 253404 253898
rect 252804 218218 252986 218454
rect 253222 218218 253404 218454
rect 252804 218134 253404 218218
rect 252804 217898 252986 218134
rect 253222 217898 253404 218134
rect 252804 182454 253404 217898
rect 252804 182218 252986 182454
rect 253222 182218 253404 182454
rect 252804 182134 253404 182218
rect 252804 181898 252986 182134
rect 253222 181898 253404 182134
rect 252804 146454 253404 181898
rect 252804 146218 252986 146454
rect 253222 146218 253404 146454
rect 252804 146134 253404 146218
rect 252804 145898 252986 146134
rect 253222 145898 253404 146134
rect 252804 110454 253404 145898
rect 252804 110218 252986 110454
rect 253222 110218 253404 110454
rect 252804 110134 253404 110218
rect 252804 109898 252986 110134
rect 253222 109898 253404 110134
rect 252804 74454 253404 109898
rect 252804 74218 252986 74454
rect 253222 74218 253404 74454
rect 252804 74134 253404 74218
rect 252804 73898 252986 74134
rect 253222 73898 253404 74134
rect 252804 38454 253404 73898
rect 252804 38218 252986 38454
rect 253222 38218 253404 38454
rect 252804 38134 253404 38218
rect 252804 37898 252986 38134
rect 253222 37898 253404 38134
rect 252804 2454 253404 37898
rect 252804 2218 252986 2454
rect 253222 2218 253404 2454
rect 252804 2134 253404 2218
rect 252804 1898 252986 2134
rect 253222 1898 253404 2134
rect 252804 -346 253404 1898
rect 252804 -582 252986 -346
rect 253222 -582 253404 -346
rect 252804 -666 253404 -582
rect 252804 -902 252986 -666
rect 253222 -902 253404 -666
rect 252804 -1844 253404 -902
rect 256404 258054 257004 293498
rect 256404 257818 256586 258054
rect 256822 257818 257004 258054
rect 256404 257734 257004 257818
rect 256404 257498 256586 257734
rect 256822 257498 257004 257734
rect 256404 222054 257004 257498
rect 256404 221818 256586 222054
rect 256822 221818 257004 222054
rect 256404 221734 257004 221818
rect 256404 221498 256586 221734
rect 256822 221498 257004 221734
rect 256404 186054 257004 221498
rect 256404 185818 256586 186054
rect 256822 185818 257004 186054
rect 256404 185734 257004 185818
rect 256404 185498 256586 185734
rect 256822 185498 257004 185734
rect 256404 150054 257004 185498
rect 256404 149818 256586 150054
rect 256822 149818 257004 150054
rect 256404 149734 257004 149818
rect 256404 149498 256586 149734
rect 256822 149498 257004 149734
rect 256404 114054 257004 149498
rect 256404 113818 256586 114054
rect 256822 113818 257004 114054
rect 256404 113734 257004 113818
rect 256404 113498 256586 113734
rect 256822 113498 257004 113734
rect 256404 78054 257004 113498
rect 256404 77818 256586 78054
rect 256822 77818 257004 78054
rect 256404 77734 257004 77818
rect 256404 77498 256586 77734
rect 256822 77498 257004 77734
rect 256404 42054 257004 77498
rect 256404 41818 256586 42054
rect 256822 41818 257004 42054
rect 256404 41734 257004 41818
rect 256404 41498 256586 41734
rect 256822 41498 257004 41734
rect 256404 6054 257004 41498
rect 256404 5818 256586 6054
rect 256822 5818 257004 6054
rect 256404 5734 257004 5818
rect 256404 5498 256586 5734
rect 256822 5498 257004 5734
rect 256404 -2186 257004 5498
rect 256404 -2422 256586 -2186
rect 256822 -2422 257004 -2186
rect 256404 -2506 257004 -2422
rect 256404 -2742 256586 -2506
rect 256822 -2742 257004 -2506
rect 256404 -3684 257004 -2742
rect 260004 693654 260604 707962
rect 260004 693418 260186 693654
rect 260422 693418 260604 693654
rect 260004 693334 260604 693418
rect 260004 693098 260186 693334
rect 260422 693098 260604 693334
rect 260004 657654 260604 693098
rect 260004 657418 260186 657654
rect 260422 657418 260604 657654
rect 260004 657334 260604 657418
rect 260004 657098 260186 657334
rect 260422 657098 260604 657334
rect 260004 621654 260604 657098
rect 260004 621418 260186 621654
rect 260422 621418 260604 621654
rect 260004 621334 260604 621418
rect 260004 621098 260186 621334
rect 260422 621098 260604 621334
rect 260004 585654 260604 621098
rect 260004 585418 260186 585654
rect 260422 585418 260604 585654
rect 260004 585334 260604 585418
rect 260004 585098 260186 585334
rect 260422 585098 260604 585334
rect 260004 549654 260604 585098
rect 260004 549418 260186 549654
rect 260422 549418 260604 549654
rect 260004 549334 260604 549418
rect 260004 549098 260186 549334
rect 260422 549098 260604 549334
rect 260004 513654 260604 549098
rect 260004 513418 260186 513654
rect 260422 513418 260604 513654
rect 260004 513334 260604 513418
rect 260004 513098 260186 513334
rect 260422 513098 260604 513334
rect 260004 477654 260604 513098
rect 260004 477418 260186 477654
rect 260422 477418 260604 477654
rect 260004 477334 260604 477418
rect 260004 477098 260186 477334
rect 260422 477098 260604 477334
rect 260004 441654 260604 477098
rect 260004 441418 260186 441654
rect 260422 441418 260604 441654
rect 260004 441334 260604 441418
rect 260004 441098 260186 441334
rect 260422 441098 260604 441334
rect 260004 405654 260604 441098
rect 260004 405418 260186 405654
rect 260422 405418 260604 405654
rect 260004 405334 260604 405418
rect 260004 405098 260186 405334
rect 260422 405098 260604 405334
rect 260004 369654 260604 405098
rect 260004 369418 260186 369654
rect 260422 369418 260604 369654
rect 260004 369334 260604 369418
rect 260004 369098 260186 369334
rect 260422 369098 260604 369334
rect 260004 333654 260604 369098
rect 260004 333418 260186 333654
rect 260422 333418 260604 333654
rect 260004 333334 260604 333418
rect 260004 333098 260186 333334
rect 260422 333098 260604 333334
rect 260004 297654 260604 333098
rect 260004 297418 260186 297654
rect 260422 297418 260604 297654
rect 260004 297334 260604 297418
rect 260004 297098 260186 297334
rect 260422 297098 260604 297334
rect 260004 261654 260604 297098
rect 260004 261418 260186 261654
rect 260422 261418 260604 261654
rect 260004 261334 260604 261418
rect 260004 261098 260186 261334
rect 260422 261098 260604 261334
rect 260004 225654 260604 261098
rect 260004 225418 260186 225654
rect 260422 225418 260604 225654
rect 260004 225334 260604 225418
rect 260004 225098 260186 225334
rect 260422 225098 260604 225334
rect 260004 189654 260604 225098
rect 260004 189418 260186 189654
rect 260422 189418 260604 189654
rect 260004 189334 260604 189418
rect 260004 189098 260186 189334
rect 260422 189098 260604 189334
rect 260004 153654 260604 189098
rect 260004 153418 260186 153654
rect 260422 153418 260604 153654
rect 260004 153334 260604 153418
rect 260004 153098 260186 153334
rect 260422 153098 260604 153334
rect 260004 117654 260604 153098
rect 260004 117418 260186 117654
rect 260422 117418 260604 117654
rect 260004 117334 260604 117418
rect 260004 117098 260186 117334
rect 260422 117098 260604 117334
rect 260004 81654 260604 117098
rect 260004 81418 260186 81654
rect 260422 81418 260604 81654
rect 260004 81334 260604 81418
rect 260004 81098 260186 81334
rect 260422 81098 260604 81334
rect 260004 45654 260604 81098
rect 260004 45418 260186 45654
rect 260422 45418 260604 45654
rect 260004 45334 260604 45418
rect 260004 45098 260186 45334
rect 260422 45098 260604 45334
rect 260004 9654 260604 45098
rect 260004 9418 260186 9654
rect 260422 9418 260604 9654
rect 260004 9334 260604 9418
rect 260004 9098 260186 9334
rect 260422 9098 260604 9334
rect 260004 -4026 260604 9098
rect 260004 -4262 260186 -4026
rect 260422 -4262 260604 -4026
rect 260004 -4346 260604 -4262
rect 260004 -4582 260186 -4346
rect 260422 -4582 260604 -4346
rect 260004 -5524 260604 -4582
rect 263604 697254 264204 709802
rect 281604 711278 282204 711300
rect 281604 711042 281786 711278
rect 282022 711042 282204 711278
rect 281604 710958 282204 711042
rect 281604 710722 281786 710958
rect 282022 710722 282204 710958
rect 278004 709438 278604 709460
rect 278004 709202 278186 709438
rect 278422 709202 278604 709438
rect 278004 709118 278604 709202
rect 278004 708882 278186 709118
rect 278422 708882 278604 709118
rect 274404 707598 275004 707620
rect 274404 707362 274586 707598
rect 274822 707362 275004 707598
rect 274404 707278 275004 707362
rect 274404 707042 274586 707278
rect 274822 707042 275004 707278
rect 263604 697018 263786 697254
rect 264022 697018 264204 697254
rect 263604 696934 264204 697018
rect 263604 696698 263786 696934
rect 264022 696698 264204 696934
rect 263604 661254 264204 696698
rect 263604 661018 263786 661254
rect 264022 661018 264204 661254
rect 263604 660934 264204 661018
rect 263604 660698 263786 660934
rect 264022 660698 264204 660934
rect 263604 625254 264204 660698
rect 263604 625018 263786 625254
rect 264022 625018 264204 625254
rect 263604 624934 264204 625018
rect 263604 624698 263786 624934
rect 264022 624698 264204 624934
rect 263604 589254 264204 624698
rect 263604 589018 263786 589254
rect 264022 589018 264204 589254
rect 263604 588934 264204 589018
rect 263604 588698 263786 588934
rect 264022 588698 264204 588934
rect 263604 553254 264204 588698
rect 263604 553018 263786 553254
rect 264022 553018 264204 553254
rect 263604 552934 264204 553018
rect 263604 552698 263786 552934
rect 264022 552698 264204 552934
rect 263604 517254 264204 552698
rect 263604 517018 263786 517254
rect 264022 517018 264204 517254
rect 263604 516934 264204 517018
rect 263604 516698 263786 516934
rect 264022 516698 264204 516934
rect 263604 481254 264204 516698
rect 263604 481018 263786 481254
rect 264022 481018 264204 481254
rect 263604 480934 264204 481018
rect 263604 480698 263786 480934
rect 264022 480698 264204 480934
rect 263604 445254 264204 480698
rect 263604 445018 263786 445254
rect 264022 445018 264204 445254
rect 263604 444934 264204 445018
rect 263604 444698 263786 444934
rect 264022 444698 264204 444934
rect 263604 409254 264204 444698
rect 263604 409018 263786 409254
rect 264022 409018 264204 409254
rect 263604 408934 264204 409018
rect 263604 408698 263786 408934
rect 264022 408698 264204 408934
rect 263604 373254 264204 408698
rect 263604 373018 263786 373254
rect 264022 373018 264204 373254
rect 263604 372934 264204 373018
rect 263604 372698 263786 372934
rect 264022 372698 264204 372934
rect 263604 337254 264204 372698
rect 263604 337018 263786 337254
rect 264022 337018 264204 337254
rect 263604 336934 264204 337018
rect 263604 336698 263786 336934
rect 264022 336698 264204 336934
rect 263604 301254 264204 336698
rect 263604 301018 263786 301254
rect 264022 301018 264204 301254
rect 263604 300934 264204 301018
rect 263604 300698 263786 300934
rect 264022 300698 264204 300934
rect 263604 265254 264204 300698
rect 263604 265018 263786 265254
rect 264022 265018 264204 265254
rect 263604 264934 264204 265018
rect 263604 264698 263786 264934
rect 264022 264698 264204 264934
rect 263604 229254 264204 264698
rect 263604 229018 263786 229254
rect 264022 229018 264204 229254
rect 263604 228934 264204 229018
rect 263604 228698 263786 228934
rect 264022 228698 264204 228934
rect 263604 193254 264204 228698
rect 263604 193018 263786 193254
rect 264022 193018 264204 193254
rect 263604 192934 264204 193018
rect 263604 192698 263786 192934
rect 264022 192698 264204 192934
rect 263604 157254 264204 192698
rect 263604 157018 263786 157254
rect 264022 157018 264204 157254
rect 263604 156934 264204 157018
rect 263604 156698 263786 156934
rect 264022 156698 264204 156934
rect 263604 121254 264204 156698
rect 263604 121018 263786 121254
rect 264022 121018 264204 121254
rect 263604 120934 264204 121018
rect 263604 120698 263786 120934
rect 264022 120698 264204 120934
rect 263604 85254 264204 120698
rect 263604 85018 263786 85254
rect 264022 85018 264204 85254
rect 263604 84934 264204 85018
rect 263604 84698 263786 84934
rect 264022 84698 264204 84934
rect 263604 49254 264204 84698
rect 263604 49018 263786 49254
rect 264022 49018 264204 49254
rect 263604 48934 264204 49018
rect 263604 48698 263786 48934
rect 264022 48698 264204 48934
rect 263604 13254 264204 48698
rect 263604 13018 263786 13254
rect 264022 13018 264204 13254
rect 263604 12934 264204 13018
rect 263604 12698 263786 12934
rect 264022 12698 264204 12934
rect 245604 -7022 245786 -6786
rect 246022 -7022 246204 -6786
rect 245604 -7106 246204 -7022
rect 245604 -7342 245786 -7106
rect 246022 -7342 246204 -7106
rect 245604 -7364 246204 -7342
rect 263604 -5866 264204 12698
rect 270804 705758 271404 705780
rect 270804 705522 270986 705758
rect 271222 705522 271404 705758
rect 270804 705438 271404 705522
rect 270804 705202 270986 705438
rect 271222 705202 271404 705438
rect 270804 668454 271404 705202
rect 270804 668218 270986 668454
rect 271222 668218 271404 668454
rect 270804 668134 271404 668218
rect 270804 667898 270986 668134
rect 271222 667898 271404 668134
rect 270804 632454 271404 667898
rect 270804 632218 270986 632454
rect 271222 632218 271404 632454
rect 270804 632134 271404 632218
rect 270804 631898 270986 632134
rect 271222 631898 271404 632134
rect 270804 596454 271404 631898
rect 270804 596218 270986 596454
rect 271222 596218 271404 596454
rect 270804 596134 271404 596218
rect 270804 595898 270986 596134
rect 271222 595898 271404 596134
rect 270804 560454 271404 595898
rect 270804 560218 270986 560454
rect 271222 560218 271404 560454
rect 270804 560134 271404 560218
rect 270804 559898 270986 560134
rect 271222 559898 271404 560134
rect 270804 524454 271404 559898
rect 270804 524218 270986 524454
rect 271222 524218 271404 524454
rect 270804 524134 271404 524218
rect 270804 523898 270986 524134
rect 271222 523898 271404 524134
rect 270804 488454 271404 523898
rect 270804 488218 270986 488454
rect 271222 488218 271404 488454
rect 270804 488134 271404 488218
rect 270804 487898 270986 488134
rect 271222 487898 271404 488134
rect 270804 452454 271404 487898
rect 270804 452218 270986 452454
rect 271222 452218 271404 452454
rect 270804 452134 271404 452218
rect 270804 451898 270986 452134
rect 271222 451898 271404 452134
rect 270804 416454 271404 451898
rect 270804 416218 270986 416454
rect 271222 416218 271404 416454
rect 270804 416134 271404 416218
rect 270804 415898 270986 416134
rect 271222 415898 271404 416134
rect 270804 380454 271404 415898
rect 270804 380218 270986 380454
rect 271222 380218 271404 380454
rect 270804 380134 271404 380218
rect 270804 379898 270986 380134
rect 271222 379898 271404 380134
rect 270804 344454 271404 379898
rect 270804 344218 270986 344454
rect 271222 344218 271404 344454
rect 270804 344134 271404 344218
rect 270804 343898 270986 344134
rect 271222 343898 271404 344134
rect 270804 308454 271404 343898
rect 270804 308218 270986 308454
rect 271222 308218 271404 308454
rect 270804 308134 271404 308218
rect 270804 307898 270986 308134
rect 271222 307898 271404 308134
rect 270804 272454 271404 307898
rect 270804 272218 270986 272454
rect 271222 272218 271404 272454
rect 270804 272134 271404 272218
rect 270804 271898 270986 272134
rect 271222 271898 271404 272134
rect 270804 236454 271404 271898
rect 270804 236218 270986 236454
rect 271222 236218 271404 236454
rect 270804 236134 271404 236218
rect 270804 235898 270986 236134
rect 271222 235898 271404 236134
rect 270804 200454 271404 235898
rect 270804 200218 270986 200454
rect 271222 200218 271404 200454
rect 270804 200134 271404 200218
rect 270804 199898 270986 200134
rect 271222 199898 271404 200134
rect 270804 164454 271404 199898
rect 270804 164218 270986 164454
rect 271222 164218 271404 164454
rect 270804 164134 271404 164218
rect 270804 163898 270986 164134
rect 271222 163898 271404 164134
rect 270804 128454 271404 163898
rect 270804 128218 270986 128454
rect 271222 128218 271404 128454
rect 270804 128134 271404 128218
rect 270804 127898 270986 128134
rect 271222 127898 271404 128134
rect 270804 92454 271404 127898
rect 270804 92218 270986 92454
rect 271222 92218 271404 92454
rect 270804 92134 271404 92218
rect 270804 91898 270986 92134
rect 271222 91898 271404 92134
rect 270804 56454 271404 91898
rect 270804 56218 270986 56454
rect 271222 56218 271404 56454
rect 270804 56134 271404 56218
rect 270804 55898 270986 56134
rect 271222 55898 271404 56134
rect 270804 20454 271404 55898
rect 270804 20218 270986 20454
rect 271222 20218 271404 20454
rect 270804 20134 271404 20218
rect 270804 19898 270986 20134
rect 271222 19898 271404 20134
rect 270804 -1266 271404 19898
rect 270804 -1502 270986 -1266
rect 271222 -1502 271404 -1266
rect 270804 -1586 271404 -1502
rect 270804 -1822 270986 -1586
rect 271222 -1822 271404 -1586
rect 270804 -1844 271404 -1822
rect 274404 672054 275004 707042
rect 274404 671818 274586 672054
rect 274822 671818 275004 672054
rect 274404 671734 275004 671818
rect 274404 671498 274586 671734
rect 274822 671498 275004 671734
rect 274404 636054 275004 671498
rect 274404 635818 274586 636054
rect 274822 635818 275004 636054
rect 274404 635734 275004 635818
rect 274404 635498 274586 635734
rect 274822 635498 275004 635734
rect 274404 600054 275004 635498
rect 274404 599818 274586 600054
rect 274822 599818 275004 600054
rect 274404 599734 275004 599818
rect 274404 599498 274586 599734
rect 274822 599498 275004 599734
rect 274404 564054 275004 599498
rect 274404 563818 274586 564054
rect 274822 563818 275004 564054
rect 274404 563734 275004 563818
rect 274404 563498 274586 563734
rect 274822 563498 275004 563734
rect 274404 528054 275004 563498
rect 274404 527818 274586 528054
rect 274822 527818 275004 528054
rect 274404 527734 275004 527818
rect 274404 527498 274586 527734
rect 274822 527498 275004 527734
rect 274404 492054 275004 527498
rect 274404 491818 274586 492054
rect 274822 491818 275004 492054
rect 274404 491734 275004 491818
rect 274404 491498 274586 491734
rect 274822 491498 275004 491734
rect 274404 456054 275004 491498
rect 274404 455818 274586 456054
rect 274822 455818 275004 456054
rect 274404 455734 275004 455818
rect 274404 455498 274586 455734
rect 274822 455498 275004 455734
rect 274404 420054 275004 455498
rect 274404 419818 274586 420054
rect 274822 419818 275004 420054
rect 274404 419734 275004 419818
rect 274404 419498 274586 419734
rect 274822 419498 275004 419734
rect 274404 384054 275004 419498
rect 278004 675654 278604 708882
rect 278004 675418 278186 675654
rect 278422 675418 278604 675654
rect 278004 675334 278604 675418
rect 278004 675098 278186 675334
rect 278422 675098 278604 675334
rect 278004 639654 278604 675098
rect 278004 639418 278186 639654
rect 278422 639418 278604 639654
rect 278004 639334 278604 639418
rect 278004 639098 278186 639334
rect 278422 639098 278604 639334
rect 278004 603654 278604 639098
rect 278004 603418 278186 603654
rect 278422 603418 278604 603654
rect 278004 603334 278604 603418
rect 278004 603098 278186 603334
rect 278422 603098 278604 603334
rect 278004 567654 278604 603098
rect 278004 567418 278186 567654
rect 278422 567418 278604 567654
rect 278004 567334 278604 567418
rect 278004 567098 278186 567334
rect 278422 567098 278604 567334
rect 278004 531654 278604 567098
rect 278004 531418 278186 531654
rect 278422 531418 278604 531654
rect 278004 531334 278604 531418
rect 278004 531098 278186 531334
rect 278422 531098 278604 531334
rect 278004 495654 278604 531098
rect 278004 495418 278186 495654
rect 278422 495418 278604 495654
rect 278004 495334 278604 495418
rect 278004 495098 278186 495334
rect 278422 495098 278604 495334
rect 278004 459654 278604 495098
rect 278004 459418 278186 459654
rect 278422 459418 278604 459654
rect 278004 459334 278604 459418
rect 278004 459098 278186 459334
rect 278422 459098 278604 459334
rect 278004 423654 278604 459098
rect 278004 423418 278186 423654
rect 278422 423418 278604 423654
rect 278004 423334 278604 423418
rect 278004 423098 278186 423334
rect 278422 423098 278604 423334
rect 276795 399396 276861 399397
rect 276795 399332 276796 399396
rect 276860 399332 276861 399396
rect 276795 399331 276861 399332
rect 276798 398717 276858 399331
rect 276795 398716 276861 398717
rect 276795 398652 276796 398716
rect 276860 398652 276861 398716
rect 276795 398651 276861 398652
rect 274404 383818 274586 384054
rect 274822 383818 275004 384054
rect 274404 383734 275004 383818
rect 274404 383498 274586 383734
rect 274822 383498 275004 383734
rect 274404 348054 275004 383498
rect 274404 347818 274586 348054
rect 274822 347818 275004 348054
rect 274404 347734 275004 347818
rect 274404 347498 274586 347734
rect 274822 347498 275004 347734
rect 274404 312054 275004 347498
rect 274404 311818 274586 312054
rect 274822 311818 275004 312054
rect 274404 311734 275004 311818
rect 274404 311498 274586 311734
rect 274822 311498 275004 311734
rect 274404 276054 275004 311498
rect 274404 275818 274586 276054
rect 274822 275818 275004 276054
rect 274404 275734 275004 275818
rect 274404 275498 274586 275734
rect 274822 275498 275004 275734
rect 274404 240054 275004 275498
rect 274404 239818 274586 240054
rect 274822 239818 275004 240054
rect 274404 239734 275004 239818
rect 274404 239498 274586 239734
rect 274822 239498 275004 239734
rect 274404 204054 275004 239498
rect 274404 203818 274586 204054
rect 274822 203818 275004 204054
rect 274404 203734 275004 203818
rect 274404 203498 274586 203734
rect 274822 203498 275004 203734
rect 274404 168054 275004 203498
rect 274404 167818 274586 168054
rect 274822 167818 275004 168054
rect 274404 167734 275004 167818
rect 274404 167498 274586 167734
rect 274822 167498 275004 167734
rect 274404 132054 275004 167498
rect 274404 131818 274586 132054
rect 274822 131818 275004 132054
rect 274404 131734 275004 131818
rect 274404 131498 274586 131734
rect 274822 131498 275004 131734
rect 274404 96054 275004 131498
rect 274404 95818 274586 96054
rect 274822 95818 275004 96054
rect 274404 95734 275004 95818
rect 274404 95498 274586 95734
rect 274822 95498 275004 95734
rect 274404 60054 275004 95498
rect 274404 59818 274586 60054
rect 274822 59818 275004 60054
rect 274404 59734 275004 59818
rect 274404 59498 274586 59734
rect 274822 59498 275004 59734
rect 274404 24054 275004 59498
rect 274404 23818 274586 24054
rect 274822 23818 275004 24054
rect 274404 23734 275004 23818
rect 274404 23498 274586 23734
rect 274822 23498 275004 23734
rect 274404 -3106 275004 23498
rect 274404 -3342 274586 -3106
rect 274822 -3342 275004 -3106
rect 274404 -3426 275004 -3342
rect 274404 -3662 274586 -3426
rect 274822 -3662 275004 -3426
rect 274404 -3684 275004 -3662
rect 278004 387654 278604 423098
rect 278004 387418 278186 387654
rect 278422 387418 278604 387654
rect 278004 387334 278604 387418
rect 278004 387098 278186 387334
rect 278422 387098 278604 387334
rect 278004 351654 278604 387098
rect 278004 351418 278186 351654
rect 278422 351418 278604 351654
rect 278004 351334 278604 351418
rect 278004 351098 278186 351334
rect 278422 351098 278604 351334
rect 278004 315654 278604 351098
rect 278004 315418 278186 315654
rect 278422 315418 278604 315654
rect 278004 315334 278604 315418
rect 278004 315098 278186 315334
rect 278422 315098 278604 315334
rect 278004 279654 278604 315098
rect 278004 279418 278186 279654
rect 278422 279418 278604 279654
rect 278004 279334 278604 279418
rect 278004 279098 278186 279334
rect 278422 279098 278604 279334
rect 278004 243654 278604 279098
rect 278004 243418 278186 243654
rect 278422 243418 278604 243654
rect 278004 243334 278604 243418
rect 278004 243098 278186 243334
rect 278422 243098 278604 243334
rect 278004 207654 278604 243098
rect 278004 207418 278186 207654
rect 278422 207418 278604 207654
rect 278004 207334 278604 207418
rect 278004 207098 278186 207334
rect 278422 207098 278604 207334
rect 278004 171654 278604 207098
rect 278004 171418 278186 171654
rect 278422 171418 278604 171654
rect 278004 171334 278604 171418
rect 278004 171098 278186 171334
rect 278422 171098 278604 171334
rect 278004 135654 278604 171098
rect 278004 135418 278186 135654
rect 278422 135418 278604 135654
rect 278004 135334 278604 135418
rect 278004 135098 278186 135334
rect 278422 135098 278604 135334
rect 278004 99654 278604 135098
rect 278004 99418 278186 99654
rect 278422 99418 278604 99654
rect 278004 99334 278604 99418
rect 278004 99098 278186 99334
rect 278422 99098 278604 99334
rect 278004 63654 278604 99098
rect 278004 63418 278186 63654
rect 278422 63418 278604 63654
rect 278004 63334 278604 63418
rect 278004 63098 278186 63334
rect 278422 63098 278604 63334
rect 278004 27654 278604 63098
rect 278004 27418 278186 27654
rect 278422 27418 278604 27654
rect 278004 27334 278604 27418
rect 278004 27098 278186 27334
rect 278422 27098 278604 27334
rect 278004 -4946 278604 27098
rect 278004 -5182 278186 -4946
rect 278422 -5182 278604 -4946
rect 278004 -5266 278604 -5182
rect 278004 -5502 278186 -5266
rect 278422 -5502 278604 -5266
rect 278004 -5524 278604 -5502
rect 281604 679254 282204 710722
rect 299604 710358 300204 711300
rect 299604 710122 299786 710358
rect 300022 710122 300204 710358
rect 299604 710038 300204 710122
rect 299604 709802 299786 710038
rect 300022 709802 300204 710038
rect 296004 708518 296604 709460
rect 296004 708282 296186 708518
rect 296422 708282 296604 708518
rect 296004 708198 296604 708282
rect 296004 707962 296186 708198
rect 296422 707962 296604 708198
rect 292404 706678 293004 707620
rect 292404 706442 292586 706678
rect 292822 706442 293004 706678
rect 292404 706358 293004 706442
rect 292404 706122 292586 706358
rect 292822 706122 293004 706358
rect 281604 679018 281786 679254
rect 282022 679018 282204 679254
rect 281604 678934 282204 679018
rect 281604 678698 281786 678934
rect 282022 678698 282204 678934
rect 281604 643254 282204 678698
rect 281604 643018 281786 643254
rect 282022 643018 282204 643254
rect 281604 642934 282204 643018
rect 281604 642698 281786 642934
rect 282022 642698 282204 642934
rect 281604 607254 282204 642698
rect 281604 607018 281786 607254
rect 282022 607018 282204 607254
rect 281604 606934 282204 607018
rect 281604 606698 281786 606934
rect 282022 606698 282204 606934
rect 281604 571254 282204 606698
rect 281604 571018 281786 571254
rect 282022 571018 282204 571254
rect 281604 570934 282204 571018
rect 281604 570698 281786 570934
rect 282022 570698 282204 570934
rect 281604 535254 282204 570698
rect 281604 535018 281786 535254
rect 282022 535018 282204 535254
rect 281604 534934 282204 535018
rect 281604 534698 281786 534934
rect 282022 534698 282204 534934
rect 281604 499254 282204 534698
rect 281604 499018 281786 499254
rect 282022 499018 282204 499254
rect 281604 498934 282204 499018
rect 281604 498698 281786 498934
rect 282022 498698 282204 498934
rect 281604 463254 282204 498698
rect 281604 463018 281786 463254
rect 282022 463018 282204 463254
rect 281604 462934 282204 463018
rect 281604 462698 281786 462934
rect 282022 462698 282204 462934
rect 281604 427254 282204 462698
rect 281604 427018 281786 427254
rect 282022 427018 282204 427254
rect 281604 426934 282204 427018
rect 281604 426698 281786 426934
rect 282022 426698 282204 426934
rect 281604 391254 282204 426698
rect 288804 704838 289404 705780
rect 288804 704602 288986 704838
rect 289222 704602 289404 704838
rect 288804 704518 289404 704602
rect 288804 704282 288986 704518
rect 289222 704282 289404 704518
rect 288804 686454 289404 704282
rect 288804 686218 288986 686454
rect 289222 686218 289404 686454
rect 288804 686134 289404 686218
rect 288804 685898 288986 686134
rect 289222 685898 289404 686134
rect 288804 650454 289404 685898
rect 288804 650218 288986 650454
rect 289222 650218 289404 650454
rect 288804 650134 289404 650218
rect 288804 649898 288986 650134
rect 289222 649898 289404 650134
rect 288804 614454 289404 649898
rect 288804 614218 288986 614454
rect 289222 614218 289404 614454
rect 288804 614134 289404 614218
rect 288804 613898 288986 614134
rect 289222 613898 289404 614134
rect 288804 578454 289404 613898
rect 288804 578218 288986 578454
rect 289222 578218 289404 578454
rect 288804 578134 289404 578218
rect 288804 577898 288986 578134
rect 289222 577898 289404 578134
rect 288804 542454 289404 577898
rect 288804 542218 288986 542454
rect 289222 542218 289404 542454
rect 288804 542134 289404 542218
rect 288804 541898 288986 542134
rect 289222 541898 289404 542134
rect 288804 506454 289404 541898
rect 288804 506218 288986 506454
rect 289222 506218 289404 506454
rect 288804 506134 289404 506218
rect 288804 505898 288986 506134
rect 289222 505898 289404 506134
rect 288804 470454 289404 505898
rect 288804 470218 288986 470454
rect 289222 470218 289404 470454
rect 288804 470134 289404 470218
rect 288804 469898 288986 470134
rect 289222 469898 289404 470134
rect 288804 434454 289404 469898
rect 288804 434218 288986 434454
rect 289222 434218 289404 434454
rect 288804 434134 289404 434218
rect 288804 433898 288986 434134
rect 289222 433898 289404 434134
rect 282867 399396 282933 399397
rect 282867 399332 282868 399396
rect 282932 399332 282933 399396
rect 282867 399331 282933 399332
rect 284339 399396 284405 399397
rect 284339 399332 284340 399396
rect 284404 399332 284405 399396
rect 284339 399331 284405 399332
rect 285627 399396 285693 399397
rect 285627 399332 285628 399396
rect 285692 399332 285693 399396
rect 285627 399331 285693 399332
rect 287283 399396 287349 399397
rect 287283 399332 287284 399396
rect 287348 399332 287349 399396
rect 287283 399331 287349 399332
rect 287835 399396 287901 399397
rect 287835 399332 287836 399396
rect 287900 399332 287901 399396
rect 287835 399331 287901 399332
rect 281604 391018 281786 391254
rect 282022 391018 282204 391254
rect 281604 390934 282204 391018
rect 281604 390698 281786 390934
rect 282022 390698 282204 390934
rect 281604 355254 282204 390698
rect 281604 355018 281786 355254
rect 282022 355018 282204 355254
rect 281604 354934 282204 355018
rect 281604 354698 281786 354934
rect 282022 354698 282204 354934
rect 281604 319254 282204 354698
rect 281604 319018 281786 319254
rect 282022 319018 282204 319254
rect 281604 318934 282204 319018
rect 281604 318698 281786 318934
rect 282022 318698 282204 318934
rect 281604 283254 282204 318698
rect 281604 283018 281786 283254
rect 282022 283018 282204 283254
rect 281604 282934 282204 283018
rect 281604 282698 281786 282934
rect 282022 282698 282204 282934
rect 281604 247254 282204 282698
rect 281604 247018 281786 247254
rect 282022 247018 282204 247254
rect 281604 246934 282204 247018
rect 281604 246698 281786 246934
rect 282022 246698 282204 246934
rect 281604 211254 282204 246698
rect 281604 211018 281786 211254
rect 282022 211018 282204 211254
rect 281604 210934 282204 211018
rect 281604 210698 281786 210934
rect 282022 210698 282204 210934
rect 281604 175254 282204 210698
rect 282870 194581 282930 399331
rect 284342 398037 284402 399331
rect 284339 398036 284405 398037
rect 284339 397972 284340 398036
rect 284404 397972 284405 398036
rect 284339 397971 284405 397972
rect 282867 194580 282933 194581
rect 282867 194516 282868 194580
rect 282932 194516 282933 194580
rect 282867 194515 282933 194516
rect 281604 175018 281786 175254
rect 282022 175018 282204 175254
rect 281604 174934 282204 175018
rect 281604 174698 281786 174934
rect 282022 174698 282204 174934
rect 281604 139254 282204 174698
rect 281604 139018 281786 139254
rect 282022 139018 282204 139254
rect 281604 138934 282204 139018
rect 281604 138698 281786 138934
rect 282022 138698 282204 138934
rect 281604 103254 282204 138698
rect 285630 109037 285690 399331
rect 287286 398309 287346 399331
rect 287283 398308 287349 398309
rect 287283 398244 287284 398308
rect 287348 398244 287349 398308
rect 287283 398243 287349 398244
rect 287838 398173 287898 399331
rect 288804 398454 289404 433898
rect 288804 398218 288986 398454
rect 289222 398218 289404 398454
rect 287835 398172 287901 398173
rect 287835 398108 287836 398172
rect 287900 398108 287901 398172
rect 287835 398107 287901 398108
rect 288804 398134 289404 398218
rect 288804 397898 288986 398134
rect 289222 397898 289404 398134
rect 288804 362454 289404 397898
rect 288804 362218 288986 362454
rect 289222 362218 289404 362454
rect 288804 362134 289404 362218
rect 288804 361898 288986 362134
rect 289222 361898 289404 362134
rect 288804 326454 289404 361898
rect 288804 326218 288986 326454
rect 289222 326218 289404 326454
rect 288804 326134 289404 326218
rect 288804 325898 288986 326134
rect 289222 325898 289404 326134
rect 288804 290454 289404 325898
rect 288804 290218 288986 290454
rect 289222 290218 289404 290454
rect 288804 290134 289404 290218
rect 288804 289898 288986 290134
rect 289222 289898 289404 290134
rect 288804 254454 289404 289898
rect 288804 254218 288986 254454
rect 289222 254218 289404 254454
rect 288804 254134 289404 254218
rect 288804 253898 288986 254134
rect 289222 253898 289404 254134
rect 288804 218454 289404 253898
rect 288804 218218 288986 218454
rect 289222 218218 289404 218454
rect 288804 218134 289404 218218
rect 288804 217898 288986 218134
rect 289222 217898 289404 218134
rect 288804 182454 289404 217898
rect 288804 182218 288986 182454
rect 289222 182218 289404 182454
rect 288804 182134 289404 182218
rect 288804 181898 288986 182134
rect 289222 181898 289404 182134
rect 288804 146454 289404 181898
rect 288804 146218 288986 146454
rect 289222 146218 289404 146454
rect 288804 146134 289404 146218
rect 288804 145898 288986 146134
rect 289222 145898 289404 146134
rect 288804 110454 289404 145898
rect 288804 110218 288986 110454
rect 289222 110218 289404 110454
rect 288804 110134 289404 110218
rect 288804 109898 288986 110134
rect 289222 109898 289404 110134
rect 285627 109036 285693 109037
rect 285627 108972 285628 109036
rect 285692 108972 285693 109036
rect 285627 108971 285693 108972
rect 281604 103018 281786 103254
rect 282022 103018 282204 103254
rect 281604 102934 282204 103018
rect 281604 102698 281786 102934
rect 282022 102698 282204 102934
rect 281604 67254 282204 102698
rect 281604 67018 281786 67254
rect 282022 67018 282204 67254
rect 281604 66934 282204 67018
rect 281604 66698 281786 66934
rect 282022 66698 282204 66934
rect 281604 31254 282204 66698
rect 281604 31018 281786 31254
rect 282022 31018 282204 31254
rect 281604 30934 282204 31018
rect 281604 30698 281786 30934
rect 282022 30698 282204 30934
rect 263604 -6102 263786 -5866
rect 264022 -6102 264204 -5866
rect 263604 -6186 264204 -6102
rect 263604 -6422 263786 -6186
rect 264022 -6422 264204 -6186
rect 263604 -7364 264204 -6422
rect 281604 -6786 282204 30698
rect 288804 74454 289404 109898
rect 288804 74218 288986 74454
rect 289222 74218 289404 74454
rect 288804 74134 289404 74218
rect 288804 73898 288986 74134
rect 289222 73898 289404 74134
rect 288804 38454 289404 73898
rect 288804 38218 288986 38454
rect 289222 38218 289404 38454
rect 288804 38134 289404 38218
rect 288804 37898 288986 38134
rect 289222 37898 289404 38134
rect 288804 2454 289404 37898
rect 288804 2218 288986 2454
rect 289222 2218 289404 2454
rect 288804 2134 289404 2218
rect 288804 1898 288986 2134
rect 289222 1898 289404 2134
rect 288804 -346 289404 1898
rect 288804 -582 288986 -346
rect 289222 -582 289404 -346
rect 288804 -666 289404 -582
rect 288804 -902 288986 -666
rect 289222 -902 289404 -666
rect 288804 -1844 289404 -902
rect 292404 690054 293004 706122
rect 292404 689818 292586 690054
rect 292822 689818 293004 690054
rect 292404 689734 293004 689818
rect 292404 689498 292586 689734
rect 292822 689498 293004 689734
rect 292404 654054 293004 689498
rect 292404 653818 292586 654054
rect 292822 653818 293004 654054
rect 292404 653734 293004 653818
rect 292404 653498 292586 653734
rect 292822 653498 293004 653734
rect 292404 618054 293004 653498
rect 292404 617818 292586 618054
rect 292822 617818 293004 618054
rect 292404 617734 293004 617818
rect 292404 617498 292586 617734
rect 292822 617498 293004 617734
rect 292404 582054 293004 617498
rect 292404 581818 292586 582054
rect 292822 581818 293004 582054
rect 292404 581734 293004 581818
rect 292404 581498 292586 581734
rect 292822 581498 293004 581734
rect 292404 546054 293004 581498
rect 292404 545818 292586 546054
rect 292822 545818 293004 546054
rect 292404 545734 293004 545818
rect 292404 545498 292586 545734
rect 292822 545498 293004 545734
rect 292404 510054 293004 545498
rect 292404 509818 292586 510054
rect 292822 509818 293004 510054
rect 292404 509734 293004 509818
rect 292404 509498 292586 509734
rect 292822 509498 293004 509734
rect 292404 474054 293004 509498
rect 292404 473818 292586 474054
rect 292822 473818 293004 474054
rect 292404 473734 293004 473818
rect 292404 473498 292586 473734
rect 292822 473498 293004 473734
rect 292404 438054 293004 473498
rect 292404 437818 292586 438054
rect 292822 437818 293004 438054
rect 292404 437734 293004 437818
rect 292404 437498 292586 437734
rect 292822 437498 293004 437734
rect 292404 402054 293004 437498
rect 292404 401818 292586 402054
rect 292822 401818 293004 402054
rect 292404 401734 293004 401818
rect 292404 401498 292586 401734
rect 292822 401498 293004 401734
rect 292404 366054 293004 401498
rect 292404 365818 292586 366054
rect 292822 365818 293004 366054
rect 292404 365734 293004 365818
rect 292404 365498 292586 365734
rect 292822 365498 293004 365734
rect 292404 330054 293004 365498
rect 292404 329818 292586 330054
rect 292822 329818 293004 330054
rect 292404 329734 293004 329818
rect 292404 329498 292586 329734
rect 292822 329498 293004 329734
rect 292404 294054 293004 329498
rect 292404 293818 292586 294054
rect 292822 293818 293004 294054
rect 292404 293734 293004 293818
rect 292404 293498 292586 293734
rect 292822 293498 293004 293734
rect 292404 258054 293004 293498
rect 292404 257818 292586 258054
rect 292822 257818 293004 258054
rect 292404 257734 293004 257818
rect 292404 257498 292586 257734
rect 292822 257498 293004 257734
rect 292404 222054 293004 257498
rect 292404 221818 292586 222054
rect 292822 221818 293004 222054
rect 292404 221734 293004 221818
rect 292404 221498 292586 221734
rect 292822 221498 293004 221734
rect 292404 186054 293004 221498
rect 292404 185818 292586 186054
rect 292822 185818 293004 186054
rect 292404 185734 293004 185818
rect 292404 185498 292586 185734
rect 292822 185498 293004 185734
rect 292404 150054 293004 185498
rect 292404 149818 292586 150054
rect 292822 149818 293004 150054
rect 292404 149734 293004 149818
rect 292404 149498 292586 149734
rect 292822 149498 293004 149734
rect 292404 114054 293004 149498
rect 292404 113818 292586 114054
rect 292822 113818 293004 114054
rect 292404 113734 293004 113818
rect 292404 113498 292586 113734
rect 292822 113498 293004 113734
rect 292404 78054 293004 113498
rect 292404 77818 292586 78054
rect 292822 77818 293004 78054
rect 292404 77734 293004 77818
rect 292404 77498 292586 77734
rect 292822 77498 293004 77734
rect 292404 42054 293004 77498
rect 292404 41818 292586 42054
rect 292822 41818 293004 42054
rect 292404 41734 293004 41818
rect 292404 41498 292586 41734
rect 292822 41498 293004 41734
rect 292404 6054 293004 41498
rect 292404 5818 292586 6054
rect 292822 5818 293004 6054
rect 292404 5734 293004 5818
rect 292404 5498 292586 5734
rect 292822 5498 293004 5734
rect 292404 -2186 293004 5498
rect 292404 -2422 292586 -2186
rect 292822 -2422 293004 -2186
rect 292404 -2506 293004 -2422
rect 292404 -2742 292586 -2506
rect 292822 -2742 293004 -2506
rect 292404 -3684 293004 -2742
rect 296004 693654 296604 707962
rect 296004 693418 296186 693654
rect 296422 693418 296604 693654
rect 296004 693334 296604 693418
rect 296004 693098 296186 693334
rect 296422 693098 296604 693334
rect 296004 657654 296604 693098
rect 296004 657418 296186 657654
rect 296422 657418 296604 657654
rect 296004 657334 296604 657418
rect 296004 657098 296186 657334
rect 296422 657098 296604 657334
rect 296004 621654 296604 657098
rect 296004 621418 296186 621654
rect 296422 621418 296604 621654
rect 296004 621334 296604 621418
rect 296004 621098 296186 621334
rect 296422 621098 296604 621334
rect 296004 585654 296604 621098
rect 296004 585418 296186 585654
rect 296422 585418 296604 585654
rect 296004 585334 296604 585418
rect 296004 585098 296186 585334
rect 296422 585098 296604 585334
rect 296004 549654 296604 585098
rect 296004 549418 296186 549654
rect 296422 549418 296604 549654
rect 296004 549334 296604 549418
rect 296004 549098 296186 549334
rect 296422 549098 296604 549334
rect 296004 513654 296604 549098
rect 296004 513418 296186 513654
rect 296422 513418 296604 513654
rect 296004 513334 296604 513418
rect 296004 513098 296186 513334
rect 296422 513098 296604 513334
rect 296004 477654 296604 513098
rect 296004 477418 296186 477654
rect 296422 477418 296604 477654
rect 296004 477334 296604 477418
rect 296004 477098 296186 477334
rect 296422 477098 296604 477334
rect 296004 441654 296604 477098
rect 296004 441418 296186 441654
rect 296422 441418 296604 441654
rect 296004 441334 296604 441418
rect 296004 441098 296186 441334
rect 296422 441098 296604 441334
rect 296004 405654 296604 441098
rect 296004 405418 296186 405654
rect 296422 405418 296604 405654
rect 296004 405334 296604 405418
rect 296004 405098 296186 405334
rect 296422 405098 296604 405334
rect 296004 369654 296604 405098
rect 296004 369418 296186 369654
rect 296422 369418 296604 369654
rect 296004 369334 296604 369418
rect 296004 369098 296186 369334
rect 296422 369098 296604 369334
rect 296004 333654 296604 369098
rect 296004 333418 296186 333654
rect 296422 333418 296604 333654
rect 296004 333334 296604 333418
rect 296004 333098 296186 333334
rect 296422 333098 296604 333334
rect 296004 297654 296604 333098
rect 296004 297418 296186 297654
rect 296422 297418 296604 297654
rect 296004 297334 296604 297418
rect 296004 297098 296186 297334
rect 296422 297098 296604 297334
rect 296004 261654 296604 297098
rect 296004 261418 296186 261654
rect 296422 261418 296604 261654
rect 296004 261334 296604 261418
rect 296004 261098 296186 261334
rect 296422 261098 296604 261334
rect 296004 225654 296604 261098
rect 296004 225418 296186 225654
rect 296422 225418 296604 225654
rect 296004 225334 296604 225418
rect 296004 225098 296186 225334
rect 296422 225098 296604 225334
rect 296004 189654 296604 225098
rect 296004 189418 296186 189654
rect 296422 189418 296604 189654
rect 296004 189334 296604 189418
rect 296004 189098 296186 189334
rect 296422 189098 296604 189334
rect 296004 153654 296604 189098
rect 296004 153418 296186 153654
rect 296422 153418 296604 153654
rect 296004 153334 296604 153418
rect 296004 153098 296186 153334
rect 296422 153098 296604 153334
rect 296004 117654 296604 153098
rect 296004 117418 296186 117654
rect 296422 117418 296604 117654
rect 296004 117334 296604 117418
rect 296004 117098 296186 117334
rect 296422 117098 296604 117334
rect 296004 81654 296604 117098
rect 296004 81418 296186 81654
rect 296422 81418 296604 81654
rect 296004 81334 296604 81418
rect 296004 81098 296186 81334
rect 296422 81098 296604 81334
rect 296004 45654 296604 81098
rect 296004 45418 296186 45654
rect 296422 45418 296604 45654
rect 296004 45334 296604 45418
rect 296004 45098 296186 45334
rect 296422 45098 296604 45334
rect 296004 9654 296604 45098
rect 296004 9418 296186 9654
rect 296422 9418 296604 9654
rect 296004 9334 296604 9418
rect 296004 9098 296186 9334
rect 296422 9098 296604 9334
rect 296004 -4026 296604 9098
rect 296004 -4262 296186 -4026
rect 296422 -4262 296604 -4026
rect 296004 -4346 296604 -4262
rect 296004 -4582 296186 -4346
rect 296422 -4582 296604 -4346
rect 296004 -5524 296604 -4582
rect 299604 697254 300204 709802
rect 317604 711278 318204 711300
rect 317604 711042 317786 711278
rect 318022 711042 318204 711278
rect 317604 710958 318204 711042
rect 317604 710722 317786 710958
rect 318022 710722 318204 710958
rect 314004 709438 314604 709460
rect 314004 709202 314186 709438
rect 314422 709202 314604 709438
rect 314004 709118 314604 709202
rect 314004 708882 314186 709118
rect 314422 708882 314604 709118
rect 310404 707598 311004 707620
rect 310404 707362 310586 707598
rect 310822 707362 311004 707598
rect 310404 707278 311004 707362
rect 310404 707042 310586 707278
rect 310822 707042 311004 707278
rect 299604 697018 299786 697254
rect 300022 697018 300204 697254
rect 299604 696934 300204 697018
rect 299604 696698 299786 696934
rect 300022 696698 300204 696934
rect 299604 661254 300204 696698
rect 299604 661018 299786 661254
rect 300022 661018 300204 661254
rect 299604 660934 300204 661018
rect 299604 660698 299786 660934
rect 300022 660698 300204 660934
rect 299604 625254 300204 660698
rect 299604 625018 299786 625254
rect 300022 625018 300204 625254
rect 299604 624934 300204 625018
rect 299604 624698 299786 624934
rect 300022 624698 300204 624934
rect 299604 589254 300204 624698
rect 299604 589018 299786 589254
rect 300022 589018 300204 589254
rect 299604 588934 300204 589018
rect 299604 588698 299786 588934
rect 300022 588698 300204 588934
rect 299604 553254 300204 588698
rect 299604 553018 299786 553254
rect 300022 553018 300204 553254
rect 299604 552934 300204 553018
rect 299604 552698 299786 552934
rect 300022 552698 300204 552934
rect 299604 517254 300204 552698
rect 299604 517018 299786 517254
rect 300022 517018 300204 517254
rect 299604 516934 300204 517018
rect 299604 516698 299786 516934
rect 300022 516698 300204 516934
rect 299604 481254 300204 516698
rect 299604 481018 299786 481254
rect 300022 481018 300204 481254
rect 299604 480934 300204 481018
rect 299604 480698 299786 480934
rect 300022 480698 300204 480934
rect 299604 445254 300204 480698
rect 299604 445018 299786 445254
rect 300022 445018 300204 445254
rect 299604 444934 300204 445018
rect 299604 444698 299786 444934
rect 300022 444698 300204 444934
rect 299604 409254 300204 444698
rect 299604 409018 299786 409254
rect 300022 409018 300204 409254
rect 299604 408934 300204 409018
rect 299604 408698 299786 408934
rect 300022 408698 300204 408934
rect 299604 373254 300204 408698
rect 299604 373018 299786 373254
rect 300022 373018 300204 373254
rect 299604 372934 300204 373018
rect 299604 372698 299786 372934
rect 300022 372698 300204 372934
rect 299604 337254 300204 372698
rect 299604 337018 299786 337254
rect 300022 337018 300204 337254
rect 299604 336934 300204 337018
rect 299604 336698 299786 336934
rect 300022 336698 300204 336934
rect 299604 301254 300204 336698
rect 299604 301018 299786 301254
rect 300022 301018 300204 301254
rect 299604 300934 300204 301018
rect 299604 300698 299786 300934
rect 300022 300698 300204 300934
rect 299604 265254 300204 300698
rect 299604 265018 299786 265254
rect 300022 265018 300204 265254
rect 299604 264934 300204 265018
rect 299604 264698 299786 264934
rect 300022 264698 300204 264934
rect 299604 229254 300204 264698
rect 299604 229018 299786 229254
rect 300022 229018 300204 229254
rect 299604 228934 300204 229018
rect 299604 228698 299786 228934
rect 300022 228698 300204 228934
rect 299604 193254 300204 228698
rect 299604 193018 299786 193254
rect 300022 193018 300204 193254
rect 299604 192934 300204 193018
rect 299604 192698 299786 192934
rect 300022 192698 300204 192934
rect 299604 157254 300204 192698
rect 299604 157018 299786 157254
rect 300022 157018 300204 157254
rect 299604 156934 300204 157018
rect 299604 156698 299786 156934
rect 300022 156698 300204 156934
rect 299604 121254 300204 156698
rect 299604 121018 299786 121254
rect 300022 121018 300204 121254
rect 299604 120934 300204 121018
rect 299604 120698 299786 120934
rect 300022 120698 300204 120934
rect 299604 85254 300204 120698
rect 299604 85018 299786 85254
rect 300022 85018 300204 85254
rect 299604 84934 300204 85018
rect 299604 84698 299786 84934
rect 300022 84698 300204 84934
rect 299604 49254 300204 84698
rect 299604 49018 299786 49254
rect 300022 49018 300204 49254
rect 299604 48934 300204 49018
rect 299604 48698 299786 48934
rect 300022 48698 300204 48934
rect 299604 13254 300204 48698
rect 299604 13018 299786 13254
rect 300022 13018 300204 13254
rect 299604 12934 300204 13018
rect 299604 12698 299786 12934
rect 300022 12698 300204 12934
rect 281604 -7022 281786 -6786
rect 282022 -7022 282204 -6786
rect 281604 -7106 282204 -7022
rect 281604 -7342 281786 -7106
rect 282022 -7342 282204 -7106
rect 281604 -7364 282204 -7342
rect 299604 -5866 300204 12698
rect 306804 705758 307404 705780
rect 306804 705522 306986 705758
rect 307222 705522 307404 705758
rect 306804 705438 307404 705522
rect 306804 705202 306986 705438
rect 307222 705202 307404 705438
rect 306804 668454 307404 705202
rect 306804 668218 306986 668454
rect 307222 668218 307404 668454
rect 306804 668134 307404 668218
rect 306804 667898 306986 668134
rect 307222 667898 307404 668134
rect 306804 632454 307404 667898
rect 306804 632218 306986 632454
rect 307222 632218 307404 632454
rect 306804 632134 307404 632218
rect 306804 631898 306986 632134
rect 307222 631898 307404 632134
rect 306804 596454 307404 631898
rect 306804 596218 306986 596454
rect 307222 596218 307404 596454
rect 306804 596134 307404 596218
rect 306804 595898 306986 596134
rect 307222 595898 307404 596134
rect 306804 560454 307404 595898
rect 306804 560218 306986 560454
rect 307222 560218 307404 560454
rect 306804 560134 307404 560218
rect 306804 559898 306986 560134
rect 307222 559898 307404 560134
rect 306804 524454 307404 559898
rect 306804 524218 306986 524454
rect 307222 524218 307404 524454
rect 306804 524134 307404 524218
rect 306804 523898 306986 524134
rect 307222 523898 307404 524134
rect 306804 488454 307404 523898
rect 306804 488218 306986 488454
rect 307222 488218 307404 488454
rect 306804 488134 307404 488218
rect 306804 487898 306986 488134
rect 307222 487898 307404 488134
rect 306804 452454 307404 487898
rect 306804 452218 306986 452454
rect 307222 452218 307404 452454
rect 306804 452134 307404 452218
rect 306804 451898 306986 452134
rect 307222 451898 307404 452134
rect 306804 416454 307404 451898
rect 306804 416218 306986 416454
rect 307222 416218 307404 416454
rect 306804 416134 307404 416218
rect 306804 415898 306986 416134
rect 307222 415898 307404 416134
rect 306804 380454 307404 415898
rect 306804 380218 306986 380454
rect 307222 380218 307404 380454
rect 306804 380134 307404 380218
rect 306804 379898 306986 380134
rect 307222 379898 307404 380134
rect 306804 344454 307404 379898
rect 306804 344218 306986 344454
rect 307222 344218 307404 344454
rect 306804 344134 307404 344218
rect 306804 343898 306986 344134
rect 307222 343898 307404 344134
rect 306804 308454 307404 343898
rect 306804 308218 306986 308454
rect 307222 308218 307404 308454
rect 306804 308134 307404 308218
rect 306804 307898 306986 308134
rect 307222 307898 307404 308134
rect 306804 272454 307404 307898
rect 306804 272218 306986 272454
rect 307222 272218 307404 272454
rect 306804 272134 307404 272218
rect 306804 271898 306986 272134
rect 307222 271898 307404 272134
rect 306804 236454 307404 271898
rect 306804 236218 306986 236454
rect 307222 236218 307404 236454
rect 306804 236134 307404 236218
rect 306804 235898 306986 236134
rect 307222 235898 307404 236134
rect 306804 200454 307404 235898
rect 306804 200218 306986 200454
rect 307222 200218 307404 200454
rect 306804 200134 307404 200218
rect 306804 199898 306986 200134
rect 307222 199898 307404 200134
rect 306804 164454 307404 199898
rect 306804 164218 306986 164454
rect 307222 164218 307404 164454
rect 306804 164134 307404 164218
rect 306804 163898 306986 164134
rect 307222 163898 307404 164134
rect 306804 128454 307404 163898
rect 306804 128218 306986 128454
rect 307222 128218 307404 128454
rect 306804 128134 307404 128218
rect 306804 127898 306986 128134
rect 307222 127898 307404 128134
rect 306804 92454 307404 127898
rect 306804 92218 306986 92454
rect 307222 92218 307404 92454
rect 306804 92134 307404 92218
rect 306804 91898 306986 92134
rect 307222 91898 307404 92134
rect 306804 56454 307404 91898
rect 306804 56218 306986 56454
rect 307222 56218 307404 56454
rect 306804 56134 307404 56218
rect 306804 55898 306986 56134
rect 307222 55898 307404 56134
rect 306804 20454 307404 55898
rect 306804 20218 306986 20454
rect 307222 20218 307404 20454
rect 306804 20134 307404 20218
rect 306804 19898 306986 20134
rect 307222 19898 307404 20134
rect 306804 -1266 307404 19898
rect 306804 -1502 306986 -1266
rect 307222 -1502 307404 -1266
rect 306804 -1586 307404 -1502
rect 306804 -1822 306986 -1586
rect 307222 -1822 307404 -1586
rect 306804 -1844 307404 -1822
rect 310404 672054 311004 707042
rect 310404 671818 310586 672054
rect 310822 671818 311004 672054
rect 310404 671734 311004 671818
rect 310404 671498 310586 671734
rect 310822 671498 311004 671734
rect 310404 636054 311004 671498
rect 310404 635818 310586 636054
rect 310822 635818 311004 636054
rect 310404 635734 311004 635818
rect 310404 635498 310586 635734
rect 310822 635498 311004 635734
rect 310404 600054 311004 635498
rect 310404 599818 310586 600054
rect 310822 599818 311004 600054
rect 310404 599734 311004 599818
rect 310404 599498 310586 599734
rect 310822 599498 311004 599734
rect 310404 564054 311004 599498
rect 310404 563818 310586 564054
rect 310822 563818 311004 564054
rect 310404 563734 311004 563818
rect 310404 563498 310586 563734
rect 310822 563498 311004 563734
rect 310404 528054 311004 563498
rect 310404 527818 310586 528054
rect 310822 527818 311004 528054
rect 310404 527734 311004 527818
rect 310404 527498 310586 527734
rect 310822 527498 311004 527734
rect 310404 492054 311004 527498
rect 310404 491818 310586 492054
rect 310822 491818 311004 492054
rect 310404 491734 311004 491818
rect 310404 491498 310586 491734
rect 310822 491498 311004 491734
rect 310404 456054 311004 491498
rect 310404 455818 310586 456054
rect 310822 455818 311004 456054
rect 310404 455734 311004 455818
rect 310404 455498 310586 455734
rect 310822 455498 311004 455734
rect 310404 420054 311004 455498
rect 310404 419818 310586 420054
rect 310822 419818 311004 420054
rect 310404 419734 311004 419818
rect 310404 419498 310586 419734
rect 310822 419498 311004 419734
rect 310404 384054 311004 419498
rect 310404 383818 310586 384054
rect 310822 383818 311004 384054
rect 310404 383734 311004 383818
rect 310404 383498 310586 383734
rect 310822 383498 311004 383734
rect 310404 348054 311004 383498
rect 310404 347818 310586 348054
rect 310822 347818 311004 348054
rect 310404 347734 311004 347818
rect 310404 347498 310586 347734
rect 310822 347498 311004 347734
rect 310404 312054 311004 347498
rect 310404 311818 310586 312054
rect 310822 311818 311004 312054
rect 310404 311734 311004 311818
rect 310404 311498 310586 311734
rect 310822 311498 311004 311734
rect 310404 276054 311004 311498
rect 310404 275818 310586 276054
rect 310822 275818 311004 276054
rect 310404 275734 311004 275818
rect 310404 275498 310586 275734
rect 310822 275498 311004 275734
rect 310404 240054 311004 275498
rect 310404 239818 310586 240054
rect 310822 239818 311004 240054
rect 310404 239734 311004 239818
rect 310404 239498 310586 239734
rect 310822 239498 311004 239734
rect 310404 204054 311004 239498
rect 310404 203818 310586 204054
rect 310822 203818 311004 204054
rect 310404 203734 311004 203818
rect 310404 203498 310586 203734
rect 310822 203498 311004 203734
rect 310404 168054 311004 203498
rect 310404 167818 310586 168054
rect 310822 167818 311004 168054
rect 310404 167734 311004 167818
rect 310404 167498 310586 167734
rect 310822 167498 311004 167734
rect 310404 132054 311004 167498
rect 310404 131818 310586 132054
rect 310822 131818 311004 132054
rect 310404 131734 311004 131818
rect 310404 131498 310586 131734
rect 310822 131498 311004 131734
rect 310404 96054 311004 131498
rect 310404 95818 310586 96054
rect 310822 95818 311004 96054
rect 310404 95734 311004 95818
rect 310404 95498 310586 95734
rect 310822 95498 311004 95734
rect 310404 60054 311004 95498
rect 310404 59818 310586 60054
rect 310822 59818 311004 60054
rect 310404 59734 311004 59818
rect 310404 59498 310586 59734
rect 310822 59498 311004 59734
rect 310404 24054 311004 59498
rect 310404 23818 310586 24054
rect 310822 23818 311004 24054
rect 310404 23734 311004 23818
rect 310404 23498 310586 23734
rect 310822 23498 311004 23734
rect 310404 -3106 311004 23498
rect 310404 -3342 310586 -3106
rect 310822 -3342 311004 -3106
rect 310404 -3426 311004 -3342
rect 310404 -3662 310586 -3426
rect 310822 -3662 311004 -3426
rect 310404 -3684 311004 -3662
rect 314004 675654 314604 708882
rect 314004 675418 314186 675654
rect 314422 675418 314604 675654
rect 314004 675334 314604 675418
rect 314004 675098 314186 675334
rect 314422 675098 314604 675334
rect 314004 639654 314604 675098
rect 314004 639418 314186 639654
rect 314422 639418 314604 639654
rect 314004 639334 314604 639418
rect 314004 639098 314186 639334
rect 314422 639098 314604 639334
rect 314004 603654 314604 639098
rect 314004 603418 314186 603654
rect 314422 603418 314604 603654
rect 314004 603334 314604 603418
rect 314004 603098 314186 603334
rect 314422 603098 314604 603334
rect 314004 567654 314604 603098
rect 314004 567418 314186 567654
rect 314422 567418 314604 567654
rect 314004 567334 314604 567418
rect 314004 567098 314186 567334
rect 314422 567098 314604 567334
rect 314004 531654 314604 567098
rect 314004 531418 314186 531654
rect 314422 531418 314604 531654
rect 314004 531334 314604 531418
rect 314004 531098 314186 531334
rect 314422 531098 314604 531334
rect 314004 495654 314604 531098
rect 314004 495418 314186 495654
rect 314422 495418 314604 495654
rect 314004 495334 314604 495418
rect 314004 495098 314186 495334
rect 314422 495098 314604 495334
rect 314004 459654 314604 495098
rect 314004 459418 314186 459654
rect 314422 459418 314604 459654
rect 314004 459334 314604 459418
rect 314004 459098 314186 459334
rect 314422 459098 314604 459334
rect 314004 423654 314604 459098
rect 314004 423418 314186 423654
rect 314422 423418 314604 423654
rect 314004 423334 314604 423418
rect 314004 423098 314186 423334
rect 314422 423098 314604 423334
rect 314004 387654 314604 423098
rect 314004 387418 314186 387654
rect 314422 387418 314604 387654
rect 314004 387334 314604 387418
rect 314004 387098 314186 387334
rect 314422 387098 314604 387334
rect 314004 351654 314604 387098
rect 314004 351418 314186 351654
rect 314422 351418 314604 351654
rect 314004 351334 314604 351418
rect 314004 351098 314186 351334
rect 314422 351098 314604 351334
rect 314004 315654 314604 351098
rect 314004 315418 314186 315654
rect 314422 315418 314604 315654
rect 314004 315334 314604 315418
rect 314004 315098 314186 315334
rect 314422 315098 314604 315334
rect 314004 279654 314604 315098
rect 314004 279418 314186 279654
rect 314422 279418 314604 279654
rect 314004 279334 314604 279418
rect 314004 279098 314186 279334
rect 314422 279098 314604 279334
rect 314004 243654 314604 279098
rect 314004 243418 314186 243654
rect 314422 243418 314604 243654
rect 314004 243334 314604 243418
rect 314004 243098 314186 243334
rect 314422 243098 314604 243334
rect 314004 207654 314604 243098
rect 314004 207418 314186 207654
rect 314422 207418 314604 207654
rect 314004 207334 314604 207418
rect 314004 207098 314186 207334
rect 314422 207098 314604 207334
rect 314004 171654 314604 207098
rect 314004 171418 314186 171654
rect 314422 171418 314604 171654
rect 314004 171334 314604 171418
rect 314004 171098 314186 171334
rect 314422 171098 314604 171334
rect 314004 135654 314604 171098
rect 314004 135418 314186 135654
rect 314422 135418 314604 135654
rect 314004 135334 314604 135418
rect 314004 135098 314186 135334
rect 314422 135098 314604 135334
rect 314004 99654 314604 135098
rect 314004 99418 314186 99654
rect 314422 99418 314604 99654
rect 314004 99334 314604 99418
rect 314004 99098 314186 99334
rect 314422 99098 314604 99334
rect 314004 63654 314604 99098
rect 314004 63418 314186 63654
rect 314422 63418 314604 63654
rect 314004 63334 314604 63418
rect 314004 63098 314186 63334
rect 314422 63098 314604 63334
rect 314004 27654 314604 63098
rect 314004 27418 314186 27654
rect 314422 27418 314604 27654
rect 314004 27334 314604 27418
rect 314004 27098 314186 27334
rect 314422 27098 314604 27334
rect 314004 -4946 314604 27098
rect 314004 -5182 314186 -4946
rect 314422 -5182 314604 -4946
rect 314004 -5266 314604 -5182
rect 314004 -5502 314186 -5266
rect 314422 -5502 314604 -5266
rect 314004 -5524 314604 -5502
rect 317604 679254 318204 710722
rect 335604 710358 336204 711300
rect 335604 710122 335786 710358
rect 336022 710122 336204 710358
rect 335604 710038 336204 710122
rect 335604 709802 335786 710038
rect 336022 709802 336204 710038
rect 332004 708518 332604 709460
rect 332004 708282 332186 708518
rect 332422 708282 332604 708518
rect 332004 708198 332604 708282
rect 332004 707962 332186 708198
rect 332422 707962 332604 708198
rect 328404 706678 329004 707620
rect 328404 706442 328586 706678
rect 328822 706442 329004 706678
rect 328404 706358 329004 706442
rect 328404 706122 328586 706358
rect 328822 706122 329004 706358
rect 317604 679018 317786 679254
rect 318022 679018 318204 679254
rect 317604 678934 318204 679018
rect 317604 678698 317786 678934
rect 318022 678698 318204 678934
rect 317604 643254 318204 678698
rect 317604 643018 317786 643254
rect 318022 643018 318204 643254
rect 317604 642934 318204 643018
rect 317604 642698 317786 642934
rect 318022 642698 318204 642934
rect 317604 607254 318204 642698
rect 317604 607018 317786 607254
rect 318022 607018 318204 607254
rect 317604 606934 318204 607018
rect 317604 606698 317786 606934
rect 318022 606698 318204 606934
rect 317604 571254 318204 606698
rect 317604 571018 317786 571254
rect 318022 571018 318204 571254
rect 317604 570934 318204 571018
rect 317604 570698 317786 570934
rect 318022 570698 318204 570934
rect 317604 535254 318204 570698
rect 317604 535018 317786 535254
rect 318022 535018 318204 535254
rect 317604 534934 318204 535018
rect 317604 534698 317786 534934
rect 318022 534698 318204 534934
rect 317604 499254 318204 534698
rect 317604 499018 317786 499254
rect 318022 499018 318204 499254
rect 317604 498934 318204 499018
rect 317604 498698 317786 498934
rect 318022 498698 318204 498934
rect 317604 463254 318204 498698
rect 317604 463018 317786 463254
rect 318022 463018 318204 463254
rect 317604 462934 318204 463018
rect 317604 462698 317786 462934
rect 318022 462698 318204 462934
rect 317604 427254 318204 462698
rect 317604 427018 317786 427254
rect 318022 427018 318204 427254
rect 317604 426934 318204 427018
rect 317604 426698 317786 426934
rect 318022 426698 318204 426934
rect 317604 391254 318204 426698
rect 317604 391018 317786 391254
rect 318022 391018 318204 391254
rect 317604 390934 318204 391018
rect 317604 390698 317786 390934
rect 318022 390698 318204 390934
rect 317604 355254 318204 390698
rect 317604 355018 317786 355254
rect 318022 355018 318204 355254
rect 317604 354934 318204 355018
rect 317604 354698 317786 354934
rect 318022 354698 318204 354934
rect 317604 319254 318204 354698
rect 317604 319018 317786 319254
rect 318022 319018 318204 319254
rect 317604 318934 318204 319018
rect 317604 318698 317786 318934
rect 318022 318698 318204 318934
rect 317604 283254 318204 318698
rect 317604 283018 317786 283254
rect 318022 283018 318204 283254
rect 317604 282934 318204 283018
rect 317604 282698 317786 282934
rect 318022 282698 318204 282934
rect 317604 247254 318204 282698
rect 317604 247018 317786 247254
rect 318022 247018 318204 247254
rect 317604 246934 318204 247018
rect 317604 246698 317786 246934
rect 318022 246698 318204 246934
rect 317604 211254 318204 246698
rect 324804 704838 325404 705780
rect 324804 704602 324986 704838
rect 325222 704602 325404 704838
rect 324804 704518 325404 704602
rect 324804 704282 324986 704518
rect 325222 704282 325404 704518
rect 324804 686454 325404 704282
rect 324804 686218 324986 686454
rect 325222 686218 325404 686454
rect 324804 686134 325404 686218
rect 324804 685898 324986 686134
rect 325222 685898 325404 686134
rect 324804 650454 325404 685898
rect 324804 650218 324986 650454
rect 325222 650218 325404 650454
rect 324804 650134 325404 650218
rect 324804 649898 324986 650134
rect 325222 649898 325404 650134
rect 324804 614454 325404 649898
rect 324804 614218 324986 614454
rect 325222 614218 325404 614454
rect 324804 614134 325404 614218
rect 324804 613898 324986 614134
rect 325222 613898 325404 614134
rect 324804 578454 325404 613898
rect 324804 578218 324986 578454
rect 325222 578218 325404 578454
rect 324804 578134 325404 578218
rect 324804 577898 324986 578134
rect 325222 577898 325404 578134
rect 324804 542454 325404 577898
rect 324804 542218 324986 542454
rect 325222 542218 325404 542454
rect 324804 542134 325404 542218
rect 324804 541898 324986 542134
rect 325222 541898 325404 542134
rect 324804 506454 325404 541898
rect 324804 506218 324986 506454
rect 325222 506218 325404 506454
rect 324804 506134 325404 506218
rect 324804 505898 324986 506134
rect 325222 505898 325404 506134
rect 324804 470454 325404 505898
rect 324804 470218 324986 470454
rect 325222 470218 325404 470454
rect 324804 470134 325404 470218
rect 324804 469898 324986 470134
rect 325222 469898 325404 470134
rect 324804 434454 325404 469898
rect 324804 434218 324986 434454
rect 325222 434218 325404 434454
rect 324804 434134 325404 434218
rect 324804 433898 324986 434134
rect 325222 433898 325404 434134
rect 324804 398454 325404 433898
rect 324804 398218 324986 398454
rect 325222 398218 325404 398454
rect 324804 398134 325404 398218
rect 324804 397898 324986 398134
rect 325222 397898 325404 398134
rect 324804 362454 325404 397898
rect 324804 362218 324986 362454
rect 325222 362218 325404 362454
rect 324804 362134 325404 362218
rect 324804 361898 324986 362134
rect 325222 361898 325404 362134
rect 324804 326454 325404 361898
rect 324804 326218 324986 326454
rect 325222 326218 325404 326454
rect 324804 326134 325404 326218
rect 324804 325898 324986 326134
rect 325222 325898 325404 326134
rect 324804 290454 325404 325898
rect 324804 290218 324986 290454
rect 325222 290218 325404 290454
rect 324804 290134 325404 290218
rect 324804 289898 324986 290134
rect 325222 289898 325404 290134
rect 324804 254454 325404 289898
rect 324804 254218 324986 254454
rect 325222 254218 325404 254454
rect 324804 254134 325404 254218
rect 324804 253898 324986 254134
rect 325222 253898 325404 254134
rect 318747 227900 318813 227901
rect 318747 227836 318748 227900
rect 318812 227836 318813 227900
rect 318747 227835 318813 227836
rect 318750 227629 318810 227835
rect 318747 227628 318813 227629
rect 318747 227564 318748 227628
rect 318812 227564 318813 227628
rect 318747 227563 318813 227564
rect 317604 211018 317786 211254
rect 318022 211018 318204 211254
rect 317604 210934 318204 211018
rect 317604 210698 317786 210934
rect 318022 210698 318204 210934
rect 317604 175254 318204 210698
rect 317604 175018 317786 175254
rect 318022 175018 318204 175254
rect 317604 174934 318204 175018
rect 317604 174698 317786 174934
rect 318022 174698 318204 174934
rect 317604 139254 318204 174698
rect 317604 139018 317786 139254
rect 318022 139018 318204 139254
rect 317604 138934 318204 139018
rect 317604 138698 317786 138934
rect 318022 138698 318204 138934
rect 317604 103254 318204 138698
rect 317604 103018 317786 103254
rect 318022 103018 318204 103254
rect 317604 102934 318204 103018
rect 317604 102698 317786 102934
rect 318022 102698 318204 102934
rect 317604 67254 318204 102698
rect 324804 218454 325404 253898
rect 324804 218218 324986 218454
rect 325222 218218 325404 218454
rect 324804 218134 325404 218218
rect 324804 217898 324986 218134
rect 325222 217898 325404 218134
rect 324804 182454 325404 217898
rect 324804 182218 324986 182454
rect 325222 182218 325404 182454
rect 324804 182134 325404 182218
rect 324804 181898 324986 182134
rect 325222 181898 325404 182134
rect 324804 146454 325404 181898
rect 324804 146218 324986 146454
rect 325222 146218 325404 146454
rect 324804 146134 325404 146218
rect 324804 145898 324986 146134
rect 325222 145898 325404 146134
rect 324804 110454 325404 145898
rect 324804 110218 324986 110454
rect 325222 110218 325404 110454
rect 324804 110134 325404 110218
rect 324804 109898 324986 110134
rect 325222 109898 325404 110134
rect 318747 76124 318813 76125
rect 318747 76060 318748 76124
rect 318812 76060 318813 76124
rect 318747 76059 318813 76060
rect 318750 75853 318810 76059
rect 318747 75852 318813 75853
rect 318747 75788 318748 75852
rect 318812 75788 318813 75852
rect 318747 75787 318813 75788
rect 317604 67018 317786 67254
rect 318022 67018 318204 67254
rect 317604 66934 318204 67018
rect 317604 66698 317786 66934
rect 318022 66698 318204 66934
rect 317604 31254 318204 66698
rect 317604 31018 317786 31254
rect 318022 31018 318204 31254
rect 317604 30934 318204 31018
rect 317604 30698 317786 30934
rect 318022 30698 318204 30934
rect 299604 -6102 299786 -5866
rect 300022 -6102 300204 -5866
rect 299604 -6186 300204 -6102
rect 299604 -6422 299786 -6186
rect 300022 -6422 300204 -6186
rect 299604 -7364 300204 -6422
rect 317604 -6786 318204 30698
rect 324804 74454 325404 109898
rect 324804 74218 324986 74454
rect 325222 74218 325404 74454
rect 324804 74134 325404 74218
rect 324804 73898 324986 74134
rect 325222 73898 325404 74134
rect 324804 38454 325404 73898
rect 324804 38218 324986 38454
rect 325222 38218 325404 38454
rect 324804 38134 325404 38218
rect 324804 37898 324986 38134
rect 325222 37898 325404 38134
rect 324804 2454 325404 37898
rect 324804 2218 324986 2454
rect 325222 2218 325404 2454
rect 324804 2134 325404 2218
rect 324804 1898 324986 2134
rect 325222 1898 325404 2134
rect 324804 -346 325404 1898
rect 324804 -582 324986 -346
rect 325222 -582 325404 -346
rect 324804 -666 325404 -582
rect 324804 -902 324986 -666
rect 325222 -902 325404 -666
rect 324804 -1844 325404 -902
rect 328404 690054 329004 706122
rect 328404 689818 328586 690054
rect 328822 689818 329004 690054
rect 328404 689734 329004 689818
rect 328404 689498 328586 689734
rect 328822 689498 329004 689734
rect 328404 654054 329004 689498
rect 328404 653818 328586 654054
rect 328822 653818 329004 654054
rect 328404 653734 329004 653818
rect 328404 653498 328586 653734
rect 328822 653498 329004 653734
rect 328404 618054 329004 653498
rect 328404 617818 328586 618054
rect 328822 617818 329004 618054
rect 328404 617734 329004 617818
rect 328404 617498 328586 617734
rect 328822 617498 329004 617734
rect 328404 582054 329004 617498
rect 328404 581818 328586 582054
rect 328822 581818 329004 582054
rect 328404 581734 329004 581818
rect 328404 581498 328586 581734
rect 328822 581498 329004 581734
rect 328404 546054 329004 581498
rect 328404 545818 328586 546054
rect 328822 545818 329004 546054
rect 328404 545734 329004 545818
rect 328404 545498 328586 545734
rect 328822 545498 329004 545734
rect 328404 510054 329004 545498
rect 328404 509818 328586 510054
rect 328822 509818 329004 510054
rect 328404 509734 329004 509818
rect 328404 509498 328586 509734
rect 328822 509498 329004 509734
rect 328404 474054 329004 509498
rect 328404 473818 328586 474054
rect 328822 473818 329004 474054
rect 328404 473734 329004 473818
rect 328404 473498 328586 473734
rect 328822 473498 329004 473734
rect 328404 438054 329004 473498
rect 328404 437818 328586 438054
rect 328822 437818 329004 438054
rect 328404 437734 329004 437818
rect 328404 437498 328586 437734
rect 328822 437498 329004 437734
rect 328404 402054 329004 437498
rect 328404 401818 328586 402054
rect 328822 401818 329004 402054
rect 328404 401734 329004 401818
rect 328404 401498 328586 401734
rect 328822 401498 329004 401734
rect 328404 366054 329004 401498
rect 328404 365818 328586 366054
rect 328822 365818 329004 366054
rect 328404 365734 329004 365818
rect 328404 365498 328586 365734
rect 328822 365498 329004 365734
rect 328404 330054 329004 365498
rect 328404 329818 328586 330054
rect 328822 329818 329004 330054
rect 328404 329734 329004 329818
rect 328404 329498 328586 329734
rect 328822 329498 329004 329734
rect 328404 294054 329004 329498
rect 328404 293818 328586 294054
rect 328822 293818 329004 294054
rect 328404 293734 329004 293818
rect 328404 293498 328586 293734
rect 328822 293498 329004 293734
rect 328404 258054 329004 293498
rect 328404 257818 328586 258054
rect 328822 257818 329004 258054
rect 328404 257734 329004 257818
rect 328404 257498 328586 257734
rect 328822 257498 329004 257734
rect 328404 222054 329004 257498
rect 328404 221818 328586 222054
rect 328822 221818 329004 222054
rect 328404 221734 329004 221818
rect 328404 221498 328586 221734
rect 328822 221498 329004 221734
rect 328404 186054 329004 221498
rect 328404 185818 328586 186054
rect 328822 185818 329004 186054
rect 328404 185734 329004 185818
rect 328404 185498 328586 185734
rect 328822 185498 329004 185734
rect 328404 150054 329004 185498
rect 328404 149818 328586 150054
rect 328822 149818 329004 150054
rect 328404 149734 329004 149818
rect 328404 149498 328586 149734
rect 328822 149498 329004 149734
rect 328404 114054 329004 149498
rect 328404 113818 328586 114054
rect 328822 113818 329004 114054
rect 328404 113734 329004 113818
rect 328404 113498 328586 113734
rect 328822 113498 329004 113734
rect 328404 78054 329004 113498
rect 328404 77818 328586 78054
rect 328822 77818 329004 78054
rect 328404 77734 329004 77818
rect 328404 77498 328586 77734
rect 328822 77498 329004 77734
rect 328404 42054 329004 77498
rect 328404 41818 328586 42054
rect 328822 41818 329004 42054
rect 328404 41734 329004 41818
rect 328404 41498 328586 41734
rect 328822 41498 329004 41734
rect 328404 6054 329004 41498
rect 328404 5818 328586 6054
rect 328822 5818 329004 6054
rect 328404 5734 329004 5818
rect 328404 5498 328586 5734
rect 328822 5498 329004 5734
rect 328404 -2186 329004 5498
rect 328404 -2422 328586 -2186
rect 328822 -2422 329004 -2186
rect 328404 -2506 329004 -2422
rect 328404 -2742 328586 -2506
rect 328822 -2742 329004 -2506
rect 328404 -3684 329004 -2742
rect 332004 693654 332604 707962
rect 332004 693418 332186 693654
rect 332422 693418 332604 693654
rect 332004 693334 332604 693418
rect 332004 693098 332186 693334
rect 332422 693098 332604 693334
rect 332004 657654 332604 693098
rect 332004 657418 332186 657654
rect 332422 657418 332604 657654
rect 332004 657334 332604 657418
rect 332004 657098 332186 657334
rect 332422 657098 332604 657334
rect 332004 621654 332604 657098
rect 332004 621418 332186 621654
rect 332422 621418 332604 621654
rect 332004 621334 332604 621418
rect 332004 621098 332186 621334
rect 332422 621098 332604 621334
rect 332004 585654 332604 621098
rect 332004 585418 332186 585654
rect 332422 585418 332604 585654
rect 332004 585334 332604 585418
rect 332004 585098 332186 585334
rect 332422 585098 332604 585334
rect 332004 549654 332604 585098
rect 332004 549418 332186 549654
rect 332422 549418 332604 549654
rect 332004 549334 332604 549418
rect 332004 549098 332186 549334
rect 332422 549098 332604 549334
rect 332004 513654 332604 549098
rect 332004 513418 332186 513654
rect 332422 513418 332604 513654
rect 332004 513334 332604 513418
rect 332004 513098 332186 513334
rect 332422 513098 332604 513334
rect 332004 477654 332604 513098
rect 332004 477418 332186 477654
rect 332422 477418 332604 477654
rect 332004 477334 332604 477418
rect 332004 477098 332186 477334
rect 332422 477098 332604 477334
rect 332004 441654 332604 477098
rect 332004 441418 332186 441654
rect 332422 441418 332604 441654
rect 332004 441334 332604 441418
rect 332004 441098 332186 441334
rect 332422 441098 332604 441334
rect 332004 405654 332604 441098
rect 332004 405418 332186 405654
rect 332422 405418 332604 405654
rect 332004 405334 332604 405418
rect 332004 405098 332186 405334
rect 332422 405098 332604 405334
rect 332004 369654 332604 405098
rect 332004 369418 332186 369654
rect 332422 369418 332604 369654
rect 332004 369334 332604 369418
rect 332004 369098 332186 369334
rect 332422 369098 332604 369334
rect 332004 333654 332604 369098
rect 332004 333418 332186 333654
rect 332422 333418 332604 333654
rect 332004 333334 332604 333418
rect 332004 333098 332186 333334
rect 332422 333098 332604 333334
rect 332004 297654 332604 333098
rect 332004 297418 332186 297654
rect 332422 297418 332604 297654
rect 332004 297334 332604 297418
rect 332004 297098 332186 297334
rect 332422 297098 332604 297334
rect 332004 261654 332604 297098
rect 332004 261418 332186 261654
rect 332422 261418 332604 261654
rect 332004 261334 332604 261418
rect 332004 261098 332186 261334
rect 332422 261098 332604 261334
rect 332004 225654 332604 261098
rect 332004 225418 332186 225654
rect 332422 225418 332604 225654
rect 332004 225334 332604 225418
rect 332004 225098 332186 225334
rect 332422 225098 332604 225334
rect 332004 189654 332604 225098
rect 332004 189418 332186 189654
rect 332422 189418 332604 189654
rect 332004 189334 332604 189418
rect 332004 189098 332186 189334
rect 332422 189098 332604 189334
rect 332004 153654 332604 189098
rect 332004 153418 332186 153654
rect 332422 153418 332604 153654
rect 332004 153334 332604 153418
rect 332004 153098 332186 153334
rect 332422 153098 332604 153334
rect 332004 117654 332604 153098
rect 332004 117418 332186 117654
rect 332422 117418 332604 117654
rect 332004 117334 332604 117418
rect 332004 117098 332186 117334
rect 332422 117098 332604 117334
rect 332004 81654 332604 117098
rect 332004 81418 332186 81654
rect 332422 81418 332604 81654
rect 332004 81334 332604 81418
rect 332004 81098 332186 81334
rect 332422 81098 332604 81334
rect 332004 45654 332604 81098
rect 332004 45418 332186 45654
rect 332422 45418 332604 45654
rect 332004 45334 332604 45418
rect 332004 45098 332186 45334
rect 332422 45098 332604 45334
rect 332004 9654 332604 45098
rect 332004 9418 332186 9654
rect 332422 9418 332604 9654
rect 332004 9334 332604 9418
rect 332004 9098 332186 9334
rect 332422 9098 332604 9334
rect 332004 -4026 332604 9098
rect 332004 -4262 332186 -4026
rect 332422 -4262 332604 -4026
rect 332004 -4346 332604 -4262
rect 332004 -4582 332186 -4346
rect 332422 -4582 332604 -4346
rect 332004 -5524 332604 -4582
rect 335604 697254 336204 709802
rect 353604 711278 354204 711300
rect 353604 711042 353786 711278
rect 354022 711042 354204 711278
rect 353604 710958 354204 711042
rect 353604 710722 353786 710958
rect 354022 710722 354204 710958
rect 350004 709438 350604 709460
rect 350004 709202 350186 709438
rect 350422 709202 350604 709438
rect 350004 709118 350604 709202
rect 350004 708882 350186 709118
rect 350422 708882 350604 709118
rect 346404 707598 347004 707620
rect 346404 707362 346586 707598
rect 346822 707362 347004 707598
rect 346404 707278 347004 707362
rect 346404 707042 346586 707278
rect 346822 707042 347004 707278
rect 335604 697018 335786 697254
rect 336022 697018 336204 697254
rect 335604 696934 336204 697018
rect 335604 696698 335786 696934
rect 336022 696698 336204 696934
rect 335604 661254 336204 696698
rect 335604 661018 335786 661254
rect 336022 661018 336204 661254
rect 335604 660934 336204 661018
rect 335604 660698 335786 660934
rect 336022 660698 336204 660934
rect 335604 625254 336204 660698
rect 335604 625018 335786 625254
rect 336022 625018 336204 625254
rect 335604 624934 336204 625018
rect 335604 624698 335786 624934
rect 336022 624698 336204 624934
rect 335604 589254 336204 624698
rect 335604 589018 335786 589254
rect 336022 589018 336204 589254
rect 335604 588934 336204 589018
rect 335604 588698 335786 588934
rect 336022 588698 336204 588934
rect 335604 553254 336204 588698
rect 335604 553018 335786 553254
rect 336022 553018 336204 553254
rect 335604 552934 336204 553018
rect 335604 552698 335786 552934
rect 336022 552698 336204 552934
rect 335604 517254 336204 552698
rect 335604 517018 335786 517254
rect 336022 517018 336204 517254
rect 335604 516934 336204 517018
rect 335604 516698 335786 516934
rect 336022 516698 336204 516934
rect 335604 481254 336204 516698
rect 335604 481018 335786 481254
rect 336022 481018 336204 481254
rect 335604 480934 336204 481018
rect 335604 480698 335786 480934
rect 336022 480698 336204 480934
rect 335604 445254 336204 480698
rect 335604 445018 335786 445254
rect 336022 445018 336204 445254
rect 335604 444934 336204 445018
rect 335604 444698 335786 444934
rect 336022 444698 336204 444934
rect 335604 409254 336204 444698
rect 335604 409018 335786 409254
rect 336022 409018 336204 409254
rect 335604 408934 336204 409018
rect 335604 408698 335786 408934
rect 336022 408698 336204 408934
rect 335604 373254 336204 408698
rect 335604 373018 335786 373254
rect 336022 373018 336204 373254
rect 335604 372934 336204 373018
rect 335604 372698 335786 372934
rect 336022 372698 336204 372934
rect 335604 337254 336204 372698
rect 335604 337018 335786 337254
rect 336022 337018 336204 337254
rect 335604 336934 336204 337018
rect 335604 336698 335786 336934
rect 336022 336698 336204 336934
rect 335604 301254 336204 336698
rect 335604 301018 335786 301254
rect 336022 301018 336204 301254
rect 335604 300934 336204 301018
rect 335604 300698 335786 300934
rect 336022 300698 336204 300934
rect 335604 265254 336204 300698
rect 335604 265018 335786 265254
rect 336022 265018 336204 265254
rect 335604 264934 336204 265018
rect 335604 264698 335786 264934
rect 336022 264698 336204 264934
rect 335604 229254 336204 264698
rect 335604 229018 335786 229254
rect 336022 229018 336204 229254
rect 335604 228934 336204 229018
rect 335604 228698 335786 228934
rect 336022 228698 336204 228934
rect 335604 193254 336204 228698
rect 342804 705758 343404 705780
rect 342804 705522 342986 705758
rect 343222 705522 343404 705758
rect 342804 705438 343404 705522
rect 342804 705202 342986 705438
rect 343222 705202 343404 705438
rect 342804 668454 343404 705202
rect 342804 668218 342986 668454
rect 343222 668218 343404 668454
rect 342804 668134 343404 668218
rect 342804 667898 342986 668134
rect 343222 667898 343404 668134
rect 342804 632454 343404 667898
rect 342804 632218 342986 632454
rect 343222 632218 343404 632454
rect 342804 632134 343404 632218
rect 342804 631898 342986 632134
rect 343222 631898 343404 632134
rect 342804 596454 343404 631898
rect 342804 596218 342986 596454
rect 343222 596218 343404 596454
rect 342804 596134 343404 596218
rect 342804 595898 342986 596134
rect 343222 595898 343404 596134
rect 342804 560454 343404 595898
rect 342804 560218 342986 560454
rect 343222 560218 343404 560454
rect 342804 560134 343404 560218
rect 342804 559898 342986 560134
rect 343222 559898 343404 560134
rect 342804 524454 343404 559898
rect 342804 524218 342986 524454
rect 343222 524218 343404 524454
rect 342804 524134 343404 524218
rect 342804 523898 342986 524134
rect 343222 523898 343404 524134
rect 342804 488454 343404 523898
rect 342804 488218 342986 488454
rect 343222 488218 343404 488454
rect 342804 488134 343404 488218
rect 342804 487898 342986 488134
rect 343222 487898 343404 488134
rect 342804 452454 343404 487898
rect 342804 452218 342986 452454
rect 343222 452218 343404 452454
rect 342804 452134 343404 452218
rect 342804 451898 342986 452134
rect 343222 451898 343404 452134
rect 342804 416454 343404 451898
rect 342804 416218 342986 416454
rect 343222 416218 343404 416454
rect 342804 416134 343404 416218
rect 342804 415898 342986 416134
rect 343222 415898 343404 416134
rect 342804 380454 343404 415898
rect 342804 380218 342986 380454
rect 343222 380218 343404 380454
rect 342804 380134 343404 380218
rect 342804 379898 342986 380134
rect 343222 379898 343404 380134
rect 342804 344454 343404 379898
rect 342804 344218 342986 344454
rect 343222 344218 343404 344454
rect 342804 344134 343404 344218
rect 342804 343898 342986 344134
rect 343222 343898 343404 344134
rect 342804 308454 343404 343898
rect 342804 308218 342986 308454
rect 343222 308218 343404 308454
rect 342804 308134 343404 308218
rect 342804 307898 342986 308134
rect 343222 307898 343404 308134
rect 342804 272454 343404 307898
rect 342804 272218 342986 272454
rect 343222 272218 343404 272454
rect 342804 272134 343404 272218
rect 342804 271898 342986 272134
rect 343222 271898 343404 272134
rect 342804 236454 343404 271898
rect 342804 236218 342986 236454
rect 343222 236218 343404 236454
rect 342804 236134 343404 236218
rect 342804 235898 342986 236134
rect 343222 235898 343404 236134
rect 338067 228036 338133 228037
rect 338067 227972 338068 228036
rect 338132 227972 338133 228036
rect 338067 227971 338133 227972
rect 338070 227765 338130 227971
rect 338067 227764 338133 227765
rect 338067 227700 338068 227764
rect 338132 227700 338133 227764
rect 338067 227699 338133 227700
rect 335604 193018 335786 193254
rect 336022 193018 336204 193254
rect 335604 192934 336204 193018
rect 335604 192698 335786 192934
rect 336022 192698 336204 192934
rect 335604 157254 336204 192698
rect 335604 157018 335786 157254
rect 336022 157018 336204 157254
rect 335604 156934 336204 157018
rect 335604 156698 335786 156934
rect 336022 156698 336204 156934
rect 335604 121254 336204 156698
rect 335604 121018 335786 121254
rect 336022 121018 336204 121254
rect 335604 120934 336204 121018
rect 335604 120698 335786 120934
rect 336022 120698 336204 120934
rect 335604 85254 336204 120698
rect 335604 85018 335786 85254
rect 336022 85018 336204 85254
rect 335604 84934 336204 85018
rect 335604 84698 335786 84934
rect 336022 84698 336204 84934
rect 335604 49254 336204 84698
rect 342804 200454 343404 235898
rect 342804 200218 342986 200454
rect 343222 200218 343404 200454
rect 342804 200134 343404 200218
rect 342804 199898 342986 200134
rect 343222 199898 343404 200134
rect 342804 164454 343404 199898
rect 342804 164218 342986 164454
rect 343222 164218 343404 164454
rect 342804 164134 343404 164218
rect 342804 163898 342986 164134
rect 343222 163898 343404 164134
rect 342804 128454 343404 163898
rect 342804 128218 342986 128454
rect 343222 128218 343404 128454
rect 342804 128134 343404 128218
rect 342804 127898 342986 128134
rect 343222 127898 343404 128134
rect 342804 92454 343404 127898
rect 342804 92218 342986 92454
rect 343222 92218 343404 92454
rect 342804 92134 343404 92218
rect 342804 91898 342986 92134
rect 343222 91898 343404 92134
rect 338067 76260 338133 76261
rect 338067 76196 338068 76260
rect 338132 76196 338133 76260
rect 338067 76195 338133 76196
rect 338070 75989 338130 76195
rect 338067 75988 338133 75989
rect 338067 75924 338068 75988
rect 338132 75924 338133 75988
rect 338067 75923 338133 75924
rect 335604 49018 335786 49254
rect 336022 49018 336204 49254
rect 335604 48934 336204 49018
rect 335604 48698 335786 48934
rect 336022 48698 336204 48934
rect 335604 13254 336204 48698
rect 335604 13018 335786 13254
rect 336022 13018 336204 13254
rect 335604 12934 336204 13018
rect 335604 12698 335786 12934
rect 336022 12698 336204 12934
rect 317604 -7022 317786 -6786
rect 318022 -7022 318204 -6786
rect 317604 -7106 318204 -7022
rect 317604 -7342 317786 -7106
rect 318022 -7342 318204 -7106
rect 317604 -7364 318204 -7342
rect 335604 -5866 336204 12698
rect 342804 56454 343404 91898
rect 342804 56218 342986 56454
rect 343222 56218 343404 56454
rect 342804 56134 343404 56218
rect 342804 55898 342986 56134
rect 343222 55898 343404 56134
rect 342804 20454 343404 55898
rect 342804 20218 342986 20454
rect 343222 20218 343404 20454
rect 342804 20134 343404 20218
rect 342804 19898 342986 20134
rect 343222 19898 343404 20134
rect 342804 -1266 343404 19898
rect 342804 -1502 342986 -1266
rect 343222 -1502 343404 -1266
rect 342804 -1586 343404 -1502
rect 342804 -1822 342986 -1586
rect 343222 -1822 343404 -1586
rect 342804 -1844 343404 -1822
rect 346404 672054 347004 707042
rect 346404 671818 346586 672054
rect 346822 671818 347004 672054
rect 346404 671734 347004 671818
rect 346404 671498 346586 671734
rect 346822 671498 347004 671734
rect 346404 636054 347004 671498
rect 346404 635818 346586 636054
rect 346822 635818 347004 636054
rect 346404 635734 347004 635818
rect 346404 635498 346586 635734
rect 346822 635498 347004 635734
rect 346404 600054 347004 635498
rect 346404 599818 346586 600054
rect 346822 599818 347004 600054
rect 346404 599734 347004 599818
rect 346404 599498 346586 599734
rect 346822 599498 347004 599734
rect 346404 564054 347004 599498
rect 346404 563818 346586 564054
rect 346822 563818 347004 564054
rect 346404 563734 347004 563818
rect 346404 563498 346586 563734
rect 346822 563498 347004 563734
rect 346404 528054 347004 563498
rect 346404 527818 346586 528054
rect 346822 527818 347004 528054
rect 346404 527734 347004 527818
rect 346404 527498 346586 527734
rect 346822 527498 347004 527734
rect 346404 492054 347004 527498
rect 346404 491818 346586 492054
rect 346822 491818 347004 492054
rect 346404 491734 347004 491818
rect 346404 491498 346586 491734
rect 346822 491498 347004 491734
rect 346404 456054 347004 491498
rect 346404 455818 346586 456054
rect 346822 455818 347004 456054
rect 346404 455734 347004 455818
rect 346404 455498 346586 455734
rect 346822 455498 347004 455734
rect 346404 420054 347004 455498
rect 346404 419818 346586 420054
rect 346822 419818 347004 420054
rect 346404 419734 347004 419818
rect 346404 419498 346586 419734
rect 346822 419498 347004 419734
rect 346404 384054 347004 419498
rect 346404 383818 346586 384054
rect 346822 383818 347004 384054
rect 346404 383734 347004 383818
rect 346404 383498 346586 383734
rect 346822 383498 347004 383734
rect 346404 348054 347004 383498
rect 346404 347818 346586 348054
rect 346822 347818 347004 348054
rect 346404 347734 347004 347818
rect 346404 347498 346586 347734
rect 346822 347498 347004 347734
rect 346404 312054 347004 347498
rect 346404 311818 346586 312054
rect 346822 311818 347004 312054
rect 346404 311734 347004 311818
rect 346404 311498 346586 311734
rect 346822 311498 347004 311734
rect 346404 276054 347004 311498
rect 346404 275818 346586 276054
rect 346822 275818 347004 276054
rect 346404 275734 347004 275818
rect 346404 275498 346586 275734
rect 346822 275498 347004 275734
rect 346404 240054 347004 275498
rect 346404 239818 346586 240054
rect 346822 239818 347004 240054
rect 346404 239734 347004 239818
rect 346404 239498 346586 239734
rect 346822 239498 347004 239734
rect 346404 204054 347004 239498
rect 346404 203818 346586 204054
rect 346822 203818 347004 204054
rect 346404 203734 347004 203818
rect 346404 203498 346586 203734
rect 346822 203498 347004 203734
rect 346404 168054 347004 203498
rect 346404 167818 346586 168054
rect 346822 167818 347004 168054
rect 346404 167734 347004 167818
rect 346404 167498 346586 167734
rect 346822 167498 347004 167734
rect 346404 132054 347004 167498
rect 346404 131818 346586 132054
rect 346822 131818 347004 132054
rect 346404 131734 347004 131818
rect 346404 131498 346586 131734
rect 346822 131498 347004 131734
rect 346404 96054 347004 131498
rect 346404 95818 346586 96054
rect 346822 95818 347004 96054
rect 346404 95734 347004 95818
rect 346404 95498 346586 95734
rect 346822 95498 347004 95734
rect 346404 60054 347004 95498
rect 346404 59818 346586 60054
rect 346822 59818 347004 60054
rect 346404 59734 347004 59818
rect 346404 59498 346586 59734
rect 346822 59498 347004 59734
rect 346404 24054 347004 59498
rect 346404 23818 346586 24054
rect 346822 23818 347004 24054
rect 346404 23734 347004 23818
rect 346404 23498 346586 23734
rect 346822 23498 347004 23734
rect 346404 -3106 347004 23498
rect 346404 -3342 346586 -3106
rect 346822 -3342 347004 -3106
rect 346404 -3426 347004 -3342
rect 346404 -3662 346586 -3426
rect 346822 -3662 347004 -3426
rect 346404 -3684 347004 -3662
rect 350004 675654 350604 708882
rect 350004 675418 350186 675654
rect 350422 675418 350604 675654
rect 350004 675334 350604 675418
rect 350004 675098 350186 675334
rect 350422 675098 350604 675334
rect 350004 639654 350604 675098
rect 350004 639418 350186 639654
rect 350422 639418 350604 639654
rect 350004 639334 350604 639418
rect 350004 639098 350186 639334
rect 350422 639098 350604 639334
rect 350004 603654 350604 639098
rect 350004 603418 350186 603654
rect 350422 603418 350604 603654
rect 350004 603334 350604 603418
rect 350004 603098 350186 603334
rect 350422 603098 350604 603334
rect 350004 567654 350604 603098
rect 350004 567418 350186 567654
rect 350422 567418 350604 567654
rect 350004 567334 350604 567418
rect 350004 567098 350186 567334
rect 350422 567098 350604 567334
rect 350004 531654 350604 567098
rect 350004 531418 350186 531654
rect 350422 531418 350604 531654
rect 350004 531334 350604 531418
rect 350004 531098 350186 531334
rect 350422 531098 350604 531334
rect 350004 495654 350604 531098
rect 350004 495418 350186 495654
rect 350422 495418 350604 495654
rect 350004 495334 350604 495418
rect 350004 495098 350186 495334
rect 350422 495098 350604 495334
rect 350004 459654 350604 495098
rect 350004 459418 350186 459654
rect 350422 459418 350604 459654
rect 350004 459334 350604 459418
rect 350004 459098 350186 459334
rect 350422 459098 350604 459334
rect 350004 423654 350604 459098
rect 350004 423418 350186 423654
rect 350422 423418 350604 423654
rect 350004 423334 350604 423418
rect 350004 423098 350186 423334
rect 350422 423098 350604 423334
rect 350004 387654 350604 423098
rect 350004 387418 350186 387654
rect 350422 387418 350604 387654
rect 350004 387334 350604 387418
rect 350004 387098 350186 387334
rect 350422 387098 350604 387334
rect 350004 351654 350604 387098
rect 350004 351418 350186 351654
rect 350422 351418 350604 351654
rect 350004 351334 350604 351418
rect 350004 351098 350186 351334
rect 350422 351098 350604 351334
rect 350004 315654 350604 351098
rect 350004 315418 350186 315654
rect 350422 315418 350604 315654
rect 350004 315334 350604 315418
rect 350004 315098 350186 315334
rect 350422 315098 350604 315334
rect 350004 279654 350604 315098
rect 350004 279418 350186 279654
rect 350422 279418 350604 279654
rect 350004 279334 350604 279418
rect 350004 279098 350186 279334
rect 350422 279098 350604 279334
rect 350004 243654 350604 279098
rect 350004 243418 350186 243654
rect 350422 243418 350604 243654
rect 350004 243334 350604 243418
rect 350004 243098 350186 243334
rect 350422 243098 350604 243334
rect 350004 207654 350604 243098
rect 350004 207418 350186 207654
rect 350422 207418 350604 207654
rect 350004 207334 350604 207418
rect 350004 207098 350186 207334
rect 350422 207098 350604 207334
rect 350004 171654 350604 207098
rect 350004 171418 350186 171654
rect 350422 171418 350604 171654
rect 350004 171334 350604 171418
rect 350004 171098 350186 171334
rect 350422 171098 350604 171334
rect 350004 135654 350604 171098
rect 350004 135418 350186 135654
rect 350422 135418 350604 135654
rect 350004 135334 350604 135418
rect 350004 135098 350186 135334
rect 350422 135098 350604 135334
rect 350004 99654 350604 135098
rect 350004 99418 350186 99654
rect 350422 99418 350604 99654
rect 350004 99334 350604 99418
rect 350004 99098 350186 99334
rect 350422 99098 350604 99334
rect 350004 63654 350604 99098
rect 350004 63418 350186 63654
rect 350422 63418 350604 63654
rect 350004 63334 350604 63418
rect 350004 63098 350186 63334
rect 350422 63098 350604 63334
rect 350004 27654 350604 63098
rect 350004 27418 350186 27654
rect 350422 27418 350604 27654
rect 350004 27334 350604 27418
rect 350004 27098 350186 27334
rect 350422 27098 350604 27334
rect 350004 -4946 350604 27098
rect 350004 -5182 350186 -4946
rect 350422 -5182 350604 -4946
rect 350004 -5266 350604 -5182
rect 350004 -5502 350186 -5266
rect 350422 -5502 350604 -5266
rect 350004 -5524 350604 -5502
rect 353604 679254 354204 710722
rect 371604 710358 372204 711300
rect 371604 710122 371786 710358
rect 372022 710122 372204 710358
rect 371604 710038 372204 710122
rect 371604 709802 371786 710038
rect 372022 709802 372204 710038
rect 368004 708518 368604 709460
rect 368004 708282 368186 708518
rect 368422 708282 368604 708518
rect 368004 708198 368604 708282
rect 368004 707962 368186 708198
rect 368422 707962 368604 708198
rect 364404 706678 365004 707620
rect 364404 706442 364586 706678
rect 364822 706442 365004 706678
rect 364404 706358 365004 706442
rect 364404 706122 364586 706358
rect 364822 706122 365004 706358
rect 353604 679018 353786 679254
rect 354022 679018 354204 679254
rect 353604 678934 354204 679018
rect 353604 678698 353786 678934
rect 354022 678698 354204 678934
rect 353604 643254 354204 678698
rect 353604 643018 353786 643254
rect 354022 643018 354204 643254
rect 353604 642934 354204 643018
rect 353604 642698 353786 642934
rect 354022 642698 354204 642934
rect 353604 607254 354204 642698
rect 353604 607018 353786 607254
rect 354022 607018 354204 607254
rect 353604 606934 354204 607018
rect 353604 606698 353786 606934
rect 354022 606698 354204 606934
rect 353604 571254 354204 606698
rect 353604 571018 353786 571254
rect 354022 571018 354204 571254
rect 353604 570934 354204 571018
rect 353604 570698 353786 570934
rect 354022 570698 354204 570934
rect 353604 535254 354204 570698
rect 353604 535018 353786 535254
rect 354022 535018 354204 535254
rect 353604 534934 354204 535018
rect 353604 534698 353786 534934
rect 354022 534698 354204 534934
rect 353604 499254 354204 534698
rect 353604 499018 353786 499254
rect 354022 499018 354204 499254
rect 353604 498934 354204 499018
rect 353604 498698 353786 498934
rect 354022 498698 354204 498934
rect 353604 463254 354204 498698
rect 353604 463018 353786 463254
rect 354022 463018 354204 463254
rect 353604 462934 354204 463018
rect 353604 462698 353786 462934
rect 354022 462698 354204 462934
rect 353604 427254 354204 462698
rect 353604 427018 353786 427254
rect 354022 427018 354204 427254
rect 353604 426934 354204 427018
rect 353604 426698 353786 426934
rect 354022 426698 354204 426934
rect 353604 391254 354204 426698
rect 353604 391018 353786 391254
rect 354022 391018 354204 391254
rect 353604 390934 354204 391018
rect 353604 390698 353786 390934
rect 354022 390698 354204 390934
rect 353604 355254 354204 390698
rect 353604 355018 353786 355254
rect 354022 355018 354204 355254
rect 353604 354934 354204 355018
rect 353604 354698 353786 354934
rect 354022 354698 354204 354934
rect 353604 319254 354204 354698
rect 353604 319018 353786 319254
rect 354022 319018 354204 319254
rect 353604 318934 354204 319018
rect 353604 318698 353786 318934
rect 354022 318698 354204 318934
rect 353604 283254 354204 318698
rect 353604 283018 353786 283254
rect 354022 283018 354204 283254
rect 353604 282934 354204 283018
rect 353604 282698 353786 282934
rect 354022 282698 354204 282934
rect 353604 247254 354204 282698
rect 353604 247018 353786 247254
rect 354022 247018 354204 247254
rect 353604 246934 354204 247018
rect 353604 246698 353786 246934
rect 354022 246698 354204 246934
rect 353604 211254 354204 246698
rect 353604 211018 353786 211254
rect 354022 211018 354204 211254
rect 353604 210934 354204 211018
rect 353604 210698 353786 210934
rect 354022 210698 354204 210934
rect 353604 175254 354204 210698
rect 353604 175018 353786 175254
rect 354022 175018 354204 175254
rect 353604 174934 354204 175018
rect 353604 174698 353786 174934
rect 354022 174698 354204 174934
rect 353604 139254 354204 174698
rect 353604 139018 353786 139254
rect 354022 139018 354204 139254
rect 353604 138934 354204 139018
rect 353604 138698 353786 138934
rect 354022 138698 354204 138934
rect 353604 103254 354204 138698
rect 353604 103018 353786 103254
rect 354022 103018 354204 103254
rect 353604 102934 354204 103018
rect 353604 102698 353786 102934
rect 354022 102698 354204 102934
rect 353604 67254 354204 102698
rect 353604 67018 353786 67254
rect 354022 67018 354204 67254
rect 353604 66934 354204 67018
rect 353604 66698 353786 66934
rect 354022 66698 354204 66934
rect 353604 31254 354204 66698
rect 353604 31018 353786 31254
rect 354022 31018 354204 31254
rect 353604 30934 354204 31018
rect 353604 30698 353786 30934
rect 354022 30698 354204 30934
rect 335604 -6102 335786 -5866
rect 336022 -6102 336204 -5866
rect 335604 -6186 336204 -6102
rect 335604 -6422 335786 -6186
rect 336022 -6422 336204 -6186
rect 335604 -7364 336204 -6422
rect 353604 -6786 354204 30698
rect 360804 704838 361404 705780
rect 360804 704602 360986 704838
rect 361222 704602 361404 704838
rect 360804 704518 361404 704602
rect 360804 704282 360986 704518
rect 361222 704282 361404 704518
rect 360804 686454 361404 704282
rect 360804 686218 360986 686454
rect 361222 686218 361404 686454
rect 360804 686134 361404 686218
rect 360804 685898 360986 686134
rect 361222 685898 361404 686134
rect 360804 650454 361404 685898
rect 360804 650218 360986 650454
rect 361222 650218 361404 650454
rect 360804 650134 361404 650218
rect 360804 649898 360986 650134
rect 361222 649898 361404 650134
rect 360804 614454 361404 649898
rect 360804 614218 360986 614454
rect 361222 614218 361404 614454
rect 360804 614134 361404 614218
rect 360804 613898 360986 614134
rect 361222 613898 361404 614134
rect 360804 578454 361404 613898
rect 360804 578218 360986 578454
rect 361222 578218 361404 578454
rect 360804 578134 361404 578218
rect 360804 577898 360986 578134
rect 361222 577898 361404 578134
rect 360804 542454 361404 577898
rect 360804 542218 360986 542454
rect 361222 542218 361404 542454
rect 360804 542134 361404 542218
rect 360804 541898 360986 542134
rect 361222 541898 361404 542134
rect 360804 506454 361404 541898
rect 360804 506218 360986 506454
rect 361222 506218 361404 506454
rect 360804 506134 361404 506218
rect 360804 505898 360986 506134
rect 361222 505898 361404 506134
rect 360804 470454 361404 505898
rect 360804 470218 360986 470454
rect 361222 470218 361404 470454
rect 360804 470134 361404 470218
rect 360804 469898 360986 470134
rect 361222 469898 361404 470134
rect 360804 434454 361404 469898
rect 360804 434218 360986 434454
rect 361222 434218 361404 434454
rect 360804 434134 361404 434218
rect 360804 433898 360986 434134
rect 361222 433898 361404 434134
rect 360804 398454 361404 433898
rect 360804 398218 360986 398454
rect 361222 398218 361404 398454
rect 360804 398134 361404 398218
rect 360804 397898 360986 398134
rect 361222 397898 361404 398134
rect 360804 362454 361404 397898
rect 360804 362218 360986 362454
rect 361222 362218 361404 362454
rect 360804 362134 361404 362218
rect 360804 361898 360986 362134
rect 361222 361898 361404 362134
rect 360804 326454 361404 361898
rect 360804 326218 360986 326454
rect 361222 326218 361404 326454
rect 360804 326134 361404 326218
rect 360804 325898 360986 326134
rect 361222 325898 361404 326134
rect 360804 290454 361404 325898
rect 360804 290218 360986 290454
rect 361222 290218 361404 290454
rect 360804 290134 361404 290218
rect 360804 289898 360986 290134
rect 361222 289898 361404 290134
rect 360804 254454 361404 289898
rect 360804 254218 360986 254454
rect 361222 254218 361404 254454
rect 360804 254134 361404 254218
rect 360804 253898 360986 254134
rect 361222 253898 361404 254134
rect 360804 218454 361404 253898
rect 360804 218218 360986 218454
rect 361222 218218 361404 218454
rect 360804 218134 361404 218218
rect 360804 217898 360986 218134
rect 361222 217898 361404 218134
rect 360804 182454 361404 217898
rect 360804 182218 360986 182454
rect 361222 182218 361404 182454
rect 360804 182134 361404 182218
rect 360804 181898 360986 182134
rect 361222 181898 361404 182134
rect 360804 146454 361404 181898
rect 360804 146218 360986 146454
rect 361222 146218 361404 146454
rect 360804 146134 361404 146218
rect 360804 145898 360986 146134
rect 361222 145898 361404 146134
rect 360804 110454 361404 145898
rect 360804 110218 360986 110454
rect 361222 110218 361404 110454
rect 360804 110134 361404 110218
rect 360804 109898 360986 110134
rect 361222 109898 361404 110134
rect 360804 74454 361404 109898
rect 360804 74218 360986 74454
rect 361222 74218 361404 74454
rect 360804 74134 361404 74218
rect 360804 73898 360986 74134
rect 361222 73898 361404 74134
rect 360804 38454 361404 73898
rect 360804 38218 360986 38454
rect 361222 38218 361404 38454
rect 360804 38134 361404 38218
rect 360804 37898 360986 38134
rect 361222 37898 361404 38134
rect 360804 2454 361404 37898
rect 360804 2218 360986 2454
rect 361222 2218 361404 2454
rect 360804 2134 361404 2218
rect 360804 1898 360986 2134
rect 361222 1898 361404 2134
rect 360804 -346 361404 1898
rect 360804 -582 360986 -346
rect 361222 -582 361404 -346
rect 360804 -666 361404 -582
rect 360804 -902 360986 -666
rect 361222 -902 361404 -666
rect 360804 -1844 361404 -902
rect 364404 690054 365004 706122
rect 364404 689818 364586 690054
rect 364822 689818 365004 690054
rect 364404 689734 365004 689818
rect 364404 689498 364586 689734
rect 364822 689498 365004 689734
rect 364404 654054 365004 689498
rect 364404 653818 364586 654054
rect 364822 653818 365004 654054
rect 364404 653734 365004 653818
rect 364404 653498 364586 653734
rect 364822 653498 365004 653734
rect 364404 618054 365004 653498
rect 364404 617818 364586 618054
rect 364822 617818 365004 618054
rect 364404 617734 365004 617818
rect 364404 617498 364586 617734
rect 364822 617498 365004 617734
rect 364404 582054 365004 617498
rect 364404 581818 364586 582054
rect 364822 581818 365004 582054
rect 364404 581734 365004 581818
rect 364404 581498 364586 581734
rect 364822 581498 365004 581734
rect 364404 546054 365004 581498
rect 364404 545818 364586 546054
rect 364822 545818 365004 546054
rect 364404 545734 365004 545818
rect 364404 545498 364586 545734
rect 364822 545498 365004 545734
rect 364404 510054 365004 545498
rect 364404 509818 364586 510054
rect 364822 509818 365004 510054
rect 364404 509734 365004 509818
rect 364404 509498 364586 509734
rect 364822 509498 365004 509734
rect 364404 474054 365004 509498
rect 364404 473818 364586 474054
rect 364822 473818 365004 474054
rect 364404 473734 365004 473818
rect 364404 473498 364586 473734
rect 364822 473498 365004 473734
rect 364404 438054 365004 473498
rect 364404 437818 364586 438054
rect 364822 437818 365004 438054
rect 364404 437734 365004 437818
rect 364404 437498 364586 437734
rect 364822 437498 365004 437734
rect 364404 402054 365004 437498
rect 364404 401818 364586 402054
rect 364822 401818 365004 402054
rect 364404 401734 365004 401818
rect 364404 401498 364586 401734
rect 364822 401498 365004 401734
rect 364404 366054 365004 401498
rect 364404 365818 364586 366054
rect 364822 365818 365004 366054
rect 364404 365734 365004 365818
rect 364404 365498 364586 365734
rect 364822 365498 365004 365734
rect 364404 330054 365004 365498
rect 364404 329818 364586 330054
rect 364822 329818 365004 330054
rect 364404 329734 365004 329818
rect 364404 329498 364586 329734
rect 364822 329498 365004 329734
rect 364404 294054 365004 329498
rect 364404 293818 364586 294054
rect 364822 293818 365004 294054
rect 364404 293734 365004 293818
rect 364404 293498 364586 293734
rect 364822 293498 365004 293734
rect 364404 258054 365004 293498
rect 364404 257818 364586 258054
rect 364822 257818 365004 258054
rect 364404 257734 365004 257818
rect 364404 257498 364586 257734
rect 364822 257498 365004 257734
rect 364404 222054 365004 257498
rect 364404 221818 364586 222054
rect 364822 221818 365004 222054
rect 364404 221734 365004 221818
rect 364404 221498 364586 221734
rect 364822 221498 365004 221734
rect 364404 186054 365004 221498
rect 364404 185818 364586 186054
rect 364822 185818 365004 186054
rect 364404 185734 365004 185818
rect 364404 185498 364586 185734
rect 364822 185498 365004 185734
rect 364404 150054 365004 185498
rect 364404 149818 364586 150054
rect 364822 149818 365004 150054
rect 364404 149734 365004 149818
rect 364404 149498 364586 149734
rect 364822 149498 365004 149734
rect 364404 114054 365004 149498
rect 364404 113818 364586 114054
rect 364822 113818 365004 114054
rect 364404 113734 365004 113818
rect 364404 113498 364586 113734
rect 364822 113498 365004 113734
rect 364404 78054 365004 113498
rect 364404 77818 364586 78054
rect 364822 77818 365004 78054
rect 364404 77734 365004 77818
rect 364404 77498 364586 77734
rect 364822 77498 365004 77734
rect 364404 42054 365004 77498
rect 364404 41818 364586 42054
rect 364822 41818 365004 42054
rect 364404 41734 365004 41818
rect 364404 41498 364586 41734
rect 364822 41498 365004 41734
rect 364404 6054 365004 41498
rect 364404 5818 364586 6054
rect 364822 5818 365004 6054
rect 364404 5734 365004 5818
rect 364404 5498 364586 5734
rect 364822 5498 365004 5734
rect 364404 -2186 365004 5498
rect 364404 -2422 364586 -2186
rect 364822 -2422 365004 -2186
rect 364404 -2506 365004 -2422
rect 364404 -2742 364586 -2506
rect 364822 -2742 365004 -2506
rect 364404 -3684 365004 -2742
rect 368004 693654 368604 707962
rect 368004 693418 368186 693654
rect 368422 693418 368604 693654
rect 368004 693334 368604 693418
rect 368004 693098 368186 693334
rect 368422 693098 368604 693334
rect 368004 657654 368604 693098
rect 368004 657418 368186 657654
rect 368422 657418 368604 657654
rect 368004 657334 368604 657418
rect 368004 657098 368186 657334
rect 368422 657098 368604 657334
rect 368004 621654 368604 657098
rect 368004 621418 368186 621654
rect 368422 621418 368604 621654
rect 368004 621334 368604 621418
rect 368004 621098 368186 621334
rect 368422 621098 368604 621334
rect 368004 585654 368604 621098
rect 368004 585418 368186 585654
rect 368422 585418 368604 585654
rect 368004 585334 368604 585418
rect 368004 585098 368186 585334
rect 368422 585098 368604 585334
rect 368004 549654 368604 585098
rect 368004 549418 368186 549654
rect 368422 549418 368604 549654
rect 368004 549334 368604 549418
rect 368004 549098 368186 549334
rect 368422 549098 368604 549334
rect 368004 513654 368604 549098
rect 368004 513418 368186 513654
rect 368422 513418 368604 513654
rect 368004 513334 368604 513418
rect 368004 513098 368186 513334
rect 368422 513098 368604 513334
rect 368004 477654 368604 513098
rect 368004 477418 368186 477654
rect 368422 477418 368604 477654
rect 368004 477334 368604 477418
rect 368004 477098 368186 477334
rect 368422 477098 368604 477334
rect 368004 441654 368604 477098
rect 368004 441418 368186 441654
rect 368422 441418 368604 441654
rect 368004 441334 368604 441418
rect 368004 441098 368186 441334
rect 368422 441098 368604 441334
rect 368004 405654 368604 441098
rect 368004 405418 368186 405654
rect 368422 405418 368604 405654
rect 368004 405334 368604 405418
rect 368004 405098 368186 405334
rect 368422 405098 368604 405334
rect 368004 369654 368604 405098
rect 368004 369418 368186 369654
rect 368422 369418 368604 369654
rect 368004 369334 368604 369418
rect 368004 369098 368186 369334
rect 368422 369098 368604 369334
rect 368004 333654 368604 369098
rect 368004 333418 368186 333654
rect 368422 333418 368604 333654
rect 368004 333334 368604 333418
rect 368004 333098 368186 333334
rect 368422 333098 368604 333334
rect 368004 297654 368604 333098
rect 368004 297418 368186 297654
rect 368422 297418 368604 297654
rect 368004 297334 368604 297418
rect 368004 297098 368186 297334
rect 368422 297098 368604 297334
rect 368004 261654 368604 297098
rect 368004 261418 368186 261654
rect 368422 261418 368604 261654
rect 368004 261334 368604 261418
rect 368004 261098 368186 261334
rect 368422 261098 368604 261334
rect 368004 225654 368604 261098
rect 368004 225418 368186 225654
rect 368422 225418 368604 225654
rect 368004 225334 368604 225418
rect 368004 225098 368186 225334
rect 368422 225098 368604 225334
rect 368004 189654 368604 225098
rect 368004 189418 368186 189654
rect 368422 189418 368604 189654
rect 368004 189334 368604 189418
rect 368004 189098 368186 189334
rect 368422 189098 368604 189334
rect 368004 153654 368604 189098
rect 368004 153418 368186 153654
rect 368422 153418 368604 153654
rect 368004 153334 368604 153418
rect 368004 153098 368186 153334
rect 368422 153098 368604 153334
rect 368004 117654 368604 153098
rect 368004 117418 368186 117654
rect 368422 117418 368604 117654
rect 368004 117334 368604 117418
rect 368004 117098 368186 117334
rect 368422 117098 368604 117334
rect 368004 81654 368604 117098
rect 368004 81418 368186 81654
rect 368422 81418 368604 81654
rect 368004 81334 368604 81418
rect 368004 81098 368186 81334
rect 368422 81098 368604 81334
rect 368004 45654 368604 81098
rect 368004 45418 368186 45654
rect 368422 45418 368604 45654
rect 368004 45334 368604 45418
rect 368004 45098 368186 45334
rect 368422 45098 368604 45334
rect 368004 9654 368604 45098
rect 368004 9418 368186 9654
rect 368422 9418 368604 9654
rect 368004 9334 368604 9418
rect 368004 9098 368186 9334
rect 368422 9098 368604 9334
rect 368004 -4026 368604 9098
rect 368004 -4262 368186 -4026
rect 368422 -4262 368604 -4026
rect 368004 -4346 368604 -4262
rect 368004 -4582 368186 -4346
rect 368422 -4582 368604 -4346
rect 368004 -5524 368604 -4582
rect 371604 697254 372204 709802
rect 389604 711278 390204 711300
rect 389604 711042 389786 711278
rect 390022 711042 390204 711278
rect 389604 710958 390204 711042
rect 389604 710722 389786 710958
rect 390022 710722 390204 710958
rect 386004 709438 386604 709460
rect 386004 709202 386186 709438
rect 386422 709202 386604 709438
rect 386004 709118 386604 709202
rect 386004 708882 386186 709118
rect 386422 708882 386604 709118
rect 382404 707598 383004 707620
rect 382404 707362 382586 707598
rect 382822 707362 383004 707598
rect 382404 707278 383004 707362
rect 382404 707042 382586 707278
rect 382822 707042 383004 707278
rect 371604 697018 371786 697254
rect 372022 697018 372204 697254
rect 371604 696934 372204 697018
rect 371604 696698 371786 696934
rect 372022 696698 372204 696934
rect 371604 661254 372204 696698
rect 371604 661018 371786 661254
rect 372022 661018 372204 661254
rect 371604 660934 372204 661018
rect 371604 660698 371786 660934
rect 372022 660698 372204 660934
rect 371604 625254 372204 660698
rect 371604 625018 371786 625254
rect 372022 625018 372204 625254
rect 371604 624934 372204 625018
rect 371604 624698 371786 624934
rect 372022 624698 372204 624934
rect 371604 589254 372204 624698
rect 371604 589018 371786 589254
rect 372022 589018 372204 589254
rect 371604 588934 372204 589018
rect 371604 588698 371786 588934
rect 372022 588698 372204 588934
rect 371604 553254 372204 588698
rect 371604 553018 371786 553254
rect 372022 553018 372204 553254
rect 371604 552934 372204 553018
rect 371604 552698 371786 552934
rect 372022 552698 372204 552934
rect 371604 517254 372204 552698
rect 371604 517018 371786 517254
rect 372022 517018 372204 517254
rect 371604 516934 372204 517018
rect 371604 516698 371786 516934
rect 372022 516698 372204 516934
rect 371604 481254 372204 516698
rect 371604 481018 371786 481254
rect 372022 481018 372204 481254
rect 371604 480934 372204 481018
rect 371604 480698 371786 480934
rect 372022 480698 372204 480934
rect 371604 445254 372204 480698
rect 371604 445018 371786 445254
rect 372022 445018 372204 445254
rect 371604 444934 372204 445018
rect 371604 444698 371786 444934
rect 372022 444698 372204 444934
rect 371604 409254 372204 444698
rect 371604 409018 371786 409254
rect 372022 409018 372204 409254
rect 371604 408934 372204 409018
rect 371604 408698 371786 408934
rect 372022 408698 372204 408934
rect 371604 373254 372204 408698
rect 371604 373018 371786 373254
rect 372022 373018 372204 373254
rect 371604 372934 372204 373018
rect 371604 372698 371786 372934
rect 372022 372698 372204 372934
rect 371604 337254 372204 372698
rect 371604 337018 371786 337254
rect 372022 337018 372204 337254
rect 371604 336934 372204 337018
rect 371604 336698 371786 336934
rect 372022 336698 372204 336934
rect 371604 301254 372204 336698
rect 371604 301018 371786 301254
rect 372022 301018 372204 301254
rect 371604 300934 372204 301018
rect 371604 300698 371786 300934
rect 372022 300698 372204 300934
rect 371604 265254 372204 300698
rect 371604 265018 371786 265254
rect 372022 265018 372204 265254
rect 371604 264934 372204 265018
rect 371604 264698 371786 264934
rect 372022 264698 372204 264934
rect 371604 229254 372204 264698
rect 371604 229018 371786 229254
rect 372022 229018 372204 229254
rect 371604 228934 372204 229018
rect 371604 228698 371786 228934
rect 372022 228698 372204 228934
rect 371604 193254 372204 228698
rect 371604 193018 371786 193254
rect 372022 193018 372204 193254
rect 371604 192934 372204 193018
rect 371604 192698 371786 192934
rect 372022 192698 372204 192934
rect 371604 157254 372204 192698
rect 371604 157018 371786 157254
rect 372022 157018 372204 157254
rect 371604 156934 372204 157018
rect 371604 156698 371786 156934
rect 372022 156698 372204 156934
rect 371604 121254 372204 156698
rect 371604 121018 371786 121254
rect 372022 121018 372204 121254
rect 371604 120934 372204 121018
rect 371604 120698 371786 120934
rect 372022 120698 372204 120934
rect 371604 85254 372204 120698
rect 371604 85018 371786 85254
rect 372022 85018 372204 85254
rect 371604 84934 372204 85018
rect 371604 84698 371786 84934
rect 372022 84698 372204 84934
rect 371604 49254 372204 84698
rect 371604 49018 371786 49254
rect 372022 49018 372204 49254
rect 371604 48934 372204 49018
rect 371604 48698 371786 48934
rect 372022 48698 372204 48934
rect 371604 13254 372204 48698
rect 371604 13018 371786 13254
rect 372022 13018 372204 13254
rect 371604 12934 372204 13018
rect 371604 12698 371786 12934
rect 372022 12698 372204 12934
rect 353604 -7022 353786 -6786
rect 354022 -7022 354204 -6786
rect 353604 -7106 354204 -7022
rect 353604 -7342 353786 -7106
rect 354022 -7342 354204 -7106
rect 353604 -7364 354204 -7342
rect 371604 -5866 372204 12698
rect 378804 705758 379404 705780
rect 378804 705522 378986 705758
rect 379222 705522 379404 705758
rect 378804 705438 379404 705522
rect 378804 705202 378986 705438
rect 379222 705202 379404 705438
rect 378804 668454 379404 705202
rect 378804 668218 378986 668454
rect 379222 668218 379404 668454
rect 378804 668134 379404 668218
rect 378804 667898 378986 668134
rect 379222 667898 379404 668134
rect 378804 632454 379404 667898
rect 378804 632218 378986 632454
rect 379222 632218 379404 632454
rect 378804 632134 379404 632218
rect 378804 631898 378986 632134
rect 379222 631898 379404 632134
rect 378804 596454 379404 631898
rect 378804 596218 378986 596454
rect 379222 596218 379404 596454
rect 378804 596134 379404 596218
rect 378804 595898 378986 596134
rect 379222 595898 379404 596134
rect 378804 560454 379404 595898
rect 378804 560218 378986 560454
rect 379222 560218 379404 560454
rect 378804 560134 379404 560218
rect 378804 559898 378986 560134
rect 379222 559898 379404 560134
rect 378804 524454 379404 559898
rect 378804 524218 378986 524454
rect 379222 524218 379404 524454
rect 378804 524134 379404 524218
rect 378804 523898 378986 524134
rect 379222 523898 379404 524134
rect 378804 488454 379404 523898
rect 378804 488218 378986 488454
rect 379222 488218 379404 488454
rect 378804 488134 379404 488218
rect 378804 487898 378986 488134
rect 379222 487898 379404 488134
rect 378804 452454 379404 487898
rect 378804 452218 378986 452454
rect 379222 452218 379404 452454
rect 378804 452134 379404 452218
rect 378804 451898 378986 452134
rect 379222 451898 379404 452134
rect 378804 416454 379404 451898
rect 378804 416218 378986 416454
rect 379222 416218 379404 416454
rect 378804 416134 379404 416218
rect 378804 415898 378986 416134
rect 379222 415898 379404 416134
rect 378804 380454 379404 415898
rect 378804 380218 378986 380454
rect 379222 380218 379404 380454
rect 378804 380134 379404 380218
rect 378804 379898 378986 380134
rect 379222 379898 379404 380134
rect 378804 344454 379404 379898
rect 378804 344218 378986 344454
rect 379222 344218 379404 344454
rect 378804 344134 379404 344218
rect 378804 343898 378986 344134
rect 379222 343898 379404 344134
rect 378804 308454 379404 343898
rect 378804 308218 378986 308454
rect 379222 308218 379404 308454
rect 378804 308134 379404 308218
rect 378804 307898 378986 308134
rect 379222 307898 379404 308134
rect 378804 272454 379404 307898
rect 378804 272218 378986 272454
rect 379222 272218 379404 272454
rect 378804 272134 379404 272218
rect 378804 271898 378986 272134
rect 379222 271898 379404 272134
rect 378804 236454 379404 271898
rect 378804 236218 378986 236454
rect 379222 236218 379404 236454
rect 378804 236134 379404 236218
rect 378804 235898 378986 236134
rect 379222 235898 379404 236134
rect 378804 200454 379404 235898
rect 378804 200218 378986 200454
rect 379222 200218 379404 200454
rect 378804 200134 379404 200218
rect 378804 199898 378986 200134
rect 379222 199898 379404 200134
rect 378804 164454 379404 199898
rect 378804 164218 378986 164454
rect 379222 164218 379404 164454
rect 378804 164134 379404 164218
rect 378804 163898 378986 164134
rect 379222 163898 379404 164134
rect 378804 128454 379404 163898
rect 378804 128218 378986 128454
rect 379222 128218 379404 128454
rect 378804 128134 379404 128218
rect 378804 127898 378986 128134
rect 379222 127898 379404 128134
rect 378804 92454 379404 127898
rect 378804 92218 378986 92454
rect 379222 92218 379404 92454
rect 378804 92134 379404 92218
rect 378804 91898 378986 92134
rect 379222 91898 379404 92134
rect 378804 56454 379404 91898
rect 378804 56218 378986 56454
rect 379222 56218 379404 56454
rect 378804 56134 379404 56218
rect 378804 55898 378986 56134
rect 379222 55898 379404 56134
rect 378804 20454 379404 55898
rect 378804 20218 378986 20454
rect 379222 20218 379404 20454
rect 378804 20134 379404 20218
rect 378804 19898 378986 20134
rect 379222 19898 379404 20134
rect 378804 -1266 379404 19898
rect 378804 -1502 378986 -1266
rect 379222 -1502 379404 -1266
rect 378804 -1586 379404 -1502
rect 378804 -1822 378986 -1586
rect 379222 -1822 379404 -1586
rect 378804 -1844 379404 -1822
rect 382404 672054 383004 707042
rect 382404 671818 382586 672054
rect 382822 671818 383004 672054
rect 382404 671734 383004 671818
rect 382404 671498 382586 671734
rect 382822 671498 383004 671734
rect 382404 636054 383004 671498
rect 382404 635818 382586 636054
rect 382822 635818 383004 636054
rect 382404 635734 383004 635818
rect 382404 635498 382586 635734
rect 382822 635498 383004 635734
rect 382404 600054 383004 635498
rect 382404 599818 382586 600054
rect 382822 599818 383004 600054
rect 382404 599734 383004 599818
rect 382404 599498 382586 599734
rect 382822 599498 383004 599734
rect 382404 564054 383004 599498
rect 382404 563818 382586 564054
rect 382822 563818 383004 564054
rect 382404 563734 383004 563818
rect 382404 563498 382586 563734
rect 382822 563498 383004 563734
rect 382404 528054 383004 563498
rect 382404 527818 382586 528054
rect 382822 527818 383004 528054
rect 382404 527734 383004 527818
rect 382404 527498 382586 527734
rect 382822 527498 383004 527734
rect 382404 492054 383004 527498
rect 382404 491818 382586 492054
rect 382822 491818 383004 492054
rect 382404 491734 383004 491818
rect 382404 491498 382586 491734
rect 382822 491498 383004 491734
rect 382404 456054 383004 491498
rect 382404 455818 382586 456054
rect 382822 455818 383004 456054
rect 382404 455734 383004 455818
rect 382404 455498 382586 455734
rect 382822 455498 383004 455734
rect 382404 420054 383004 455498
rect 382404 419818 382586 420054
rect 382822 419818 383004 420054
rect 382404 419734 383004 419818
rect 382404 419498 382586 419734
rect 382822 419498 383004 419734
rect 382404 384054 383004 419498
rect 382404 383818 382586 384054
rect 382822 383818 383004 384054
rect 382404 383734 383004 383818
rect 382404 383498 382586 383734
rect 382822 383498 383004 383734
rect 382404 348054 383004 383498
rect 382404 347818 382586 348054
rect 382822 347818 383004 348054
rect 382404 347734 383004 347818
rect 382404 347498 382586 347734
rect 382822 347498 383004 347734
rect 382404 312054 383004 347498
rect 382404 311818 382586 312054
rect 382822 311818 383004 312054
rect 382404 311734 383004 311818
rect 382404 311498 382586 311734
rect 382822 311498 383004 311734
rect 382404 276054 383004 311498
rect 382404 275818 382586 276054
rect 382822 275818 383004 276054
rect 382404 275734 383004 275818
rect 382404 275498 382586 275734
rect 382822 275498 383004 275734
rect 382404 240054 383004 275498
rect 382404 239818 382586 240054
rect 382822 239818 383004 240054
rect 382404 239734 383004 239818
rect 382404 239498 382586 239734
rect 382822 239498 383004 239734
rect 382404 204054 383004 239498
rect 382404 203818 382586 204054
rect 382822 203818 383004 204054
rect 382404 203734 383004 203818
rect 382404 203498 382586 203734
rect 382822 203498 383004 203734
rect 382404 168054 383004 203498
rect 382404 167818 382586 168054
rect 382822 167818 383004 168054
rect 382404 167734 383004 167818
rect 382404 167498 382586 167734
rect 382822 167498 383004 167734
rect 382404 132054 383004 167498
rect 382404 131818 382586 132054
rect 382822 131818 383004 132054
rect 382404 131734 383004 131818
rect 382404 131498 382586 131734
rect 382822 131498 383004 131734
rect 382404 96054 383004 131498
rect 382404 95818 382586 96054
rect 382822 95818 383004 96054
rect 382404 95734 383004 95818
rect 382404 95498 382586 95734
rect 382822 95498 383004 95734
rect 382404 60054 383004 95498
rect 382404 59818 382586 60054
rect 382822 59818 383004 60054
rect 382404 59734 383004 59818
rect 382404 59498 382586 59734
rect 382822 59498 383004 59734
rect 382404 24054 383004 59498
rect 382404 23818 382586 24054
rect 382822 23818 383004 24054
rect 382404 23734 383004 23818
rect 382404 23498 382586 23734
rect 382822 23498 383004 23734
rect 382404 -3106 383004 23498
rect 382404 -3342 382586 -3106
rect 382822 -3342 383004 -3106
rect 382404 -3426 383004 -3342
rect 382404 -3662 382586 -3426
rect 382822 -3662 383004 -3426
rect 382404 -3684 383004 -3662
rect 386004 675654 386604 708882
rect 386004 675418 386186 675654
rect 386422 675418 386604 675654
rect 386004 675334 386604 675418
rect 386004 675098 386186 675334
rect 386422 675098 386604 675334
rect 386004 639654 386604 675098
rect 386004 639418 386186 639654
rect 386422 639418 386604 639654
rect 386004 639334 386604 639418
rect 386004 639098 386186 639334
rect 386422 639098 386604 639334
rect 386004 603654 386604 639098
rect 386004 603418 386186 603654
rect 386422 603418 386604 603654
rect 386004 603334 386604 603418
rect 386004 603098 386186 603334
rect 386422 603098 386604 603334
rect 386004 567654 386604 603098
rect 386004 567418 386186 567654
rect 386422 567418 386604 567654
rect 386004 567334 386604 567418
rect 386004 567098 386186 567334
rect 386422 567098 386604 567334
rect 386004 531654 386604 567098
rect 386004 531418 386186 531654
rect 386422 531418 386604 531654
rect 386004 531334 386604 531418
rect 386004 531098 386186 531334
rect 386422 531098 386604 531334
rect 386004 495654 386604 531098
rect 386004 495418 386186 495654
rect 386422 495418 386604 495654
rect 386004 495334 386604 495418
rect 386004 495098 386186 495334
rect 386422 495098 386604 495334
rect 386004 459654 386604 495098
rect 386004 459418 386186 459654
rect 386422 459418 386604 459654
rect 386004 459334 386604 459418
rect 386004 459098 386186 459334
rect 386422 459098 386604 459334
rect 386004 423654 386604 459098
rect 386004 423418 386186 423654
rect 386422 423418 386604 423654
rect 386004 423334 386604 423418
rect 386004 423098 386186 423334
rect 386422 423098 386604 423334
rect 386004 387654 386604 423098
rect 386004 387418 386186 387654
rect 386422 387418 386604 387654
rect 386004 387334 386604 387418
rect 386004 387098 386186 387334
rect 386422 387098 386604 387334
rect 386004 351654 386604 387098
rect 386004 351418 386186 351654
rect 386422 351418 386604 351654
rect 386004 351334 386604 351418
rect 386004 351098 386186 351334
rect 386422 351098 386604 351334
rect 386004 315654 386604 351098
rect 386004 315418 386186 315654
rect 386422 315418 386604 315654
rect 386004 315334 386604 315418
rect 386004 315098 386186 315334
rect 386422 315098 386604 315334
rect 386004 279654 386604 315098
rect 386004 279418 386186 279654
rect 386422 279418 386604 279654
rect 386004 279334 386604 279418
rect 386004 279098 386186 279334
rect 386422 279098 386604 279334
rect 386004 243654 386604 279098
rect 386004 243418 386186 243654
rect 386422 243418 386604 243654
rect 386004 243334 386604 243418
rect 386004 243098 386186 243334
rect 386422 243098 386604 243334
rect 386004 207654 386604 243098
rect 386004 207418 386186 207654
rect 386422 207418 386604 207654
rect 386004 207334 386604 207418
rect 386004 207098 386186 207334
rect 386422 207098 386604 207334
rect 386004 171654 386604 207098
rect 386004 171418 386186 171654
rect 386422 171418 386604 171654
rect 386004 171334 386604 171418
rect 386004 171098 386186 171334
rect 386422 171098 386604 171334
rect 386004 135654 386604 171098
rect 386004 135418 386186 135654
rect 386422 135418 386604 135654
rect 386004 135334 386604 135418
rect 386004 135098 386186 135334
rect 386422 135098 386604 135334
rect 386004 99654 386604 135098
rect 386004 99418 386186 99654
rect 386422 99418 386604 99654
rect 386004 99334 386604 99418
rect 386004 99098 386186 99334
rect 386422 99098 386604 99334
rect 386004 63654 386604 99098
rect 386004 63418 386186 63654
rect 386422 63418 386604 63654
rect 386004 63334 386604 63418
rect 386004 63098 386186 63334
rect 386422 63098 386604 63334
rect 386004 27654 386604 63098
rect 386004 27418 386186 27654
rect 386422 27418 386604 27654
rect 386004 27334 386604 27418
rect 386004 27098 386186 27334
rect 386422 27098 386604 27334
rect 386004 -4946 386604 27098
rect 386004 -5182 386186 -4946
rect 386422 -5182 386604 -4946
rect 386004 -5266 386604 -5182
rect 386004 -5502 386186 -5266
rect 386422 -5502 386604 -5266
rect 386004 -5524 386604 -5502
rect 389604 679254 390204 710722
rect 407604 710358 408204 711300
rect 407604 710122 407786 710358
rect 408022 710122 408204 710358
rect 407604 710038 408204 710122
rect 407604 709802 407786 710038
rect 408022 709802 408204 710038
rect 404004 708518 404604 709460
rect 404004 708282 404186 708518
rect 404422 708282 404604 708518
rect 404004 708198 404604 708282
rect 404004 707962 404186 708198
rect 404422 707962 404604 708198
rect 400404 706678 401004 707620
rect 400404 706442 400586 706678
rect 400822 706442 401004 706678
rect 400404 706358 401004 706442
rect 400404 706122 400586 706358
rect 400822 706122 401004 706358
rect 389604 679018 389786 679254
rect 390022 679018 390204 679254
rect 389604 678934 390204 679018
rect 389604 678698 389786 678934
rect 390022 678698 390204 678934
rect 389604 643254 390204 678698
rect 389604 643018 389786 643254
rect 390022 643018 390204 643254
rect 389604 642934 390204 643018
rect 389604 642698 389786 642934
rect 390022 642698 390204 642934
rect 389604 607254 390204 642698
rect 389604 607018 389786 607254
rect 390022 607018 390204 607254
rect 389604 606934 390204 607018
rect 389604 606698 389786 606934
rect 390022 606698 390204 606934
rect 389604 571254 390204 606698
rect 389604 571018 389786 571254
rect 390022 571018 390204 571254
rect 389604 570934 390204 571018
rect 389604 570698 389786 570934
rect 390022 570698 390204 570934
rect 389604 535254 390204 570698
rect 389604 535018 389786 535254
rect 390022 535018 390204 535254
rect 389604 534934 390204 535018
rect 389604 534698 389786 534934
rect 390022 534698 390204 534934
rect 389604 499254 390204 534698
rect 389604 499018 389786 499254
rect 390022 499018 390204 499254
rect 389604 498934 390204 499018
rect 389604 498698 389786 498934
rect 390022 498698 390204 498934
rect 389604 463254 390204 498698
rect 389604 463018 389786 463254
rect 390022 463018 390204 463254
rect 389604 462934 390204 463018
rect 389604 462698 389786 462934
rect 390022 462698 390204 462934
rect 389604 427254 390204 462698
rect 389604 427018 389786 427254
rect 390022 427018 390204 427254
rect 389604 426934 390204 427018
rect 389604 426698 389786 426934
rect 390022 426698 390204 426934
rect 389604 391254 390204 426698
rect 389604 391018 389786 391254
rect 390022 391018 390204 391254
rect 389604 390934 390204 391018
rect 389604 390698 389786 390934
rect 390022 390698 390204 390934
rect 389604 355254 390204 390698
rect 389604 355018 389786 355254
rect 390022 355018 390204 355254
rect 389604 354934 390204 355018
rect 389604 354698 389786 354934
rect 390022 354698 390204 354934
rect 389604 319254 390204 354698
rect 389604 319018 389786 319254
rect 390022 319018 390204 319254
rect 389604 318934 390204 319018
rect 389604 318698 389786 318934
rect 390022 318698 390204 318934
rect 389604 283254 390204 318698
rect 389604 283018 389786 283254
rect 390022 283018 390204 283254
rect 389604 282934 390204 283018
rect 389604 282698 389786 282934
rect 390022 282698 390204 282934
rect 389604 247254 390204 282698
rect 389604 247018 389786 247254
rect 390022 247018 390204 247254
rect 389604 246934 390204 247018
rect 389604 246698 389786 246934
rect 390022 246698 390204 246934
rect 389604 211254 390204 246698
rect 389604 211018 389786 211254
rect 390022 211018 390204 211254
rect 389604 210934 390204 211018
rect 389604 210698 389786 210934
rect 390022 210698 390204 210934
rect 389604 175254 390204 210698
rect 389604 175018 389786 175254
rect 390022 175018 390204 175254
rect 389604 174934 390204 175018
rect 389604 174698 389786 174934
rect 390022 174698 390204 174934
rect 389604 139254 390204 174698
rect 389604 139018 389786 139254
rect 390022 139018 390204 139254
rect 389604 138934 390204 139018
rect 389604 138698 389786 138934
rect 390022 138698 390204 138934
rect 389604 103254 390204 138698
rect 389604 103018 389786 103254
rect 390022 103018 390204 103254
rect 389604 102934 390204 103018
rect 389604 102698 389786 102934
rect 390022 102698 390204 102934
rect 389604 67254 390204 102698
rect 389604 67018 389786 67254
rect 390022 67018 390204 67254
rect 389604 66934 390204 67018
rect 389604 66698 389786 66934
rect 390022 66698 390204 66934
rect 389604 31254 390204 66698
rect 389604 31018 389786 31254
rect 390022 31018 390204 31254
rect 389604 30934 390204 31018
rect 389604 30698 389786 30934
rect 390022 30698 390204 30934
rect 371604 -6102 371786 -5866
rect 372022 -6102 372204 -5866
rect 371604 -6186 372204 -6102
rect 371604 -6422 371786 -6186
rect 372022 -6422 372204 -6186
rect 371604 -7364 372204 -6422
rect 389604 -6786 390204 30698
rect 396804 704838 397404 705780
rect 396804 704602 396986 704838
rect 397222 704602 397404 704838
rect 396804 704518 397404 704602
rect 396804 704282 396986 704518
rect 397222 704282 397404 704518
rect 396804 686454 397404 704282
rect 396804 686218 396986 686454
rect 397222 686218 397404 686454
rect 396804 686134 397404 686218
rect 396804 685898 396986 686134
rect 397222 685898 397404 686134
rect 396804 650454 397404 685898
rect 396804 650218 396986 650454
rect 397222 650218 397404 650454
rect 396804 650134 397404 650218
rect 396804 649898 396986 650134
rect 397222 649898 397404 650134
rect 396804 614454 397404 649898
rect 396804 614218 396986 614454
rect 397222 614218 397404 614454
rect 396804 614134 397404 614218
rect 396804 613898 396986 614134
rect 397222 613898 397404 614134
rect 396804 578454 397404 613898
rect 396804 578218 396986 578454
rect 397222 578218 397404 578454
rect 396804 578134 397404 578218
rect 396804 577898 396986 578134
rect 397222 577898 397404 578134
rect 396804 542454 397404 577898
rect 396804 542218 396986 542454
rect 397222 542218 397404 542454
rect 396804 542134 397404 542218
rect 396804 541898 396986 542134
rect 397222 541898 397404 542134
rect 396804 506454 397404 541898
rect 396804 506218 396986 506454
rect 397222 506218 397404 506454
rect 396804 506134 397404 506218
rect 396804 505898 396986 506134
rect 397222 505898 397404 506134
rect 396804 470454 397404 505898
rect 396804 470218 396986 470454
rect 397222 470218 397404 470454
rect 396804 470134 397404 470218
rect 396804 469898 396986 470134
rect 397222 469898 397404 470134
rect 396804 434454 397404 469898
rect 396804 434218 396986 434454
rect 397222 434218 397404 434454
rect 396804 434134 397404 434218
rect 396804 433898 396986 434134
rect 397222 433898 397404 434134
rect 396804 398454 397404 433898
rect 396804 398218 396986 398454
rect 397222 398218 397404 398454
rect 396804 398134 397404 398218
rect 396804 397898 396986 398134
rect 397222 397898 397404 398134
rect 396804 362454 397404 397898
rect 396804 362218 396986 362454
rect 397222 362218 397404 362454
rect 396804 362134 397404 362218
rect 396804 361898 396986 362134
rect 397222 361898 397404 362134
rect 396804 326454 397404 361898
rect 396804 326218 396986 326454
rect 397222 326218 397404 326454
rect 396804 326134 397404 326218
rect 396804 325898 396986 326134
rect 397222 325898 397404 326134
rect 396804 290454 397404 325898
rect 396804 290218 396986 290454
rect 397222 290218 397404 290454
rect 396804 290134 397404 290218
rect 396804 289898 396986 290134
rect 397222 289898 397404 290134
rect 396804 254454 397404 289898
rect 396804 254218 396986 254454
rect 397222 254218 397404 254454
rect 396804 254134 397404 254218
rect 396804 253898 396986 254134
rect 397222 253898 397404 254134
rect 396804 218454 397404 253898
rect 396804 218218 396986 218454
rect 397222 218218 397404 218454
rect 396804 218134 397404 218218
rect 396804 217898 396986 218134
rect 397222 217898 397404 218134
rect 396804 182454 397404 217898
rect 396804 182218 396986 182454
rect 397222 182218 397404 182454
rect 396804 182134 397404 182218
rect 396804 181898 396986 182134
rect 397222 181898 397404 182134
rect 396804 146454 397404 181898
rect 396804 146218 396986 146454
rect 397222 146218 397404 146454
rect 396804 146134 397404 146218
rect 396804 145898 396986 146134
rect 397222 145898 397404 146134
rect 396804 110454 397404 145898
rect 396804 110218 396986 110454
rect 397222 110218 397404 110454
rect 396804 110134 397404 110218
rect 396804 109898 396986 110134
rect 397222 109898 397404 110134
rect 396804 74454 397404 109898
rect 396804 74218 396986 74454
rect 397222 74218 397404 74454
rect 396804 74134 397404 74218
rect 396804 73898 396986 74134
rect 397222 73898 397404 74134
rect 396804 38454 397404 73898
rect 396804 38218 396986 38454
rect 397222 38218 397404 38454
rect 396804 38134 397404 38218
rect 396804 37898 396986 38134
rect 397222 37898 397404 38134
rect 396804 2454 397404 37898
rect 396804 2218 396986 2454
rect 397222 2218 397404 2454
rect 396804 2134 397404 2218
rect 396804 1898 396986 2134
rect 397222 1898 397404 2134
rect 396804 -346 397404 1898
rect 396804 -582 396986 -346
rect 397222 -582 397404 -346
rect 396804 -666 397404 -582
rect 396804 -902 396986 -666
rect 397222 -902 397404 -666
rect 396804 -1844 397404 -902
rect 400404 690054 401004 706122
rect 400404 689818 400586 690054
rect 400822 689818 401004 690054
rect 400404 689734 401004 689818
rect 400404 689498 400586 689734
rect 400822 689498 401004 689734
rect 400404 654054 401004 689498
rect 400404 653818 400586 654054
rect 400822 653818 401004 654054
rect 400404 653734 401004 653818
rect 400404 653498 400586 653734
rect 400822 653498 401004 653734
rect 400404 618054 401004 653498
rect 400404 617818 400586 618054
rect 400822 617818 401004 618054
rect 400404 617734 401004 617818
rect 400404 617498 400586 617734
rect 400822 617498 401004 617734
rect 400404 582054 401004 617498
rect 400404 581818 400586 582054
rect 400822 581818 401004 582054
rect 400404 581734 401004 581818
rect 400404 581498 400586 581734
rect 400822 581498 401004 581734
rect 400404 546054 401004 581498
rect 400404 545818 400586 546054
rect 400822 545818 401004 546054
rect 400404 545734 401004 545818
rect 400404 545498 400586 545734
rect 400822 545498 401004 545734
rect 400404 510054 401004 545498
rect 400404 509818 400586 510054
rect 400822 509818 401004 510054
rect 400404 509734 401004 509818
rect 400404 509498 400586 509734
rect 400822 509498 401004 509734
rect 400404 474054 401004 509498
rect 400404 473818 400586 474054
rect 400822 473818 401004 474054
rect 400404 473734 401004 473818
rect 400404 473498 400586 473734
rect 400822 473498 401004 473734
rect 400404 438054 401004 473498
rect 400404 437818 400586 438054
rect 400822 437818 401004 438054
rect 400404 437734 401004 437818
rect 400404 437498 400586 437734
rect 400822 437498 401004 437734
rect 400404 402054 401004 437498
rect 400404 401818 400586 402054
rect 400822 401818 401004 402054
rect 400404 401734 401004 401818
rect 400404 401498 400586 401734
rect 400822 401498 401004 401734
rect 400404 366054 401004 401498
rect 400404 365818 400586 366054
rect 400822 365818 401004 366054
rect 400404 365734 401004 365818
rect 400404 365498 400586 365734
rect 400822 365498 401004 365734
rect 400404 330054 401004 365498
rect 400404 329818 400586 330054
rect 400822 329818 401004 330054
rect 400404 329734 401004 329818
rect 400404 329498 400586 329734
rect 400822 329498 401004 329734
rect 400404 294054 401004 329498
rect 400404 293818 400586 294054
rect 400822 293818 401004 294054
rect 400404 293734 401004 293818
rect 400404 293498 400586 293734
rect 400822 293498 401004 293734
rect 400404 258054 401004 293498
rect 400404 257818 400586 258054
rect 400822 257818 401004 258054
rect 400404 257734 401004 257818
rect 400404 257498 400586 257734
rect 400822 257498 401004 257734
rect 400404 222054 401004 257498
rect 400404 221818 400586 222054
rect 400822 221818 401004 222054
rect 400404 221734 401004 221818
rect 400404 221498 400586 221734
rect 400822 221498 401004 221734
rect 400404 186054 401004 221498
rect 400404 185818 400586 186054
rect 400822 185818 401004 186054
rect 400404 185734 401004 185818
rect 400404 185498 400586 185734
rect 400822 185498 401004 185734
rect 400404 150054 401004 185498
rect 400404 149818 400586 150054
rect 400822 149818 401004 150054
rect 400404 149734 401004 149818
rect 400404 149498 400586 149734
rect 400822 149498 401004 149734
rect 400404 114054 401004 149498
rect 400404 113818 400586 114054
rect 400822 113818 401004 114054
rect 400404 113734 401004 113818
rect 400404 113498 400586 113734
rect 400822 113498 401004 113734
rect 400404 78054 401004 113498
rect 400404 77818 400586 78054
rect 400822 77818 401004 78054
rect 400404 77734 401004 77818
rect 400404 77498 400586 77734
rect 400822 77498 401004 77734
rect 400404 42054 401004 77498
rect 400404 41818 400586 42054
rect 400822 41818 401004 42054
rect 400404 41734 401004 41818
rect 400404 41498 400586 41734
rect 400822 41498 401004 41734
rect 400404 6054 401004 41498
rect 400404 5818 400586 6054
rect 400822 5818 401004 6054
rect 400404 5734 401004 5818
rect 400404 5498 400586 5734
rect 400822 5498 401004 5734
rect 400404 -2186 401004 5498
rect 400404 -2422 400586 -2186
rect 400822 -2422 401004 -2186
rect 400404 -2506 401004 -2422
rect 400404 -2742 400586 -2506
rect 400822 -2742 401004 -2506
rect 400404 -3684 401004 -2742
rect 404004 693654 404604 707962
rect 404004 693418 404186 693654
rect 404422 693418 404604 693654
rect 404004 693334 404604 693418
rect 404004 693098 404186 693334
rect 404422 693098 404604 693334
rect 404004 657654 404604 693098
rect 404004 657418 404186 657654
rect 404422 657418 404604 657654
rect 404004 657334 404604 657418
rect 404004 657098 404186 657334
rect 404422 657098 404604 657334
rect 404004 621654 404604 657098
rect 404004 621418 404186 621654
rect 404422 621418 404604 621654
rect 404004 621334 404604 621418
rect 404004 621098 404186 621334
rect 404422 621098 404604 621334
rect 404004 585654 404604 621098
rect 404004 585418 404186 585654
rect 404422 585418 404604 585654
rect 404004 585334 404604 585418
rect 404004 585098 404186 585334
rect 404422 585098 404604 585334
rect 404004 549654 404604 585098
rect 404004 549418 404186 549654
rect 404422 549418 404604 549654
rect 404004 549334 404604 549418
rect 404004 549098 404186 549334
rect 404422 549098 404604 549334
rect 404004 513654 404604 549098
rect 404004 513418 404186 513654
rect 404422 513418 404604 513654
rect 404004 513334 404604 513418
rect 404004 513098 404186 513334
rect 404422 513098 404604 513334
rect 404004 477654 404604 513098
rect 404004 477418 404186 477654
rect 404422 477418 404604 477654
rect 404004 477334 404604 477418
rect 404004 477098 404186 477334
rect 404422 477098 404604 477334
rect 404004 441654 404604 477098
rect 404004 441418 404186 441654
rect 404422 441418 404604 441654
rect 404004 441334 404604 441418
rect 404004 441098 404186 441334
rect 404422 441098 404604 441334
rect 404004 405654 404604 441098
rect 404004 405418 404186 405654
rect 404422 405418 404604 405654
rect 404004 405334 404604 405418
rect 404004 405098 404186 405334
rect 404422 405098 404604 405334
rect 404004 369654 404604 405098
rect 404004 369418 404186 369654
rect 404422 369418 404604 369654
rect 404004 369334 404604 369418
rect 404004 369098 404186 369334
rect 404422 369098 404604 369334
rect 404004 333654 404604 369098
rect 404004 333418 404186 333654
rect 404422 333418 404604 333654
rect 404004 333334 404604 333418
rect 404004 333098 404186 333334
rect 404422 333098 404604 333334
rect 404004 297654 404604 333098
rect 404004 297418 404186 297654
rect 404422 297418 404604 297654
rect 404004 297334 404604 297418
rect 404004 297098 404186 297334
rect 404422 297098 404604 297334
rect 404004 261654 404604 297098
rect 404004 261418 404186 261654
rect 404422 261418 404604 261654
rect 404004 261334 404604 261418
rect 404004 261098 404186 261334
rect 404422 261098 404604 261334
rect 404004 225654 404604 261098
rect 404004 225418 404186 225654
rect 404422 225418 404604 225654
rect 404004 225334 404604 225418
rect 404004 225098 404186 225334
rect 404422 225098 404604 225334
rect 404004 189654 404604 225098
rect 404004 189418 404186 189654
rect 404422 189418 404604 189654
rect 404004 189334 404604 189418
rect 404004 189098 404186 189334
rect 404422 189098 404604 189334
rect 404004 153654 404604 189098
rect 404004 153418 404186 153654
rect 404422 153418 404604 153654
rect 404004 153334 404604 153418
rect 404004 153098 404186 153334
rect 404422 153098 404604 153334
rect 404004 117654 404604 153098
rect 404004 117418 404186 117654
rect 404422 117418 404604 117654
rect 404004 117334 404604 117418
rect 404004 117098 404186 117334
rect 404422 117098 404604 117334
rect 404004 81654 404604 117098
rect 404004 81418 404186 81654
rect 404422 81418 404604 81654
rect 404004 81334 404604 81418
rect 404004 81098 404186 81334
rect 404422 81098 404604 81334
rect 404004 45654 404604 81098
rect 404004 45418 404186 45654
rect 404422 45418 404604 45654
rect 404004 45334 404604 45418
rect 404004 45098 404186 45334
rect 404422 45098 404604 45334
rect 404004 9654 404604 45098
rect 404004 9418 404186 9654
rect 404422 9418 404604 9654
rect 404004 9334 404604 9418
rect 404004 9098 404186 9334
rect 404422 9098 404604 9334
rect 404004 -4026 404604 9098
rect 404004 -4262 404186 -4026
rect 404422 -4262 404604 -4026
rect 404004 -4346 404604 -4262
rect 404004 -4582 404186 -4346
rect 404422 -4582 404604 -4346
rect 404004 -5524 404604 -4582
rect 407604 697254 408204 709802
rect 425604 711278 426204 711300
rect 425604 711042 425786 711278
rect 426022 711042 426204 711278
rect 425604 710958 426204 711042
rect 425604 710722 425786 710958
rect 426022 710722 426204 710958
rect 422004 709438 422604 709460
rect 422004 709202 422186 709438
rect 422422 709202 422604 709438
rect 422004 709118 422604 709202
rect 422004 708882 422186 709118
rect 422422 708882 422604 709118
rect 418404 707598 419004 707620
rect 418404 707362 418586 707598
rect 418822 707362 419004 707598
rect 418404 707278 419004 707362
rect 418404 707042 418586 707278
rect 418822 707042 419004 707278
rect 407604 697018 407786 697254
rect 408022 697018 408204 697254
rect 407604 696934 408204 697018
rect 407604 696698 407786 696934
rect 408022 696698 408204 696934
rect 407604 661254 408204 696698
rect 407604 661018 407786 661254
rect 408022 661018 408204 661254
rect 407604 660934 408204 661018
rect 407604 660698 407786 660934
rect 408022 660698 408204 660934
rect 407604 625254 408204 660698
rect 407604 625018 407786 625254
rect 408022 625018 408204 625254
rect 407604 624934 408204 625018
rect 407604 624698 407786 624934
rect 408022 624698 408204 624934
rect 407604 589254 408204 624698
rect 407604 589018 407786 589254
rect 408022 589018 408204 589254
rect 407604 588934 408204 589018
rect 407604 588698 407786 588934
rect 408022 588698 408204 588934
rect 407604 553254 408204 588698
rect 407604 553018 407786 553254
rect 408022 553018 408204 553254
rect 407604 552934 408204 553018
rect 407604 552698 407786 552934
rect 408022 552698 408204 552934
rect 407604 517254 408204 552698
rect 407604 517018 407786 517254
rect 408022 517018 408204 517254
rect 407604 516934 408204 517018
rect 407604 516698 407786 516934
rect 408022 516698 408204 516934
rect 407604 481254 408204 516698
rect 407604 481018 407786 481254
rect 408022 481018 408204 481254
rect 407604 480934 408204 481018
rect 407604 480698 407786 480934
rect 408022 480698 408204 480934
rect 407604 445254 408204 480698
rect 407604 445018 407786 445254
rect 408022 445018 408204 445254
rect 407604 444934 408204 445018
rect 407604 444698 407786 444934
rect 408022 444698 408204 444934
rect 407604 409254 408204 444698
rect 407604 409018 407786 409254
rect 408022 409018 408204 409254
rect 407604 408934 408204 409018
rect 407604 408698 407786 408934
rect 408022 408698 408204 408934
rect 407604 373254 408204 408698
rect 407604 373018 407786 373254
rect 408022 373018 408204 373254
rect 407604 372934 408204 373018
rect 407604 372698 407786 372934
rect 408022 372698 408204 372934
rect 407604 337254 408204 372698
rect 407604 337018 407786 337254
rect 408022 337018 408204 337254
rect 407604 336934 408204 337018
rect 407604 336698 407786 336934
rect 408022 336698 408204 336934
rect 407604 301254 408204 336698
rect 407604 301018 407786 301254
rect 408022 301018 408204 301254
rect 407604 300934 408204 301018
rect 407604 300698 407786 300934
rect 408022 300698 408204 300934
rect 407604 265254 408204 300698
rect 407604 265018 407786 265254
rect 408022 265018 408204 265254
rect 407604 264934 408204 265018
rect 407604 264698 407786 264934
rect 408022 264698 408204 264934
rect 407604 229254 408204 264698
rect 407604 229018 407786 229254
rect 408022 229018 408204 229254
rect 407604 228934 408204 229018
rect 407604 228698 407786 228934
rect 408022 228698 408204 228934
rect 407604 193254 408204 228698
rect 407604 193018 407786 193254
rect 408022 193018 408204 193254
rect 407604 192934 408204 193018
rect 407604 192698 407786 192934
rect 408022 192698 408204 192934
rect 407604 157254 408204 192698
rect 407604 157018 407786 157254
rect 408022 157018 408204 157254
rect 407604 156934 408204 157018
rect 407604 156698 407786 156934
rect 408022 156698 408204 156934
rect 407604 121254 408204 156698
rect 407604 121018 407786 121254
rect 408022 121018 408204 121254
rect 407604 120934 408204 121018
rect 407604 120698 407786 120934
rect 408022 120698 408204 120934
rect 407604 85254 408204 120698
rect 407604 85018 407786 85254
rect 408022 85018 408204 85254
rect 407604 84934 408204 85018
rect 407604 84698 407786 84934
rect 408022 84698 408204 84934
rect 407604 49254 408204 84698
rect 407604 49018 407786 49254
rect 408022 49018 408204 49254
rect 407604 48934 408204 49018
rect 407604 48698 407786 48934
rect 408022 48698 408204 48934
rect 407604 13254 408204 48698
rect 407604 13018 407786 13254
rect 408022 13018 408204 13254
rect 407604 12934 408204 13018
rect 407604 12698 407786 12934
rect 408022 12698 408204 12934
rect 389604 -7022 389786 -6786
rect 390022 -7022 390204 -6786
rect 389604 -7106 390204 -7022
rect 389604 -7342 389786 -7106
rect 390022 -7342 390204 -7106
rect 389604 -7364 390204 -7342
rect 407604 -5866 408204 12698
rect 414804 705758 415404 705780
rect 414804 705522 414986 705758
rect 415222 705522 415404 705758
rect 414804 705438 415404 705522
rect 414804 705202 414986 705438
rect 415222 705202 415404 705438
rect 414804 668454 415404 705202
rect 414804 668218 414986 668454
rect 415222 668218 415404 668454
rect 414804 668134 415404 668218
rect 414804 667898 414986 668134
rect 415222 667898 415404 668134
rect 414804 632454 415404 667898
rect 414804 632218 414986 632454
rect 415222 632218 415404 632454
rect 414804 632134 415404 632218
rect 414804 631898 414986 632134
rect 415222 631898 415404 632134
rect 414804 596454 415404 631898
rect 414804 596218 414986 596454
rect 415222 596218 415404 596454
rect 414804 596134 415404 596218
rect 414804 595898 414986 596134
rect 415222 595898 415404 596134
rect 414804 560454 415404 595898
rect 414804 560218 414986 560454
rect 415222 560218 415404 560454
rect 414804 560134 415404 560218
rect 414804 559898 414986 560134
rect 415222 559898 415404 560134
rect 414804 524454 415404 559898
rect 414804 524218 414986 524454
rect 415222 524218 415404 524454
rect 414804 524134 415404 524218
rect 414804 523898 414986 524134
rect 415222 523898 415404 524134
rect 414804 488454 415404 523898
rect 414804 488218 414986 488454
rect 415222 488218 415404 488454
rect 414804 488134 415404 488218
rect 414804 487898 414986 488134
rect 415222 487898 415404 488134
rect 414804 452454 415404 487898
rect 414804 452218 414986 452454
rect 415222 452218 415404 452454
rect 414804 452134 415404 452218
rect 414804 451898 414986 452134
rect 415222 451898 415404 452134
rect 414804 416454 415404 451898
rect 414804 416218 414986 416454
rect 415222 416218 415404 416454
rect 414804 416134 415404 416218
rect 414804 415898 414986 416134
rect 415222 415898 415404 416134
rect 414804 380454 415404 415898
rect 414804 380218 414986 380454
rect 415222 380218 415404 380454
rect 414804 380134 415404 380218
rect 414804 379898 414986 380134
rect 415222 379898 415404 380134
rect 414804 344454 415404 379898
rect 414804 344218 414986 344454
rect 415222 344218 415404 344454
rect 414804 344134 415404 344218
rect 414804 343898 414986 344134
rect 415222 343898 415404 344134
rect 414804 308454 415404 343898
rect 414804 308218 414986 308454
rect 415222 308218 415404 308454
rect 414804 308134 415404 308218
rect 414804 307898 414986 308134
rect 415222 307898 415404 308134
rect 414804 272454 415404 307898
rect 414804 272218 414986 272454
rect 415222 272218 415404 272454
rect 414804 272134 415404 272218
rect 414804 271898 414986 272134
rect 415222 271898 415404 272134
rect 414804 236454 415404 271898
rect 414804 236218 414986 236454
rect 415222 236218 415404 236454
rect 414804 236134 415404 236218
rect 414804 235898 414986 236134
rect 415222 235898 415404 236134
rect 414804 200454 415404 235898
rect 414804 200218 414986 200454
rect 415222 200218 415404 200454
rect 414804 200134 415404 200218
rect 414804 199898 414986 200134
rect 415222 199898 415404 200134
rect 414804 164454 415404 199898
rect 414804 164218 414986 164454
rect 415222 164218 415404 164454
rect 414804 164134 415404 164218
rect 414804 163898 414986 164134
rect 415222 163898 415404 164134
rect 414804 128454 415404 163898
rect 414804 128218 414986 128454
rect 415222 128218 415404 128454
rect 414804 128134 415404 128218
rect 414804 127898 414986 128134
rect 415222 127898 415404 128134
rect 414804 92454 415404 127898
rect 414804 92218 414986 92454
rect 415222 92218 415404 92454
rect 414804 92134 415404 92218
rect 414804 91898 414986 92134
rect 415222 91898 415404 92134
rect 414804 56454 415404 91898
rect 414804 56218 414986 56454
rect 415222 56218 415404 56454
rect 414804 56134 415404 56218
rect 414804 55898 414986 56134
rect 415222 55898 415404 56134
rect 414804 20454 415404 55898
rect 414804 20218 414986 20454
rect 415222 20218 415404 20454
rect 414804 20134 415404 20218
rect 414804 19898 414986 20134
rect 415222 19898 415404 20134
rect 414804 -1266 415404 19898
rect 414804 -1502 414986 -1266
rect 415222 -1502 415404 -1266
rect 414804 -1586 415404 -1502
rect 414804 -1822 414986 -1586
rect 415222 -1822 415404 -1586
rect 414804 -1844 415404 -1822
rect 418404 672054 419004 707042
rect 418404 671818 418586 672054
rect 418822 671818 419004 672054
rect 418404 671734 419004 671818
rect 418404 671498 418586 671734
rect 418822 671498 419004 671734
rect 418404 636054 419004 671498
rect 418404 635818 418586 636054
rect 418822 635818 419004 636054
rect 418404 635734 419004 635818
rect 418404 635498 418586 635734
rect 418822 635498 419004 635734
rect 418404 600054 419004 635498
rect 418404 599818 418586 600054
rect 418822 599818 419004 600054
rect 418404 599734 419004 599818
rect 418404 599498 418586 599734
rect 418822 599498 419004 599734
rect 418404 564054 419004 599498
rect 418404 563818 418586 564054
rect 418822 563818 419004 564054
rect 418404 563734 419004 563818
rect 418404 563498 418586 563734
rect 418822 563498 419004 563734
rect 418404 528054 419004 563498
rect 418404 527818 418586 528054
rect 418822 527818 419004 528054
rect 418404 527734 419004 527818
rect 418404 527498 418586 527734
rect 418822 527498 419004 527734
rect 418404 492054 419004 527498
rect 418404 491818 418586 492054
rect 418822 491818 419004 492054
rect 418404 491734 419004 491818
rect 418404 491498 418586 491734
rect 418822 491498 419004 491734
rect 418404 456054 419004 491498
rect 418404 455818 418586 456054
rect 418822 455818 419004 456054
rect 418404 455734 419004 455818
rect 418404 455498 418586 455734
rect 418822 455498 419004 455734
rect 418404 420054 419004 455498
rect 418404 419818 418586 420054
rect 418822 419818 419004 420054
rect 418404 419734 419004 419818
rect 418404 419498 418586 419734
rect 418822 419498 419004 419734
rect 418404 384054 419004 419498
rect 418404 383818 418586 384054
rect 418822 383818 419004 384054
rect 418404 383734 419004 383818
rect 418404 383498 418586 383734
rect 418822 383498 419004 383734
rect 418404 348054 419004 383498
rect 418404 347818 418586 348054
rect 418822 347818 419004 348054
rect 418404 347734 419004 347818
rect 418404 347498 418586 347734
rect 418822 347498 419004 347734
rect 418404 312054 419004 347498
rect 418404 311818 418586 312054
rect 418822 311818 419004 312054
rect 418404 311734 419004 311818
rect 418404 311498 418586 311734
rect 418822 311498 419004 311734
rect 418404 276054 419004 311498
rect 418404 275818 418586 276054
rect 418822 275818 419004 276054
rect 418404 275734 419004 275818
rect 418404 275498 418586 275734
rect 418822 275498 419004 275734
rect 418404 240054 419004 275498
rect 418404 239818 418586 240054
rect 418822 239818 419004 240054
rect 418404 239734 419004 239818
rect 418404 239498 418586 239734
rect 418822 239498 419004 239734
rect 418404 204054 419004 239498
rect 418404 203818 418586 204054
rect 418822 203818 419004 204054
rect 418404 203734 419004 203818
rect 418404 203498 418586 203734
rect 418822 203498 419004 203734
rect 418404 168054 419004 203498
rect 418404 167818 418586 168054
rect 418822 167818 419004 168054
rect 418404 167734 419004 167818
rect 418404 167498 418586 167734
rect 418822 167498 419004 167734
rect 418404 132054 419004 167498
rect 418404 131818 418586 132054
rect 418822 131818 419004 132054
rect 418404 131734 419004 131818
rect 418404 131498 418586 131734
rect 418822 131498 419004 131734
rect 418404 96054 419004 131498
rect 418404 95818 418586 96054
rect 418822 95818 419004 96054
rect 418404 95734 419004 95818
rect 418404 95498 418586 95734
rect 418822 95498 419004 95734
rect 418404 60054 419004 95498
rect 418404 59818 418586 60054
rect 418822 59818 419004 60054
rect 418404 59734 419004 59818
rect 418404 59498 418586 59734
rect 418822 59498 419004 59734
rect 418404 24054 419004 59498
rect 418404 23818 418586 24054
rect 418822 23818 419004 24054
rect 418404 23734 419004 23818
rect 418404 23498 418586 23734
rect 418822 23498 419004 23734
rect 418404 -3106 419004 23498
rect 418404 -3342 418586 -3106
rect 418822 -3342 419004 -3106
rect 418404 -3426 419004 -3342
rect 418404 -3662 418586 -3426
rect 418822 -3662 419004 -3426
rect 418404 -3684 419004 -3662
rect 422004 675654 422604 708882
rect 422004 675418 422186 675654
rect 422422 675418 422604 675654
rect 422004 675334 422604 675418
rect 422004 675098 422186 675334
rect 422422 675098 422604 675334
rect 422004 639654 422604 675098
rect 422004 639418 422186 639654
rect 422422 639418 422604 639654
rect 422004 639334 422604 639418
rect 422004 639098 422186 639334
rect 422422 639098 422604 639334
rect 422004 603654 422604 639098
rect 422004 603418 422186 603654
rect 422422 603418 422604 603654
rect 422004 603334 422604 603418
rect 422004 603098 422186 603334
rect 422422 603098 422604 603334
rect 422004 567654 422604 603098
rect 422004 567418 422186 567654
rect 422422 567418 422604 567654
rect 422004 567334 422604 567418
rect 422004 567098 422186 567334
rect 422422 567098 422604 567334
rect 422004 531654 422604 567098
rect 422004 531418 422186 531654
rect 422422 531418 422604 531654
rect 422004 531334 422604 531418
rect 422004 531098 422186 531334
rect 422422 531098 422604 531334
rect 422004 495654 422604 531098
rect 422004 495418 422186 495654
rect 422422 495418 422604 495654
rect 422004 495334 422604 495418
rect 422004 495098 422186 495334
rect 422422 495098 422604 495334
rect 422004 459654 422604 495098
rect 422004 459418 422186 459654
rect 422422 459418 422604 459654
rect 422004 459334 422604 459418
rect 422004 459098 422186 459334
rect 422422 459098 422604 459334
rect 422004 423654 422604 459098
rect 422004 423418 422186 423654
rect 422422 423418 422604 423654
rect 422004 423334 422604 423418
rect 422004 423098 422186 423334
rect 422422 423098 422604 423334
rect 422004 387654 422604 423098
rect 422004 387418 422186 387654
rect 422422 387418 422604 387654
rect 422004 387334 422604 387418
rect 422004 387098 422186 387334
rect 422422 387098 422604 387334
rect 422004 351654 422604 387098
rect 422004 351418 422186 351654
rect 422422 351418 422604 351654
rect 422004 351334 422604 351418
rect 422004 351098 422186 351334
rect 422422 351098 422604 351334
rect 422004 315654 422604 351098
rect 422004 315418 422186 315654
rect 422422 315418 422604 315654
rect 422004 315334 422604 315418
rect 422004 315098 422186 315334
rect 422422 315098 422604 315334
rect 422004 279654 422604 315098
rect 422004 279418 422186 279654
rect 422422 279418 422604 279654
rect 422004 279334 422604 279418
rect 422004 279098 422186 279334
rect 422422 279098 422604 279334
rect 422004 243654 422604 279098
rect 422004 243418 422186 243654
rect 422422 243418 422604 243654
rect 422004 243334 422604 243418
rect 422004 243098 422186 243334
rect 422422 243098 422604 243334
rect 422004 207654 422604 243098
rect 422004 207418 422186 207654
rect 422422 207418 422604 207654
rect 422004 207334 422604 207418
rect 422004 207098 422186 207334
rect 422422 207098 422604 207334
rect 422004 171654 422604 207098
rect 422004 171418 422186 171654
rect 422422 171418 422604 171654
rect 422004 171334 422604 171418
rect 422004 171098 422186 171334
rect 422422 171098 422604 171334
rect 422004 135654 422604 171098
rect 422004 135418 422186 135654
rect 422422 135418 422604 135654
rect 422004 135334 422604 135418
rect 422004 135098 422186 135334
rect 422422 135098 422604 135334
rect 422004 99654 422604 135098
rect 422004 99418 422186 99654
rect 422422 99418 422604 99654
rect 422004 99334 422604 99418
rect 422004 99098 422186 99334
rect 422422 99098 422604 99334
rect 422004 63654 422604 99098
rect 422004 63418 422186 63654
rect 422422 63418 422604 63654
rect 422004 63334 422604 63418
rect 422004 63098 422186 63334
rect 422422 63098 422604 63334
rect 422004 27654 422604 63098
rect 422004 27418 422186 27654
rect 422422 27418 422604 27654
rect 422004 27334 422604 27418
rect 422004 27098 422186 27334
rect 422422 27098 422604 27334
rect 422004 -4946 422604 27098
rect 422004 -5182 422186 -4946
rect 422422 -5182 422604 -4946
rect 422004 -5266 422604 -5182
rect 422004 -5502 422186 -5266
rect 422422 -5502 422604 -5266
rect 422004 -5524 422604 -5502
rect 425604 679254 426204 710722
rect 443604 710358 444204 711300
rect 443604 710122 443786 710358
rect 444022 710122 444204 710358
rect 443604 710038 444204 710122
rect 443604 709802 443786 710038
rect 444022 709802 444204 710038
rect 440004 708518 440604 709460
rect 440004 708282 440186 708518
rect 440422 708282 440604 708518
rect 440004 708198 440604 708282
rect 440004 707962 440186 708198
rect 440422 707962 440604 708198
rect 436404 706678 437004 707620
rect 436404 706442 436586 706678
rect 436822 706442 437004 706678
rect 436404 706358 437004 706442
rect 436404 706122 436586 706358
rect 436822 706122 437004 706358
rect 425604 679018 425786 679254
rect 426022 679018 426204 679254
rect 425604 678934 426204 679018
rect 425604 678698 425786 678934
rect 426022 678698 426204 678934
rect 425604 643254 426204 678698
rect 425604 643018 425786 643254
rect 426022 643018 426204 643254
rect 425604 642934 426204 643018
rect 425604 642698 425786 642934
rect 426022 642698 426204 642934
rect 425604 607254 426204 642698
rect 425604 607018 425786 607254
rect 426022 607018 426204 607254
rect 425604 606934 426204 607018
rect 425604 606698 425786 606934
rect 426022 606698 426204 606934
rect 425604 571254 426204 606698
rect 425604 571018 425786 571254
rect 426022 571018 426204 571254
rect 425604 570934 426204 571018
rect 425604 570698 425786 570934
rect 426022 570698 426204 570934
rect 425604 535254 426204 570698
rect 425604 535018 425786 535254
rect 426022 535018 426204 535254
rect 425604 534934 426204 535018
rect 425604 534698 425786 534934
rect 426022 534698 426204 534934
rect 425604 499254 426204 534698
rect 425604 499018 425786 499254
rect 426022 499018 426204 499254
rect 425604 498934 426204 499018
rect 425604 498698 425786 498934
rect 426022 498698 426204 498934
rect 425604 463254 426204 498698
rect 425604 463018 425786 463254
rect 426022 463018 426204 463254
rect 425604 462934 426204 463018
rect 425604 462698 425786 462934
rect 426022 462698 426204 462934
rect 425604 427254 426204 462698
rect 425604 427018 425786 427254
rect 426022 427018 426204 427254
rect 425604 426934 426204 427018
rect 425604 426698 425786 426934
rect 426022 426698 426204 426934
rect 425604 391254 426204 426698
rect 425604 391018 425786 391254
rect 426022 391018 426204 391254
rect 425604 390934 426204 391018
rect 425604 390698 425786 390934
rect 426022 390698 426204 390934
rect 425604 355254 426204 390698
rect 425604 355018 425786 355254
rect 426022 355018 426204 355254
rect 425604 354934 426204 355018
rect 425604 354698 425786 354934
rect 426022 354698 426204 354934
rect 425604 319254 426204 354698
rect 425604 319018 425786 319254
rect 426022 319018 426204 319254
rect 425604 318934 426204 319018
rect 425604 318698 425786 318934
rect 426022 318698 426204 318934
rect 425604 283254 426204 318698
rect 425604 283018 425786 283254
rect 426022 283018 426204 283254
rect 425604 282934 426204 283018
rect 425604 282698 425786 282934
rect 426022 282698 426204 282934
rect 425604 247254 426204 282698
rect 425604 247018 425786 247254
rect 426022 247018 426204 247254
rect 425604 246934 426204 247018
rect 425604 246698 425786 246934
rect 426022 246698 426204 246934
rect 425604 211254 426204 246698
rect 425604 211018 425786 211254
rect 426022 211018 426204 211254
rect 425604 210934 426204 211018
rect 425604 210698 425786 210934
rect 426022 210698 426204 210934
rect 425604 175254 426204 210698
rect 425604 175018 425786 175254
rect 426022 175018 426204 175254
rect 425604 174934 426204 175018
rect 425604 174698 425786 174934
rect 426022 174698 426204 174934
rect 425604 139254 426204 174698
rect 425604 139018 425786 139254
rect 426022 139018 426204 139254
rect 425604 138934 426204 139018
rect 425604 138698 425786 138934
rect 426022 138698 426204 138934
rect 425604 103254 426204 138698
rect 425604 103018 425786 103254
rect 426022 103018 426204 103254
rect 425604 102934 426204 103018
rect 425604 102698 425786 102934
rect 426022 102698 426204 102934
rect 425604 67254 426204 102698
rect 425604 67018 425786 67254
rect 426022 67018 426204 67254
rect 425604 66934 426204 67018
rect 425604 66698 425786 66934
rect 426022 66698 426204 66934
rect 425604 31254 426204 66698
rect 425604 31018 425786 31254
rect 426022 31018 426204 31254
rect 425604 30934 426204 31018
rect 425604 30698 425786 30934
rect 426022 30698 426204 30934
rect 407604 -6102 407786 -5866
rect 408022 -6102 408204 -5866
rect 407604 -6186 408204 -6102
rect 407604 -6422 407786 -6186
rect 408022 -6422 408204 -6186
rect 407604 -7364 408204 -6422
rect 425604 -6786 426204 30698
rect 432804 704838 433404 705780
rect 432804 704602 432986 704838
rect 433222 704602 433404 704838
rect 432804 704518 433404 704602
rect 432804 704282 432986 704518
rect 433222 704282 433404 704518
rect 432804 686454 433404 704282
rect 432804 686218 432986 686454
rect 433222 686218 433404 686454
rect 432804 686134 433404 686218
rect 432804 685898 432986 686134
rect 433222 685898 433404 686134
rect 432804 650454 433404 685898
rect 432804 650218 432986 650454
rect 433222 650218 433404 650454
rect 432804 650134 433404 650218
rect 432804 649898 432986 650134
rect 433222 649898 433404 650134
rect 432804 614454 433404 649898
rect 432804 614218 432986 614454
rect 433222 614218 433404 614454
rect 432804 614134 433404 614218
rect 432804 613898 432986 614134
rect 433222 613898 433404 614134
rect 432804 578454 433404 613898
rect 432804 578218 432986 578454
rect 433222 578218 433404 578454
rect 432804 578134 433404 578218
rect 432804 577898 432986 578134
rect 433222 577898 433404 578134
rect 432804 542454 433404 577898
rect 432804 542218 432986 542454
rect 433222 542218 433404 542454
rect 432804 542134 433404 542218
rect 432804 541898 432986 542134
rect 433222 541898 433404 542134
rect 432804 506454 433404 541898
rect 432804 506218 432986 506454
rect 433222 506218 433404 506454
rect 432804 506134 433404 506218
rect 432804 505898 432986 506134
rect 433222 505898 433404 506134
rect 432804 470454 433404 505898
rect 432804 470218 432986 470454
rect 433222 470218 433404 470454
rect 432804 470134 433404 470218
rect 432804 469898 432986 470134
rect 433222 469898 433404 470134
rect 432804 434454 433404 469898
rect 432804 434218 432986 434454
rect 433222 434218 433404 434454
rect 432804 434134 433404 434218
rect 432804 433898 432986 434134
rect 433222 433898 433404 434134
rect 432804 398454 433404 433898
rect 432804 398218 432986 398454
rect 433222 398218 433404 398454
rect 432804 398134 433404 398218
rect 432804 397898 432986 398134
rect 433222 397898 433404 398134
rect 432804 362454 433404 397898
rect 432804 362218 432986 362454
rect 433222 362218 433404 362454
rect 432804 362134 433404 362218
rect 432804 361898 432986 362134
rect 433222 361898 433404 362134
rect 432804 326454 433404 361898
rect 432804 326218 432986 326454
rect 433222 326218 433404 326454
rect 432804 326134 433404 326218
rect 432804 325898 432986 326134
rect 433222 325898 433404 326134
rect 432804 290454 433404 325898
rect 432804 290218 432986 290454
rect 433222 290218 433404 290454
rect 432804 290134 433404 290218
rect 432804 289898 432986 290134
rect 433222 289898 433404 290134
rect 432804 254454 433404 289898
rect 432804 254218 432986 254454
rect 433222 254218 433404 254454
rect 432804 254134 433404 254218
rect 432804 253898 432986 254134
rect 433222 253898 433404 254134
rect 432804 218454 433404 253898
rect 432804 218218 432986 218454
rect 433222 218218 433404 218454
rect 432804 218134 433404 218218
rect 432804 217898 432986 218134
rect 433222 217898 433404 218134
rect 432804 182454 433404 217898
rect 432804 182218 432986 182454
rect 433222 182218 433404 182454
rect 432804 182134 433404 182218
rect 432804 181898 432986 182134
rect 433222 181898 433404 182134
rect 432804 146454 433404 181898
rect 432804 146218 432986 146454
rect 433222 146218 433404 146454
rect 432804 146134 433404 146218
rect 432804 145898 432986 146134
rect 433222 145898 433404 146134
rect 432804 110454 433404 145898
rect 432804 110218 432986 110454
rect 433222 110218 433404 110454
rect 432804 110134 433404 110218
rect 432804 109898 432986 110134
rect 433222 109898 433404 110134
rect 432804 74454 433404 109898
rect 432804 74218 432986 74454
rect 433222 74218 433404 74454
rect 432804 74134 433404 74218
rect 432804 73898 432986 74134
rect 433222 73898 433404 74134
rect 432804 38454 433404 73898
rect 432804 38218 432986 38454
rect 433222 38218 433404 38454
rect 432804 38134 433404 38218
rect 432804 37898 432986 38134
rect 433222 37898 433404 38134
rect 432804 2454 433404 37898
rect 432804 2218 432986 2454
rect 433222 2218 433404 2454
rect 432804 2134 433404 2218
rect 432804 1898 432986 2134
rect 433222 1898 433404 2134
rect 432804 -346 433404 1898
rect 432804 -582 432986 -346
rect 433222 -582 433404 -346
rect 432804 -666 433404 -582
rect 432804 -902 432986 -666
rect 433222 -902 433404 -666
rect 432804 -1844 433404 -902
rect 436404 690054 437004 706122
rect 436404 689818 436586 690054
rect 436822 689818 437004 690054
rect 436404 689734 437004 689818
rect 436404 689498 436586 689734
rect 436822 689498 437004 689734
rect 436404 654054 437004 689498
rect 436404 653818 436586 654054
rect 436822 653818 437004 654054
rect 436404 653734 437004 653818
rect 436404 653498 436586 653734
rect 436822 653498 437004 653734
rect 436404 618054 437004 653498
rect 436404 617818 436586 618054
rect 436822 617818 437004 618054
rect 436404 617734 437004 617818
rect 436404 617498 436586 617734
rect 436822 617498 437004 617734
rect 436404 582054 437004 617498
rect 436404 581818 436586 582054
rect 436822 581818 437004 582054
rect 436404 581734 437004 581818
rect 436404 581498 436586 581734
rect 436822 581498 437004 581734
rect 436404 546054 437004 581498
rect 436404 545818 436586 546054
rect 436822 545818 437004 546054
rect 436404 545734 437004 545818
rect 436404 545498 436586 545734
rect 436822 545498 437004 545734
rect 436404 510054 437004 545498
rect 436404 509818 436586 510054
rect 436822 509818 437004 510054
rect 436404 509734 437004 509818
rect 436404 509498 436586 509734
rect 436822 509498 437004 509734
rect 436404 474054 437004 509498
rect 436404 473818 436586 474054
rect 436822 473818 437004 474054
rect 436404 473734 437004 473818
rect 436404 473498 436586 473734
rect 436822 473498 437004 473734
rect 436404 438054 437004 473498
rect 436404 437818 436586 438054
rect 436822 437818 437004 438054
rect 436404 437734 437004 437818
rect 436404 437498 436586 437734
rect 436822 437498 437004 437734
rect 436404 402054 437004 437498
rect 436404 401818 436586 402054
rect 436822 401818 437004 402054
rect 436404 401734 437004 401818
rect 436404 401498 436586 401734
rect 436822 401498 437004 401734
rect 436404 366054 437004 401498
rect 436404 365818 436586 366054
rect 436822 365818 437004 366054
rect 436404 365734 437004 365818
rect 436404 365498 436586 365734
rect 436822 365498 437004 365734
rect 436404 330054 437004 365498
rect 436404 329818 436586 330054
rect 436822 329818 437004 330054
rect 436404 329734 437004 329818
rect 436404 329498 436586 329734
rect 436822 329498 437004 329734
rect 436404 294054 437004 329498
rect 436404 293818 436586 294054
rect 436822 293818 437004 294054
rect 436404 293734 437004 293818
rect 436404 293498 436586 293734
rect 436822 293498 437004 293734
rect 436404 258054 437004 293498
rect 436404 257818 436586 258054
rect 436822 257818 437004 258054
rect 436404 257734 437004 257818
rect 436404 257498 436586 257734
rect 436822 257498 437004 257734
rect 436404 222054 437004 257498
rect 436404 221818 436586 222054
rect 436822 221818 437004 222054
rect 436404 221734 437004 221818
rect 436404 221498 436586 221734
rect 436822 221498 437004 221734
rect 436404 186054 437004 221498
rect 436404 185818 436586 186054
rect 436822 185818 437004 186054
rect 436404 185734 437004 185818
rect 436404 185498 436586 185734
rect 436822 185498 437004 185734
rect 436404 150054 437004 185498
rect 436404 149818 436586 150054
rect 436822 149818 437004 150054
rect 436404 149734 437004 149818
rect 436404 149498 436586 149734
rect 436822 149498 437004 149734
rect 436404 114054 437004 149498
rect 436404 113818 436586 114054
rect 436822 113818 437004 114054
rect 436404 113734 437004 113818
rect 436404 113498 436586 113734
rect 436822 113498 437004 113734
rect 436404 78054 437004 113498
rect 436404 77818 436586 78054
rect 436822 77818 437004 78054
rect 436404 77734 437004 77818
rect 436404 77498 436586 77734
rect 436822 77498 437004 77734
rect 436404 42054 437004 77498
rect 436404 41818 436586 42054
rect 436822 41818 437004 42054
rect 436404 41734 437004 41818
rect 436404 41498 436586 41734
rect 436822 41498 437004 41734
rect 436404 6054 437004 41498
rect 436404 5818 436586 6054
rect 436822 5818 437004 6054
rect 436404 5734 437004 5818
rect 436404 5498 436586 5734
rect 436822 5498 437004 5734
rect 436404 -2186 437004 5498
rect 436404 -2422 436586 -2186
rect 436822 -2422 437004 -2186
rect 436404 -2506 437004 -2422
rect 436404 -2742 436586 -2506
rect 436822 -2742 437004 -2506
rect 436404 -3684 437004 -2742
rect 440004 693654 440604 707962
rect 440004 693418 440186 693654
rect 440422 693418 440604 693654
rect 440004 693334 440604 693418
rect 440004 693098 440186 693334
rect 440422 693098 440604 693334
rect 440004 657654 440604 693098
rect 440004 657418 440186 657654
rect 440422 657418 440604 657654
rect 440004 657334 440604 657418
rect 440004 657098 440186 657334
rect 440422 657098 440604 657334
rect 440004 621654 440604 657098
rect 440004 621418 440186 621654
rect 440422 621418 440604 621654
rect 440004 621334 440604 621418
rect 440004 621098 440186 621334
rect 440422 621098 440604 621334
rect 440004 585654 440604 621098
rect 440004 585418 440186 585654
rect 440422 585418 440604 585654
rect 440004 585334 440604 585418
rect 440004 585098 440186 585334
rect 440422 585098 440604 585334
rect 440004 549654 440604 585098
rect 440004 549418 440186 549654
rect 440422 549418 440604 549654
rect 440004 549334 440604 549418
rect 440004 549098 440186 549334
rect 440422 549098 440604 549334
rect 440004 513654 440604 549098
rect 440004 513418 440186 513654
rect 440422 513418 440604 513654
rect 440004 513334 440604 513418
rect 440004 513098 440186 513334
rect 440422 513098 440604 513334
rect 440004 477654 440604 513098
rect 440004 477418 440186 477654
rect 440422 477418 440604 477654
rect 440004 477334 440604 477418
rect 440004 477098 440186 477334
rect 440422 477098 440604 477334
rect 440004 441654 440604 477098
rect 440004 441418 440186 441654
rect 440422 441418 440604 441654
rect 440004 441334 440604 441418
rect 440004 441098 440186 441334
rect 440422 441098 440604 441334
rect 440004 405654 440604 441098
rect 440004 405418 440186 405654
rect 440422 405418 440604 405654
rect 440004 405334 440604 405418
rect 440004 405098 440186 405334
rect 440422 405098 440604 405334
rect 440004 369654 440604 405098
rect 440004 369418 440186 369654
rect 440422 369418 440604 369654
rect 440004 369334 440604 369418
rect 440004 369098 440186 369334
rect 440422 369098 440604 369334
rect 440004 333654 440604 369098
rect 440004 333418 440186 333654
rect 440422 333418 440604 333654
rect 440004 333334 440604 333418
rect 440004 333098 440186 333334
rect 440422 333098 440604 333334
rect 440004 297654 440604 333098
rect 440004 297418 440186 297654
rect 440422 297418 440604 297654
rect 440004 297334 440604 297418
rect 440004 297098 440186 297334
rect 440422 297098 440604 297334
rect 440004 261654 440604 297098
rect 440004 261418 440186 261654
rect 440422 261418 440604 261654
rect 440004 261334 440604 261418
rect 440004 261098 440186 261334
rect 440422 261098 440604 261334
rect 440004 225654 440604 261098
rect 440004 225418 440186 225654
rect 440422 225418 440604 225654
rect 440004 225334 440604 225418
rect 440004 225098 440186 225334
rect 440422 225098 440604 225334
rect 440004 189654 440604 225098
rect 440004 189418 440186 189654
rect 440422 189418 440604 189654
rect 440004 189334 440604 189418
rect 440004 189098 440186 189334
rect 440422 189098 440604 189334
rect 440004 153654 440604 189098
rect 440004 153418 440186 153654
rect 440422 153418 440604 153654
rect 440004 153334 440604 153418
rect 440004 153098 440186 153334
rect 440422 153098 440604 153334
rect 440004 117654 440604 153098
rect 440004 117418 440186 117654
rect 440422 117418 440604 117654
rect 440004 117334 440604 117418
rect 440004 117098 440186 117334
rect 440422 117098 440604 117334
rect 440004 81654 440604 117098
rect 440004 81418 440186 81654
rect 440422 81418 440604 81654
rect 440004 81334 440604 81418
rect 440004 81098 440186 81334
rect 440422 81098 440604 81334
rect 440004 45654 440604 81098
rect 440004 45418 440186 45654
rect 440422 45418 440604 45654
rect 440004 45334 440604 45418
rect 440004 45098 440186 45334
rect 440422 45098 440604 45334
rect 440004 9654 440604 45098
rect 440004 9418 440186 9654
rect 440422 9418 440604 9654
rect 440004 9334 440604 9418
rect 440004 9098 440186 9334
rect 440422 9098 440604 9334
rect 440004 -4026 440604 9098
rect 440004 -4262 440186 -4026
rect 440422 -4262 440604 -4026
rect 440004 -4346 440604 -4262
rect 440004 -4582 440186 -4346
rect 440422 -4582 440604 -4346
rect 440004 -5524 440604 -4582
rect 443604 697254 444204 709802
rect 461604 711278 462204 711300
rect 461604 711042 461786 711278
rect 462022 711042 462204 711278
rect 461604 710958 462204 711042
rect 461604 710722 461786 710958
rect 462022 710722 462204 710958
rect 458004 709438 458604 709460
rect 458004 709202 458186 709438
rect 458422 709202 458604 709438
rect 458004 709118 458604 709202
rect 458004 708882 458186 709118
rect 458422 708882 458604 709118
rect 454404 707598 455004 707620
rect 454404 707362 454586 707598
rect 454822 707362 455004 707598
rect 454404 707278 455004 707362
rect 454404 707042 454586 707278
rect 454822 707042 455004 707278
rect 443604 697018 443786 697254
rect 444022 697018 444204 697254
rect 443604 696934 444204 697018
rect 443604 696698 443786 696934
rect 444022 696698 444204 696934
rect 443604 661254 444204 696698
rect 443604 661018 443786 661254
rect 444022 661018 444204 661254
rect 443604 660934 444204 661018
rect 443604 660698 443786 660934
rect 444022 660698 444204 660934
rect 443604 625254 444204 660698
rect 443604 625018 443786 625254
rect 444022 625018 444204 625254
rect 443604 624934 444204 625018
rect 443604 624698 443786 624934
rect 444022 624698 444204 624934
rect 443604 589254 444204 624698
rect 443604 589018 443786 589254
rect 444022 589018 444204 589254
rect 443604 588934 444204 589018
rect 443604 588698 443786 588934
rect 444022 588698 444204 588934
rect 443604 553254 444204 588698
rect 443604 553018 443786 553254
rect 444022 553018 444204 553254
rect 443604 552934 444204 553018
rect 443604 552698 443786 552934
rect 444022 552698 444204 552934
rect 443604 517254 444204 552698
rect 443604 517018 443786 517254
rect 444022 517018 444204 517254
rect 443604 516934 444204 517018
rect 443604 516698 443786 516934
rect 444022 516698 444204 516934
rect 443604 481254 444204 516698
rect 443604 481018 443786 481254
rect 444022 481018 444204 481254
rect 443604 480934 444204 481018
rect 443604 480698 443786 480934
rect 444022 480698 444204 480934
rect 443604 445254 444204 480698
rect 443604 445018 443786 445254
rect 444022 445018 444204 445254
rect 443604 444934 444204 445018
rect 443604 444698 443786 444934
rect 444022 444698 444204 444934
rect 443604 409254 444204 444698
rect 443604 409018 443786 409254
rect 444022 409018 444204 409254
rect 443604 408934 444204 409018
rect 443604 408698 443786 408934
rect 444022 408698 444204 408934
rect 443604 373254 444204 408698
rect 443604 373018 443786 373254
rect 444022 373018 444204 373254
rect 443604 372934 444204 373018
rect 443604 372698 443786 372934
rect 444022 372698 444204 372934
rect 443604 337254 444204 372698
rect 443604 337018 443786 337254
rect 444022 337018 444204 337254
rect 443604 336934 444204 337018
rect 443604 336698 443786 336934
rect 444022 336698 444204 336934
rect 443604 301254 444204 336698
rect 443604 301018 443786 301254
rect 444022 301018 444204 301254
rect 443604 300934 444204 301018
rect 443604 300698 443786 300934
rect 444022 300698 444204 300934
rect 443604 265254 444204 300698
rect 443604 265018 443786 265254
rect 444022 265018 444204 265254
rect 443604 264934 444204 265018
rect 443604 264698 443786 264934
rect 444022 264698 444204 264934
rect 443604 229254 444204 264698
rect 443604 229018 443786 229254
rect 444022 229018 444204 229254
rect 443604 228934 444204 229018
rect 443604 228698 443786 228934
rect 444022 228698 444204 228934
rect 443604 193254 444204 228698
rect 443604 193018 443786 193254
rect 444022 193018 444204 193254
rect 443604 192934 444204 193018
rect 443604 192698 443786 192934
rect 444022 192698 444204 192934
rect 443604 157254 444204 192698
rect 443604 157018 443786 157254
rect 444022 157018 444204 157254
rect 443604 156934 444204 157018
rect 443604 156698 443786 156934
rect 444022 156698 444204 156934
rect 443604 121254 444204 156698
rect 443604 121018 443786 121254
rect 444022 121018 444204 121254
rect 443604 120934 444204 121018
rect 443604 120698 443786 120934
rect 444022 120698 444204 120934
rect 443604 85254 444204 120698
rect 443604 85018 443786 85254
rect 444022 85018 444204 85254
rect 443604 84934 444204 85018
rect 443604 84698 443786 84934
rect 444022 84698 444204 84934
rect 443604 49254 444204 84698
rect 443604 49018 443786 49254
rect 444022 49018 444204 49254
rect 443604 48934 444204 49018
rect 443604 48698 443786 48934
rect 444022 48698 444204 48934
rect 443604 13254 444204 48698
rect 443604 13018 443786 13254
rect 444022 13018 444204 13254
rect 443604 12934 444204 13018
rect 443604 12698 443786 12934
rect 444022 12698 444204 12934
rect 425604 -7022 425786 -6786
rect 426022 -7022 426204 -6786
rect 425604 -7106 426204 -7022
rect 425604 -7342 425786 -7106
rect 426022 -7342 426204 -7106
rect 425604 -7364 426204 -7342
rect 443604 -5866 444204 12698
rect 450804 705758 451404 705780
rect 450804 705522 450986 705758
rect 451222 705522 451404 705758
rect 450804 705438 451404 705522
rect 450804 705202 450986 705438
rect 451222 705202 451404 705438
rect 450804 668454 451404 705202
rect 450804 668218 450986 668454
rect 451222 668218 451404 668454
rect 450804 668134 451404 668218
rect 450804 667898 450986 668134
rect 451222 667898 451404 668134
rect 450804 632454 451404 667898
rect 450804 632218 450986 632454
rect 451222 632218 451404 632454
rect 450804 632134 451404 632218
rect 450804 631898 450986 632134
rect 451222 631898 451404 632134
rect 450804 596454 451404 631898
rect 450804 596218 450986 596454
rect 451222 596218 451404 596454
rect 450804 596134 451404 596218
rect 450804 595898 450986 596134
rect 451222 595898 451404 596134
rect 450804 560454 451404 595898
rect 450804 560218 450986 560454
rect 451222 560218 451404 560454
rect 450804 560134 451404 560218
rect 450804 559898 450986 560134
rect 451222 559898 451404 560134
rect 450804 524454 451404 559898
rect 450804 524218 450986 524454
rect 451222 524218 451404 524454
rect 450804 524134 451404 524218
rect 450804 523898 450986 524134
rect 451222 523898 451404 524134
rect 450804 488454 451404 523898
rect 450804 488218 450986 488454
rect 451222 488218 451404 488454
rect 450804 488134 451404 488218
rect 450804 487898 450986 488134
rect 451222 487898 451404 488134
rect 450804 452454 451404 487898
rect 450804 452218 450986 452454
rect 451222 452218 451404 452454
rect 450804 452134 451404 452218
rect 450804 451898 450986 452134
rect 451222 451898 451404 452134
rect 450804 416454 451404 451898
rect 450804 416218 450986 416454
rect 451222 416218 451404 416454
rect 450804 416134 451404 416218
rect 450804 415898 450986 416134
rect 451222 415898 451404 416134
rect 450804 380454 451404 415898
rect 450804 380218 450986 380454
rect 451222 380218 451404 380454
rect 450804 380134 451404 380218
rect 450804 379898 450986 380134
rect 451222 379898 451404 380134
rect 450804 344454 451404 379898
rect 450804 344218 450986 344454
rect 451222 344218 451404 344454
rect 450804 344134 451404 344218
rect 450804 343898 450986 344134
rect 451222 343898 451404 344134
rect 450804 308454 451404 343898
rect 450804 308218 450986 308454
rect 451222 308218 451404 308454
rect 450804 308134 451404 308218
rect 450804 307898 450986 308134
rect 451222 307898 451404 308134
rect 450804 272454 451404 307898
rect 450804 272218 450986 272454
rect 451222 272218 451404 272454
rect 450804 272134 451404 272218
rect 450804 271898 450986 272134
rect 451222 271898 451404 272134
rect 450804 236454 451404 271898
rect 450804 236218 450986 236454
rect 451222 236218 451404 236454
rect 450804 236134 451404 236218
rect 450804 235898 450986 236134
rect 451222 235898 451404 236134
rect 450804 200454 451404 235898
rect 450804 200218 450986 200454
rect 451222 200218 451404 200454
rect 450804 200134 451404 200218
rect 450804 199898 450986 200134
rect 451222 199898 451404 200134
rect 450804 164454 451404 199898
rect 450804 164218 450986 164454
rect 451222 164218 451404 164454
rect 450804 164134 451404 164218
rect 450804 163898 450986 164134
rect 451222 163898 451404 164134
rect 450804 128454 451404 163898
rect 450804 128218 450986 128454
rect 451222 128218 451404 128454
rect 450804 128134 451404 128218
rect 450804 127898 450986 128134
rect 451222 127898 451404 128134
rect 450804 92454 451404 127898
rect 450804 92218 450986 92454
rect 451222 92218 451404 92454
rect 450804 92134 451404 92218
rect 450804 91898 450986 92134
rect 451222 91898 451404 92134
rect 450804 56454 451404 91898
rect 450804 56218 450986 56454
rect 451222 56218 451404 56454
rect 450804 56134 451404 56218
rect 450804 55898 450986 56134
rect 451222 55898 451404 56134
rect 450804 20454 451404 55898
rect 450804 20218 450986 20454
rect 451222 20218 451404 20454
rect 450804 20134 451404 20218
rect 450804 19898 450986 20134
rect 451222 19898 451404 20134
rect 450804 -1266 451404 19898
rect 450804 -1502 450986 -1266
rect 451222 -1502 451404 -1266
rect 450804 -1586 451404 -1502
rect 450804 -1822 450986 -1586
rect 451222 -1822 451404 -1586
rect 450804 -1844 451404 -1822
rect 454404 672054 455004 707042
rect 454404 671818 454586 672054
rect 454822 671818 455004 672054
rect 454404 671734 455004 671818
rect 454404 671498 454586 671734
rect 454822 671498 455004 671734
rect 454404 636054 455004 671498
rect 454404 635818 454586 636054
rect 454822 635818 455004 636054
rect 454404 635734 455004 635818
rect 454404 635498 454586 635734
rect 454822 635498 455004 635734
rect 454404 600054 455004 635498
rect 454404 599818 454586 600054
rect 454822 599818 455004 600054
rect 454404 599734 455004 599818
rect 454404 599498 454586 599734
rect 454822 599498 455004 599734
rect 454404 564054 455004 599498
rect 454404 563818 454586 564054
rect 454822 563818 455004 564054
rect 454404 563734 455004 563818
rect 454404 563498 454586 563734
rect 454822 563498 455004 563734
rect 454404 528054 455004 563498
rect 454404 527818 454586 528054
rect 454822 527818 455004 528054
rect 454404 527734 455004 527818
rect 454404 527498 454586 527734
rect 454822 527498 455004 527734
rect 454404 492054 455004 527498
rect 454404 491818 454586 492054
rect 454822 491818 455004 492054
rect 454404 491734 455004 491818
rect 454404 491498 454586 491734
rect 454822 491498 455004 491734
rect 454404 456054 455004 491498
rect 454404 455818 454586 456054
rect 454822 455818 455004 456054
rect 454404 455734 455004 455818
rect 454404 455498 454586 455734
rect 454822 455498 455004 455734
rect 454404 420054 455004 455498
rect 454404 419818 454586 420054
rect 454822 419818 455004 420054
rect 454404 419734 455004 419818
rect 454404 419498 454586 419734
rect 454822 419498 455004 419734
rect 454404 384054 455004 419498
rect 454404 383818 454586 384054
rect 454822 383818 455004 384054
rect 454404 383734 455004 383818
rect 454404 383498 454586 383734
rect 454822 383498 455004 383734
rect 454404 348054 455004 383498
rect 454404 347818 454586 348054
rect 454822 347818 455004 348054
rect 454404 347734 455004 347818
rect 454404 347498 454586 347734
rect 454822 347498 455004 347734
rect 454404 312054 455004 347498
rect 454404 311818 454586 312054
rect 454822 311818 455004 312054
rect 454404 311734 455004 311818
rect 454404 311498 454586 311734
rect 454822 311498 455004 311734
rect 454404 276054 455004 311498
rect 454404 275818 454586 276054
rect 454822 275818 455004 276054
rect 454404 275734 455004 275818
rect 454404 275498 454586 275734
rect 454822 275498 455004 275734
rect 454404 240054 455004 275498
rect 454404 239818 454586 240054
rect 454822 239818 455004 240054
rect 454404 239734 455004 239818
rect 454404 239498 454586 239734
rect 454822 239498 455004 239734
rect 454404 204054 455004 239498
rect 454404 203818 454586 204054
rect 454822 203818 455004 204054
rect 454404 203734 455004 203818
rect 454404 203498 454586 203734
rect 454822 203498 455004 203734
rect 454404 168054 455004 203498
rect 454404 167818 454586 168054
rect 454822 167818 455004 168054
rect 454404 167734 455004 167818
rect 454404 167498 454586 167734
rect 454822 167498 455004 167734
rect 454404 132054 455004 167498
rect 454404 131818 454586 132054
rect 454822 131818 455004 132054
rect 454404 131734 455004 131818
rect 454404 131498 454586 131734
rect 454822 131498 455004 131734
rect 454404 96054 455004 131498
rect 454404 95818 454586 96054
rect 454822 95818 455004 96054
rect 454404 95734 455004 95818
rect 454404 95498 454586 95734
rect 454822 95498 455004 95734
rect 454404 60054 455004 95498
rect 454404 59818 454586 60054
rect 454822 59818 455004 60054
rect 454404 59734 455004 59818
rect 454404 59498 454586 59734
rect 454822 59498 455004 59734
rect 454404 24054 455004 59498
rect 454404 23818 454586 24054
rect 454822 23818 455004 24054
rect 454404 23734 455004 23818
rect 454404 23498 454586 23734
rect 454822 23498 455004 23734
rect 454404 -3106 455004 23498
rect 454404 -3342 454586 -3106
rect 454822 -3342 455004 -3106
rect 454404 -3426 455004 -3342
rect 454404 -3662 454586 -3426
rect 454822 -3662 455004 -3426
rect 454404 -3684 455004 -3662
rect 458004 675654 458604 708882
rect 458004 675418 458186 675654
rect 458422 675418 458604 675654
rect 458004 675334 458604 675418
rect 458004 675098 458186 675334
rect 458422 675098 458604 675334
rect 458004 639654 458604 675098
rect 458004 639418 458186 639654
rect 458422 639418 458604 639654
rect 458004 639334 458604 639418
rect 458004 639098 458186 639334
rect 458422 639098 458604 639334
rect 458004 603654 458604 639098
rect 458004 603418 458186 603654
rect 458422 603418 458604 603654
rect 458004 603334 458604 603418
rect 458004 603098 458186 603334
rect 458422 603098 458604 603334
rect 458004 567654 458604 603098
rect 458004 567418 458186 567654
rect 458422 567418 458604 567654
rect 458004 567334 458604 567418
rect 458004 567098 458186 567334
rect 458422 567098 458604 567334
rect 458004 531654 458604 567098
rect 458004 531418 458186 531654
rect 458422 531418 458604 531654
rect 458004 531334 458604 531418
rect 458004 531098 458186 531334
rect 458422 531098 458604 531334
rect 458004 495654 458604 531098
rect 458004 495418 458186 495654
rect 458422 495418 458604 495654
rect 458004 495334 458604 495418
rect 458004 495098 458186 495334
rect 458422 495098 458604 495334
rect 458004 459654 458604 495098
rect 458004 459418 458186 459654
rect 458422 459418 458604 459654
rect 458004 459334 458604 459418
rect 458004 459098 458186 459334
rect 458422 459098 458604 459334
rect 458004 423654 458604 459098
rect 458004 423418 458186 423654
rect 458422 423418 458604 423654
rect 458004 423334 458604 423418
rect 458004 423098 458186 423334
rect 458422 423098 458604 423334
rect 458004 387654 458604 423098
rect 458004 387418 458186 387654
rect 458422 387418 458604 387654
rect 458004 387334 458604 387418
rect 458004 387098 458186 387334
rect 458422 387098 458604 387334
rect 458004 351654 458604 387098
rect 458004 351418 458186 351654
rect 458422 351418 458604 351654
rect 458004 351334 458604 351418
rect 458004 351098 458186 351334
rect 458422 351098 458604 351334
rect 458004 315654 458604 351098
rect 458004 315418 458186 315654
rect 458422 315418 458604 315654
rect 458004 315334 458604 315418
rect 458004 315098 458186 315334
rect 458422 315098 458604 315334
rect 458004 279654 458604 315098
rect 458004 279418 458186 279654
rect 458422 279418 458604 279654
rect 458004 279334 458604 279418
rect 458004 279098 458186 279334
rect 458422 279098 458604 279334
rect 458004 243654 458604 279098
rect 458004 243418 458186 243654
rect 458422 243418 458604 243654
rect 458004 243334 458604 243418
rect 458004 243098 458186 243334
rect 458422 243098 458604 243334
rect 458004 207654 458604 243098
rect 458004 207418 458186 207654
rect 458422 207418 458604 207654
rect 458004 207334 458604 207418
rect 458004 207098 458186 207334
rect 458422 207098 458604 207334
rect 458004 171654 458604 207098
rect 458004 171418 458186 171654
rect 458422 171418 458604 171654
rect 458004 171334 458604 171418
rect 458004 171098 458186 171334
rect 458422 171098 458604 171334
rect 458004 135654 458604 171098
rect 458004 135418 458186 135654
rect 458422 135418 458604 135654
rect 458004 135334 458604 135418
rect 458004 135098 458186 135334
rect 458422 135098 458604 135334
rect 458004 99654 458604 135098
rect 458004 99418 458186 99654
rect 458422 99418 458604 99654
rect 458004 99334 458604 99418
rect 458004 99098 458186 99334
rect 458422 99098 458604 99334
rect 458004 63654 458604 99098
rect 458004 63418 458186 63654
rect 458422 63418 458604 63654
rect 458004 63334 458604 63418
rect 458004 63098 458186 63334
rect 458422 63098 458604 63334
rect 458004 27654 458604 63098
rect 458004 27418 458186 27654
rect 458422 27418 458604 27654
rect 458004 27334 458604 27418
rect 458004 27098 458186 27334
rect 458422 27098 458604 27334
rect 458004 -4946 458604 27098
rect 458004 -5182 458186 -4946
rect 458422 -5182 458604 -4946
rect 458004 -5266 458604 -5182
rect 458004 -5502 458186 -5266
rect 458422 -5502 458604 -5266
rect 458004 -5524 458604 -5502
rect 461604 679254 462204 710722
rect 479604 710358 480204 711300
rect 479604 710122 479786 710358
rect 480022 710122 480204 710358
rect 479604 710038 480204 710122
rect 479604 709802 479786 710038
rect 480022 709802 480204 710038
rect 476004 708518 476604 709460
rect 476004 708282 476186 708518
rect 476422 708282 476604 708518
rect 476004 708198 476604 708282
rect 476004 707962 476186 708198
rect 476422 707962 476604 708198
rect 472404 706678 473004 707620
rect 472404 706442 472586 706678
rect 472822 706442 473004 706678
rect 472404 706358 473004 706442
rect 472404 706122 472586 706358
rect 472822 706122 473004 706358
rect 461604 679018 461786 679254
rect 462022 679018 462204 679254
rect 461604 678934 462204 679018
rect 461604 678698 461786 678934
rect 462022 678698 462204 678934
rect 461604 643254 462204 678698
rect 461604 643018 461786 643254
rect 462022 643018 462204 643254
rect 461604 642934 462204 643018
rect 461604 642698 461786 642934
rect 462022 642698 462204 642934
rect 461604 607254 462204 642698
rect 461604 607018 461786 607254
rect 462022 607018 462204 607254
rect 461604 606934 462204 607018
rect 461604 606698 461786 606934
rect 462022 606698 462204 606934
rect 461604 571254 462204 606698
rect 461604 571018 461786 571254
rect 462022 571018 462204 571254
rect 461604 570934 462204 571018
rect 461604 570698 461786 570934
rect 462022 570698 462204 570934
rect 461604 535254 462204 570698
rect 461604 535018 461786 535254
rect 462022 535018 462204 535254
rect 461604 534934 462204 535018
rect 461604 534698 461786 534934
rect 462022 534698 462204 534934
rect 461604 499254 462204 534698
rect 461604 499018 461786 499254
rect 462022 499018 462204 499254
rect 461604 498934 462204 499018
rect 461604 498698 461786 498934
rect 462022 498698 462204 498934
rect 461604 463254 462204 498698
rect 461604 463018 461786 463254
rect 462022 463018 462204 463254
rect 461604 462934 462204 463018
rect 461604 462698 461786 462934
rect 462022 462698 462204 462934
rect 461604 427254 462204 462698
rect 461604 427018 461786 427254
rect 462022 427018 462204 427254
rect 461604 426934 462204 427018
rect 461604 426698 461786 426934
rect 462022 426698 462204 426934
rect 461604 391254 462204 426698
rect 461604 391018 461786 391254
rect 462022 391018 462204 391254
rect 461604 390934 462204 391018
rect 461604 390698 461786 390934
rect 462022 390698 462204 390934
rect 461604 355254 462204 390698
rect 461604 355018 461786 355254
rect 462022 355018 462204 355254
rect 461604 354934 462204 355018
rect 461604 354698 461786 354934
rect 462022 354698 462204 354934
rect 461604 319254 462204 354698
rect 461604 319018 461786 319254
rect 462022 319018 462204 319254
rect 461604 318934 462204 319018
rect 461604 318698 461786 318934
rect 462022 318698 462204 318934
rect 461604 283254 462204 318698
rect 461604 283018 461786 283254
rect 462022 283018 462204 283254
rect 461604 282934 462204 283018
rect 461604 282698 461786 282934
rect 462022 282698 462204 282934
rect 461604 247254 462204 282698
rect 461604 247018 461786 247254
rect 462022 247018 462204 247254
rect 461604 246934 462204 247018
rect 461604 246698 461786 246934
rect 462022 246698 462204 246934
rect 461604 211254 462204 246698
rect 461604 211018 461786 211254
rect 462022 211018 462204 211254
rect 461604 210934 462204 211018
rect 461604 210698 461786 210934
rect 462022 210698 462204 210934
rect 461604 175254 462204 210698
rect 461604 175018 461786 175254
rect 462022 175018 462204 175254
rect 461604 174934 462204 175018
rect 461604 174698 461786 174934
rect 462022 174698 462204 174934
rect 461604 139254 462204 174698
rect 461604 139018 461786 139254
rect 462022 139018 462204 139254
rect 461604 138934 462204 139018
rect 461604 138698 461786 138934
rect 462022 138698 462204 138934
rect 461604 103254 462204 138698
rect 461604 103018 461786 103254
rect 462022 103018 462204 103254
rect 461604 102934 462204 103018
rect 461604 102698 461786 102934
rect 462022 102698 462204 102934
rect 461604 67254 462204 102698
rect 461604 67018 461786 67254
rect 462022 67018 462204 67254
rect 461604 66934 462204 67018
rect 461604 66698 461786 66934
rect 462022 66698 462204 66934
rect 461604 31254 462204 66698
rect 461604 31018 461786 31254
rect 462022 31018 462204 31254
rect 461604 30934 462204 31018
rect 461604 30698 461786 30934
rect 462022 30698 462204 30934
rect 443604 -6102 443786 -5866
rect 444022 -6102 444204 -5866
rect 443604 -6186 444204 -6102
rect 443604 -6422 443786 -6186
rect 444022 -6422 444204 -6186
rect 443604 -7364 444204 -6422
rect 461604 -6786 462204 30698
rect 468804 704838 469404 705780
rect 468804 704602 468986 704838
rect 469222 704602 469404 704838
rect 468804 704518 469404 704602
rect 468804 704282 468986 704518
rect 469222 704282 469404 704518
rect 468804 686454 469404 704282
rect 468804 686218 468986 686454
rect 469222 686218 469404 686454
rect 468804 686134 469404 686218
rect 468804 685898 468986 686134
rect 469222 685898 469404 686134
rect 468804 650454 469404 685898
rect 468804 650218 468986 650454
rect 469222 650218 469404 650454
rect 468804 650134 469404 650218
rect 468804 649898 468986 650134
rect 469222 649898 469404 650134
rect 468804 614454 469404 649898
rect 468804 614218 468986 614454
rect 469222 614218 469404 614454
rect 468804 614134 469404 614218
rect 468804 613898 468986 614134
rect 469222 613898 469404 614134
rect 468804 578454 469404 613898
rect 468804 578218 468986 578454
rect 469222 578218 469404 578454
rect 468804 578134 469404 578218
rect 468804 577898 468986 578134
rect 469222 577898 469404 578134
rect 468804 542454 469404 577898
rect 468804 542218 468986 542454
rect 469222 542218 469404 542454
rect 468804 542134 469404 542218
rect 468804 541898 468986 542134
rect 469222 541898 469404 542134
rect 468804 506454 469404 541898
rect 468804 506218 468986 506454
rect 469222 506218 469404 506454
rect 468804 506134 469404 506218
rect 468804 505898 468986 506134
rect 469222 505898 469404 506134
rect 468804 470454 469404 505898
rect 468804 470218 468986 470454
rect 469222 470218 469404 470454
rect 468804 470134 469404 470218
rect 468804 469898 468986 470134
rect 469222 469898 469404 470134
rect 468804 434454 469404 469898
rect 468804 434218 468986 434454
rect 469222 434218 469404 434454
rect 468804 434134 469404 434218
rect 468804 433898 468986 434134
rect 469222 433898 469404 434134
rect 468804 398454 469404 433898
rect 468804 398218 468986 398454
rect 469222 398218 469404 398454
rect 468804 398134 469404 398218
rect 468804 397898 468986 398134
rect 469222 397898 469404 398134
rect 468804 362454 469404 397898
rect 468804 362218 468986 362454
rect 469222 362218 469404 362454
rect 468804 362134 469404 362218
rect 468804 361898 468986 362134
rect 469222 361898 469404 362134
rect 468804 326454 469404 361898
rect 468804 326218 468986 326454
rect 469222 326218 469404 326454
rect 468804 326134 469404 326218
rect 468804 325898 468986 326134
rect 469222 325898 469404 326134
rect 468804 290454 469404 325898
rect 468804 290218 468986 290454
rect 469222 290218 469404 290454
rect 468804 290134 469404 290218
rect 468804 289898 468986 290134
rect 469222 289898 469404 290134
rect 468804 254454 469404 289898
rect 468804 254218 468986 254454
rect 469222 254218 469404 254454
rect 468804 254134 469404 254218
rect 468804 253898 468986 254134
rect 469222 253898 469404 254134
rect 468804 218454 469404 253898
rect 468804 218218 468986 218454
rect 469222 218218 469404 218454
rect 468804 218134 469404 218218
rect 468804 217898 468986 218134
rect 469222 217898 469404 218134
rect 468804 182454 469404 217898
rect 468804 182218 468986 182454
rect 469222 182218 469404 182454
rect 468804 182134 469404 182218
rect 468804 181898 468986 182134
rect 469222 181898 469404 182134
rect 468804 146454 469404 181898
rect 468804 146218 468986 146454
rect 469222 146218 469404 146454
rect 468804 146134 469404 146218
rect 468804 145898 468986 146134
rect 469222 145898 469404 146134
rect 468804 110454 469404 145898
rect 468804 110218 468986 110454
rect 469222 110218 469404 110454
rect 468804 110134 469404 110218
rect 468804 109898 468986 110134
rect 469222 109898 469404 110134
rect 468804 74454 469404 109898
rect 468804 74218 468986 74454
rect 469222 74218 469404 74454
rect 468804 74134 469404 74218
rect 468804 73898 468986 74134
rect 469222 73898 469404 74134
rect 468804 38454 469404 73898
rect 468804 38218 468986 38454
rect 469222 38218 469404 38454
rect 468804 38134 469404 38218
rect 468804 37898 468986 38134
rect 469222 37898 469404 38134
rect 468804 2454 469404 37898
rect 468804 2218 468986 2454
rect 469222 2218 469404 2454
rect 468804 2134 469404 2218
rect 468804 1898 468986 2134
rect 469222 1898 469404 2134
rect 468804 -346 469404 1898
rect 468804 -582 468986 -346
rect 469222 -582 469404 -346
rect 468804 -666 469404 -582
rect 468804 -902 468986 -666
rect 469222 -902 469404 -666
rect 468804 -1844 469404 -902
rect 472404 690054 473004 706122
rect 472404 689818 472586 690054
rect 472822 689818 473004 690054
rect 472404 689734 473004 689818
rect 472404 689498 472586 689734
rect 472822 689498 473004 689734
rect 472404 654054 473004 689498
rect 472404 653818 472586 654054
rect 472822 653818 473004 654054
rect 472404 653734 473004 653818
rect 472404 653498 472586 653734
rect 472822 653498 473004 653734
rect 472404 618054 473004 653498
rect 472404 617818 472586 618054
rect 472822 617818 473004 618054
rect 472404 617734 473004 617818
rect 472404 617498 472586 617734
rect 472822 617498 473004 617734
rect 472404 582054 473004 617498
rect 472404 581818 472586 582054
rect 472822 581818 473004 582054
rect 472404 581734 473004 581818
rect 472404 581498 472586 581734
rect 472822 581498 473004 581734
rect 472404 546054 473004 581498
rect 472404 545818 472586 546054
rect 472822 545818 473004 546054
rect 472404 545734 473004 545818
rect 472404 545498 472586 545734
rect 472822 545498 473004 545734
rect 472404 510054 473004 545498
rect 472404 509818 472586 510054
rect 472822 509818 473004 510054
rect 472404 509734 473004 509818
rect 472404 509498 472586 509734
rect 472822 509498 473004 509734
rect 472404 474054 473004 509498
rect 472404 473818 472586 474054
rect 472822 473818 473004 474054
rect 472404 473734 473004 473818
rect 472404 473498 472586 473734
rect 472822 473498 473004 473734
rect 472404 438054 473004 473498
rect 472404 437818 472586 438054
rect 472822 437818 473004 438054
rect 472404 437734 473004 437818
rect 472404 437498 472586 437734
rect 472822 437498 473004 437734
rect 472404 402054 473004 437498
rect 472404 401818 472586 402054
rect 472822 401818 473004 402054
rect 472404 401734 473004 401818
rect 472404 401498 472586 401734
rect 472822 401498 473004 401734
rect 472404 366054 473004 401498
rect 472404 365818 472586 366054
rect 472822 365818 473004 366054
rect 472404 365734 473004 365818
rect 472404 365498 472586 365734
rect 472822 365498 473004 365734
rect 472404 330054 473004 365498
rect 472404 329818 472586 330054
rect 472822 329818 473004 330054
rect 472404 329734 473004 329818
rect 472404 329498 472586 329734
rect 472822 329498 473004 329734
rect 472404 294054 473004 329498
rect 472404 293818 472586 294054
rect 472822 293818 473004 294054
rect 472404 293734 473004 293818
rect 472404 293498 472586 293734
rect 472822 293498 473004 293734
rect 472404 258054 473004 293498
rect 472404 257818 472586 258054
rect 472822 257818 473004 258054
rect 472404 257734 473004 257818
rect 472404 257498 472586 257734
rect 472822 257498 473004 257734
rect 472404 222054 473004 257498
rect 472404 221818 472586 222054
rect 472822 221818 473004 222054
rect 472404 221734 473004 221818
rect 472404 221498 472586 221734
rect 472822 221498 473004 221734
rect 472404 186054 473004 221498
rect 472404 185818 472586 186054
rect 472822 185818 473004 186054
rect 472404 185734 473004 185818
rect 472404 185498 472586 185734
rect 472822 185498 473004 185734
rect 472404 150054 473004 185498
rect 472404 149818 472586 150054
rect 472822 149818 473004 150054
rect 472404 149734 473004 149818
rect 472404 149498 472586 149734
rect 472822 149498 473004 149734
rect 472404 114054 473004 149498
rect 472404 113818 472586 114054
rect 472822 113818 473004 114054
rect 472404 113734 473004 113818
rect 472404 113498 472586 113734
rect 472822 113498 473004 113734
rect 472404 78054 473004 113498
rect 472404 77818 472586 78054
rect 472822 77818 473004 78054
rect 472404 77734 473004 77818
rect 472404 77498 472586 77734
rect 472822 77498 473004 77734
rect 472404 42054 473004 77498
rect 472404 41818 472586 42054
rect 472822 41818 473004 42054
rect 472404 41734 473004 41818
rect 472404 41498 472586 41734
rect 472822 41498 473004 41734
rect 472404 6054 473004 41498
rect 472404 5818 472586 6054
rect 472822 5818 473004 6054
rect 472404 5734 473004 5818
rect 472404 5498 472586 5734
rect 472822 5498 473004 5734
rect 472404 -2186 473004 5498
rect 472404 -2422 472586 -2186
rect 472822 -2422 473004 -2186
rect 472404 -2506 473004 -2422
rect 472404 -2742 472586 -2506
rect 472822 -2742 473004 -2506
rect 472404 -3684 473004 -2742
rect 476004 693654 476604 707962
rect 476004 693418 476186 693654
rect 476422 693418 476604 693654
rect 476004 693334 476604 693418
rect 476004 693098 476186 693334
rect 476422 693098 476604 693334
rect 476004 657654 476604 693098
rect 476004 657418 476186 657654
rect 476422 657418 476604 657654
rect 476004 657334 476604 657418
rect 476004 657098 476186 657334
rect 476422 657098 476604 657334
rect 476004 621654 476604 657098
rect 476004 621418 476186 621654
rect 476422 621418 476604 621654
rect 476004 621334 476604 621418
rect 476004 621098 476186 621334
rect 476422 621098 476604 621334
rect 476004 585654 476604 621098
rect 476004 585418 476186 585654
rect 476422 585418 476604 585654
rect 476004 585334 476604 585418
rect 476004 585098 476186 585334
rect 476422 585098 476604 585334
rect 476004 549654 476604 585098
rect 476004 549418 476186 549654
rect 476422 549418 476604 549654
rect 476004 549334 476604 549418
rect 476004 549098 476186 549334
rect 476422 549098 476604 549334
rect 476004 513654 476604 549098
rect 476004 513418 476186 513654
rect 476422 513418 476604 513654
rect 476004 513334 476604 513418
rect 476004 513098 476186 513334
rect 476422 513098 476604 513334
rect 476004 477654 476604 513098
rect 476004 477418 476186 477654
rect 476422 477418 476604 477654
rect 476004 477334 476604 477418
rect 476004 477098 476186 477334
rect 476422 477098 476604 477334
rect 476004 441654 476604 477098
rect 476004 441418 476186 441654
rect 476422 441418 476604 441654
rect 476004 441334 476604 441418
rect 476004 441098 476186 441334
rect 476422 441098 476604 441334
rect 476004 405654 476604 441098
rect 476004 405418 476186 405654
rect 476422 405418 476604 405654
rect 476004 405334 476604 405418
rect 476004 405098 476186 405334
rect 476422 405098 476604 405334
rect 476004 369654 476604 405098
rect 476004 369418 476186 369654
rect 476422 369418 476604 369654
rect 476004 369334 476604 369418
rect 476004 369098 476186 369334
rect 476422 369098 476604 369334
rect 476004 333654 476604 369098
rect 476004 333418 476186 333654
rect 476422 333418 476604 333654
rect 476004 333334 476604 333418
rect 476004 333098 476186 333334
rect 476422 333098 476604 333334
rect 476004 297654 476604 333098
rect 476004 297418 476186 297654
rect 476422 297418 476604 297654
rect 476004 297334 476604 297418
rect 476004 297098 476186 297334
rect 476422 297098 476604 297334
rect 476004 261654 476604 297098
rect 476004 261418 476186 261654
rect 476422 261418 476604 261654
rect 476004 261334 476604 261418
rect 476004 261098 476186 261334
rect 476422 261098 476604 261334
rect 476004 225654 476604 261098
rect 476004 225418 476186 225654
rect 476422 225418 476604 225654
rect 476004 225334 476604 225418
rect 476004 225098 476186 225334
rect 476422 225098 476604 225334
rect 476004 189654 476604 225098
rect 476004 189418 476186 189654
rect 476422 189418 476604 189654
rect 476004 189334 476604 189418
rect 476004 189098 476186 189334
rect 476422 189098 476604 189334
rect 476004 153654 476604 189098
rect 476004 153418 476186 153654
rect 476422 153418 476604 153654
rect 476004 153334 476604 153418
rect 476004 153098 476186 153334
rect 476422 153098 476604 153334
rect 476004 117654 476604 153098
rect 476004 117418 476186 117654
rect 476422 117418 476604 117654
rect 476004 117334 476604 117418
rect 476004 117098 476186 117334
rect 476422 117098 476604 117334
rect 476004 81654 476604 117098
rect 476004 81418 476186 81654
rect 476422 81418 476604 81654
rect 476004 81334 476604 81418
rect 476004 81098 476186 81334
rect 476422 81098 476604 81334
rect 476004 45654 476604 81098
rect 476004 45418 476186 45654
rect 476422 45418 476604 45654
rect 476004 45334 476604 45418
rect 476004 45098 476186 45334
rect 476422 45098 476604 45334
rect 476004 9654 476604 45098
rect 476004 9418 476186 9654
rect 476422 9418 476604 9654
rect 476004 9334 476604 9418
rect 476004 9098 476186 9334
rect 476422 9098 476604 9334
rect 476004 -4026 476604 9098
rect 476004 -4262 476186 -4026
rect 476422 -4262 476604 -4026
rect 476004 -4346 476604 -4262
rect 476004 -4582 476186 -4346
rect 476422 -4582 476604 -4346
rect 476004 -5524 476604 -4582
rect 479604 697254 480204 709802
rect 497604 711278 498204 711300
rect 497604 711042 497786 711278
rect 498022 711042 498204 711278
rect 497604 710958 498204 711042
rect 497604 710722 497786 710958
rect 498022 710722 498204 710958
rect 494004 709438 494604 709460
rect 494004 709202 494186 709438
rect 494422 709202 494604 709438
rect 494004 709118 494604 709202
rect 494004 708882 494186 709118
rect 494422 708882 494604 709118
rect 490404 707598 491004 707620
rect 490404 707362 490586 707598
rect 490822 707362 491004 707598
rect 490404 707278 491004 707362
rect 490404 707042 490586 707278
rect 490822 707042 491004 707278
rect 479604 697018 479786 697254
rect 480022 697018 480204 697254
rect 479604 696934 480204 697018
rect 479604 696698 479786 696934
rect 480022 696698 480204 696934
rect 479604 661254 480204 696698
rect 479604 661018 479786 661254
rect 480022 661018 480204 661254
rect 479604 660934 480204 661018
rect 479604 660698 479786 660934
rect 480022 660698 480204 660934
rect 479604 625254 480204 660698
rect 479604 625018 479786 625254
rect 480022 625018 480204 625254
rect 479604 624934 480204 625018
rect 479604 624698 479786 624934
rect 480022 624698 480204 624934
rect 479604 589254 480204 624698
rect 479604 589018 479786 589254
rect 480022 589018 480204 589254
rect 479604 588934 480204 589018
rect 479604 588698 479786 588934
rect 480022 588698 480204 588934
rect 479604 553254 480204 588698
rect 479604 553018 479786 553254
rect 480022 553018 480204 553254
rect 479604 552934 480204 553018
rect 479604 552698 479786 552934
rect 480022 552698 480204 552934
rect 479604 517254 480204 552698
rect 479604 517018 479786 517254
rect 480022 517018 480204 517254
rect 479604 516934 480204 517018
rect 479604 516698 479786 516934
rect 480022 516698 480204 516934
rect 479604 481254 480204 516698
rect 479604 481018 479786 481254
rect 480022 481018 480204 481254
rect 479604 480934 480204 481018
rect 479604 480698 479786 480934
rect 480022 480698 480204 480934
rect 479604 445254 480204 480698
rect 479604 445018 479786 445254
rect 480022 445018 480204 445254
rect 479604 444934 480204 445018
rect 479604 444698 479786 444934
rect 480022 444698 480204 444934
rect 479604 409254 480204 444698
rect 479604 409018 479786 409254
rect 480022 409018 480204 409254
rect 479604 408934 480204 409018
rect 479604 408698 479786 408934
rect 480022 408698 480204 408934
rect 479604 373254 480204 408698
rect 479604 373018 479786 373254
rect 480022 373018 480204 373254
rect 479604 372934 480204 373018
rect 479604 372698 479786 372934
rect 480022 372698 480204 372934
rect 479604 337254 480204 372698
rect 479604 337018 479786 337254
rect 480022 337018 480204 337254
rect 479604 336934 480204 337018
rect 479604 336698 479786 336934
rect 480022 336698 480204 336934
rect 479604 301254 480204 336698
rect 479604 301018 479786 301254
rect 480022 301018 480204 301254
rect 479604 300934 480204 301018
rect 479604 300698 479786 300934
rect 480022 300698 480204 300934
rect 479604 265254 480204 300698
rect 479604 265018 479786 265254
rect 480022 265018 480204 265254
rect 479604 264934 480204 265018
rect 479604 264698 479786 264934
rect 480022 264698 480204 264934
rect 479604 229254 480204 264698
rect 479604 229018 479786 229254
rect 480022 229018 480204 229254
rect 479604 228934 480204 229018
rect 479604 228698 479786 228934
rect 480022 228698 480204 228934
rect 479604 193254 480204 228698
rect 479604 193018 479786 193254
rect 480022 193018 480204 193254
rect 479604 192934 480204 193018
rect 479604 192698 479786 192934
rect 480022 192698 480204 192934
rect 479604 157254 480204 192698
rect 479604 157018 479786 157254
rect 480022 157018 480204 157254
rect 479604 156934 480204 157018
rect 479604 156698 479786 156934
rect 480022 156698 480204 156934
rect 479604 121254 480204 156698
rect 479604 121018 479786 121254
rect 480022 121018 480204 121254
rect 479604 120934 480204 121018
rect 479604 120698 479786 120934
rect 480022 120698 480204 120934
rect 479604 85254 480204 120698
rect 479604 85018 479786 85254
rect 480022 85018 480204 85254
rect 479604 84934 480204 85018
rect 479604 84698 479786 84934
rect 480022 84698 480204 84934
rect 479604 49254 480204 84698
rect 479604 49018 479786 49254
rect 480022 49018 480204 49254
rect 479604 48934 480204 49018
rect 479604 48698 479786 48934
rect 480022 48698 480204 48934
rect 479604 13254 480204 48698
rect 479604 13018 479786 13254
rect 480022 13018 480204 13254
rect 479604 12934 480204 13018
rect 479604 12698 479786 12934
rect 480022 12698 480204 12934
rect 461604 -7022 461786 -6786
rect 462022 -7022 462204 -6786
rect 461604 -7106 462204 -7022
rect 461604 -7342 461786 -7106
rect 462022 -7342 462204 -7106
rect 461604 -7364 462204 -7342
rect 479604 -5866 480204 12698
rect 486804 705758 487404 705780
rect 486804 705522 486986 705758
rect 487222 705522 487404 705758
rect 486804 705438 487404 705522
rect 486804 705202 486986 705438
rect 487222 705202 487404 705438
rect 486804 668454 487404 705202
rect 486804 668218 486986 668454
rect 487222 668218 487404 668454
rect 486804 668134 487404 668218
rect 486804 667898 486986 668134
rect 487222 667898 487404 668134
rect 486804 632454 487404 667898
rect 486804 632218 486986 632454
rect 487222 632218 487404 632454
rect 486804 632134 487404 632218
rect 486804 631898 486986 632134
rect 487222 631898 487404 632134
rect 486804 596454 487404 631898
rect 486804 596218 486986 596454
rect 487222 596218 487404 596454
rect 486804 596134 487404 596218
rect 486804 595898 486986 596134
rect 487222 595898 487404 596134
rect 486804 560454 487404 595898
rect 486804 560218 486986 560454
rect 487222 560218 487404 560454
rect 486804 560134 487404 560218
rect 486804 559898 486986 560134
rect 487222 559898 487404 560134
rect 486804 524454 487404 559898
rect 486804 524218 486986 524454
rect 487222 524218 487404 524454
rect 486804 524134 487404 524218
rect 486804 523898 486986 524134
rect 487222 523898 487404 524134
rect 486804 488454 487404 523898
rect 486804 488218 486986 488454
rect 487222 488218 487404 488454
rect 486804 488134 487404 488218
rect 486804 487898 486986 488134
rect 487222 487898 487404 488134
rect 486804 452454 487404 487898
rect 486804 452218 486986 452454
rect 487222 452218 487404 452454
rect 486804 452134 487404 452218
rect 486804 451898 486986 452134
rect 487222 451898 487404 452134
rect 486804 416454 487404 451898
rect 486804 416218 486986 416454
rect 487222 416218 487404 416454
rect 486804 416134 487404 416218
rect 486804 415898 486986 416134
rect 487222 415898 487404 416134
rect 486804 380454 487404 415898
rect 486804 380218 486986 380454
rect 487222 380218 487404 380454
rect 486804 380134 487404 380218
rect 486804 379898 486986 380134
rect 487222 379898 487404 380134
rect 486804 344454 487404 379898
rect 486804 344218 486986 344454
rect 487222 344218 487404 344454
rect 486804 344134 487404 344218
rect 486804 343898 486986 344134
rect 487222 343898 487404 344134
rect 486804 308454 487404 343898
rect 486804 308218 486986 308454
rect 487222 308218 487404 308454
rect 486804 308134 487404 308218
rect 486804 307898 486986 308134
rect 487222 307898 487404 308134
rect 486804 272454 487404 307898
rect 486804 272218 486986 272454
rect 487222 272218 487404 272454
rect 486804 272134 487404 272218
rect 486804 271898 486986 272134
rect 487222 271898 487404 272134
rect 486804 236454 487404 271898
rect 486804 236218 486986 236454
rect 487222 236218 487404 236454
rect 486804 236134 487404 236218
rect 486804 235898 486986 236134
rect 487222 235898 487404 236134
rect 486804 200454 487404 235898
rect 486804 200218 486986 200454
rect 487222 200218 487404 200454
rect 486804 200134 487404 200218
rect 486804 199898 486986 200134
rect 487222 199898 487404 200134
rect 486804 164454 487404 199898
rect 486804 164218 486986 164454
rect 487222 164218 487404 164454
rect 486804 164134 487404 164218
rect 486804 163898 486986 164134
rect 487222 163898 487404 164134
rect 486804 128454 487404 163898
rect 486804 128218 486986 128454
rect 487222 128218 487404 128454
rect 486804 128134 487404 128218
rect 486804 127898 486986 128134
rect 487222 127898 487404 128134
rect 486804 92454 487404 127898
rect 486804 92218 486986 92454
rect 487222 92218 487404 92454
rect 486804 92134 487404 92218
rect 486804 91898 486986 92134
rect 487222 91898 487404 92134
rect 486804 56454 487404 91898
rect 486804 56218 486986 56454
rect 487222 56218 487404 56454
rect 486804 56134 487404 56218
rect 486804 55898 486986 56134
rect 487222 55898 487404 56134
rect 486804 20454 487404 55898
rect 486804 20218 486986 20454
rect 487222 20218 487404 20454
rect 486804 20134 487404 20218
rect 486804 19898 486986 20134
rect 487222 19898 487404 20134
rect 486804 -1266 487404 19898
rect 486804 -1502 486986 -1266
rect 487222 -1502 487404 -1266
rect 486804 -1586 487404 -1502
rect 486804 -1822 486986 -1586
rect 487222 -1822 487404 -1586
rect 486804 -1844 487404 -1822
rect 490404 672054 491004 707042
rect 490404 671818 490586 672054
rect 490822 671818 491004 672054
rect 490404 671734 491004 671818
rect 490404 671498 490586 671734
rect 490822 671498 491004 671734
rect 490404 636054 491004 671498
rect 490404 635818 490586 636054
rect 490822 635818 491004 636054
rect 490404 635734 491004 635818
rect 490404 635498 490586 635734
rect 490822 635498 491004 635734
rect 490404 600054 491004 635498
rect 490404 599818 490586 600054
rect 490822 599818 491004 600054
rect 490404 599734 491004 599818
rect 490404 599498 490586 599734
rect 490822 599498 491004 599734
rect 490404 564054 491004 599498
rect 490404 563818 490586 564054
rect 490822 563818 491004 564054
rect 490404 563734 491004 563818
rect 490404 563498 490586 563734
rect 490822 563498 491004 563734
rect 490404 528054 491004 563498
rect 490404 527818 490586 528054
rect 490822 527818 491004 528054
rect 490404 527734 491004 527818
rect 490404 527498 490586 527734
rect 490822 527498 491004 527734
rect 490404 492054 491004 527498
rect 490404 491818 490586 492054
rect 490822 491818 491004 492054
rect 490404 491734 491004 491818
rect 490404 491498 490586 491734
rect 490822 491498 491004 491734
rect 490404 456054 491004 491498
rect 490404 455818 490586 456054
rect 490822 455818 491004 456054
rect 490404 455734 491004 455818
rect 490404 455498 490586 455734
rect 490822 455498 491004 455734
rect 490404 420054 491004 455498
rect 490404 419818 490586 420054
rect 490822 419818 491004 420054
rect 490404 419734 491004 419818
rect 490404 419498 490586 419734
rect 490822 419498 491004 419734
rect 490404 384054 491004 419498
rect 490404 383818 490586 384054
rect 490822 383818 491004 384054
rect 490404 383734 491004 383818
rect 490404 383498 490586 383734
rect 490822 383498 491004 383734
rect 490404 348054 491004 383498
rect 490404 347818 490586 348054
rect 490822 347818 491004 348054
rect 490404 347734 491004 347818
rect 490404 347498 490586 347734
rect 490822 347498 491004 347734
rect 490404 312054 491004 347498
rect 490404 311818 490586 312054
rect 490822 311818 491004 312054
rect 490404 311734 491004 311818
rect 490404 311498 490586 311734
rect 490822 311498 491004 311734
rect 490404 276054 491004 311498
rect 490404 275818 490586 276054
rect 490822 275818 491004 276054
rect 490404 275734 491004 275818
rect 490404 275498 490586 275734
rect 490822 275498 491004 275734
rect 490404 240054 491004 275498
rect 490404 239818 490586 240054
rect 490822 239818 491004 240054
rect 490404 239734 491004 239818
rect 490404 239498 490586 239734
rect 490822 239498 491004 239734
rect 490404 204054 491004 239498
rect 490404 203818 490586 204054
rect 490822 203818 491004 204054
rect 490404 203734 491004 203818
rect 490404 203498 490586 203734
rect 490822 203498 491004 203734
rect 490404 168054 491004 203498
rect 490404 167818 490586 168054
rect 490822 167818 491004 168054
rect 490404 167734 491004 167818
rect 490404 167498 490586 167734
rect 490822 167498 491004 167734
rect 490404 132054 491004 167498
rect 490404 131818 490586 132054
rect 490822 131818 491004 132054
rect 490404 131734 491004 131818
rect 490404 131498 490586 131734
rect 490822 131498 491004 131734
rect 490404 96054 491004 131498
rect 490404 95818 490586 96054
rect 490822 95818 491004 96054
rect 490404 95734 491004 95818
rect 490404 95498 490586 95734
rect 490822 95498 491004 95734
rect 490404 60054 491004 95498
rect 494004 675654 494604 708882
rect 494004 675418 494186 675654
rect 494422 675418 494604 675654
rect 494004 675334 494604 675418
rect 494004 675098 494186 675334
rect 494422 675098 494604 675334
rect 494004 639654 494604 675098
rect 494004 639418 494186 639654
rect 494422 639418 494604 639654
rect 494004 639334 494604 639418
rect 494004 639098 494186 639334
rect 494422 639098 494604 639334
rect 494004 603654 494604 639098
rect 494004 603418 494186 603654
rect 494422 603418 494604 603654
rect 494004 603334 494604 603418
rect 494004 603098 494186 603334
rect 494422 603098 494604 603334
rect 494004 567654 494604 603098
rect 494004 567418 494186 567654
rect 494422 567418 494604 567654
rect 494004 567334 494604 567418
rect 494004 567098 494186 567334
rect 494422 567098 494604 567334
rect 494004 531654 494604 567098
rect 494004 531418 494186 531654
rect 494422 531418 494604 531654
rect 494004 531334 494604 531418
rect 494004 531098 494186 531334
rect 494422 531098 494604 531334
rect 494004 495654 494604 531098
rect 494004 495418 494186 495654
rect 494422 495418 494604 495654
rect 494004 495334 494604 495418
rect 494004 495098 494186 495334
rect 494422 495098 494604 495334
rect 494004 459654 494604 495098
rect 494004 459418 494186 459654
rect 494422 459418 494604 459654
rect 494004 459334 494604 459418
rect 494004 459098 494186 459334
rect 494422 459098 494604 459334
rect 494004 423654 494604 459098
rect 494004 423418 494186 423654
rect 494422 423418 494604 423654
rect 494004 423334 494604 423418
rect 494004 423098 494186 423334
rect 494422 423098 494604 423334
rect 494004 387654 494604 423098
rect 494004 387418 494186 387654
rect 494422 387418 494604 387654
rect 494004 387334 494604 387418
rect 494004 387098 494186 387334
rect 494422 387098 494604 387334
rect 494004 351654 494604 387098
rect 494004 351418 494186 351654
rect 494422 351418 494604 351654
rect 494004 351334 494604 351418
rect 494004 351098 494186 351334
rect 494422 351098 494604 351334
rect 494004 315654 494604 351098
rect 494004 315418 494186 315654
rect 494422 315418 494604 315654
rect 494004 315334 494604 315418
rect 494004 315098 494186 315334
rect 494422 315098 494604 315334
rect 494004 279654 494604 315098
rect 494004 279418 494186 279654
rect 494422 279418 494604 279654
rect 494004 279334 494604 279418
rect 494004 279098 494186 279334
rect 494422 279098 494604 279334
rect 494004 243654 494604 279098
rect 494004 243418 494186 243654
rect 494422 243418 494604 243654
rect 494004 243334 494604 243418
rect 494004 243098 494186 243334
rect 494422 243098 494604 243334
rect 494004 207654 494604 243098
rect 494004 207418 494186 207654
rect 494422 207418 494604 207654
rect 494004 207334 494604 207418
rect 494004 207098 494186 207334
rect 494422 207098 494604 207334
rect 494004 171654 494604 207098
rect 494004 171418 494186 171654
rect 494422 171418 494604 171654
rect 494004 171334 494604 171418
rect 494004 171098 494186 171334
rect 494422 171098 494604 171334
rect 494004 135654 494604 171098
rect 494004 135418 494186 135654
rect 494422 135418 494604 135654
rect 494004 135334 494604 135418
rect 494004 135098 494186 135334
rect 494422 135098 494604 135334
rect 494004 99654 494604 135098
rect 494004 99418 494186 99654
rect 494422 99418 494604 99654
rect 494004 99334 494604 99418
rect 494004 99098 494186 99334
rect 494422 99098 494604 99334
rect 492627 76124 492693 76125
rect 492627 76060 492628 76124
rect 492692 76060 492693 76124
rect 492627 76059 492693 76060
rect 492630 75853 492690 76059
rect 492627 75852 492693 75853
rect 492627 75788 492628 75852
rect 492692 75788 492693 75852
rect 492627 75787 492693 75788
rect 490404 59818 490586 60054
rect 490822 59818 491004 60054
rect 490404 59734 491004 59818
rect 490404 59498 490586 59734
rect 490822 59498 491004 59734
rect 490404 24054 491004 59498
rect 490404 23818 490586 24054
rect 490822 23818 491004 24054
rect 490404 23734 491004 23818
rect 490404 23498 490586 23734
rect 490822 23498 491004 23734
rect 490404 -3106 491004 23498
rect 490404 -3342 490586 -3106
rect 490822 -3342 491004 -3106
rect 490404 -3426 491004 -3342
rect 490404 -3662 490586 -3426
rect 490822 -3662 491004 -3426
rect 490404 -3684 491004 -3662
rect 494004 63654 494604 99098
rect 494004 63418 494186 63654
rect 494422 63418 494604 63654
rect 494004 63334 494604 63418
rect 494004 63098 494186 63334
rect 494422 63098 494604 63334
rect 494004 27654 494604 63098
rect 494004 27418 494186 27654
rect 494422 27418 494604 27654
rect 494004 27334 494604 27418
rect 494004 27098 494186 27334
rect 494422 27098 494604 27334
rect 494004 -4946 494604 27098
rect 494004 -5182 494186 -4946
rect 494422 -5182 494604 -4946
rect 494004 -5266 494604 -5182
rect 494004 -5502 494186 -5266
rect 494422 -5502 494604 -5266
rect 494004 -5524 494604 -5502
rect 497604 679254 498204 710722
rect 515604 710358 516204 711300
rect 515604 710122 515786 710358
rect 516022 710122 516204 710358
rect 515604 710038 516204 710122
rect 515604 709802 515786 710038
rect 516022 709802 516204 710038
rect 512004 708518 512604 709460
rect 512004 708282 512186 708518
rect 512422 708282 512604 708518
rect 512004 708198 512604 708282
rect 512004 707962 512186 708198
rect 512422 707962 512604 708198
rect 508404 706678 509004 707620
rect 508404 706442 508586 706678
rect 508822 706442 509004 706678
rect 508404 706358 509004 706442
rect 508404 706122 508586 706358
rect 508822 706122 509004 706358
rect 497604 679018 497786 679254
rect 498022 679018 498204 679254
rect 497604 678934 498204 679018
rect 497604 678698 497786 678934
rect 498022 678698 498204 678934
rect 497604 643254 498204 678698
rect 497604 643018 497786 643254
rect 498022 643018 498204 643254
rect 497604 642934 498204 643018
rect 497604 642698 497786 642934
rect 498022 642698 498204 642934
rect 497604 607254 498204 642698
rect 497604 607018 497786 607254
rect 498022 607018 498204 607254
rect 497604 606934 498204 607018
rect 497604 606698 497786 606934
rect 498022 606698 498204 606934
rect 497604 571254 498204 606698
rect 497604 571018 497786 571254
rect 498022 571018 498204 571254
rect 497604 570934 498204 571018
rect 497604 570698 497786 570934
rect 498022 570698 498204 570934
rect 497604 535254 498204 570698
rect 497604 535018 497786 535254
rect 498022 535018 498204 535254
rect 497604 534934 498204 535018
rect 497604 534698 497786 534934
rect 498022 534698 498204 534934
rect 497604 499254 498204 534698
rect 497604 499018 497786 499254
rect 498022 499018 498204 499254
rect 497604 498934 498204 499018
rect 497604 498698 497786 498934
rect 498022 498698 498204 498934
rect 497604 463254 498204 498698
rect 497604 463018 497786 463254
rect 498022 463018 498204 463254
rect 497604 462934 498204 463018
rect 497604 462698 497786 462934
rect 498022 462698 498204 462934
rect 497604 427254 498204 462698
rect 497604 427018 497786 427254
rect 498022 427018 498204 427254
rect 497604 426934 498204 427018
rect 497604 426698 497786 426934
rect 498022 426698 498204 426934
rect 497604 391254 498204 426698
rect 497604 391018 497786 391254
rect 498022 391018 498204 391254
rect 497604 390934 498204 391018
rect 497604 390698 497786 390934
rect 498022 390698 498204 390934
rect 497604 355254 498204 390698
rect 497604 355018 497786 355254
rect 498022 355018 498204 355254
rect 497604 354934 498204 355018
rect 497604 354698 497786 354934
rect 498022 354698 498204 354934
rect 497604 319254 498204 354698
rect 497604 319018 497786 319254
rect 498022 319018 498204 319254
rect 497604 318934 498204 319018
rect 497604 318698 497786 318934
rect 498022 318698 498204 318934
rect 497604 283254 498204 318698
rect 497604 283018 497786 283254
rect 498022 283018 498204 283254
rect 497604 282934 498204 283018
rect 497604 282698 497786 282934
rect 498022 282698 498204 282934
rect 497604 247254 498204 282698
rect 497604 247018 497786 247254
rect 498022 247018 498204 247254
rect 497604 246934 498204 247018
rect 497604 246698 497786 246934
rect 498022 246698 498204 246934
rect 497604 211254 498204 246698
rect 497604 211018 497786 211254
rect 498022 211018 498204 211254
rect 497604 210934 498204 211018
rect 497604 210698 497786 210934
rect 498022 210698 498204 210934
rect 497604 175254 498204 210698
rect 497604 175018 497786 175254
rect 498022 175018 498204 175254
rect 497604 174934 498204 175018
rect 497604 174698 497786 174934
rect 498022 174698 498204 174934
rect 497604 139254 498204 174698
rect 497604 139018 497786 139254
rect 498022 139018 498204 139254
rect 497604 138934 498204 139018
rect 497604 138698 497786 138934
rect 498022 138698 498204 138934
rect 497604 103254 498204 138698
rect 497604 103018 497786 103254
rect 498022 103018 498204 103254
rect 497604 102934 498204 103018
rect 497604 102698 497786 102934
rect 498022 102698 498204 102934
rect 497604 67254 498204 102698
rect 497604 67018 497786 67254
rect 498022 67018 498204 67254
rect 497604 66934 498204 67018
rect 497604 66698 497786 66934
rect 498022 66698 498204 66934
rect 497604 31254 498204 66698
rect 497604 31018 497786 31254
rect 498022 31018 498204 31254
rect 497604 30934 498204 31018
rect 497604 30698 497786 30934
rect 498022 30698 498204 30934
rect 479604 -6102 479786 -5866
rect 480022 -6102 480204 -5866
rect 479604 -6186 480204 -6102
rect 479604 -6422 479786 -6186
rect 480022 -6422 480204 -6186
rect 479604 -7364 480204 -6422
rect 497604 -6786 498204 30698
rect 504804 704838 505404 705780
rect 504804 704602 504986 704838
rect 505222 704602 505404 704838
rect 504804 704518 505404 704602
rect 504804 704282 504986 704518
rect 505222 704282 505404 704518
rect 504804 686454 505404 704282
rect 504804 686218 504986 686454
rect 505222 686218 505404 686454
rect 504804 686134 505404 686218
rect 504804 685898 504986 686134
rect 505222 685898 505404 686134
rect 504804 650454 505404 685898
rect 504804 650218 504986 650454
rect 505222 650218 505404 650454
rect 504804 650134 505404 650218
rect 504804 649898 504986 650134
rect 505222 649898 505404 650134
rect 504804 614454 505404 649898
rect 504804 614218 504986 614454
rect 505222 614218 505404 614454
rect 504804 614134 505404 614218
rect 504804 613898 504986 614134
rect 505222 613898 505404 614134
rect 504804 578454 505404 613898
rect 504804 578218 504986 578454
rect 505222 578218 505404 578454
rect 504804 578134 505404 578218
rect 504804 577898 504986 578134
rect 505222 577898 505404 578134
rect 504804 542454 505404 577898
rect 504804 542218 504986 542454
rect 505222 542218 505404 542454
rect 504804 542134 505404 542218
rect 504804 541898 504986 542134
rect 505222 541898 505404 542134
rect 504804 506454 505404 541898
rect 504804 506218 504986 506454
rect 505222 506218 505404 506454
rect 504804 506134 505404 506218
rect 504804 505898 504986 506134
rect 505222 505898 505404 506134
rect 504804 470454 505404 505898
rect 504804 470218 504986 470454
rect 505222 470218 505404 470454
rect 504804 470134 505404 470218
rect 504804 469898 504986 470134
rect 505222 469898 505404 470134
rect 504804 434454 505404 469898
rect 504804 434218 504986 434454
rect 505222 434218 505404 434454
rect 504804 434134 505404 434218
rect 504804 433898 504986 434134
rect 505222 433898 505404 434134
rect 504804 398454 505404 433898
rect 504804 398218 504986 398454
rect 505222 398218 505404 398454
rect 504804 398134 505404 398218
rect 504804 397898 504986 398134
rect 505222 397898 505404 398134
rect 504804 362454 505404 397898
rect 504804 362218 504986 362454
rect 505222 362218 505404 362454
rect 504804 362134 505404 362218
rect 504804 361898 504986 362134
rect 505222 361898 505404 362134
rect 504804 326454 505404 361898
rect 504804 326218 504986 326454
rect 505222 326218 505404 326454
rect 504804 326134 505404 326218
rect 504804 325898 504986 326134
rect 505222 325898 505404 326134
rect 504804 290454 505404 325898
rect 504804 290218 504986 290454
rect 505222 290218 505404 290454
rect 504804 290134 505404 290218
rect 504804 289898 504986 290134
rect 505222 289898 505404 290134
rect 504804 254454 505404 289898
rect 504804 254218 504986 254454
rect 505222 254218 505404 254454
rect 504804 254134 505404 254218
rect 504804 253898 504986 254134
rect 505222 253898 505404 254134
rect 504804 218454 505404 253898
rect 504804 218218 504986 218454
rect 505222 218218 505404 218454
rect 504804 218134 505404 218218
rect 504804 217898 504986 218134
rect 505222 217898 505404 218134
rect 504804 182454 505404 217898
rect 504804 182218 504986 182454
rect 505222 182218 505404 182454
rect 504804 182134 505404 182218
rect 504804 181898 504986 182134
rect 505222 181898 505404 182134
rect 504804 146454 505404 181898
rect 504804 146218 504986 146454
rect 505222 146218 505404 146454
rect 504804 146134 505404 146218
rect 504804 145898 504986 146134
rect 505222 145898 505404 146134
rect 504804 110454 505404 145898
rect 504804 110218 504986 110454
rect 505222 110218 505404 110454
rect 504804 110134 505404 110218
rect 504804 109898 504986 110134
rect 505222 109898 505404 110134
rect 504804 74454 505404 109898
rect 504804 74218 504986 74454
rect 505222 74218 505404 74454
rect 504804 74134 505404 74218
rect 504804 73898 504986 74134
rect 505222 73898 505404 74134
rect 504804 38454 505404 73898
rect 504804 38218 504986 38454
rect 505222 38218 505404 38454
rect 504804 38134 505404 38218
rect 504804 37898 504986 38134
rect 505222 37898 505404 38134
rect 504804 2454 505404 37898
rect 504804 2218 504986 2454
rect 505222 2218 505404 2454
rect 504804 2134 505404 2218
rect 504804 1898 504986 2134
rect 505222 1898 505404 2134
rect 504804 -346 505404 1898
rect 504804 -582 504986 -346
rect 505222 -582 505404 -346
rect 504804 -666 505404 -582
rect 504804 -902 504986 -666
rect 505222 -902 505404 -666
rect 504804 -1844 505404 -902
rect 508404 690054 509004 706122
rect 508404 689818 508586 690054
rect 508822 689818 509004 690054
rect 508404 689734 509004 689818
rect 508404 689498 508586 689734
rect 508822 689498 509004 689734
rect 508404 654054 509004 689498
rect 508404 653818 508586 654054
rect 508822 653818 509004 654054
rect 508404 653734 509004 653818
rect 508404 653498 508586 653734
rect 508822 653498 509004 653734
rect 508404 618054 509004 653498
rect 508404 617818 508586 618054
rect 508822 617818 509004 618054
rect 508404 617734 509004 617818
rect 508404 617498 508586 617734
rect 508822 617498 509004 617734
rect 508404 582054 509004 617498
rect 508404 581818 508586 582054
rect 508822 581818 509004 582054
rect 508404 581734 509004 581818
rect 508404 581498 508586 581734
rect 508822 581498 509004 581734
rect 508404 546054 509004 581498
rect 508404 545818 508586 546054
rect 508822 545818 509004 546054
rect 508404 545734 509004 545818
rect 508404 545498 508586 545734
rect 508822 545498 509004 545734
rect 508404 510054 509004 545498
rect 508404 509818 508586 510054
rect 508822 509818 509004 510054
rect 508404 509734 509004 509818
rect 508404 509498 508586 509734
rect 508822 509498 509004 509734
rect 508404 474054 509004 509498
rect 508404 473818 508586 474054
rect 508822 473818 509004 474054
rect 508404 473734 509004 473818
rect 508404 473498 508586 473734
rect 508822 473498 509004 473734
rect 508404 438054 509004 473498
rect 508404 437818 508586 438054
rect 508822 437818 509004 438054
rect 508404 437734 509004 437818
rect 508404 437498 508586 437734
rect 508822 437498 509004 437734
rect 508404 402054 509004 437498
rect 508404 401818 508586 402054
rect 508822 401818 509004 402054
rect 508404 401734 509004 401818
rect 508404 401498 508586 401734
rect 508822 401498 509004 401734
rect 508404 366054 509004 401498
rect 508404 365818 508586 366054
rect 508822 365818 509004 366054
rect 508404 365734 509004 365818
rect 508404 365498 508586 365734
rect 508822 365498 509004 365734
rect 508404 330054 509004 365498
rect 508404 329818 508586 330054
rect 508822 329818 509004 330054
rect 508404 329734 509004 329818
rect 508404 329498 508586 329734
rect 508822 329498 509004 329734
rect 508404 294054 509004 329498
rect 508404 293818 508586 294054
rect 508822 293818 509004 294054
rect 508404 293734 509004 293818
rect 508404 293498 508586 293734
rect 508822 293498 509004 293734
rect 508404 258054 509004 293498
rect 508404 257818 508586 258054
rect 508822 257818 509004 258054
rect 508404 257734 509004 257818
rect 508404 257498 508586 257734
rect 508822 257498 509004 257734
rect 508404 222054 509004 257498
rect 508404 221818 508586 222054
rect 508822 221818 509004 222054
rect 508404 221734 509004 221818
rect 508404 221498 508586 221734
rect 508822 221498 509004 221734
rect 508404 186054 509004 221498
rect 508404 185818 508586 186054
rect 508822 185818 509004 186054
rect 508404 185734 509004 185818
rect 508404 185498 508586 185734
rect 508822 185498 509004 185734
rect 508404 150054 509004 185498
rect 508404 149818 508586 150054
rect 508822 149818 509004 150054
rect 508404 149734 509004 149818
rect 508404 149498 508586 149734
rect 508822 149498 509004 149734
rect 508404 114054 509004 149498
rect 508404 113818 508586 114054
rect 508822 113818 509004 114054
rect 508404 113734 509004 113818
rect 508404 113498 508586 113734
rect 508822 113498 509004 113734
rect 508404 78054 509004 113498
rect 508404 77818 508586 78054
rect 508822 77818 509004 78054
rect 508404 77734 509004 77818
rect 508404 77498 508586 77734
rect 508822 77498 509004 77734
rect 508404 42054 509004 77498
rect 508404 41818 508586 42054
rect 508822 41818 509004 42054
rect 508404 41734 509004 41818
rect 508404 41498 508586 41734
rect 508822 41498 509004 41734
rect 508404 6054 509004 41498
rect 508404 5818 508586 6054
rect 508822 5818 509004 6054
rect 508404 5734 509004 5818
rect 508404 5498 508586 5734
rect 508822 5498 509004 5734
rect 508404 -2186 509004 5498
rect 508404 -2422 508586 -2186
rect 508822 -2422 509004 -2186
rect 508404 -2506 509004 -2422
rect 508404 -2742 508586 -2506
rect 508822 -2742 509004 -2506
rect 508404 -3684 509004 -2742
rect 512004 693654 512604 707962
rect 512004 693418 512186 693654
rect 512422 693418 512604 693654
rect 512004 693334 512604 693418
rect 512004 693098 512186 693334
rect 512422 693098 512604 693334
rect 512004 657654 512604 693098
rect 512004 657418 512186 657654
rect 512422 657418 512604 657654
rect 512004 657334 512604 657418
rect 512004 657098 512186 657334
rect 512422 657098 512604 657334
rect 512004 621654 512604 657098
rect 512004 621418 512186 621654
rect 512422 621418 512604 621654
rect 512004 621334 512604 621418
rect 512004 621098 512186 621334
rect 512422 621098 512604 621334
rect 512004 585654 512604 621098
rect 512004 585418 512186 585654
rect 512422 585418 512604 585654
rect 512004 585334 512604 585418
rect 512004 585098 512186 585334
rect 512422 585098 512604 585334
rect 512004 549654 512604 585098
rect 512004 549418 512186 549654
rect 512422 549418 512604 549654
rect 512004 549334 512604 549418
rect 512004 549098 512186 549334
rect 512422 549098 512604 549334
rect 512004 513654 512604 549098
rect 512004 513418 512186 513654
rect 512422 513418 512604 513654
rect 512004 513334 512604 513418
rect 512004 513098 512186 513334
rect 512422 513098 512604 513334
rect 512004 477654 512604 513098
rect 512004 477418 512186 477654
rect 512422 477418 512604 477654
rect 512004 477334 512604 477418
rect 512004 477098 512186 477334
rect 512422 477098 512604 477334
rect 512004 441654 512604 477098
rect 512004 441418 512186 441654
rect 512422 441418 512604 441654
rect 512004 441334 512604 441418
rect 512004 441098 512186 441334
rect 512422 441098 512604 441334
rect 512004 405654 512604 441098
rect 512004 405418 512186 405654
rect 512422 405418 512604 405654
rect 512004 405334 512604 405418
rect 512004 405098 512186 405334
rect 512422 405098 512604 405334
rect 512004 369654 512604 405098
rect 512004 369418 512186 369654
rect 512422 369418 512604 369654
rect 512004 369334 512604 369418
rect 512004 369098 512186 369334
rect 512422 369098 512604 369334
rect 512004 333654 512604 369098
rect 512004 333418 512186 333654
rect 512422 333418 512604 333654
rect 512004 333334 512604 333418
rect 512004 333098 512186 333334
rect 512422 333098 512604 333334
rect 512004 297654 512604 333098
rect 512004 297418 512186 297654
rect 512422 297418 512604 297654
rect 512004 297334 512604 297418
rect 512004 297098 512186 297334
rect 512422 297098 512604 297334
rect 512004 261654 512604 297098
rect 512004 261418 512186 261654
rect 512422 261418 512604 261654
rect 512004 261334 512604 261418
rect 512004 261098 512186 261334
rect 512422 261098 512604 261334
rect 512004 225654 512604 261098
rect 512004 225418 512186 225654
rect 512422 225418 512604 225654
rect 512004 225334 512604 225418
rect 512004 225098 512186 225334
rect 512422 225098 512604 225334
rect 512004 189654 512604 225098
rect 512004 189418 512186 189654
rect 512422 189418 512604 189654
rect 512004 189334 512604 189418
rect 512004 189098 512186 189334
rect 512422 189098 512604 189334
rect 512004 153654 512604 189098
rect 512004 153418 512186 153654
rect 512422 153418 512604 153654
rect 512004 153334 512604 153418
rect 512004 153098 512186 153334
rect 512422 153098 512604 153334
rect 512004 117654 512604 153098
rect 512004 117418 512186 117654
rect 512422 117418 512604 117654
rect 512004 117334 512604 117418
rect 512004 117098 512186 117334
rect 512422 117098 512604 117334
rect 512004 81654 512604 117098
rect 512004 81418 512186 81654
rect 512422 81418 512604 81654
rect 512004 81334 512604 81418
rect 512004 81098 512186 81334
rect 512422 81098 512604 81334
rect 512004 45654 512604 81098
rect 512004 45418 512186 45654
rect 512422 45418 512604 45654
rect 512004 45334 512604 45418
rect 512004 45098 512186 45334
rect 512422 45098 512604 45334
rect 512004 9654 512604 45098
rect 512004 9418 512186 9654
rect 512422 9418 512604 9654
rect 512004 9334 512604 9418
rect 512004 9098 512186 9334
rect 512422 9098 512604 9334
rect 512004 -4026 512604 9098
rect 512004 -4262 512186 -4026
rect 512422 -4262 512604 -4026
rect 512004 -4346 512604 -4262
rect 512004 -4582 512186 -4346
rect 512422 -4582 512604 -4346
rect 512004 -5524 512604 -4582
rect 515604 697254 516204 709802
rect 533604 711278 534204 711300
rect 533604 711042 533786 711278
rect 534022 711042 534204 711278
rect 533604 710958 534204 711042
rect 533604 710722 533786 710958
rect 534022 710722 534204 710958
rect 530004 709438 530604 709460
rect 530004 709202 530186 709438
rect 530422 709202 530604 709438
rect 530004 709118 530604 709202
rect 530004 708882 530186 709118
rect 530422 708882 530604 709118
rect 526404 707598 527004 707620
rect 526404 707362 526586 707598
rect 526822 707362 527004 707598
rect 526404 707278 527004 707362
rect 526404 707042 526586 707278
rect 526822 707042 527004 707278
rect 515604 697018 515786 697254
rect 516022 697018 516204 697254
rect 515604 696934 516204 697018
rect 515604 696698 515786 696934
rect 516022 696698 516204 696934
rect 515604 661254 516204 696698
rect 515604 661018 515786 661254
rect 516022 661018 516204 661254
rect 515604 660934 516204 661018
rect 515604 660698 515786 660934
rect 516022 660698 516204 660934
rect 515604 625254 516204 660698
rect 515604 625018 515786 625254
rect 516022 625018 516204 625254
rect 515604 624934 516204 625018
rect 515604 624698 515786 624934
rect 516022 624698 516204 624934
rect 515604 589254 516204 624698
rect 515604 589018 515786 589254
rect 516022 589018 516204 589254
rect 515604 588934 516204 589018
rect 515604 588698 515786 588934
rect 516022 588698 516204 588934
rect 515604 553254 516204 588698
rect 515604 553018 515786 553254
rect 516022 553018 516204 553254
rect 515604 552934 516204 553018
rect 515604 552698 515786 552934
rect 516022 552698 516204 552934
rect 515604 517254 516204 552698
rect 515604 517018 515786 517254
rect 516022 517018 516204 517254
rect 515604 516934 516204 517018
rect 515604 516698 515786 516934
rect 516022 516698 516204 516934
rect 515604 481254 516204 516698
rect 515604 481018 515786 481254
rect 516022 481018 516204 481254
rect 515604 480934 516204 481018
rect 515604 480698 515786 480934
rect 516022 480698 516204 480934
rect 515604 445254 516204 480698
rect 515604 445018 515786 445254
rect 516022 445018 516204 445254
rect 515604 444934 516204 445018
rect 515604 444698 515786 444934
rect 516022 444698 516204 444934
rect 515604 409254 516204 444698
rect 515604 409018 515786 409254
rect 516022 409018 516204 409254
rect 515604 408934 516204 409018
rect 515604 408698 515786 408934
rect 516022 408698 516204 408934
rect 515604 373254 516204 408698
rect 515604 373018 515786 373254
rect 516022 373018 516204 373254
rect 515604 372934 516204 373018
rect 515604 372698 515786 372934
rect 516022 372698 516204 372934
rect 515604 337254 516204 372698
rect 515604 337018 515786 337254
rect 516022 337018 516204 337254
rect 515604 336934 516204 337018
rect 515604 336698 515786 336934
rect 516022 336698 516204 336934
rect 515604 301254 516204 336698
rect 515604 301018 515786 301254
rect 516022 301018 516204 301254
rect 515604 300934 516204 301018
rect 515604 300698 515786 300934
rect 516022 300698 516204 300934
rect 515604 265254 516204 300698
rect 515604 265018 515786 265254
rect 516022 265018 516204 265254
rect 515604 264934 516204 265018
rect 515604 264698 515786 264934
rect 516022 264698 516204 264934
rect 515604 229254 516204 264698
rect 515604 229018 515786 229254
rect 516022 229018 516204 229254
rect 515604 228934 516204 229018
rect 515604 228698 515786 228934
rect 516022 228698 516204 228934
rect 515604 193254 516204 228698
rect 515604 193018 515786 193254
rect 516022 193018 516204 193254
rect 515604 192934 516204 193018
rect 515604 192698 515786 192934
rect 516022 192698 516204 192934
rect 515604 157254 516204 192698
rect 515604 157018 515786 157254
rect 516022 157018 516204 157254
rect 515604 156934 516204 157018
rect 515604 156698 515786 156934
rect 516022 156698 516204 156934
rect 515604 121254 516204 156698
rect 515604 121018 515786 121254
rect 516022 121018 516204 121254
rect 515604 120934 516204 121018
rect 515604 120698 515786 120934
rect 516022 120698 516204 120934
rect 515604 85254 516204 120698
rect 515604 85018 515786 85254
rect 516022 85018 516204 85254
rect 515604 84934 516204 85018
rect 515604 84698 515786 84934
rect 516022 84698 516204 84934
rect 515604 49254 516204 84698
rect 515604 49018 515786 49254
rect 516022 49018 516204 49254
rect 515604 48934 516204 49018
rect 515604 48698 515786 48934
rect 516022 48698 516204 48934
rect 515604 13254 516204 48698
rect 515604 13018 515786 13254
rect 516022 13018 516204 13254
rect 515604 12934 516204 13018
rect 515604 12698 515786 12934
rect 516022 12698 516204 12934
rect 497604 -7022 497786 -6786
rect 498022 -7022 498204 -6786
rect 497604 -7106 498204 -7022
rect 497604 -7342 497786 -7106
rect 498022 -7342 498204 -7106
rect 497604 -7364 498204 -7342
rect 515604 -5866 516204 12698
rect 522804 705758 523404 705780
rect 522804 705522 522986 705758
rect 523222 705522 523404 705758
rect 522804 705438 523404 705522
rect 522804 705202 522986 705438
rect 523222 705202 523404 705438
rect 522804 668454 523404 705202
rect 522804 668218 522986 668454
rect 523222 668218 523404 668454
rect 522804 668134 523404 668218
rect 522804 667898 522986 668134
rect 523222 667898 523404 668134
rect 522804 632454 523404 667898
rect 522804 632218 522986 632454
rect 523222 632218 523404 632454
rect 522804 632134 523404 632218
rect 522804 631898 522986 632134
rect 523222 631898 523404 632134
rect 522804 596454 523404 631898
rect 522804 596218 522986 596454
rect 523222 596218 523404 596454
rect 522804 596134 523404 596218
rect 522804 595898 522986 596134
rect 523222 595898 523404 596134
rect 522804 560454 523404 595898
rect 522804 560218 522986 560454
rect 523222 560218 523404 560454
rect 522804 560134 523404 560218
rect 522804 559898 522986 560134
rect 523222 559898 523404 560134
rect 522804 524454 523404 559898
rect 522804 524218 522986 524454
rect 523222 524218 523404 524454
rect 522804 524134 523404 524218
rect 522804 523898 522986 524134
rect 523222 523898 523404 524134
rect 522804 488454 523404 523898
rect 522804 488218 522986 488454
rect 523222 488218 523404 488454
rect 522804 488134 523404 488218
rect 522804 487898 522986 488134
rect 523222 487898 523404 488134
rect 522804 452454 523404 487898
rect 522804 452218 522986 452454
rect 523222 452218 523404 452454
rect 522804 452134 523404 452218
rect 522804 451898 522986 452134
rect 523222 451898 523404 452134
rect 522804 416454 523404 451898
rect 522804 416218 522986 416454
rect 523222 416218 523404 416454
rect 522804 416134 523404 416218
rect 522804 415898 522986 416134
rect 523222 415898 523404 416134
rect 522804 380454 523404 415898
rect 522804 380218 522986 380454
rect 523222 380218 523404 380454
rect 522804 380134 523404 380218
rect 522804 379898 522986 380134
rect 523222 379898 523404 380134
rect 522804 344454 523404 379898
rect 522804 344218 522986 344454
rect 523222 344218 523404 344454
rect 522804 344134 523404 344218
rect 522804 343898 522986 344134
rect 523222 343898 523404 344134
rect 522804 308454 523404 343898
rect 522804 308218 522986 308454
rect 523222 308218 523404 308454
rect 522804 308134 523404 308218
rect 522804 307898 522986 308134
rect 523222 307898 523404 308134
rect 522804 272454 523404 307898
rect 522804 272218 522986 272454
rect 523222 272218 523404 272454
rect 522804 272134 523404 272218
rect 522804 271898 522986 272134
rect 523222 271898 523404 272134
rect 522804 236454 523404 271898
rect 522804 236218 522986 236454
rect 523222 236218 523404 236454
rect 522804 236134 523404 236218
rect 522804 235898 522986 236134
rect 523222 235898 523404 236134
rect 522804 200454 523404 235898
rect 522804 200218 522986 200454
rect 523222 200218 523404 200454
rect 522804 200134 523404 200218
rect 522804 199898 522986 200134
rect 523222 199898 523404 200134
rect 522804 164454 523404 199898
rect 522804 164218 522986 164454
rect 523222 164218 523404 164454
rect 522804 164134 523404 164218
rect 522804 163898 522986 164134
rect 523222 163898 523404 164134
rect 522804 128454 523404 163898
rect 522804 128218 522986 128454
rect 523222 128218 523404 128454
rect 522804 128134 523404 128218
rect 522804 127898 522986 128134
rect 523222 127898 523404 128134
rect 522804 92454 523404 127898
rect 522804 92218 522986 92454
rect 523222 92218 523404 92454
rect 522804 92134 523404 92218
rect 522804 91898 522986 92134
rect 523222 91898 523404 92134
rect 522804 56454 523404 91898
rect 522804 56218 522986 56454
rect 523222 56218 523404 56454
rect 522804 56134 523404 56218
rect 522804 55898 522986 56134
rect 523222 55898 523404 56134
rect 522804 20454 523404 55898
rect 522804 20218 522986 20454
rect 523222 20218 523404 20454
rect 522804 20134 523404 20218
rect 522804 19898 522986 20134
rect 523222 19898 523404 20134
rect 522804 -1266 523404 19898
rect 522804 -1502 522986 -1266
rect 523222 -1502 523404 -1266
rect 522804 -1586 523404 -1502
rect 522804 -1822 522986 -1586
rect 523222 -1822 523404 -1586
rect 522804 -1844 523404 -1822
rect 526404 672054 527004 707042
rect 526404 671818 526586 672054
rect 526822 671818 527004 672054
rect 526404 671734 527004 671818
rect 526404 671498 526586 671734
rect 526822 671498 527004 671734
rect 526404 636054 527004 671498
rect 526404 635818 526586 636054
rect 526822 635818 527004 636054
rect 526404 635734 527004 635818
rect 526404 635498 526586 635734
rect 526822 635498 527004 635734
rect 526404 600054 527004 635498
rect 526404 599818 526586 600054
rect 526822 599818 527004 600054
rect 526404 599734 527004 599818
rect 526404 599498 526586 599734
rect 526822 599498 527004 599734
rect 526404 564054 527004 599498
rect 526404 563818 526586 564054
rect 526822 563818 527004 564054
rect 526404 563734 527004 563818
rect 526404 563498 526586 563734
rect 526822 563498 527004 563734
rect 526404 528054 527004 563498
rect 526404 527818 526586 528054
rect 526822 527818 527004 528054
rect 526404 527734 527004 527818
rect 526404 527498 526586 527734
rect 526822 527498 527004 527734
rect 526404 492054 527004 527498
rect 526404 491818 526586 492054
rect 526822 491818 527004 492054
rect 526404 491734 527004 491818
rect 526404 491498 526586 491734
rect 526822 491498 527004 491734
rect 526404 456054 527004 491498
rect 526404 455818 526586 456054
rect 526822 455818 527004 456054
rect 526404 455734 527004 455818
rect 526404 455498 526586 455734
rect 526822 455498 527004 455734
rect 526404 420054 527004 455498
rect 526404 419818 526586 420054
rect 526822 419818 527004 420054
rect 526404 419734 527004 419818
rect 526404 419498 526586 419734
rect 526822 419498 527004 419734
rect 526404 384054 527004 419498
rect 526404 383818 526586 384054
rect 526822 383818 527004 384054
rect 526404 383734 527004 383818
rect 526404 383498 526586 383734
rect 526822 383498 527004 383734
rect 526404 348054 527004 383498
rect 526404 347818 526586 348054
rect 526822 347818 527004 348054
rect 526404 347734 527004 347818
rect 526404 347498 526586 347734
rect 526822 347498 527004 347734
rect 526404 312054 527004 347498
rect 526404 311818 526586 312054
rect 526822 311818 527004 312054
rect 526404 311734 527004 311818
rect 526404 311498 526586 311734
rect 526822 311498 527004 311734
rect 526404 276054 527004 311498
rect 526404 275818 526586 276054
rect 526822 275818 527004 276054
rect 526404 275734 527004 275818
rect 526404 275498 526586 275734
rect 526822 275498 527004 275734
rect 526404 240054 527004 275498
rect 526404 239818 526586 240054
rect 526822 239818 527004 240054
rect 526404 239734 527004 239818
rect 526404 239498 526586 239734
rect 526822 239498 527004 239734
rect 526404 204054 527004 239498
rect 526404 203818 526586 204054
rect 526822 203818 527004 204054
rect 526404 203734 527004 203818
rect 526404 203498 526586 203734
rect 526822 203498 527004 203734
rect 526404 168054 527004 203498
rect 526404 167818 526586 168054
rect 526822 167818 527004 168054
rect 526404 167734 527004 167818
rect 526404 167498 526586 167734
rect 526822 167498 527004 167734
rect 526404 132054 527004 167498
rect 526404 131818 526586 132054
rect 526822 131818 527004 132054
rect 526404 131734 527004 131818
rect 526404 131498 526586 131734
rect 526822 131498 527004 131734
rect 526404 96054 527004 131498
rect 526404 95818 526586 96054
rect 526822 95818 527004 96054
rect 526404 95734 527004 95818
rect 526404 95498 526586 95734
rect 526822 95498 527004 95734
rect 526404 60054 527004 95498
rect 526404 59818 526586 60054
rect 526822 59818 527004 60054
rect 526404 59734 527004 59818
rect 526404 59498 526586 59734
rect 526822 59498 527004 59734
rect 526404 24054 527004 59498
rect 526404 23818 526586 24054
rect 526822 23818 527004 24054
rect 526404 23734 527004 23818
rect 526404 23498 526586 23734
rect 526822 23498 527004 23734
rect 526404 -3106 527004 23498
rect 526404 -3342 526586 -3106
rect 526822 -3342 527004 -3106
rect 526404 -3426 527004 -3342
rect 526404 -3662 526586 -3426
rect 526822 -3662 527004 -3426
rect 526404 -3684 527004 -3662
rect 530004 675654 530604 708882
rect 530004 675418 530186 675654
rect 530422 675418 530604 675654
rect 530004 675334 530604 675418
rect 530004 675098 530186 675334
rect 530422 675098 530604 675334
rect 530004 639654 530604 675098
rect 530004 639418 530186 639654
rect 530422 639418 530604 639654
rect 530004 639334 530604 639418
rect 530004 639098 530186 639334
rect 530422 639098 530604 639334
rect 530004 603654 530604 639098
rect 530004 603418 530186 603654
rect 530422 603418 530604 603654
rect 530004 603334 530604 603418
rect 530004 603098 530186 603334
rect 530422 603098 530604 603334
rect 530004 567654 530604 603098
rect 530004 567418 530186 567654
rect 530422 567418 530604 567654
rect 530004 567334 530604 567418
rect 530004 567098 530186 567334
rect 530422 567098 530604 567334
rect 530004 531654 530604 567098
rect 530004 531418 530186 531654
rect 530422 531418 530604 531654
rect 530004 531334 530604 531418
rect 530004 531098 530186 531334
rect 530422 531098 530604 531334
rect 530004 495654 530604 531098
rect 530004 495418 530186 495654
rect 530422 495418 530604 495654
rect 530004 495334 530604 495418
rect 530004 495098 530186 495334
rect 530422 495098 530604 495334
rect 530004 459654 530604 495098
rect 530004 459418 530186 459654
rect 530422 459418 530604 459654
rect 530004 459334 530604 459418
rect 530004 459098 530186 459334
rect 530422 459098 530604 459334
rect 530004 423654 530604 459098
rect 530004 423418 530186 423654
rect 530422 423418 530604 423654
rect 530004 423334 530604 423418
rect 530004 423098 530186 423334
rect 530422 423098 530604 423334
rect 530004 387654 530604 423098
rect 530004 387418 530186 387654
rect 530422 387418 530604 387654
rect 530004 387334 530604 387418
rect 530004 387098 530186 387334
rect 530422 387098 530604 387334
rect 530004 351654 530604 387098
rect 530004 351418 530186 351654
rect 530422 351418 530604 351654
rect 530004 351334 530604 351418
rect 530004 351098 530186 351334
rect 530422 351098 530604 351334
rect 530004 315654 530604 351098
rect 530004 315418 530186 315654
rect 530422 315418 530604 315654
rect 530004 315334 530604 315418
rect 530004 315098 530186 315334
rect 530422 315098 530604 315334
rect 530004 279654 530604 315098
rect 530004 279418 530186 279654
rect 530422 279418 530604 279654
rect 530004 279334 530604 279418
rect 530004 279098 530186 279334
rect 530422 279098 530604 279334
rect 530004 243654 530604 279098
rect 530004 243418 530186 243654
rect 530422 243418 530604 243654
rect 530004 243334 530604 243418
rect 530004 243098 530186 243334
rect 530422 243098 530604 243334
rect 530004 207654 530604 243098
rect 530004 207418 530186 207654
rect 530422 207418 530604 207654
rect 530004 207334 530604 207418
rect 530004 207098 530186 207334
rect 530422 207098 530604 207334
rect 530004 171654 530604 207098
rect 530004 171418 530186 171654
rect 530422 171418 530604 171654
rect 530004 171334 530604 171418
rect 530004 171098 530186 171334
rect 530422 171098 530604 171334
rect 530004 135654 530604 171098
rect 530004 135418 530186 135654
rect 530422 135418 530604 135654
rect 530004 135334 530604 135418
rect 530004 135098 530186 135334
rect 530422 135098 530604 135334
rect 530004 99654 530604 135098
rect 530004 99418 530186 99654
rect 530422 99418 530604 99654
rect 530004 99334 530604 99418
rect 530004 99098 530186 99334
rect 530422 99098 530604 99334
rect 530004 63654 530604 99098
rect 530004 63418 530186 63654
rect 530422 63418 530604 63654
rect 530004 63334 530604 63418
rect 530004 63098 530186 63334
rect 530422 63098 530604 63334
rect 530004 27654 530604 63098
rect 530004 27418 530186 27654
rect 530422 27418 530604 27654
rect 530004 27334 530604 27418
rect 530004 27098 530186 27334
rect 530422 27098 530604 27334
rect 530004 -4946 530604 27098
rect 530004 -5182 530186 -4946
rect 530422 -5182 530604 -4946
rect 530004 -5266 530604 -5182
rect 530004 -5502 530186 -5266
rect 530422 -5502 530604 -5266
rect 530004 -5524 530604 -5502
rect 533604 679254 534204 710722
rect 551604 710358 552204 711300
rect 551604 710122 551786 710358
rect 552022 710122 552204 710358
rect 551604 710038 552204 710122
rect 551604 709802 551786 710038
rect 552022 709802 552204 710038
rect 548004 708518 548604 709460
rect 548004 708282 548186 708518
rect 548422 708282 548604 708518
rect 548004 708198 548604 708282
rect 548004 707962 548186 708198
rect 548422 707962 548604 708198
rect 544404 706678 545004 707620
rect 544404 706442 544586 706678
rect 544822 706442 545004 706678
rect 544404 706358 545004 706442
rect 544404 706122 544586 706358
rect 544822 706122 545004 706358
rect 533604 679018 533786 679254
rect 534022 679018 534204 679254
rect 533604 678934 534204 679018
rect 533604 678698 533786 678934
rect 534022 678698 534204 678934
rect 533604 643254 534204 678698
rect 533604 643018 533786 643254
rect 534022 643018 534204 643254
rect 533604 642934 534204 643018
rect 533604 642698 533786 642934
rect 534022 642698 534204 642934
rect 533604 607254 534204 642698
rect 533604 607018 533786 607254
rect 534022 607018 534204 607254
rect 533604 606934 534204 607018
rect 533604 606698 533786 606934
rect 534022 606698 534204 606934
rect 533604 571254 534204 606698
rect 533604 571018 533786 571254
rect 534022 571018 534204 571254
rect 533604 570934 534204 571018
rect 533604 570698 533786 570934
rect 534022 570698 534204 570934
rect 533604 535254 534204 570698
rect 533604 535018 533786 535254
rect 534022 535018 534204 535254
rect 533604 534934 534204 535018
rect 533604 534698 533786 534934
rect 534022 534698 534204 534934
rect 533604 499254 534204 534698
rect 533604 499018 533786 499254
rect 534022 499018 534204 499254
rect 533604 498934 534204 499018
rect 533604 498698 533786 498934
rect 534022 498698 534204 498934
rect 533604 463254 534204 498698
rect 533604 463018 533786 463254
rect 534022 463018 534204 463254
rect 533604 462934 534204 463018
rect 533604 462698 533786 462934
rect 534022 462698 534204 462934
rect 533604 427254 534204 462698
rect 533604 427018 533786 427254
rect 534022 427018 534204 427254
rect 533604 426934 534204 427018
rect 533604 426698 533786 426934
rect 534022 426698 534204 426934
rect 533604 391254 534204 426698
rect 533604 391018 533786 391254
rect 534022 391018 534204 391254
rect 533604 390934 534204 391018
rect 533604 390698 533786 390934
rect 534022 390698 534204 390934
rect 533604 355254 534204 390698
rect 533604 355018 533786 355254
rect 534022 355018 534204 355254
rect 533604 354934 534204 355018
rect 533604 354698 533786 354934
rect 534022 354698 534204 354934
rect 533604 319254 534204 354698
rect 533604 319018 533786 319254
rect 534022 319018 534204 319254
rect 533604 318934 534204 319018
rect 533604 318698 533786 318934
rect 534022 318698 534204 318934
rect 533604 283254 534204 318698
rect 533604 283018 533786 283254
rect 534022 283018 534204 283254
rect 533604 282934 534204 283018
rect 533604 282698 533786 282934
rect 534022 282698 534204 282934
rect 533604 247254 534204 282698
rect 533604 247018 533786 247254
rect 534022 247018 534204 247254
rect 533604 246934 534204 247018
rect 533604 246698 533786 246934
rect 534022 246698 534204 246934
rect 533604 211254 534204 246698
rect 533604 211018 533786 211254
rect 534022 211018 534204 211254
rect 533604 210934 534204 211018
rect 533604 210698 533786 210934
rect 534022 210698 534204 210934
rect 533604 175254 534204 210698
rect 533604 175018 533786 175254
rect 534022 175018 534204 175254
rect 533604 174934 534204 175018
rect 533604 174698 533786 174934
rect 534022 174698 534204 174934
rect 533604 139254 534204 174698
rect 533604 139018 533786 139254
rect 534022 139018 534204 139254
rect 533604 138934 534204 139018
rect 533604 138698 533786 138934
rect 534022 138698 534204 138934
rect 533604 103254 534204 138698
rect 533604 103018 533786 103254
rect 534022 103018 534204 103254
rect 533604 102934 534204 103018
rect 533604 102698 533786 102934
rect 534022 102698 534204 102934
rect 533604 67254 534204 102698
rect 533604 67018 533786 67254
rect 534022 67018 534204 67254
rect 533604 66934 534204 67018
rect 533604 66698 533786 66934
rect 534022 66698 534204 66934
rect 533604 31254 534204 66698
rect 533604 31018 533786 31254
rect 534022 31018 534204 31254
rect 533604 30934 534204 31018
rect 533604 30698 533786 30934
rect 534022 30698 534204 30934
rect 515604 -6102 515786 -5866
rect 516022 -6102 516204 -5866
rect 515604 -6186 516204 -6102
rect 515604 -6422 515786 -6186
rect 516022 -6422 516204 -6186
rect 515604 -7364 516204 -6422
rect 533604 -6786 534204 30698
rect 540804 704838 541404 705780
rect 540804 704602 540986 704838
rect 541222 704602 541404 704838
rect 540804 704518 541404 704602
rect 540804 704282 540986 704518
rect 541222 704282 541404 704518
rect 540804 686454 541404 704282
rect 540804 686218 540986 686454
rect 541222 686218 541404 686454
rect 540804 686134 541404 686218
rect 540804 685898 540986 686134
rect 541222 685898 541404 686134
rect 540804 650454 541404 685898
rect 540804 650218 540986 650454
rect 541222 650218 541404 650454
rect 540804 650134 541404 650218
rect 540804 649898 540986 650134
rect 541222 649898 541404 650134
rect 540804 614454 541404 649898
rect 540804 614218 540986 614454
rect 541222 614218 541404 614454
rect 540804 614134 541404 614218
rect 540804 613898 540986 614134
rect 541222 613898 541404 614134
rect 540804 578454 541404 613898
rect 540804 578218 540986 578454
rect 541222 578218 541404 578454
rect 540804 578134 541404 578218
rect 540804 577898 540986 578134
rect 541222 577898 541404 578134
rect 540804 542454 541404 577898
rect 540804 542218 540986 542454
rect 541222 542218 541404 542454
rect 540804 542134 541404 542218
rect 540804 541898 540986 542134
rect 541222 541898 541404 542134
rect 540804 506454 541404 541898
rect 540804 506218 540986 506454
rect 541222 506218 541404 506454
rect 540804 506134 541404 506218
rect 540804 505898 540986 506134
rect 541222 505898 541404 506134
rect 540804 470454 541404 505898
rect 540804 470218 540986 470454
rect 541222 470218 541404 470454
rect 540804 470134 541404 470218
rect 540804 469898 540986 470134
rect 541222 469898 541404 470134
rect 540804 434454 541404 469898
rect 540804 434218 540986 434454
rect 541222 434218 541404 434454
rect 540804 434134 541404 434218
rect 540804 433898 540986 434134
rect 541222 433898 541404 434134
rect 540804 398454 541404 433898
rect 540804 398218 540986 398454
rect 541222 398218 541404 398454
rect 540804 398134 541404 398218
rect 540804 397898 540986 398134
rect 541222 397898 541404 398134
rect 540804 362454 541404 397898
rect 540804 362218 540986 362454
rect 541222 362218 541404 362454
rect 540804 362134 541404 362218
rect 540804 361898 540986 362134
rect 541222 361898 541404 362134
rect 540804 326454 541404 361898
rect 540804 326218 540986 326454
rect 541222 326218 541404 326454
rect 540804 326134 541404 326218
rect 540804 325898 540986 326134
rect 541222 325898 541404 326134
rect 540804 290454 541404 325898
rect 540804 290218 540986 290454
rect 541222 290218 541404 290454
rect 540804 290134 541404 290218
rect 540804 289898 540986 290134
rect 541222 289898 541404 290134
rect 540804 254454 541404 289898
rect 540804 254218 540986 254454
rect 541222 254218 541404 254454
rect 540804 254134 541404 254218
rect 540804 253898 540986 254134
rect 541222 253898 541404 254134
rect 540804 218454 541404 253898
rect 540804 218218 540986 218454
rect 541222 218218 541404 218454
rect 540804 218134 541404 218218
rect 540804 217898 540986 218134
rect 541222 217898 541404 218134
rect 540804 182454 541404 217898
rect 540804 182218 540986 182454
rect 541222 182218 541404 182454
rect 540804 182134 541404 182218
rect 540804 181898 540986 182134
rect 541222 181898 541404 182134
rect 540804 146454 541404 181898
rect 540804 146218 540986 146454
rect 541222 146218 541404 146454
rect 540804 146134 541404 146218
rect 540804 145898 540986 146134
rect 541222 145898 541404 146134
rect 540804 110454 541404 145898
rect 540804 110218 540986 110454
rect 541222 110218 541404 110454
rect 540804 110134 541404 110218
rect 540804 109898 540986 110134
rect 541222 109898 541404 110134
rect 540804 74454 541404 109898
rect 540804 74218 540986 74454
rect 541222 74218 541404 74454
rect 540804 74134 541404 74218
rect 540804 73898 540986 74134
rect 541222 73898 541404 74134
rect 540804 38454 541404 73898
rect 540804 38218 540986 38454
rect 541222 38218 541404 38454
rect 540804 38134 541404 38218
rect 540804 37898 540986 38134
rect 541222 37898 541404 38134
rect 540804 2454 541404 37898
rect 540804 2218 540986 2454
rect 541222 2218 541404 2454
rect 540804 2134 541404 2218
rect 540804 1898 540986 2134
rect 541222 1898 541404 2134
rect 540804 -346 541404 1898
rect 540804 -582 540986 -346
rect 541222 -582 541404 -346
rect 540804 -666 541404 -582
rect 540804 -902 540986 -666
rect 541222 -902 541404 -666
rect 540804 -1844 541404 -902
rect 544404 690054 545004 706122
rect 544404 689818 544586 690054
rect 544822 689818 545004 690054
rect 544404 689734 545004 689818
rect 544404 689498 544586 689734
rect 544822 689498 545004 689734
rect 544404 654054 545004 689498
rect 544404 653818 544586 654054
rect 544822 653818 545004 654054
rect 544404 653734 545004 653818
rect 544404 653498 544586 653734
rect 544822 653498 545004 653734
rect 544404 618054 545004 653498
rect 544404 617818 544586 618054
rect 544822 617818 545004 618054
rect 544404 617734 545004 617818
rect 544404 617498 544586 617734
rect 544822 617498 545004 617734
rect 544404 582054 545004 617498
rect 544404 581818 544586 582054
rect 544822 581818 545004 582054
rect 544404 581734 545004 581818
rect 544404 581498 544586 581734
rect 544822 581498 545004 581734
rect 544404 546054 545004 581498
rect 544404 545818 544586 546054
rect 544822 545818 545004 546054
rect 544404 545734 545004 545818
rect 544404 545498 544586 545734
rect 544822 545498 545004 545734
rect 544404 510054 545004 545498
rect 544404 509818 544586 510054
rect 544822 509818 545004 510054
rect 544404 509734 545004 509818
rect 544404 509498 544586 509734
rect 544822 509498 545004 509734
rect 544404 474054 545004 509498
rect 544404 473818 544586 474054
rect 544822 473818 545004 474054
rect 544404 473734 545004 473818
rect 544404 473498 544586 473734
rect 544822 473498 545004 473734
rect 544404 438054 545004 473498
rect 544404 437818 544586 438054
rect 544822 437818 545004 438054
rect 544404 437734 545004 437818
rect 544404 437498 544586 437734
rect 544822 437498 545004 437734
rect 544404 402054 545004 437498
rect 544404 401818 544586 402054
rect 544822 401818 545004 402054
rect 544404 401734 545004 401818
rect 544404 401498 544586 401734
rect 544822 401498 545004 401734
rect 544404 366054 545004 401498
rect 544404 365818 544586 366054
rect 544822 365818 545004 366054
rect 544404 365734 545004 365818
rect 544404 365498 544586 365734
rect 544822 365498 545004 365734
rect 544404 330054 545004 365498
rect 544404 329818 544586 330054
rect 544822 329818 545004 330054
rect 544404 329734 545004 329818
rect 544404 329498 544586 329734
rect 544822 329498 545004 329734
rect 544404 294054 545004 329498
rect 544404 293818 544586 294054
rect 544822 293818 545004 294054
rect 544404 293734 545004 293818
rect 544404 293498 544586 293734
rect 544822 293498 545004 293734
rect 544404 258054 545004 293498
rect 544404 257818 544586 258054
rect 544822 257818 545004 258054
rect 544404 257734 545004 257818
rect 544404 257498 544586 257734
rect 544822 257498 545004 257734
rect 544404 222054 545004 257498
rect 544404 221818 544586 222054
rect 544822 221818 545004 222054
rect 544404 221734 545004 221818
rect 544404 221498 544586 221734
rect 544822 221498 545004 221734
rect 544404 186054 545004 221498
rect 544404 185818 544586 186054
rect 544822 185818 545004 186054
rect 544404 185734 545004 185818
rect 544404 185498 544586 185734
rect 544822 185498 545004 185734
rect 544404 150054 545004 185498
rect 544404 149818 544586 150054
rect 544822 149818 545004 150054
rect 544404 149734 545004 149818
rect 544404 149498 544586 149734
rect 544822 149498 545004 149734
rect 544404 114054 545004 149498
rect 544404 113818 544586 114054
rect 544822 113818 545004 114054
rect 544404 113734 545004 113818
rect 544404 113498 544586 113734
rect 544822 113498 545004 113734
rect 544404 78054 545004 113498
rect 544404 77818 544586 78054
rect 544822 77818 545004 78054
rect 544404 77734 545004 77818
rect 544404 77498 544586 77734
rect 544822 77498 545004 77734
rect 544404 42054 545004 77498
rect 544404 41818 544586 42054
rect 544822 41818 545004 42054
rect 544404 41734 545004 41818
rect 544404 41498 544586 41734
rect 544822 41498 545004 41734
rect 544404 6054 545004 41498
rect 544404 5818 544586 6054
rect 544822 5818 545004 6054
rect 544404 5734 545004 5818
rect 544404 5498 544586 5734
rect 544822 5498 545004 5734
rect 544404 -2186 545004 5498
rect 544404 -2422 544586 -2186
rect 544822 -2422 545004 -2186
rect 544404 -2506 545004 -2422
rect 544404 -2742 544586 -2506
rect 544822 -2742 545004 -2506
rect 544404 -3684 545004 -2742
rect 548004 693654 548604 707962
rect 548004 693418 548186 693654
rect 548422 693418 548604 693654
rect 548004 693334 548604 693418
rect 548004 693098 548186 693334
rect 548422 693098 548604 693334
rect 548004 657654 548604 693098
rect 548004 657418 548186 657654
rect 548422 657418 548604 657654
rect 548004 657334 548604 657418
rect 548004 657098 548186 657334
rect 548422 657098 548604 657334
rect 548004 621654 548604 657098
rect 548004 621418 548186 621654
rect 548422 621418 548604 621654
rect 548004 621334 548604 621418
rect 548004 621098 548186 621334
rect 548422 621098 548604 621334
rect 548004 585654 548604 621098
rect 548004 585418 548186 585654
rect 548422 585418 548604 585654
rect 548004 585334 548604 585418
rect 548004 585098 548186 585334
rect 548422 585098 548604 585334
rect 548004 549654 548604 585098
rect 548004 549418 548186 549654
rect 548422 549418 548604 549654
rect 548004 549334 548604 549418
rect 548004 549098 548186 549334
rect 548422 549098 548604 549334
rect 548004 513654 548604 549098
rect 548004 513418 548186 513654
rect 548422 513418 548604 513654
rect 548004 513334 548604 513418
rect 548004 513098 548186 513334
rect 548422 513098 548604 513334
rect 548004 477654 548604 513098
rect 548004 477418 548186 477654
rect 548422 477418 548604 477654
rect 548004 477334 548604 477418
rect 548004 477098 548186 477334
rect 548422 477098 548604 477334
rect 548004 441654 548604 477098
rect 548004 441418 548186 441654
rect 548422 441418 548604 441654
rect 548004 441334 548604 441418
rect 548004 441098 548186 441334
rect 548422 441098 548604 441334
rect 548004 405654 548604 441098
rect 548004 405418 548186 405654
rect 548422 405418 548604 405654
rect 548004 405334 548604 405418
rect 548004 405098 548186 405334
rect 548422 405098 548604 405334
rect 548004 369654 548604 405098
rect 548004 369418 548186 369654
rect 548422 369418 548604 369654
rect 548004 369334 548604 369418
rect 548004 369098 548186 369334
rect 548422 369098 548604 369334
rect 548004 333654 548604 369098
rect 548004 333418 548186 333654
rect 548422 333418 548604 333654
rect 548004 333334 548604 333418
rect 548004 333098 548186 333334
rect 548422 333098 548604 333334
rect 548004 297654 548604 333098
rect 548004 297418 548186 297654
rect 548422 297418 548604 297654
rect 548004 297334 548604 297418
rect 548004 297098 548186 297334
rect 548422 297098 548604 297334
rect 548004 261654 548604 297098
rect 548004 261418 548186 261654
rect 548422 261418 548604 261654
rect 548004 261334 548604 261418
rect 548004 261098 548186 261334
rect 548422 261098 548604 261334
rect 548004 225654 548604 261098
rect 548004 225418 548186 225654
rect 548422 225418 548604 225654
rect 548004 225334 548604 225418
rect 548004 225098 548186 225334
rect 548422 225098 548604 225334
rect 548004 189654 548604 225098
rect 548004 189418 548186 189654
rect 548422 189418 548604 189654
rect 548004 189334 548604 189418
rect 548004 189098 548186 189334
rect 548422 189098 548604 189334
rect 548004 153654 548604 189098
rect 548004 153418 548186 153654
rect 548422 153418 548604 153654
rect 548004 153334 548604 153418
rect 548004 153098 548186 153334
rect 548422 153098 548604 153334
rect 548004 117654 548604 153098
rect 548004 117418 548186 117654
rect 548422 117418 548604 117654
rect 548004 117334 548604 117418
rect 548004 117098 548186 117334
rect 548422 117098 548604 117334
rect 548004 81654 548604 117098
rect 548004 81418 548186 81654
rect 548422 81418 548604 81654
rect 548004 81334 548604 81418
rect 548004 81098 548186 81334
rect 548422 81098 548604 81334
rect 548004 45654 548604 81098
rect 548004 45418 548186 45654
rect 548422 45418 548604 45654
rect 548004 45334 548604 45418
rect 548004 45098 548186 45334
rect 548422 45098 548604 45334
rect 548004 9654 548604 45098
rect 548004 9418 548186 9654
rect 548422 9418 548604 9654
rect 548004 9334 548604 9418
rect 548004 9098 548186 9334
rect 548422 9098 548604 9334
rect 548004 -4026 548604 9098
rect 548004 -4262 548186 -4026
rect 548422 -4262 548604 -4026
rect 548004 -4346 548604 -4262
rect 548004 -4582 548186 -4346
rect 548422 -4582 548604 -4346
rect 548004 -5524 548604 -4582
rect 551604 697254 552204 709802
rect 569604 711278 570204 711300
rect 569604 711042 569786 711278
rect 570022 711042 570204 711278
rect 569604 710958 570204 711042
rect 569604 710722 569786 710958
rect 570022 710722 570204 710958
rect 566004 709438 566604 709460
rect 566004 709202 566186 709438
rect 566422 709202 566604 709438
rect 566004 709118 566604 709202
rect 566004 708882 566186 709118
rect 566422 708882 566604 709118
rect 562404 707598 563004 707620
rect 562404 707362 562586 707598
rect 562822 707362 563004 707598
rect 562404 707278 563004 707362
rect 562404 707042 562586 707278
rect 562822 707042 563004 707278
rect 551604 697018 551786 697254
rect 552022 697018 552204 697254
rect 551604 696934 552204 697018
rect 551604 696698 551786 696934
rect 552022 696698 552204 696934
rect 551604 661254 552204 696698
rect 551604 661018 551786 661254
rect 552022 661018 552204 661254
rect 551604 660934 552204 661018
rect 551604 660698 551786 660934
rect 552022 660698 552204 660934
rect 551604 625254 552204 660698
rect 551604 625018 551786 625254
rect 552022 625018 552204 625254
rect 551604 624934 552204 625018
rect 551604 624698 551786 624934
rect 552022 624698 552204 624934
rect 551604 589254 552204 624698
rect 551604 589018 551786 589254
rect 552022 589018 552204 589254
rect 551604 588934 552204 589018
rect 551604 588698 551786 588934
rect 552022 588698 552204 588934
rect 551604 553254 552204 588698
rect 551604 553018 551786 553254
rect 552022 553018 552204 553254
rect 551604 552934 552204 553018
rect 551604 552698 551786 552934
rect 552022 552698 552204 552934
rect 551604 517254 552204 552698
rect 551604 517018 551786 517254
rect 552022 517018 552204 517254
rect 551604 516934 552204 517018
rect 551604 516698 551786 516934
rect 552022 516698 552204 516934
rect 551604 481254 552204 516698
rect 551604 481018 551786 481254
rect 552022 481018 552204 481254
rect 551604 480934 552204 481018
rect 551604 480698 551786 480934
rect 552022 480698 552204 480934
rect 551604 445254 552204 480698
rect 551604 445018 551786 445254
rect 552022 445018 552204 445254
rect 551604 444934 552204 445018
rect 551604 444698 551786 444934
rect 552022 444698 552204 444934
rect 551604 409254 552204 444698
rect 551604 409018 551786 409254
rect 552022 409018 552204 409254
rect 551604 408934 552204 409018
rect 551604 408698 551786 408934
rect 552022 408698 552204 408934
rect 551604 373254 552204 408698
rect 551604 373018 551786 373254
rect 552022 373018 552204 373254
rect 551604 372934 552204 373018
rect 551604 372698 551786 372934
rect 552022 372698 552204 372934
rect 551604 337254 552204 372698
rect 551604 337018 551786 337254
rect 552022 337018 552204 337254
rect 551604 336934 552204 337018
rect 551604 336698 551786 336934
rect 552022 336698 552204 336934
rect 551604 301254 552204 336698
rect 551604 301018 551786 301254
rect 552022 301018 552204 301254
rect 551604 300934 552204 301018
rect 551604 300698 551786 300934
rect 552022 300698 552204 300934
rect 551604 265254 552204 300698
rect 551604 265018 551786 265254
rect 552022 265018 552204 265254
rect 551604 264934 552204 265018
rect 551604 264698 551786 264934
rect 552022 264698 552204 264934
rect 551604 229254 552204 264698
rect 551604 229018 551786 229254
rect 552022 229018 552204 229254
rect 551604 228934 552204 229018
rect 551604 228698 551786 228934
rect 552022 228698 552204 228934
rect 551604 193254 552204 228698
rect 551604 193018 551786 193254
rect 552022 193018 552204 193254
rect 551604 192934 552204 193018
rect 551604 192698 551786 192934
rect 552022 192698 552204 192934
rect 551604 157254 552204 192698
rect 551604 157018 551786 157254
rect 552022 157018 552204 157254
rect 551604 156934 552204 157018
rect 551604 156698 551786 156934
rect 552022 156698 552204 156934
rect 551604 121254 552204 156698
rect 551604 121018 551786 121254
rect 552022 121018 552204 121254
rect 551604 120934 552204 121018
rect 551604 120698 551786 120934
rect 552022 120698 552204 120934
rect 551604 85254 552204 120698
rect 551604 85018 551786 85254
rect 552022 85018 552204 85254
rect 551604 84934 552204 85018
rect 551604 84698 551786 84934
rect 552022 84698 552204 84934
rect 551604 49254 552204 84698
rect 551604 49018 551786 49254
rect 552022 49018 552204 49254
rect 551604 48934 552204 49018
rect 551604 48698 551786 48934
rect 552022 48698 552204 48934
rect 551604 13254 552204 48698
rect 551604 13018 551786 13254
rect 552022 13018 552204 13254
rect 551604 12934 552204 13018
rect 551604 12698 551786 12934
rect 552022 12698 552204 12934
rect 533604 -7022 533786 -6786
rect 534022 -7022 534204 -6786
rect 533604 -7106 534204 -7022
rect 533604 -7342 533786 -7106
rect 534022 -7342 534204 -7106
rect 533604 -7364 534204 -7342
rect 551604 -5866 552204 12698
rect 558804 705758 559404 705780
rect 558804 705522 558986 705758
rect 559222 705522 559404 705758
rect 558804 705438 559404 705522
rect 558804 705202 558986 705438
rect 559222 705202 559404 705438
rect 558804 668454 559404 705202
rect 558804 668218 558986 668454
rect 559222 668218 559404 668454
rect 558804 668134 559404 668218
rect 558804 667898 558986 668134
rect 559222 667898 559404 668134
rect 558804 632454 559404 667898
rect 558804 632218 558986 632454
rect 559222 632218 559404 632454
rect 558804 632134 559404 632218
rect 558804 631898 558986 632134
rect 559222 631898 559404 632134
rect 558804 596454 559404 631898
rect 558804 596218 558986 596454
rect 559222 596218 559404 596454
rect 558804 596134 559404 596218
rect 558804 595898 558986 596134
rect 559222 595898 559404 596134
rect 558804 560454 559404 595898
rect 558804 560218 558986 560454
rect 559222 560218 559404 560454
rect 558804 560134 559404 560218
rect 558804 559898 558986 560134
rect 559222 559898 559404 560134
rect 558804 524454 559404 559898
rect 558804 524218 558986 524454
rect 559222 524218 559404 524454
rect 558804 524134 559404 524218
rect 558804 523898 558986 524134
rect 559222 523898 559404 524134
rect 558804 488454 559404 523898
rect 558804 488218 558986 488454
rect 559222 488218 559404 488454
rect 558804 488134 559404 488218
rect 558804 487898 558986 488134
rect 559222 487898 559404 488134
rect 558804 452454 559404 487898
rect 558804 452218 558986 452454
rect 559222 452218 559404 452454
rect 558804 452134 559404 452218
rect 558804 451898 558986 452134
rect 559222 451898 559404 452134
rect 558804 416454 559404 451898
rect 558804 416218 558986 416454
rect 559222 416218 559404 416454
rect 558804 416134 559404 416218
rect 558804 415898 558986 416134
rect 559222 415898 559404 416134
rect 558804 380454 559404 415898
rect 558804 380218 558986 380454
rect 559222 380218 559404 380454
rect 558804 380134 559404 380218
rect 558804 379898 558986 380134
rect 559222 379898 559404 380134
rect 558804 344454 559404 379898
rect 558804 344218 558986 344454
rect 559222 344218 559404 344454
rect 558804 344134 559404 344218
rect 558804 343898 558986 344134
rect 559222 343898 559404 344134
rect 558804 308454 559404 343898
rect 558804 308218 558986 308454
rect 559222 308218 559404 308454
rect 558804 308134 559404 308218
rect 558804 307898 558986 308134
rect 559222 307898 559404 308134
rect 558804 272454 559404 307898
rect 558804 272218 558986 272454
rect 559222 272218 559404 272454
rect 558804 272134 559404 272218
rect 558804 271898 558986 272134
rect 559222 271898 559404 272134
rect 558804 236454 559404 271898
rect 558804 236218 558986 236454
rect 559222 236218 559404 236454
rect 558804 236134 559404 236218
rect 558804 235898 558986 236134
rect 559222 235898 559404 236134
rect 558804 200454 559404 235898
rect 558804 200218 558986 200454
rect 559222 200218 559404 200454
rect 558804 200134 559404 200218
rect 558804 199898 558986 200134
rect 559222 199898 559404 200134
rect 558804 164454 559404 199898
rect 558804 164218 558986 164454
rect 559222 164218 559404 164454
rect 558804 164134 559404 164218
rect 558804 163898 558986 164134
rect 559222 163898 559404 164134
rect 558804 128454 559404 163898
rect 558804 128218 558986 128454
rect 559222 128218 559404 128454
rect 558804 128134 559404 128218
rect 558804 127898 558986 128134
rect 559222 127898 559404 128134
rect 558804 92454 559404 127898
rect 558804 92218 558986 92454
rect 559222 92218 559404 92454
rect 558804 92134 559404 92218
rect 558804 91898 558986 92134
rect 559222 91898 559404 92134
rect 558804 56454 559404 91898
rect 558804 56218 558986 56454
rect 559222 56218 559404 56454
rect 558804 56134 559404 56218
rect 558804 55898 558986 56134
rect 559222 55898 559404 56134
rect 558804 20454 559404 55898
rect 558804 20218 558986 20454
rect 559222 20218 559404 20454
rect 558804 20134 559404 20218
rect 558804 19898 558986 20134
rect 559222 19898 559404 20134
rect 558804 -1266 559404 19898
rect 558804 -1502 558986 -1266
rect 559222 -1502 559404 -1266
rect 558804 -1586 559404 -1502
rect 558804 -1822 558986 -1586
rect 559222 -1822 559404 -1586
rect 558804 -1844 559404 -1822
rect 562404 672054 563004 707042
rect 562404 671818 562586 672054
rect 562822 671818 563004 672054
rect 562404 671734 563004 671818
rect 562404 671498 562586 671734
rect 562822 671498 563004 671734
rect 562404 636054 563004 671498
rect 562404 635818 562586 636054
rect 562822 635818 563004 636054
rect 562404 635734 563004 635818
rect 562404 635498 562586 635734
rect 562822 635498 563004 635734
rect 562404 600054 563004 635498
rect 562404 599818 562586 600054
rect 562822 599818 563004 600054
rect 562404 599734 563004 599818
rect 562404 599498 562586 599734
rect 562822 599498 563004 599734
rect 562404 564054 563004 599498
rect 562404 563818 562586 564054
rect 562822 563818 563004 564054
rect 562404 563734 563004 563818
rect 562404 563498 562586 563734
rect 562822 563498 563004 563734
rect 562404 528054 563004 563498
rect 562404 527818 562586 528054
rect 562822 527818 563004 528054
rect 562404 527734 563004 527818
rect 562404 527498 562586 527734
rect 562822 527498 563004 527734
rect 562404 492054 563004 527498
rect 562404 491818 562586 492054
rect 562822 491818 563004 492054
rect 562404 491734 563004 491818
rect 562404 491498 562586 491734
rect 562822 491498 563004 491734
rect 562404 456054 563004 491498
rect 562404 455818 562586 456054
rect 562822 455818 563004 456054
rect 562404 455734 563004 455818
rect 562404 455498 562586 455734
rect 562822 455498 563004 455734
rect 562404 420054 563004 455498
rect 562404 419818 562586 420054
rect 562822 419818 563004 420054
rect 562404 419734 563004 419818
rect 562404 419498 562586 419734
rect 562822 419498 563004 419734
rect 562404 384054 563004 419498
rect 562404 383818 562586 384054
rect 562822 383818 563004 384054
rect 562404 383734 563004 383818
rect 562404 383498 562586 383734
rect 562822 383498 563004 383734
rect 562404 348054 563004 383498
rect 562404 347818 562586 348054
rect 562822 347818 563004 348054
rect 562404 347734 563004 347818
rect 562404 347498 562586 347734
rect 562822 347498 563004 347734
rect 562404 312054 563004 347498
rect 562404 311818 562586 312054
rect 562822 311818 563004 312054
rect 562404 311734 563004 311818
rect 562404 311498 562586 311734
rect 562822 311498 563004 311734
rect 562404 276054 563004 311498
rect 562404 275818 562586 276054
rect 562822 275818 563004 276054
rect 562404 275734 563004 275818
rect 562404 275498 562586 275734
rect 562822 275498 563004 275734
rect 562404 240054 563004 275498
rect 562404 239818 562586 240054
rect 562822 239818 563004 240054
rect 562404 239734 563004 239818
rect 562404 239498 562586 239734
rect 562822 239498 563004 239734
rect 562404 204054 563004 239498
rect 562404 203818 562586 204054
rect 562822 203818 563004 204054
rect 562404 203734 563004 203818
rect 562404 203498 562586 203734
rect 562822 203498 563004 203734
rect 562404 168054 563004 203498
rect 562404 167818 562586 168054
rect 562822 167818 563004 168054
rect 562404 167734 563004 167818
rect 562404 167498 562586 167734
rect 562822 167498 563004 167734
rect 562404 132054 563004 167498
rect 562404 131818 562586 132054
rect 562822 131818 563004 132054
rect 562404 131734 563004 131818
rect 562404 131498 562586 131734
rect 562822 131498 563004 131734
rect 562404 96054 563004 131498
rect 562404 95818 562586 96054
rect 562822 95818 563004 96054
rect 562404 95734 563004 95818
rect 562404 95498 562586 95734
rect 562822 95498 563004 95734
rect 562404 60054 563004 95498
rect 562404 59818 562586 60054
rect 562822 59818 563004 60054
rect 562404 59734 563004 59818
rect 562404 59498 562586 59734
rect 562822 59498 563004 59734
rect 562404 24054 563004 59498
rect 562404 23818 562586 24054
rect 562822 23818 563004 24054
rect 562404 23734 563004 23818
rect 562404 23498 562586 23734
rect 562822 23498 563004 23734
rect 562404 -3106 563004 23498
rect 562404 -3342 562586 -3106
rect 562822 -3342 563004 -3106
rect 562404 -3426 563004 -3342
rect 562404 -3662 562586 -3426
rect 562822 -3662 563004 -3426
rect 562404 -3684 563004 -3662
rect 566004 675654 566604 708882
rect 566004 675418 566186 675654
rect 566422 675418 566604 675654
rect 566004 675334 566604 675418
rect 566004 675098 566186 675334
rect 566422 675098 566604 675334
rect 566004 639654 566604 675098
rect 566004 639418 566186 639654
rect 566422 639418 566604 639654
rect 566004 639334 566604 639418
rect 566004 639098 566186 639334
rect 566422 639098 566604 639334
rect 566004 603654 566604 639098
rect 566004 603418 566186 603654
rect 566422 603418 566604 603654
rect 566004 603334 566604 603418
rect 566004 603098 566186 603334
rect 566422 603098 566604 603334
rect 566004 567654 566604 603098
rect 566004 567418 566186 567654
rect 566422 567418 566604 567654
rect 566004 567334 566604 567418
rect 566004 567098 566186 567334
rect 566422 567098 566604 567334
rect 566004 531654 566604 567098
rect 566004 531418 566186 531654
rect 566422 531418 566604 531654
rect 566004 531334 566604 531418
rect 566004 531098 566186 531334
rect 566422 531098 566604 531334
rect 566004 495654 566604 531098
rect 566004 495418 566186 495654
rect 566422 495418 566604 495654
rect 566004 495334 566604 495418
rect 566004 495098 566186 495334
rect 566422 495098 566604 495334
rect 566004 459654 566604 495098
rect 566004 459418 566186 459654
rect 566422 459418 566604 459654
rect 566004 459334 566604 459418
rect 566004 459098 566186 459334
rect 566422 459098 566604 459334
rect 566004 423654 566604 459098
rect 566004 423418 566186 423654
rect 566422 423418 566604 423654
rect 566004 423334 566604 423418
rect 566004 423098 566186 423334
rect 566422 423098 566604 423334
rect 566004 387654 566604 423098
rect 566004 387418 566186 387654
rect 566422 387418 566604 387654
rect 566004 387334 566604 387418
rect 566004 387098 566186 387334
rect 566422 387098 566604 387334
rect 566004 351654 566604 387098
rect 566004 351418 566186 351654
rect 566422 351418 566604 351654
rect 566004 351334 566604 351418
rect 566004 351098 566186 351334
rect 566422 351098 566604 351334
rect 566004 315654 566604 351098
rect 566004 315418 566186 315654
rect 566422 315418 566604 315654
rect 566004 315334 566604 315418
rect 566004 315098 566186 315334
rect 566422 315098 566604 315334
rect 566004 279654 566604 315098
rect 566004 279418 566186 279654
rect 566422 279418 566604 279654
rect 566004 279334 566604 279418
rect 566004 279098 566186 279334
rect 566422 279098 566604 279334
rect 566004 243654 566604 279098
rect 566004 243418 566186 243654
rect 566422 243418 566604 243654
rect 566004 243334 566604 243418
rect 566004 243098 566186 243334
rect 566422 243098 566604 243334
rect 566004 207654 566604 243098
rect 566004 207418 566186 207654
rect 566422 207418 566604 207654
rect 566004 207334 566604 207418
rect 566004 207098 566186 207334
rect 566422 207098 566604 207334
rect 566004 171654 566604 207098
rect 566004 171418 566186 171654
rect 566422 171418 566604 171654
rect 566004 171334 566604 171418
rect 566004 171098 566186 171334
rect 566422 171098 566604 171334
rect 566004 135654 566604 171098
rect 566004 135418 566186 135654
rect 566422 135418 566604 135654
rect 566004 135334 566604 135418
rect 566004 135098 566186 135334
rect 566422 135098 566604 135334
rect 566004 99654 566604 135098
rect 566004 99418 566186 99654
rect 566422 99418 566604 99654
rect 566004 99334 566604 99418
rect 566004 99098 566186 99334
rect 566422 99098 566604 99334
rect 566004 63654 566604 99098
rect 566004 63418 566186 63654
rect 566422 63418 566604 63654
rect 566004 63334 566604 63418
rect 566004 63098 566186 63334
rect 566422 63098 566604 63334
rect 566004 27654 566604 63098
rect 566004 27418 566186 27654
rect 566422 27418 566604 27654
rect 566004 27334 566604 27418
rect 566004 27098 566186 27334
rect 566422 27098 566604 27334
rect 566004 -4946 566604 27098
rect 566004 -5182 566186 -4946
rect 566422 -5182 566604 -4946
rect 566004 -5266 566604 -5182
rect 566004 -5502 566186 -5266
rect 566422 -5502 566604 -5266
rect 566004 -5524 566604 -5502
rect 569604 679254 570204 710722
rect 591760 711278 592360 711300
rect 591760 711042 591942 711278
rect 592178 711042 592360 711278
rect 591760 710958 592360 711042
rect 591760 710722 591942 710958
rect 592178 710722 592360 710958
rect 590840 710358 591440 710380
rect 590840 710122 591022 710358
rect 591258 710122 591440 710358
rect 590840 710038 591440 710122
rect 590840 709802 591022 710038
rect 591258 709802 591440 710038
rect 589920 709438 590520 709460
rect 589920 709202 590102 709438
rect 590338 709202 590520 709438
rect 589920 709118 590520 709202
rect 589920 708882 590102 709118
rect 590338 708882 590520 709118
rect 589000 708518 589600 708540
rect 589000 708282 589182 708518
rect 589418 708282 589600 708518
rect 589000 708198 589600 708282
rect 589000 707962 589182 708198
rect 589418 707962 589600 708198
rect 580404 706678 581004 707620
rect 588080 707598 588680 707620
rect 588080 707362 588262 707598
rect 588498 707362 588680 707598
rect 588080 707278 588680 707362
rect 588080 707042 588262 707278
rect 588498 707042 588680 707278
rect 580404 706442 580586 706678
rect 580822 706442 581004 706678
rect 580404 706358 581004 706442
rect 580404 706122 580586 706358
rect 580822 706122 581004 706358
rect 569604 679018 569786 679254
rect 570022 679018 570204 679254
rect 569604 678934 570204 679018
rect 569604 678698 569786 678934
rect 570022 678698 570204 678934
rect 569604 643254 570204 678698
rect 569604 643018 569786 643254
rect 570022 643018 570204 643254
rect 569604 642934 570204 643018
rect 569604 642698 569786 642934
rect 570022 642698 570204 642934
rect 569604 607254 570204 642698
rect 569604 607018 569786 607254
rect 570022 607018 570204 607254
rect 569604 606934 570204 607018
rect 569604 606698 569786 606934
rect 570022 606698 570204 606934
rect 569604 571254 570204 606698
rect 569604 571018 569786 571254
rect 570022 571018 570204 571254
rect 569604 570934 570204 571018
rect 569604 570698 569786 570934
rect 570022 570698 570204 570934
rect 569604 535254 570204 570698
rect 569604 535018 569786 535254
rect 570022 535018 570204 535254
rect 569604 534934 570204 535018
rect 569604 534698 569786 534934
rect 570022 534698 570204 534934
rect 569604 499254 570204 534698
rect 569604 499018 569786 499254
rect 570022 499018 570204 499254
rect 569604 498934 570204 499018
rect 569604 498698 569786 498934
rect 570022 498698 570204 498934
rect 569604 463254 570204 498698
rect 569604 463018 569786 463254
rect 570022 463018 570204 463254
rect 569604 462934 570204 463018
rect 569604 462698 569786 462934
rect 570022 462698 570204 462934
rect 569604 427254 570204 462698
rect 569604 427018 569786 427254
rect 570022 427018 570204 427254
rect 569604 426934 570204 427018
rect 569604 426698 569786 426934
rect 570022 426698 570204 426934
rect 569604 391254 570204 426698
rect 569604 391018 569786 391254
rect 570022 391018 570204 391254
rect 569604 390934 570204 391018
rect 569604 390698 569786 390934
rect 570022 390698 570204 390934
rect 569604 355254 570204 390698
rect 569604 355018 569786 355254
rect 570022 355018 570204 355254
rect 569604 354934 570204 355018
rect 569604 354698 569786 354934
rect 570022 354698 570204 354934
rect 569604 319254 570204 354698
rect 569604 319018 569786 319254
rect 570022 319018 570204 319254
rect 569604 318934 570204 319018
rect 569604 318698 569786 318934
rect 570022 318698 570204 318934
rect 569604 283254 570204 318698
rect 569604 283018 569786 283254
rect 570022 283018 570204 283254
rect 569604 282934 570204 283018
rect 569604 282698 569786 282934
rect 570022 282698 570204 282934
rect 569604 247254 570204 282698
rect 569604 247018 569786 247254
rect 570022 247018 570204 247254
rect 569604 246934 570204 247018
rect 569604 246698 569786 246934
rect 570022 246698 570204 246934
rect 569604 211254 570204 246698
rect 569604 211018 569786 211254
rect 570022 211018 570204 211254
rect 569604 210934 570204 211018
rect 569604 210698 569786 210934
rect 570022 210698 570204 210934
rect 569604 175254 570204 210698
rect 569604 175018 569786 175254
rect 570022 175018 570204 175254
rect 569604 174934 570204 175018
rect 569604 174698 569786 174934
rect 570022 174698 570204 174934
rect 569604 139254 570204 174698
rect 569604 139018 569786 139254
rect 570022 139018 570204 139254
rect 569604 138934 570204 139018
rect 569604 138698 569786 138934
rect 570022 138698 570204 138934
rect 569604 103254 570204 138698
rect 569604 103018 569786 103254
rect 570022 103018 570204 103254
rect 569604 102934 570204 103018
rect 569604 102698 569786 102934
rect 570022 102698 570204 102934
rect 569604 67254 570204 102698
rect 569604 67018 569786 67254
rect 570022 67018 570204 67254
rect 569604 66934 570204 67018
rect 569604 66698 569786 66934
rect 570022 66698 570204 66934
rect 569604 31254 570204 66698
rect 569604 31018 569786 31254
rect 570022 31018 570204 31254
rect 569604 30934 570204 31018
rect 569604 30698 569786 30934
rect 570022 30698 570204 30934
rect 551604 -6102 551786 -5866
rect 552022 -6102 552204 -5866
rect 551604 -6186 552204 -6102
rect 551604 -6422 551786 -6186
rect 552022 -6422 552204 -6186
rect 551604 -7364 552204 -6422
rect 569604 -6786 570204 30698
rect 576804 704838 577404 705780
rect 576804 704602 576986 704838
rect 577222 704602 577404 704838
rect 576804 704518 577404 704602
rect 576804 704282 576986 704518
rect 577222 704282 577404 704518
rect 576804 686454 577404 704282
rect 576804 686218 576986 686454
rect 577222 686218 577404 686454
rect 576804 686134 577404 686218
rect 576804 685898 576986 686134
rect 577222 685898 577404 686134
rect 576804 650454 577404 685898
rect 576804 650218 576986 650454
rect 577222 650218 577404 650454
rect 576804 650134 577404 650218
rect 576804 649898 576986 650134
rect 577222 649898 577404 650134
rect 576804 614454 577404 649898
rect 576804 614218 576986 614454
rect 577222 614218 577404 614454
rect 576804 614134 577404 614218
rect 576804 613898 576986 614134
rect 577222 613898 577404 614134
rect 576804 578454 577404 613898
rect 576804 578218 576986 578454
rect 577222 578218 577404 578454
rect 576804 578134 577404 578218
rect 576804 577898 576986 578134
rect 577222 577898 577404 578134
rect 576804 542454 577404 577898
rect 576804 542218 576986 542454
rect 577222 542218 577404 542454
rect 576804 542134 577404 542218
rect 576804 541898 576986 542134
rect 577222 541898 577404 542134
rect 576804 506454 577404 541898
rect 576804 506218 576986 506454
rect 577222 506218 577404 506454
rect 576804 506134 577404 506218
rect 576804 505898 576986 506134
rect 577222 505898 577404 506134
rect 576804 470454 577404 505898
rect 576804 470218 576986 470454
rect 577222 470218 577404 470454
rect 576804 470134 577404 470218
rect 576804 469898 576986 470134
rect 577222 469898 577404 470134
rect 576804 434454 577404 469898
rect 576804 434218 576986 434454
rect 577222 434218 577404 434454
rect 576804 434134 577404 434218
rect 576804 433898 576986 434134
rect 577222 433898 577404 434134
rect 576804 398454 577404 433898
rect 576804 398218 576986 398454
rect 577222 398218 577404 398454
rect 576804 398134 577404 398218
rect 576804 397898 576986 398134
rect 577222 397898 577404 398134
rect 576804 362454 577404 397898
rect 576804 362218 576986 362454
rect 577222 362218 577404 362454
rect 576804 362134 577404 362218
rect 576804 361898 576986 362134
rect 577222 361898 577404 362134
rect 576804 326454 577404 361898
rect 576804 326218 576986 326454
rect 577222 326218 577404 326454
rect 576804 326134 577404 326218
rect 576804 325898 576986 326134
rect 577222 325898 577404 326134
rect 576804 290454 577404 325898
rect 576804 290218 576986 290454
rect 577222 290218 577404 290454
rect 576804 290134 577404 290218
rect 576804 289898 576986 290134
rect 577222 289898 577404 290134
rect 576804 254454 577404 289898
rect 576804 254218 576986 254454
rect 577222 254218 577404 254454
rect 576804 254134 577404 254218
rect 576804 253898 576986 254134
rect 577222 253898 577404 254134
rect 576804 218454 577404 253898
rect 576804 218218 576986 218454
rect 577222 218218 577404 218454
rect 576804 218134 577404 218218
rect 576804 217898 576986 218134
rect 577222 217898 577404 218134
rect 576804 182454 577404 217898
rect 576804 182218 576986 182454
rect 577222 182218 577404 182454
rect 576804 182134 577404 182218
rect 576804 181898 576986 182134
rect 577222 181898 577404 182134
rect 576804 146454 577404 181898
rect 576804 146218 576986 146454
rect 577222 146218 577404 146454
rect 576804 146134 577404 146218
rect 576804 145898 576986 146134
rect 577222 145898 577404 146134
rect 576804 110454 577404 145898
rect 576804 110218 576986 110454
rect 577222 110218 577404 110454
rect 576804 110134 577404 110218
rect 576804 109898 576986 110134
rect 577222 109898 577404 110134
rect 576804 74454 577404 109898
rect 576804 74218 576986 74454
rect 577222 74218 577404 74454
rect 576804 74134 577404 74218
rect 576804 73898 576986 74134
rect 577222 73898 577404 74134
rect 576804 38454 577404 73898
rect 576804 38218 576986 38454
rect 577222 38218 577404 38454
rect 576804 38134 577404 38218
rect 576804 37898 576986 38134
rect 577222 37898 577404 38134
rect 576804 2454 577404 37898
rect 576804 2218 576986 2454
rect 577222 2218 577404 2454
rect 576804 2134 577404 2218
rect 576804 1898 576986 2134
rect 577222 1898 577404 2134
rect 576804 -346 577404 1898
rect 576804 -582 576986 -346
rect 577222 -582 577404 -346
rect 576804 -666 577404 -582
rect 576804 -902 576986 -666
rect 577222 -902 577404 -666
rect 576804 -1844 577404 -902
rect 580404 690054 581004 706122
rect 587160 706678 587760 706700
rect 587160 706442 587342 706678
rect 587578 706442 587760 706678
rect 587160 706358 587760 706442
rect 587160 706122 587342 706358
rect 587578 706122 587760 706358
rect 586240 705758 586840 705780
rect 586240 705522 586422 705758
rect 586658 705522 586840 705758
rect 586240 705438 586840 705522
rect 586240 705202 586422 705438
rect 586658 705202 586840 705438
rect 580404 689818 580586 690054
rect 580822 689818 581004 690054
rect 580404 689734 581004 689818
rect 580404 689498 580586 689734
rect 580822 689498 581004 689734
rect 580404 654054 581004 689498
rect 580404 653818 580586 654054
rect 580822 653818 581004 654054
rect 580404 653734 581004 653818
rect 580404 653498 580586 653734
rect 580822 653498 581004 653734
rect 580404 618054 581004 653498
rect 580404 617818 580586 618054
rect 580822 617818 581004 618054
rect 580404 617734 581004 617818
rect 580404 617498 580586 617734
rect 580822 617498 581004 617734
rect 580404 582054 581004 617498
rect 580404 581818 580586 582054
rect 580822 581818 581004 582054
rect 580404 581734 581004 581818
rect 580404 581498 580586 581734
rect 580822 581498 581004 581734
rect 580404 546054 581004 581498
rect 580404 545818 580586 546054
rect 580822 545818 581004 546054
rect 580404 545734 581004 545818
rect 580404 545498 580586 545734
rect 580822 545498 581004 545734
rect 580404 510054 581004 545498
rect 580404 509818 580586 510054
rect 580822 509818 581004 510054
rect 580404 509734 581004 509818
rect 580404 509498 580586 509734
rect 580822 509498 581004 509734
rect 580404 474054 581004 509498
rect 580404 473818 580586 474054
rect 580822 473818 581004 474054
rect 580404 473734 581004 473818
rect 580404 473498 580586 473734
rect 580822 473498 581004 473734
rect 580404 438054 581004 473498
rect 580404 437818 580586 438054
rect 580822 437818 581004 438054
rect 580404 437734 581004 437818
rect 580404 437498 580586 437734
rect 580822 437498 581004 437734
rect 580404 402054 581004 437498
rect 580404 401818 580586 402054
rect 580822 401818 581004 402054
rect 580404 401734 581004 401818
rect 580404 401498 580586 401734
rect 580822 401498 581004 401734
rect 580404 366054 581004 401498
rect 580404 365818 580586 366054
rect 580822 365818 581004 366054
rect 580404 365734 581004 365818
rect 580404 365498 580586 365734
rect 580822 365498 581004 365734
rect 580404 330054 581004 365498
rect 580404 329818 580586 330054
rect 580822 329818 581004 330054
rect 580404 329734 581004 329818
rect 580404 329498 580586 329734
rect 580822 329498 581004 329734
rect 580404 294054 581004 329498
rect 580404 293818 580586 294054
rect 580822 293818 581004 294054
rect 580404 293734 581004 293818
rect 580404 293498 580586 293734
rect 580822 293498 581004 293734
rect 580404 258054 581004 293498
rect 580404 257818 580586 258054
rect 580822 257818 581004 258054
rect 580404 257734 581004 257818
rect 580404 257498 580586 257734
rect 580822 257498 581004 257734
rect 580404 222054 581004 257498
rect 580404 221818 580586 222054
rect 580822 221818 581004 222054
rect 580404 221734 581004 221818
rect 580404 221498 580586 221734
rect 580822 221498 581004 221734
rect 580404 186054 581004 221498
rect 580404 185818 580586 186054
rect 580822 185818 581004 186054
rect 580404 185734 581004 185818
rect 580404 185498 580586 185734
rect 580822 185498 581004 185734
rect 580404 150054 581004 185498
rect 580404 149818 580586 150054
rect 580822 149818 581004 150054
rect 580404 149734 581004 149818
rect 580404 149498 580586 149734
rect 580822 149498 581004 149734
rect 580404 114054 581004 149498
rect 580404 113818 580586 114054
rect 580822 113818 581004 114054
rect 580404 113734 581004 113818
rect 580404 113498 580586 113734
rect 580822 113498 581004 113734
rect 580404 78054 581004 113498
rect 580404 77818 580586 78054
rect 580822 77818 581004 78054
rect 580404 77734 581004 77818
rect 580404 77498 580586 77734
rect 580822 77498 581004 77734
rect 580404 42054 581004 77498
rect 580404 41818 580586 42054
rect 580822 41818 581004 42054
rect 580404 41734 581004 41818
rect 580404 41498 580586 41734
rect 580822 41498 581004 41734
rect 580404 6054 581004 41498
rect 580404 5818 580586 6054
rect 580822 5818 581004 6054
rect 580404 5734 581004 5818
rect 580404 5498 580586 5734
rect 580822 5498 581004 5734
rect 580404 -2186 581004 5498
rect 585320 704838 585920 704860
rect 585320 704602 585502 704838
rect 585738 704602 585920 704838
rect 585320 704518 585920 704602
rect 585320 704282 585502 704518
rect 585738 704282 585920 704518
rect 585320 686454 585920 704282
rect 585320 686218 585502 686454
rect 585738 686218 585920 686454
rect 585320 686134 585920 686218
rect 585320 685898 585502 686134
rect 585738 685898 585920 686134
rect 585320 650454 585920 685898
rect 585320 650218 585502 650454
rect 585738 650218 585920 650454
rect 585320 650134 585920 650218
rect 585320 649898 585502 650134
rect 585738 649898 585920 650134
rect 585320 614454 585920 649898
rect 585320 614218 585502 614454
rect 585738 614218 585920 614454
rect 585320 614134 585920 614218
rect 585320 613898 585502 614134
rect 585738 613898 585920 614134
rect 585320 578454 585920 613898
rect 585320 578218 585502 578454
rect 585738 578218 585920 578454
rect 585320 578134 585920 578218
rect 585320 577898 585502 578134
rect 585738 577898 585920 578134
rect 585320 542454 585920 577898
rect 585320 542218 585502 542454
rect 585738 542218 585920 542454
rect 585320 542134 585920 542218
rect 585320 541898 585502 542134
rect 585738 541898 585920 542134
rect 585320 506454 585920 541898
rect 585320 506218 585502 506454
rect 585738 506218 585920 506454
rect 585320 506134 585920 506218
rect 585320 505898 585502 506134
rect 585738 505898 585920 506134
rect 585320 470454 585920 505898
rect 585320 470218 585502 470454
rect 585738 470218 585920 470454
rect 585320 470134 585920 470218
rect 585320 469898 585502 470134
rect 585738 469898 585920 470134
rect 585320 434454 585920 469898
rect 585320 434218 585502 434454
rect 585738 434218 585920 434454
rect 585320 434134 585920 434218
rect 585320 433898 585502 434134
rect 585738 433898 585920 434134
rect 585320 398454 585920 433898
rect 585320 398218 585502 398454
rect 585738 398218 585920 398454
rect 585320 398134 585920 398218
rect 585320 397898 585502 398134
rect 585738 397898 585920 398134
rect 585320 362454 585920 397898
rect 585320 362218 585502 362454
rect 585738 362218 585920 362454
rect 585320 362134 585920 362218
rect 585320 361898 585502 362134
rect 585738 361898 585920 362134
rect 585320 326454 585920 361898
rect 585320 326218 585502 326454
rect 585738 326218 585920 326454
rect 585320 326134 585920 326218
rect 585320 325898 585502 326134
rect 585738 325898 585920 326134
rect 585320 290454 585920 325898
rect 585320 290218 585502 290454
rect 585738 290218 585920 290454
rect 585320 290134 585920 290218
rect 585320 289898 585502 290134
rect 585738 289898 585920 290134
rect 585320 254454 585920 289898
rect 585320 254218 585502 254454
rect 585738 254218 585920 254454
rect 585320 254134 585920 254218
rect 585320 253898 585502 254134
rect 585738 253898 585920 254134
rect 585320 218454 585920 253898
rect 585320 218218 585502 218454
rect 585738 218218 585920 218454
rect 585320 218134 585920 218218
rect 585320 217898 585502 218134
rect 585738 217898 585920 218134
rect 585320 182454 585920 217898
rect 585320 182218 585502 182454
rect 585738 182218 585920 182454
rect 585320 182134 585920 182218
rect 585320 181898 585502 182134
rect 585738 181898 585920 182134
rect 585320 146454 585920 181898
rect 585320 146218 585502 146454
rect 585738 146218 585920 146454
rect 585320 146134 585920 146218
rect 585320 145898 585502 146134
rect 585738 145898 585920 146134
rect 585320 110454 585920 145898
rect 585320 110218 585502 110454
rect 585738 110218 585920 110454
rect 585320 110134 585920 110218
rect 585320 109898 585502 110134
rect 585738 109898 585920 110134
rect 585320 74454 585920 109898
rect 585320 74218 585502 74454
rect 585738 74218 585920 74454
rect 585320 74134 585920 74218
rect 585320 73898 585502 74134
rect 585738 73898 585920 74134
rect 585320 38454 585920 73898
rect 585320 38218 585502 38454
rect 585738 38218 585920 38454
rect 585320 38134 585920 38218
rect 585320 37898 585502 38134
rect 585738 37898 585920 38134
rect 585320 2454 585920 37898
rect 585320 2218 585502 2454
rect 585738 2218 585920 2454
rect 585320 2134 585920 2218
rect 585320 1898 585502 2134
rect 585738 1898 585920 2134
rect 585320 -346 585920 1898
rect 585320 -582 585502 -346
rect 585738 -582 585920 -346
rect 585320 -666 585920 -582
rect 585320 -902 585502 -666
rect 585738 -902 585920 -666
rect 585320 -924 585920 -902
rect 586240 668454 586840 705202
rect 586240 668218 586422 668454
rect 586658 668218 586840 668454
rect 586240 668134 586840 668218
rect 586240 667898 586422 668134
rect 586658 667898 586840 668134
rect 586240 632454 586840 667898
rect 586240 632218 586422 632454
rect 586658 632218 586840 632454
rect 586240 632134 586840 632218
rect 586240 631898 586422 632134
rect 586658 631898 586840 632134
rect 586240 596454 586840 631898
rect 586240 596218 586422 596454
rect 586658 596218 586840 596454
rect 586240 596134 586840 596218
rect 586240 595898 586422 596134
rect 586658 595898 586840 596134
rect 586240 560454 586840 595898
rect 586240 560218 586422 560454
rect 586658 560218 586840 560454
rect 586240 560134 586840 560218
rect 586240 559898 586422 560134
rect 586658 559898 586840 560134
rect 586240 524454 586840 559898
rect 586240 524218 586422 524454
rect 586658 524218 586840 524454
rect 586240 524134 586840 524218
rect 586240 523898 586422 524134
rect 586658 523898 586840 524134
rect 586240 488454 586840 523898
rect 586240 488218 586422 488454
rect 586658 488218 586840 488454
rect 586240 488134 586840 488218
rect 586240 487898 586422 488134
rect 586658 487898 586840 488134
rect 586240 452454 586840 487898
rect 586240 452218 586422 452454
rect 586658 452218 586840 452454
rect 586240 452134 586840 452218
rect 586240 451898 586422 452134
rect 586658 451898 586840 452134
rect 586240 416454 586840 451898
rect 586240 416218 586422 416454
rect 586658 416218 586840 416454
rect 586240 416134 586840 416218
rect 586240 415898 586422 416134
rect 586658 415898 586840 416134
rect 586240 380454 586840 415898
rect 586240 380218 586422 380454
rect 586658 380218 586840 380454
rect 586240 380134 586840 380218
rect 586240 379898 586422 380134
rect 586658 379898 586840 380134
rect 586240 344454 586840 379898
rect 586240 344218 586422 344454
rect 586658 344218 586840 344454
rect 586240 344134 586840 344218
rect 586240 343898 586422 344134
rect 586658 343898 586840 344134
rect 586240 308454 586840 343898
rect 586240 308218 586422 308454
rect 586658 308218 586840 308454
rect 586240 308134 586840 308218
rect 586240 307898 586422 308134
rect 586658 307898 586840 308134
rect 586240 272454 586840 307898
rect 586240 272218 586422 272454
rect 586658 272218 586840 272454
rect 586240 272134 586840 272218
rect 586240 271898 586422 272134
rect 586658 271898 586840 272134
rect 586240 236454 586840 271898
rect 586240 236218 586422 236454
rect 586658 236218 586840 236454
rect 586240 236134 586840 236218
rect 586240 235898 586422 236134
rect 586658 235898 586840 236134
rect 586240 200454 586840 235898
rect 586240 200218 586422 200454
rect 586658 200218 586840 200454
rect 586240 200134 586840 200218
rect 586240 199898 586422 200134
rect 586658 199898 586840 200134
rect 586240 164454 586840 199898
rect 586240 164218 586422 164454
rect 586658 164218 586840 164454
rect 586240 164134 586840 164218
rect 586240 163898 586422 164134
rect 586658 163898 586840 164134
rect 586240 128454 586840 163898
rect 586240 128218 586422 128454
rect 586658 128218 586840 128454
rect 586240 128134 586840 128218
rect 586240 127898 586422 128134
rect 586658 127898 586840 128134
rect 586240 92454 586840 127898
rect 586240 92218 586422 92454
rect 586658 92218 586840 92454
rect 586240 92134 586840 92218
rect 586240 91898 586422 92134
rect 586658 91898 586840 92134
rect 586240 56454 586840 91898
rect 586240 56218 586422 56454
rect 586658 56218 586840 56454
rect 586240 56134 586840 56218
rect 586240 55898 586422 56134
rect 586658 55898 586840 56134
rect 586240 20454 586840 55898
rect 586240 20218 586422 20454
rect 586658 20218 586840 20454
rect 586240 20134 586840 20218
rect 586240 19898 586422 20134
rect 586658 19898 586840 20134
rect 586240 -1266 586840 19898
rect 586240 -1502 586422 -1266
rect 586658 -1502 586840 -1266
rect 586240 -1586 586840 -1502
rect 586240 -1822 586422 -1586
rect 586658 -1822 586840 -1586
rect 586240 -1844 586840 -1822
rect 587160 690054 587760 706122
rect 587160 689818 587342 690054
rect 587578 689818 587760 690054
rect 587160 689734 587760 689818
rect 587160 689498 587342 689734
rect 587578 689498 587760 689734
rect 587160 654054 587760 689498
rect 587160 653818 587342 654054
rect 587578 653818 587760 654054
rect 587160 653734 587760 653818
rect 587160 653498 587342 653734
rect 587578 653498 587760 653734
rect 587160 618054 587760 653498
rect 587160 617818 587342 618054
rect 587578 617818 587760 618054
rect 587160 617734 587760 617818
rect 587160 617498 587342 617734
rect 587578 617498 587760 617734
rect 587160 582054 587760 617498
rect 587160 581818 587342 582054
rect 587578 581818 587760 582054
rect 587160 581734 587760 581818
rect 587160 581498 587342 581734
rect 587578 581498 587760 581734
rect 587160 546054 587760 581498
rect 587160 545818 587342 546054
rect 587578 545818 587760 546054
rect 587160 545734 587760 545818
rect 587160 545498 587342 545734
rect 587578 545498 587760 545734
rect 587160 510054 587760 545498
rect 587160 509818 587342 510054
rect 587578 509818 587760 510054
rect 587160 509734 587760 509818
rect 587160 509498 587342 509734
rect 587578 509498 587760 509734
rect 587160 474054 587760 509498
rect 587160 473818 587342 474054
rect 587578 473818 587760 474054
rect 587160 473734 587760 473818
rect 587160 473498 587342 473734
rect 587578 473498 587760 473734
rect 587160 438054 587760 473498
rect 587160 437818 587342 438054
rect 587578 437818 587760 438054
rect 587160 437734 587760 437818
rect 587160 437498 587342 437734
rect 587578 437498 587760 437734
rect 587160 402054 587760 437498
rect 587160 401818 587342 402054
rect 587578 401818 587760 402054
rect 587160 401734 587760 401818
rect 587160 401498 587342 401734
rect 587578 401498 587760 401734
rect 587160 366054 587760 401498
rect 587160 365818 587342 366054
rect 587578 365818 587760 366054
rect 587160 365734 587760 365818
rect 587160 365498 587342 365734
rect 587578 365498 587760 365734
rect 587160 330054 587760 365498
rect 587160 329818 587342 330054
rect 587578 329818 587760 330054
rect 587160 329734 587760 329818
rect 587160 329498 587342 329734
rect 587578 329498 587760 329734
rect 587160 294054 587760 329498
rect 587160 293818 587342 294054
rect 587578 293818 587760 294054
rect 587160 293734 587760 293818
rect 587160 293498 587342 293734
rect 587578 293498 587760 293734
rect 587160 258054 587760 293498
rect 587160 257818 587342 258054
rect 587578 257818 587760 258054
rect 587160 257734 587760 257818
rect 587160 257498 587342 257734
rect 587578 257498 587760 257734
rect 587160 222054 587760 257498
rect 587160 221818 587342 222054
rect 587578 221818 587760 222054
rect 587160 221734 587760 221818
rect 587160 221498 587342 221734
rect 587578 221498 587760 221734
rect 587160 186054 587760 221498
rect 587160 185818 587342 186054
rect 587578 185818 587760 186054
rect 587160 185734 587760 185818
rect 587160 185498 587342 185734
rect 587578 185498 587760 185734
rect 587160 150054 587760 185498
rect 587160 149818 587342 150054
rect 587578 149818 587760 150054
rect 587160 149734 587760 149818
rect 587160 149498 587342 149734
rect 587578 149498 587760 149734
rect 587160 114054 587760 149498
rect 587160 113818 587342 114054
rect 587578 113818 587760 114054
rect 587160 113734 587760 113818
rect 587160 113498 587342 113734
rect 587578 113498 587760 113734
rect 587160 78054 587760 113498
rect 587160 77818 587342 78054
rect 587578 77818 587760 78054
rect 587160 77734 587760 77818
rect 587160 77498 587342 77734
rect 587578 77498 587760 77734
rect 587160 42054 587760 77498
rect 587160 41818 587342 42054
rect 587578 41818 587760 42054
rect 587160 41734 587760 41818
rect 587160 41498 587342 41734
rect 587578 41498 587760 41734
rect 587160 6054 587760 41498
rect 587160 5818 587342 6054
rect 587578 5818 587760 6054
rect 587160 5734 587760 5818
rect 587160 5498 587342 5734
rect 587578 5498 587760 5734
rect 580404 -2422 580586 -2186
rect 580822 -2422 581004 -2186
rect 580404 -2506 581004 -2422
rect 580404 -2742 580586 -2506
rect 580822 -2742 581004 -2506
rect 580404 -3684 581004 -2742
rect 587160 -2186 587760 5498
rect 587160 -2422 587342 -2186
rect 587578 -2422 587760 -2186
rect 587160 -2506 587760 -2422
rect 587160 -2742 587342 -2506
rect 587578 -2742 587760 -2506
rect 587160 -2764 587760 -2742
rect 588080 672054 588680 707042
rect 588080 671818 588262 672054
rect 588498 671818 588680 672054
rect 588080 671734 588680 671818
rect 588080 671498 588262 671734
rect 588498 671498 588680 671734
rect 588080 636054 588680 671498
rect 588080 635818 588262 636054
rect 588498 635818 588680 636054
rect 588080 635734 588680 635818
rect 588080 635498 588262 635734
rect 588498 635498 588680 635734
rect 588080 600054 588680 635498
rect 588080 599818 588262 600054
rect 588498 599818 588680 600054
rect 588080 599734 588680 599818
rect 588080 599498 588262 599734
rect 588498 599498 588680 599734
rect 588080 564054 588680 599498
rect 588080 563818 588262 564054
rect 588498 563818 588680 564054
rect 588080 563734 588680 563818
rect 588080 563498 588262 563734
rect 588498 563498 588680 563734
rect 588080 528054 588680 563498
rect 588080 527818 588262 528054
rect 588498 527818 588680 528054
rect 588080 527734 588680 527818
rect 588080 527498 588262 527734
rect 588498 527498 588680 527734
rect 588080 492054 588680 527498
rect 588080 491818 588262 492054
rect 588498 491818 588680 492054
rect 588080 491734 588680 491818
rect 588080 491498 588262 491734
rect 588498 491498 588680 491734
rect 588080 456054 588680 491498
rect 588080 455818 588262 456054
rect 588498 455818 588680 456054
rect 588080 455734 588680 455818
rect 588080 455498 588262 455734
rect 588498 455498 588680 455734
rect 588080 420054 588680 455498
rect 588080 419818 588262 420054
rect 588498 419818 588680 420054
rect 588080 419734 588680 419818
rect 588080 419498 588262 419734
rect 588498 419498 588680 419734
rect 588080 384054 588680 419498
rect 588080 383818 588262 384054
rect 588498 383818 588680 384054
rect 588080 383734 588680 383818
rect 588080 383498 588262 383734
rect 588498 383498 588680 383734
rect 588080 348054 588680 383498
rect 588080 347818 588262 348054
rect 588498 347818 588680 348054
rect 588080 347734 588680 347818
rect 588080 347498 588262 347734
rect 588498 347498 588680 347734
rect 588080 312054 588680 347498
rect 588080 311818 588262 312054
rect 588498 311818 588680 312054
rect 588080 311734 588680 311818
rect 588080 311498 588262 311734
rect 588498 311498 588680 311734
rect 588080 276054 588680 311498
rect 588080 275818 588262 276054
rect 588498 275818 588680 276054
rect 588080 275734 588680 275818
rect 588080 275498 588262 275734
rect 588498 275498 588680 275734
rect 588080 240054 588680 275498
rect 588080 239818 588262 240054
rect 588498 239818 588680 240054
rect 588080 239734 588680 239818
rect 588080 239498 588262 239734
rect 588498 239498 588680 239734
rect 588080 204054 588680 239498
rect 588080 203818 588262 204054
rect 588498 203818 588680 204054
rect 588080 203734 588680 203818
rect 588080 203498 588262 203734
rect 588498 203498 588680 203734
rect 588080 168054 588680 203498
rect 588080 167818 588262 168054
rect 588498 167818 588680 168054
rect 588080 167734 588680 167818
rect 588080 167498 588262 167734
rect 588498 167498 588680 167734
rect 588080 132054 588680 167498
rect 588080 131818 588262 132054
rect 588498 131818 588680 132054
rect 588080 131734 588680 131818
rect 588080 131498 588262 131734
rect 588498 131498 588680 131734
rect 588080 96054 588680 131498
rect 588080 95818 588262 96054
rect 588498 95818 588680 96054
rect 588080 95734 588680 95818
rect 588080 95498 588262 95734
rect 588498 95498 588680 95734
rect 588080 60054 588680 95498
rect 588080 59818 588262 60054
rect 588498 59818 588680 60054
rect 588080 59734 588680 59818
rect 588080 59498 588262 59734
rect 588498 59498 588680 59734
rect 588080 24054 588680 59498
rect 588080 23818 588262 24054
rect 588498 23818 588680 24054
rect 588080 23734 588680 23818
rect 588080 23498 588262 23734
rect 588498 23498 588680 23734
rect 588080 -3106 588680 23498
rect 588080 -3342 588262 -3106
rect 588498 -3342 588680 -3106
rect 588080 -3426 588680 -3342
rect 588080 -3662 588262 -3426
rect 588498 -3662 588680 -3426
rect 588080 -3684 588680 -3662
rect 589000 693654 589600 707962
rect 589000 693418 589182 693654
rect 589418 693418 589600 693654
rect 589000 693334 589600 693418
rect 589000 693098 589182 693334
rect 589418 693098 589600 693334
rect 589000 657654 589600 693098
rect 589000 657418 589182 657654
rect 589418 657418 589600 657654
rect 589000 657334 589600 657418
rect 589000 657098 589182 657334
rect 589418 657098 589600 657334
rect 589000 621654 589600 657098
rect 589000 621418 589182 621654
rect 589418 621418 589600 621654
rect 589000 621334 589600 621418
rect 589000 621098 589182 621334
rect 589418 621098 589600 621334
rect 589000 585654 589600 621098
rect 589000 585418 589182 585654
rect 589418 585418 589600 585654
rect 589000 585334 589600 585418
rect 589000 585098 589182 585334
rect 589418 585098 589600 585334
rect 589000 549654 589600 585098
rect 589000 549418 589182 549654
rect 589418 549418 589600 549654
rect 589000 549334 589600 549418
rect 589000 549098 589182 549334
rect 589418 549098 589600 549334
rect 589000 513654 589600 549098
rect 589000 513418 589182 513654
rect 589418 513418 589600 513654
rect 589000 513334 589600 513418
rect 589000 513098 589182 513334
rect 589418 513098 589600 513334
rect 589000 477654 589600 513098
rect 589000 477418 589182 477654
rect 589418 477418 589600 477654
rect 589000 477334 589600 477418
rect 589000 477098 589182 477334
rect 589418 477098 589600 477334
rect 589000 441654 589600 477098
rect 589000 441418 589182 441654
rect 589418 441418 589600 441654
rect 589000 441334 589600 441418
rect 589000 441098 589182 441334
rect 589418 441098 589600 441334
rect 589000 405654 589600 441098
rect 589000 405418 589182 405654
rect 589418 405418 589600 405654
rect 589000 405334 589600 405418
rect 589000 405098 589182 405334
rect 589418 405098 589600 405334
rect 589000 369654 589600 405098
rect 589000 369418 589182 369654
rect 589418 369418 589600 369654
rect 589000 369334 589600 369418
rect 589000 369098 589182 369334
rect 589418 369098 589600 369334
rect 589000 333654 589600 369098
rect 589000 333418 589182 333654
rect 589418 333418 589600 333654
rect 589000 333334 589600 333418
rect 589000 333098 589182 333334
rect 589418 333098 589600 333334
rect 589000 297654 589600 333098
rect 589000 297418 589182 297654
rect 589418 297418 589600 297654
rect 589000 297334 589600 297418
rect 589000 297098 589182 297334
rect 589418 297098 589600 297334
rect 589000 261654 589600 297098
rect 589000 261418 589182 261654
rect 589418 261418 589600 261654
rect 589000 261334 589600 261418
rect 589000 261098 589182 261334
rect 589418 261098 589600 261334
rect 589000 225654 589600 261098
rect 589000 225418 589182 225654
rect 589418 225418 589600 225654
rect 589000 225334 589600 225418
rect 589000 225098 589182 225334
rect 589418 225098 589600 225334
rect 589000 189654 589600 225098
rect 589000 189418 589182 189654
rect 589418 189418 589600 189654
rect 589000 189334 589600 189418
rect 589000 189098 589182 189334
rect 589418 189098 589600 189334
rect 589000 153654 589600 189098
rect 589000 153418 589182 153654
rect 589418 153418 589600 153654
rect 589000 153334 589600 153418
rect 589000 153098 589182 153334
rect 589418 153098 589600 153334
rect 589000 117654 589600 153098
rect 589000 117418 589182 117654
rect 589418 117418 589600 117654
rect 589000 117334 589600 117418
rect 589000 117098 589182 117334
rect 589418 117098 589600 117334
rect 589000 81654 589600 117098
rect 589000 81418 589182 81654
rect 589418 81418 589600 81654
rect 589000 81334 589600 81418
rect 589000 81098 589182 81334
rect 589418 81098 589600 81334
rect 589000 45654 589600 81098
rect 589000 45418 589182 45654
rect 589418 45418 589600 45654
rect 589000 45334 589600 45418
rect 589000 45098 589182 45334
rect 589418 45098 589600 45334
rect 589000 9654 589600 45098
rect 589000 9418 589182 9654
rect 589418 9418 589600 9654
rect 589000 9334 589600 9418
rect 589000 9098 589182 9334
rect 589418 9098 589600 9334
rect 589000 -4026 589600 9098
rect 589000 -4262 589182 -4026
rect 589418 -4262 589600 -4026
rect 589000 -4346 589600 -4262
rect 589000 -4582 589182 -4346
rect 589418 -4582 589600 -4346
rect 589000 -4604 589600 -4582
rect 589920 675654 590520 708882
rect 589920 675418 590102 675654
rect 590338 675418 590520 675654
rect 589920 675334 590520 675418
rect 589920 675098 590102 675334
rect 590338 675098 590520 675334
rect 589920 639654 590520 675098
rect 589920 639418 590102 639654
rect 590338 639418 590520 639654
rect 589920 639334 590520 639418
rect 589920 639098 590102 639334
rect 590338 639098 590520 639334
rect 589920 603654 590520 639098
rect 589920 603418 590102 603654
rect 590338 603418 590520 603654
rect 589920 603334 590520 603418
rect 589920 603098 590102 603334
rect 590338 603098 590520 603334
rect 589920 567654 590520 603098
rect 589920 567418 590102 567654
rect 590338 567418 590520 567654
rect 589920 567334 590520 567418
rect 589920 567098 590102 567334
rect 590338 567098 590520 567334
rect 589920 531654 590520 567098
rect 589920 531418 590102 531654
rect 590338 531418 590520 531654
rect 589920 531334 590520 531418
rect 589920 531098 590102 531334
rect 590338 531098 590520 531334
rect 589920 495654 590520 531098
rect 589920 495418 590102 495654
rect 590338 495418 590520 495654
rect 589920 495334 590520 495418
rect 589920 495098 590102 495334
rect 590338 495098 590520 495334
rect 589920 459654 590520 495098
rect 589920 459418 590102 459654
rect 590338 459418 590520 459654
rect 589920 459334 590520 459418
rect 589920 459098 590102 459334
rect 590338 459098 590520 459334
rect 589920 423654 590520 459098
rect 589920 423418 590102 423654
rect 590338 423418 590520 423654
rect 589920 423334 590520 423418
rect 589920 423098 590102 423334
rect 590338 423098 590520 423334
rect 589920 387654 590520 423098
rect 589920 387418 590102 387654
rect 590338 387418 590520 387654
rect 589920 387334 590520 387418
rect 589920 387098 590102 387334
rect 590338 387098 590520 387334
rect 589920 351654 590520 387098
rect 589920 351418 590102 351654
rect 590338 351418 590520 351654
rect 589920 351334 590520 351418
rect 589920 351098 590102 351334
rect 590338 351098 590520 351334
rect 589920 315654 590520 351098
rect 589920 315418 590102 315654
rect 590338 315418 590520 315654
rect 589920 315334 590520 315418
rect 589920 315098 590102 315334
rect 590338 315098 590520 315334
rect 589920 279654 590520 315098
rect 589920 279418 590102 279654
rect 590338 279418 590520 279654
rect 589920 279334 590520 279418
rect 589920 279098 590102 279334
rect 590338 279098 590520 279334
rect 589920 243654 590520 279098
rect 589920 243418 590102 243654
rect 590338 243418 590520 243654
rect 589920 243334 590520 243418
rect 589920 243098 590102 243334
rect 590338 243098 590520 243334
rect 589920 207654 590520 243098
rect 589920 207418 590102 207654
rect 590338 207418 590520 207654
rect 589920 207334 590520 207418
rect 589920 207098 590102 207334
rect 590338 207098 590520 207334
rect 589920 171654 590520 207098
rect 589920 171418 590102 171654
rect 590338 171418 590520 171654
rect 589920 171334 590520 171418
rect 589920 171098 590102 171334
rect 590338 171098 590520 171334
rect 589920 135654 590520 171098
rect 589920 135418 590102 135654
rect 590338 135418 590520 135654
rect 589920 135334 590520 135418
rect 589920 135098 590102 135334
rect 590338 135098 590520 135334
rect 589920 99654 590520 135098
rect 589920 99418 590102 99654
rect 590338 99418 590520 99654
rect 589920 99334 590520 99418
rect 589920 99098 590102 99334
rect 590338 99098 590520 99334
rect 589920 63654 590520 99098
rect 589920 63418 590102 63654
rect 590338 63418 590520 63654
rect 589920 63334 590520 63418
rect 589920 63098 590102 63334
rect 590338 63098 590520 63334
rect 589920 27654 590520 63098
rect 589920 27418 590102 27654
rect 590338 27418 590520 27654
rect 589920 27334 590520 27418
rect 589920 27098 590102 27334
rect 590338 27098 590520 27334
rect 589920 -4946 590520 27098
rect 589920 -5182 590102 -4946
rect 590338 -5182 590520 -4946
rect 589920 -5266 590520 -5182
rect 589920 -5502 590102 -5266
rect 590338 -5502 590520 -5266
rect 589920 -5524 590520 -5502
rect 590840 697254 591440 709802
rect 590840 697018 591022 697254
rect 591258 697018 591440 697254
rect 590840 696934 591440 697018
rect 590840 696698 591022 696934
rect 591258 696698 591440 696934
rect 590840 661254 591440 696698
rect 590840 661018 591022 661254
rect 591258 661018 591440 661254
rect 590840 660934 591440 661018
rect 590840 660698 591022 660934
rect 591258 660698 591440 660934
rect 590840 625254 591440 660698
rect 590840 625018 591022 625254
rect 591258 625018 591440 625254
rect 590840 624934 591440 625018
rect 590840 624698 591022 624934
rect 591258 624698 591440 624934
rect 590840 589254 591440 624698
rect 590840 589018 591022 589254
rect 591258 589018 591440 589254
rect 590840 588934 591440 589018
rect 590840 588698 591022 588934
rect 591258 588698 591440 588934
rect 590840 553254 591440 588698
rect 590840 553018 591022 553254
rect 591258 553018 591440 553254
rect 590840 552934 591440 553018
rect 590840 552698 591022 552934
rect 591258 552698 591440 552934
rect 590840 517254 591440 552698
rect 590840 517018 591022 517254
rect 591258 517018 591440 517254
rect 590840 516934 591440 517018
rect 590840 516698 591022 516934
rect 591258 516698 591440 516934
rect 590840 481254 591440 516698
rect 590840 481018 591022 481254
rect 591258 481018 591440 481254
rect 590840 480934 591440 481018
rect 590840 480698 591022 480934
rect 591258 480698 591440 480934
rect 590840 445254 591440 480698
rect 590840 445018 591022 445254
rect 591258 445018 591440 445254
rect 590840 444934 591440 445018
rect 590840 444698 591022 444934
rect 591258 444698 591440 444934
rect 590840 409254 591440 444698
rect 590840 409018 591022 409254
rect 591258 409018 591440 409254
rect 590840 408934 591440 409018
rect 590840 408698 591022 408934
rect 591258 408698 591440 408934
rect 590840 373254 591440 408698
rect 590840 373018 591022 373254
rect 591258 373018 591440 373254
rect 590840 372934 591440 373018
rect 590840 372698 591022 372934
rect 591258 372698 591440 372934
rect 590840 337254 591440 372698
rect 590840 337018 591022 337254
rect 591258 337018 591440 337254
rect 590840 336934 591440 337018
rect 590840 336698 591022 336934
rect 591258 336698 591440 336934
rect 590840 301254 591440 336698
rect 590840 301018 591022 301254
rect 591258 301018 591440 301254
rect 590840 300934 591440 301018
rect 590840 300698 591022 300934
rect 591258 300698 591440 300934
rect 590840 265254 591440 300698
rect 590840 265018 591022 265254
rect 591258 265018 591440 265254
rect 590840 264934 591440 265018
rect 590840 264698 591022 264934
rect 591258 264698 591440 264934
rect 590840 229254 591440 264698
rect 590840 229018 591022 229254
rect 591258 229018 591440 229254
rect 590840 228934 591440 229018
rect 590840 228698 591022 228934
rect 591258 228698 591440 228934
rect 590840 193254 591440 228698
rect 590840 193018 591022 193254
rect 591258 193018 591440 193254
rect 590840 192934 591440 193018
rect 590840 192698 591022 192934
rect 591258 192698 591440 192934
rect 590840 157254 591440 192698
rect 590840 157018 591022 157254
rect 591258 157018 591440 157254
rect 590840 156934 591440 157018
rect 590840 156698 591022 156934
rect 591258 156698 591440 156934
rect 590840 121254 591440 156698
rect 590840 121018 591022 121254
rect 591258 121018 591440 121254
rect 590840 120934 591440 121018
rect 590840 120698 591022 120934
rect 591258 120698 591440 120934
rect 590840 85254 591440 120698
rect 590840 85018 591022 85254
rect 591258 85018 591440 85254
rect 590840 84934 591440 85018
rect 590840 84698 591022 84934
rect 591258 84698 591440 84934
rect 590840 49254 591440 84698
rect 590840 49018 591022 49254
rect 591258 49018 591440 49254
rect 590840 48934 591440 49018
rect 590840 48698 591022 48934
rect 591258 48698 591440 48934
rect 590840 13254 591440 48698
rect 590840 13018 591022 13254
rect 591258 13018 591440 13254
rect 590840 12934 591440 13018
rect 590840 12698 591022 12934
rect 591258 12698 591440 12934
rect 590840 -5866 591440 12698
rect 590840 -6102 591022 -5866
rect 591258 -6102 591440 -5866
rect 590840 -6186 591440 -6102
rect 590840 -6422 591022 -6186
rect 591258 -6422 591440 -6186
rect 590840 -6444 591440 -6422
rect 591760 679254 592360 710722
rect 591760 679018 591942 679254
rect 592178 679018 592360 679254
rect 591760 678934 592360 679018
rect 591760 678698 591942 678934
rect 592178 678698 592360 678934
rect 591760 643254 592360 678698
rect 591760 643018 591942 643254
rect 592178 643018 592360 643254
rect 591760 642934 592360 643018
rect 591760 642698 591942 642934
rect 592178 642698 592360 642934
rect 591760 607254 592360 642698
rect 591760 607018 591942 607254
rect 592178 607018 592360 607254
rect 591760 606934 592360 607018
rect 591760 606698 591942 606934
rect 592178 606698 592360 606934
rect 591760 571254 592360 606698
rect 591760 571018 591942 571254
rect 592178 571018 592360 571254
rect 591760 570934 592360 571018
rect 591760 570698 591942 570934
rect 592178 570698 592360 570934
rect 591760 535254 592360 570698
rect 591760 535018 591942 535254
rect 592178 535018 592360 535254
rect 591760 534934 592360 535018
rect 591760 534698 591942 534934
rect 592178 534698 592360 534934
rect 591760 499254 592360 534698
rect 591760 499018 591942 499254
rect 592178 499018 592360 499254
rect 591760 498934 592360 499018
rect 591760 498698 591942 498934
rect 592178 498698 592360 498934
rect 591760 463254 592360 498698
rect 591760 463018 591942 463254
rect 592178 463018 592360 463254
rect 591760 462934 592360 463018
rect 591760 462698 591942 462934
rect 592178 462698 592360 462934
rect 591760 427254 592360 462698
rect 591760 427018 591942 427254
rect 592178 427018 592360 427254
rect 591760 426934 592360 427018
rect 591760 426698 591942 426934
rect 592178 426698 592360 426934
rect 591760 391254 592360 426698
rect 591760 391018 591942 391254
rect 592178 391018 592360 391254
rect 591760 390934 592360 391018
rect 591760 390698 591942 390934
rect 592178 390698 592360 390934
rect 591760 355254 592360 390698
rect 591760 355018 591942 355254
rect 592178 355018 592360 355254
rect 591760 354934 592360 355018
rect 591760 354698 591942 354934
rect 592178 354698 592360 354934
rect 591760 319254 592360 354698
rect 591760 319018 591942 319254
rect 592178 319018 592360 319254
rect 591760 318934 592360 319018
rect 591760 318698 591942 318934
rect 592178 318698 592360 318934
rect 591760 283254 592360 318698
rect 591760 283018 591942 283254
rect 592178 283018 592360 283254
rect 591760 282934 592360 283018
rect 591760 282698 591942 282934
rect 592178 282698 592360 282934
rect 591760 247254 592360 282698
rect 591760 247018 591942 247254
rect 592178 247018 592360 247254
rect 591760 246934 592360 247018
rect 591760 246698 591942 246934
rect 592178 246698 592360 246934
rect 591760 211254 592360 246698
rect 591760 211018 591942 211254
rect 592178 211018 592360 211254
rect 591760 210934 592360 211018
rect 591760 210698 591942 210934
rect 592178 210698 592360 210934
rect 591760 175254 592360 210698
rect 591760 175018 591942 175254
rect 592178 175018 592360 175254
rect 591760 174934 592360 175018
rect 591760 174698 591942 174934
rect 592178 174698 592360 174934
rect 591760 139254 592360 174698
rect 591760 139018 591942 139254
rect 592178 139018 592360 139254
rect 591760 138934 592360 139018
rect 591760 138698 591942 138934
rect 592178 138698 592360 138934
rect 591760 103254 592360 138698
rect 591760 103018 591942 103254
rect 592178 103018 592360 103254
rect 591760 102934 592360 103018
rect 591760 102698 591942 102934
rect 592178 102698 592360 102934
rect 591760 67254 592360 102698
rect 591760 67018 591942 67254
rect 592178 67018 592360 67254
rect 591760 66934 592360 67018
rect 591760 66698 591942 66934
rect 592178 66698 592360 66934
rect 591760 31254 592360 66698
rect 591760 31018 591942 31254
rect 592178 31018 592360 31254
rect 591760 30934 592360 31018
rect 591760 30698 591942 30934
rect 592178 30698 592360 30934
rect 569604 -7022 569786 -6786
rect 570022 -7022 570204 -6786
rect 569604 -7106 570204 -7022
rect 569604 -7342 569786 -7106
rect 570022 -7342 570204 -7106
rect 569604 -7364 570204 -7342
rect 591760 -6786 592360 30698
rect 591760 -7022 591942 -6786
rect 592178 -7022 592360 -6786
rect 591760 -7106 592360 -7022
rect 591760 -7342 591942 -7106
rect 592178 -7342 592360 -7106
rect 591760 -7364 592360 -7342
<< via4 >>
rect -8254 711042 -8018 711278
rect -8254 710722 -8018 710958
rect -8254 679018 -8018 679254
rect -8254 678698 -8018 678934
rect -8254 643018 -8018 643254
rect -8254 642698 -8018 642934
rect -8254 607018 -8018 607254
rect -8254 606698 -8018 606934
rect -8254 571018 -8018 571254
rect -8254 570698 -8018 570934
rect -8254 535018 -8018 535254
rect -8254 534698 -8018 534934
rect -8254 499018 -8018 499254
rect -8254 498698 -8018 498934
rect -8254 463018 -8018 463254
rect -8254 462698 -8018 462934
rect -8254 427018 -8018 427254
rect -8254 426698 -8018 426934
rect -8254 391018 -8018 391254
rect -8254 390698 -8018 390934
rect -8254 355018 -8018 355254
rect -8254 354698 -8018 354934
rect -8254 319018 -8018 319254
rect -8254 318698 -8018 318934
rect -8254 283018 -8018 283254
rect -8254 282698 -8018 282934
rect -8254 247018 -8018 247254
rect -8254 246698 -8018 246934
rect -8254 211018 -8018 211254
rect -8254 210698 -8018 210934
rect -8254 175018 -8018 175254
rect -8254 174698 -8018 174934
rect -8254 139018 -8018 139254
rect -8254 138698 -8018 138934
rect -8254 103018 -8018 103254
rect -8254 102698 -8018 102934
rect -8254 67018 -8018 67254
rect -8254 66698 -8018 66934
rect -8254 31018 -8018 31254
rect -8254 30698 -8018 30934
rect -7334 710122 -7098 710358
rect -7334 709802 -7098 710038
rect 11786 710122 12022 710358
rect 11786 709802 12022 710038
rect -7334 697018 -7098 697254
rect -7334 696698 -7098 696934
rect -7334 661018 -7098 661254
rect -7334 660698 -7098 660934
rect -7334 625018 -7098 625254
rect -7334 624698 -7098 624934
rect -7334 589018 -7098 589254
rect -7334 588698 -7098 588934
rect -7334 553018 -7098 553254
rect -7334 552698 -7098 552934
rect -7334 517018 -7098 517254
rect -7334 516698 -7098 516934
rect -7334 481018 -7098 481254
rect -7334 480698 -7098 480934
rect -7334 445018 -7098 445254
rect -7334 444698 -7098 444934
rect -7334 409018 -7098 409254
rect -7334 408698 -7098 408934
rect -7334 373018 -7098 373254
rect -7334 372698 -7098 372934
rect -7334 337018 -7098 337254
rect -7334 336698 -7098 336934
rect -7334 301018 -7098 301254
rect -7334 300698 -7098 300934
rect -7334 265018 -7098 265254
rect -7334 264698 -7098 264934
rect -7334 229018 -7098 229254
rect -7334 228698 -7098 228934
rect -7334 193018 -7098 193254
rect -7334 192698 -7098 192934
rect -7334 157018 -7098 157254
rect -7334 156698 -7098 156934
rect -7334 121018 -7098 121254
rect -7334 120698 -7098 120934
rect -7334 85018 -7098 85254
rect -7334 84698 -7098 84934
rect -7334 49018 -7098 49254
rect -7334 48698 -7098 48934
rect -7334 13018 -7098 13254
rect -7334 12698 -7098 12934
rect -6414 709202 -6178 709438
rect -6414 708882 -6178 709118
rect -6414 675418 -6178 675654
rect -6414 675098 -6178 675334
rect -6414 639418 -6178 639654
rect -6414 639098 -6178 639334
rect -6414 603418 -6178 603654
rect -6414 603098 -6178 603334
rect -6414 567418 -6178 567654
rect -6414 567098 -6178 567334
rect -6414 531418 -6178 531654
rect -6414 531098 -6178 531334
rect -6414 495418 -6178 495654
rect -6414 495098 -6178 495334
rect -6414 459418 -6178 459654
rect -6414 459098 -6178 459334
rect -6414 423418 -6178 423654
rect -6414 423098 -6178 423334
rect -6414 387418 -6178 387654
rect -6414 387098 -6178 387334
rect -6414 351418 -6178 351654
rect -6414 351098 -6178 351334
rect -6414 315418 -6178 315654
rect -6414 315098 -6178 315334
rect -6414 279418 -6178 279654
rect -6414 279098 -6178 279334
rect -6414 243418 -6178 243654
rect -6414 243098 -6178 243334
rect -6414 207418 -6178 207654
rect -6414 207098 -6178 207334
rect -6414 171418 -6178 171654
rect -6414 171098 -6178 171334
rect -6414 135418 -6178 135654
rect -6414 135098 -6178 135334
rect -6414 99418 -6178 99654
rect -6414 99098 -6178 99334
rect -6414 63418 -6178 63654
rect -6414 63098 -6178 63334
rect -6414 27418 -6178 27654
rect -6414 27098 -6178 27334
rect -5494 708282 -5258 708518
rect -5494 707962 -5258 708198
rect 8186 708282 8422 708518
rect 8186 707962 8422 708198
rect -5494 693418 -5258 693654
rect -5494 693098 -5258 693334
rect -5494 657418 -5258 657654
rect -5494 657098 -5258 657334
rect -5494 621418 -5258 621654
rect -5494 621098 -5258 621334
rect -5494 585418 -5258 585654
rect -5494 585098 -5258 585334
rect -5494 549418 -5258 549654
rect -5494 549098 -5258 549334
rect -5494 513418 -5258 513654
rect -5494 513098 -5258 513334
rect -5494 477418 -5258 477654
rect -5494 477098 -5258 477334
rect -5494 441418 -5258 441654
rect -5494 441098 -5258 441334
rect -5494 405418 -5258 405654
rect -5494 405098 -5258 405334
rect -5494 369418 -5258 369654
rect -5494 369098 -5258 369334
rect -5494 333418 -5258 333654
rect -5494 333098 -5258 333334
rect -5494 297418 -5258 297654
rect -5494 297098 -5258 297334
rect -5494 261418 -5258 261654
rect -5494 261098 -5258 261334
rect -5494 225418 -5258 225654
rect -5494 225098 -5258 225334
rect -5494 189418 -5258 189654
rect -5494 189098 -5258 189334
rect -5494 153418 -5258 153654
rect -5494 153098 -5258 153334
rect -5494 117418 -5258 117654
rect -5494 117098 -5258 117334
rect -5494 81418 -5258 81654
rect -5494 81098 -5258 81334
rect -5494 45418 -5258 45654
rect -5494 45098 -5258 45334
rect -5494 9418 -5258 9654
rect -5494 9098 -5258 9334
rect -4574 707362 -4338 707598
rect -4574 707042 -4338 707278
rect -4574 671818 -4338 672054
rect -4574 671498 -4338 671734
rect -4574 635818 -4338 636054
rect -4574 635498 -4338 635734
rect -4574 599818 -4338 600054
rect -4574 599498 -4338 599734
rect -4574 563818 -4338 564054
rect -4574 563498 -4338 563734
rect -4574 527818 -4338 528054
rect -4574 527498 -4338 527734
rect -4574 491818 -4338 492054
rect -4574 491498 -4338 491734
rect -4574 455818 -4338 456054
rect -4574 455498 -4338 455734
rect -4574 419818 -4338 420054
rect -4574 419498 -4338 419734
rect -4574 383818 -4338 384054
rect -4574 383498 -4338 383734
rect -4574 347818 -4338 348054
rect -4574 347498 -4338 347734
rect -4574 311818 -4338 312054
rect -4574 311498 -4338 311734
rect -4574 275818 -4338 276054
rect -4574 275498 -4338 275734
rect -4574 239818 -4338 240054
rect -4574 239498 -4338 239734
rect -4574 203818 -4338 204054
rect -4574 203498 -4338 203734
rect -4574 167818 -4338 168054
rect -4574 167498 -4338 167734
rect -4574 131818 -4338 132054
rect -4574 131498 -4338 131734
rect -4574 95818 -4338 96054
rect -4574 95498 -4338 95734
rect -4574 59818 -4338 60054
rect -4574 59498 -4338 59734
rect -4574 23818 -4338 24054
rect -4574 23498 -4338 23734
rect -3654 706442 -3418 706678
rect -3654 706122 -3418 706358
rect 4586 706442 4822 706678
rect 4586 706122 4822 706358
rect -3654 689818 -3418 690054
rect -3654 689498 -3418 689734
rect -3654 653818 -3418 654054
rect -3654 653498 -3418 653734
rect -3654 617818 -3418 618054
rect -3654 617498 -3418 617734
rect -3654 581818 -3418 582054
rect -3654 581498 -3418 581734
rect -3654 545818 -3418 546054
rect -3654 545498 -3418 545734
rect -3654 509818 -3418 510054
rect -3654 509498 -3418 509734
rect -3654 473818 -3418 474054
rect -3654 473498 -3418 473734
rect -3654 437818 -3418 438054
rect -3654 437498 -3418 437734
rect -3654 401818 -3418 402054
rect -3654 401498 -3418 401734
rect -3654 365818 -3418 366054
rect -3654 365498 -3418 365734
rect -3654 329818 -3418 330054
rect -3654 329498 -3418 329734
rect -3654 293818 -3418 294054
rect -3654 293498 -3418 293734
rect -3654 257818 -3418 258054
rect -3654 257498 -3418 257734
rect -3654 221818 -3418 222054
rect -3654 221498 -3418 221734
rect -3654 185818 -3418 186054
rect -3654 185498 -3418 185734
rect -3654 149818 -3418 150054
rect -3654 149498 -3418 149734
rect -3654 113818 -3418 114054
rect -3654 113498 -3418 113734
rect -3654 77818 -3418 78054
rect -3654 77498 -3418 77734
rect -3654 41818 -3418 42054
rect -3654 41498 -3418 41734
rect -3654 5818 -3418 6054
rect -3654 5498 -3418 5734
rect -2734 705522 -2498 705758
rect -2734 705202 -2498 705438
rect -2734 668218 -2498 668454
rect -2734 667898 -2498 668134
rect -2734 632218 -2498 632454
rect -2734 631898 -2498 632134
rect -2734 596218 -2498 596454
rect -2734 595898 -2498 596134
rect -2734 560218 -2498 560454
rect -2734 559898 -2498 560134
rect -2734 524218 -2498 524454
rect -2734 523898 -2498 524134
rect -2734 488218 -2498 488454
rect -2734 487898 -2498 488134
rect -2734 452218 -2498 452454
rect -2734 451898 -2498 452134
rect -2734 416218 -2498 416454
rect -2734 415898 -2498 416134
rect -2734 380218 -2498 380454
rect -2734 379898 -2498 380134
rect -2734 344218 -2498 344454
rect -2734 343898 -2498 344134
rect -2734 308218 -2498 308454
rect -2734 307898 -2498 308134
rect -2734 272218 -2498 272454
rect -2734 271898 -2498 272134
rect -2734 236218 -2498 236454
rect -2734 235898 -2498 236134
rect -2734 200218 -2498 200454
rect -2734 199898 -2498 200134
rect -2734 164218 -2498 164454
rect -2734 163898 -2498 164134
rect -2734 128218 -2498 128454
rect -2734 127898 -2498 128134
rect -2734 92218 -2498 92454
rect -2734 91898 -2498 92134
rect -2734 56218 -2498 56454
rect -2734 55898 -2498 56134
rect -2734 20218 -2498 20454
rect -2734 19898 -2498 20134
rect -1814 704602 -1578 704838
rect -1814 704282 -1578 704518
rect -1814 686218 -1578 686454
rect -1814 685898 -1578 686134
rect -1814 650218 -1578 650454
rect -1814 649898 -1578 650134
rect -1814 614218 -1578 614454
rect -1814 613898 -1578 614134
rect -1814 578218 -1578 578454
rect -1814 577898 -1578 578134
rect -1814 542218 -1578 542454
rect -1814 541898 -1578 542134
rect -1814 506218 -1578 506454
rect -1814 505898 -1578 506134
rect -1814 470218 -1578 470454
rect -1814 469898 -1578 470134
rect -1814 434218 -1578 434454
rect -1814 433898 -1578 434134
rect -1814 398218 -1578 398454
rect -1814 397898 -1578 398134
rect -1814 362218 -1578 362454
rect -1814 361898 -1578 362134
rect -1814 326218 -1578 326454
rect -1814 325898 -1578 326134
rect -1814 290218 -1578 290454
rect -1814 289898 -1578 290134
rect -1814 254218 -1578 254454
rect -1814 253898 -1578 254134
rect -1814 218218 -1578 218454
rect -1814 217898 -1578 218134
rect -1814 182218 -1578 182454
rect -1814 181898 -1578 182134
rect -1814 146218 -1578 146454
rect -1814 145898 -1578 146134
rect -1814 110218 -1578 110454
rect -1814 109898 -1578 110134
rect -1814 74218 -1578 74454
rect -1814 73898 -1578 74134
rect -1814 38218 -1578 38454
rect -1814 37898 -1578 38134
rect -1814 2218 -1578 2454
rect -1814 1898 -1578 2134
rect -1814 -582 -1578 -346
rect -1814 -902 -1578 -666
rect 986 704602 1222 704838
rect 986 704282 1222 704518
rect 986 686218 1222 686454
rect 986 685898 1222 686134
rect 986 650218 1222 650454
rect 986 649898 1222 650134
rect 986 614218 1222 614454
rect 986 613898 1222 614134
rect 986 578218 1222 578454
rect 986 577898 1222 578134
rect 986 542218 1222 542454
rect 986 541898 1222 542134
rect 986 506218 1222 506454
rect 986 505898 1222 506134
rect 986 470218 1222 470454
rect 986 469898 1222 470134
rect 986 434218 1222 434454
rect 986 433898 1222 434134
rect 986 398218 1222 398454
rect 986 397898 1222 398134
rect 986 362218 1222 362454
rect 986 361898 1222 362134
rect 986 326218 1222 326454
rect 986 325898 1222 326134
rect 986 290218 1222 290454
rect 986 289898 1222 290134
rect 986 254218 1222 254454
rect 986 253898 1222 254134
rect 986 218218 1222 218454
rect 986 217898 1222 218134
rect 986 182218 1222 182454
rect 986 181898 1222 182134
rect 986 146218 1222 146454
rect 986 145898 1222 146134
rect 986 110218 1222 110454
rect 986 109898 1222 110134
rect 986 74218 1222 74454
rect 986 73898 1222 74134
rect 986 38218 1222 38454
rect 986 37898 1222 38134
rect 986 2218 1222 2454
rect 986 1898 1222 2134
rect 986 -582 1222 -346
rect 986 -902 1222 -666
rect -2734 -1502 -2498 -1266
rect -2734 -1822 -2498 -1586
rect 4586 689818 4822 690054
rect 4586 689498 4822 689734
rect 4586 653818 4822 654054
rect 4586 653498 4822 653734
rect 4586 617818 4822 618054
rect 4586 617498 4822 617734
rect 4586 581818 4822 582054
rect 4586 581498 4822 581734
rect 4586 545818 4822 546054
rect 4586 545498 4822 545734
rect 4586 509818 4822 510054
rect 4586 509498 4822 509734
rect 4586 473818 4822 474054
rect 4586 473498 4822 473734
rect 4586 437818 4822 438054
rect 4586 437498 4822 437734
rect 4586 401818 4822 402054
rect 4586 401498 4822 401734
rect 4586 365818 4822 366054
rect 4586 365498 4822 365734
rect 4586 329818 4822 330054
rect 4586 329498 4822 329734
rect 4586 293818 4822 294054
rect 4586 293498 4822 293734
rect 4586 257818 4822 258054
rect 4586 257498 4822 257734
rect 4586 221818 4822 222054
rect 4586 221498 4822 221734
rect 4586 185818 4822 186054
rect 4586 185498 4822 185734
rect 4586 149818 4822 150054
rect 4586 149498 4822 149734
rect 4586 113818 4822 114054
rect 4586 113498 4822 113734
rect 4586 77818 4822 78054
rect 4586 77498 4822 77734
rect 4586 41818 4822 42054
rect 4586 41498 4822 41734
rect 4586 5818 4822 6054
rect 4586 5498 4822 5734
rect -3654 -2422 -3418 -2186
rect -3654 -2742 -3418 -2506
rect 4586 -2422 4822 -2186
rect 4586 -2742 4822 -2506
rect -4574 -3342 -4338 -3106
rect -4574 -3662 -4338 -3426
rect 8186 693418 8422 693654
rect 8186 693098 8422 693334
rect 8186 657418 8422 657654
rect 8186 657098 8422 657334
rect 8186 621418 8422 621654
rect 8186 621098 8422 621334
rect 8186 585418 8422 585654
rect 8186 585098 8422 585334
rect 8186 549418 8422 549654
rect 8186 549098 8422 549334
rect 8186 513418 8422 513654
rect 8186 513098 8422 513334
rect 8186 477418 8422 477654
rect 8186 477098 8422 477334
rect 8186 441418 8422 441654
rect 8186 441098 8422 441334
rect 8186 405418 8422 405654
rect 8186 405098 8422 405334
rect 8186 369418 8422 369654
rect 8186 369098 8422 369334
rect 8186 333418 8422 333654
rect 8186 333098 8422 333334
rect 8186 297418 8422 297654
rect 8186 297098 8422 297334
rect 8186 261418 8422 261654
rect 8186 261098 8422 261334
rect 8186 225418 8422 225654
rect 8186 225098 8422 225334
rect 8186 189418 8422 189654
rect 8186 189098 8422 189334
rect 8186 153418 8422 153654
rect 8186 153098 8422 153334
rect 8186 117418 8422 117654
rect 8186 117098 8422 117334
rect 8186 81418 8422 81654
rect 8186 81098 8422 81334
rect 8186 45418 8422 45654
rect 8186 45098 8422 45334
rect 8186 9418 8422 9654
rect 8186 9098 8422 9334
rect -5494 -4262 -5258 -4026
rect -5494 -4582 -5258 -4346
rect 8186 -4262 8422 -4026
rect 8186 -4582 8422 -4346
rect -6414 -5182 -6178 -4946
rect -6414 -5502 -6178 -5266
rect 29786 711042 30022 711278
rect 29786 710722 30022 710958
rect 26186 709202 26422 709438
rect 26186 708882 26422 709118
rect 22586 707362 22822 707598
rect 22586 707042 22822 707278
rect 11786 697018 12022 697254
rect 11786 696698 12022 696934
rect 11786 661018 12022 661254
rect 11786 660698 12022 660934
rect 11786 625018 12022 625254
rect 11786 624698 12022 624934
rect 11786 589018 12022 589254
rect 11786 588698 12022 588934
rect 11786 553018 12022 553254
rect 11786 552698 12022 552934
rect 11786 517018 12022 517254
rect 11786 516698 12022 516934
rect 11786 481018 12022 481254
rect 11786 480698 12022 480934
rect 11786 445018 12022 445254
rect 11786 444698 12022 444934
rect 11786 409018 12022 409254
rect 11786 408698 12022 408934
rect 11786 373018 12022 373254
rect 11786 372698 12022 372934
rect 11786 337018 12022 337254
rect 11786 336698 12022 336934
rect 11786 301018 12022 301254
rect 11786 300698 12022 300934
rect 11786 265018 12022 265254
rect 11786 264698 12022 264934
rect 11786 229018 12022 229254
rect 11786 228698 12022 228934
rect 11786 193018 12022 193254
rect 11786 192698 12022 192934
rect 11786 157018 12022 157254
rect 11786 156698 12022 156934
rect 11786 121018 12022 121254
rect 11786 120698 12022 120934
rect 11786 85018 12022 85254
rect 11786 84698 12022 84934
rect 11786 49018 12022 49254
rect 11786 48698 12022 48934
rect 11786 13018 12022 13254
rect 11786 12698 12022 12934
rect -7334 -6102 -7098 -5866
rect -7334 -6422 -7098 -6186
rect 18986 705522 19222 705758
rect 18986 705202 19222 705438
rect 18986 668218 19222 668454
rect 18986 667898 19222 668134
rect 18986 632218 19222 632454
rect 18986 631898 19222 632134
rect 18986 596218 19222 596454
rect 18986 595898 19222 596134
rect 18986 560218 19222 560454
rect 18986 559898 19222 560134
rect 18986 524218 19222 524454
rect 18986 523898 19222 524134
rect 18986 488218 19222 488454
rect 18986 487898 19222 488134
rect 18986 452218 19222 452454
rect 18986 451898 19222 452134
rect 18986 416218 19222 416454
rect 18986 415898 19222 416134
rect 18986 380218 19222 380454
rect 18986 379898 19222 380134
rect 18986 344218 19222 344454
rect 18986 343898 19222 344134
rect 18986 308218 19222 308454
rect 18986 307898 19222 308134
rect 18986 272218 19222 272454
rect 18986 271898 19222 272134
rect 18986 236218 19222 236454
rect 18986 235898 19222 236134
rect 18986 200218 19222 200454
rect 18986 199898 19222 200134
rect 18986 164218 19222 164454
rect 18986 163898 19222 164134
rect 18986 128218 19222 128454
rect 18986 127898 19222 128134
rect 18986 92218 19222 92454
rect 18986 91898 19222 92134
rect 18986 56218 19222 56454
rect 18986 55898 19222 56134
rect 18986 20218 19222 20454
rect 18986 19898 19222 20134
rect 18986 -1502 19222 -1266
rect 18986 -1822 19222 -1586
rect 22586 671818 22822 672054
rect 22586 671498 22822 671734
rect 22586 635818 22822 636054
rect 22586 635498 22822 635734
rect 22586 599818 22822 600054
rect 22586 599498 22822 599734
rect 22586 563818 22822 564054
rect 22586 563498 22822 563734
rect 22586 527818 22822 528054
rect 22586 527498 22822 527734
rect 22586 491818 22822 492054
rect 22586 491498 22822 491734
rect 22586 455818 22822 456054
rect 22586 455498 22822 455734
rect 22586 419818 22822 420054
rect 22586 419498 22822 419734
rect 22586 383818 22822 384054
rect 22586 383498 22822 383734
rect 22586 347818 22822 348054
rect 22586 347498 22822 347734
rect 22586 311818 22822 312054
rect 22586 311498 22822 311734
rect 22586 275818 22822 276054
rect 22586 275498 22822 275734
rect 22586 239818 22822 240054
rect 22586 239498 22822 239734
rect 22586 203818 22822 204054
rect 22586 203498 22822 203734
rect 22586 167818 22822 168054
rect 22586 167498 22822 167734
rect 22586 131818 22822 132054
rect 22586 131498 22822 131734
rect 22586 95818 22822 96054
rect 22586 95498 22822 95734
rect 22586 59818 22822 60054
rect 22586 59498 22822 59734
rect 22586 23818 22822 24054
rect 22586 23498 22822 23734
rect 22586 -3342 22822 -3106
rect 22586 -3662 22822 -3426
rect 26186 675418 26422 675654
rect 26186 675098 26422 675334
rect 26186 639418 26422 639654
rect 26186 639098 26422 639334
rect 26186 603418 26422 603654
rect 26186 603098 26422 603334
rect 26186 567418 26422 567654
rect 26186 567098 26422 567334
rect 26186 531418 26422 531654
rect 26186 531098 26422 531334
rect 26186 495418 26422 495654
rect 26186 495098 26422 495334
rect 26186 459418 26422 459654
rect 26186 459098 26422 459334
rect 26186 423418 26422 423654
rect 26186 423098 26422 423334
rect 26186 387418 26422 387654
rect 26186 387098 26422 387334
rect 26186 351418 26422 351654
rect 26186 351098 26422 351334
rect 26186 315418 26422 315654
rect 26186 315098 26422 315334
rect 26186 279418 26422 279654
rect 26186 279098 26422 279334
rect 26186 243418 26422 243654
rect 26186 243098 26422 243334
rect 26186 207418 26422 207654
rect 26186 207098 26422 207334
rect 26186 171418 26422 171654
rect 26186 171098 26422 171334
rect 26186 135418 26422 135654
rect 26186 135098 26422 135334
rect 26186 99418 26422 99654
rect 26186 99098 26422 99334
rect 26186 63418 26422 63654
rect 26186 63098 26422 63334
rect 26186 27418 26422 27654
rect 26186 27098 26422 27334
rect 26186 -5182 26422 -4946
rect 26186 -5502 26422 -5266
rect 47786 710122 48022 710358
rect 47786 709802 48022 710038
rect 44186 708282 44422 708518
rect 44186 707962 44422 708198
rect 40586 706442 40822 706678
rect 40586 706122 40822 706358
rect 29786 679018 30022 679254
rect 29786 678698 30022 678934
rect 29786 643018 30022 643254
rect 29786 642698 30022 642934
rect 29786 607018 30022 607254
rect 29786 606698 30022 606934
rect 29786 571018 30022 571254
rect 29786 570698 30022 570934
rect 29786 535018 30022 535254
rect 29786 534698 30022 534934
rect 29786 499018 30022 499254
rect 29786 498698 30022 498934
rect 29786 463018 30022 463254
rect 29786 462698 30022 462934
rect 29786 427018 30022 427254
rect 29786 426698 30022 426934
rect 29786 391018 30022 391254
rect 29786 390698 30022 390934
rect 29786 355018 30022 355254
rect 29786 354698 30022 354934
rect 29786 319018 30022 319254
rect 29786 318698 30022 318934
rect 29786 283018 30022 283254
rect 29786 282698 30022 282934
rect 29786 247018 30022 247254
rect 29786 246698 30022 246934
rect 29786 211018 30022 211254
rect 29786 210698 30022 210934
rect 29786 175018 30022 175254
rect 29786 174698 30022 174934
rect 29786 139018 30022 139254
rect 29786 138698 30022 138934
rect 29786 103018 30022 103254
rect 29786 102698 30022 102934
rect 29786 67018 30022 67254
rect 29786 66698 30022 66934
rect 29786 31018 30022 31254
rect 29786 30698 30022 30934
rect 11786 -6102 12022 -5866
rect 11786 -6422 12022 -6186
rect -8254 -7022 -8018 -6786
rect -8254 -7342 -8018 -7106
rect 36986 704602 37222 704838
rect 36986 704282 37222 704518
rect 36986 686218 37222 686454
rect 36986 685898 37222 686134
rect 36986 650218 37222 650454
rect 36986 649898 37222 650134
rect 36986 614218 37222 614454
rect 36986 613898 37222 614134
rect 36986 578218 37222 578454
rect 36986 577898 37222 578134
rect 36986 542218 37222 542454
rect 36986 541898 37222 542134
rect 36986 506218 37222 506454
rect 36986 505898 37222 506134
rect 36986 470218 37222 470454
rect 36986 469898 37222 470134
rect 36986 434218 37222 434454
rect 36986 433898 37222 434134
rect 36986 398218 37222 398454
rect 36986 397898 37222 398134
rect 36986 362218 37222 362454
rect 36986 361898 37222 362134
rect 36986 326218 37222 326454
rect 36986 325898 37222 326134
rect 36986 290218 37222 290454
rect 36986 289898 37222 290134
rect 36986 254218 37222 254454
rect 36986 253898 37222 254134
rect 36986 218218 37222 218454
rect 36986 217898 37222 218134
rect 36986 182218 37222 182454
rect 36986 181898 37222 182134
rect 36986 146218 37222 146454
rect 36986 145898 37222 146134
rect 36986 110218 37222 110454
rect 36986 109898 37222 110134
rect 36986 74218 37222 74454
rect 36986 73898 37222 74134
rect 36986 38218 37222 38454
rect 36986 37898 37222 38134
rect 36986 2218 37222 2454
rect 36986 1898 37222 2134
rect 36986 -582 37222 -346
rect 36986 -902 37222 -666
rect 40586 689818 40822 690054
rect 40586 689498 40822 689734
rect 40586 653818 40822 654054
rect 40586 653498 40822 653734
rect 40586 617818 40822 618054
rect 40586 617498 40822 617734
rect 40586 581818 40822 582054
rect 40586 581498 40822 581734
rect 40586 545818 40822 546054
rect 40586 545498 40822 545734
rect 40586 509818 40822 510054
rect 40586 509498 40822 509734
rect 40586 473818 40822 474054
rect 40586 473498 40822 473734
rect 40586 437818 40822 438054
rect 40586 437498 40822 437734
rect 40586 401818 40822 402054
rect 40586 401498 40822 401734
rect 40586 365818 40822 366054
rect 40586 365498 40822 365734
rect 40586 329818 40822 330054
rect 40586 329498 40822 329734
rect 40586 293818 40822 294054
rect 40586 293498 40822 293734
rect 40586 257818 40822 258054
rect 40586 257498 40822 257734
rect 40586 221818 40822 222054
rect 40586 221498 40822 221734
rect 40586 185818 40822 186054
rect 40586 185498 40822 185734
rect 40586 149818 40822 150054
rect 40586 149498 40822 149734
rect 40586 113818 40822 114054
rect 40586 113498 40822 113734
rect 40586 77818 40822 78054
rect 40586 77498 40822 77734
rect 40586 41818 40822 42054
rect 40586 41498 40822 41734
rect 40586 5818 40822 6054
rect 40586 5498 40822 5734
rect 40586 -2422 40822 -2186
rect 40586 -2742 40822 -2506
rect 44186 693418 44422 693654
rect 44186 693098 44422 693334
rect 44186 657418 44422 657654
rect 44186 657098 44422 657334
rect 44186 621418 44422 621654
rect 44186 621098 44422 621334
rect 44186 585418 44422 585654
rect 44186 585098 44422 585334
rect 44186 549418 44422 549654
rect 44186 549098 44422 549334
rect 44186 513418 44422 513654
rect 44186 513098 44422 513334
rect 44186 477418 44422 477654
rect 44186 477098 44422 477334
rect 44186 441418 44422 441654
rect 44186 441098 44422 441334
rect 44186 405418 44422 405654
rect 44186 405098 44422 405334
rect 44186 369418 44422 369654
rect 44186 369098 44422 369334
rect 44186 333418 44422 333654
rect 44186 333098 44422 333334
rect 44186 297418 44422 297654
rect 44186 297098 44422 297334
rect 44186 261418 44422 261654
rect 44186 261098 44422 261334
rect 44186 225418 44422 225654
rect 44186 225098 44422 225334
rect 44186 189418 44422 189654
rect 44186 189098 44422 189334
rect 44186 153418 44422 153654
rect 44186 153098 44422 153334
rect 44186 117418 44422 117654
rect 44186 117098 44422 117334
rect 44186 81418 44422 81654
rect 44186 81098 44422 81334
rect 44186 45418 44422 45654
rect 44186 45098 44422 45334
rect 44186 9418 44422 9654
rect 44186 9098 44422 9334
rect 44186 -4262 44422 -4026
rect 44186 -4582 44422 -4346
rect 65786 711042 66022 711278
rect 65786 710722 66022 710958
rect 62186 709202 62422 709438
rect 62186 708882 62422 709118
rect 58586 707362 58822 707598
rect 58586 707042 58822 707278
rect 47786 697018 48022 697254
rect 47786 696698 48022 696934
rect 47786 661018 48022 661254
rect 47786 660698 48022 660934
rect 47786 625018 48022 625254
rect 47786 624698 48022 624934
rect 47786 589018 48022 589254
rect 47786 588698 48022 588934
rect 47786 553018 48022 553254
rect 47786 552698 48022 552934
rect 47786 517018 48022 517254
rect 47786 516698 48022 516934
rect 47786 481018 48022 481254
rect 47786 480698 48022 480934
rect 47786 445018 48022 445254
rect 47786 444698 48022 444934
rect 47786 409018 48022 409254
rect 47786 408698 48022 408934
rect 47786 373018 48022 373254
rect 47786 372698 48022 372934
rect 47786 337018 48022 337254
rect 47786 336698 48022 336934
rect 47786 301018 48022 301254
rect 47786 300698 48022 300934
rect 47786 265018 48022 265254
rect 47786 264698 48022 264934
rect 47786 229018 48022 229254
rect 47786 228698 48022 228934
rect 47786 193018 48022 193254
rect 47786 192698 48022 192934
rect 47786 157018 48022 157254
rect 47786 156698 48022 156934
rect 47786 121018 48022 121254
rect 47786 120698 48022 120934
rect 47786 85018 48022 85254
rect 47786 84698 48022 84934
rect 47786 49018 48022 49254
rect 47786 48698 48022 48934
rect 47786 13018 48022 13254
rect 47786 12698 48022 12934
rect 29786 -7022 30022 -6786
rect 29786 -7342 30022 -7106
rect 54986 705522 55222 705758
rect 54986 705202 55222 705438
rect 54986 668218 55222 668454
rect 54986 667898 55222 668134
rect 54986 632218 55222 632454
rect 54986 631898 55222 632134
rect 54986 596218 55222 596454
rect 54986 595898 55222 596134
rect 54986 560218 55222 560454
rect 54986 559898 55222 560134
rect 54986 524218 55222 524454
rect 54986 523898 55222 524134
rect 54986 488218 55222 488454
rect 54986 487898 55222 488134
rect 54986 452218 55222 452454
rect 54986 451898 55222 452134
rect 54986 416218 55222 416454
rect 54986 415898 55222 416134
rect 54986 380218 55222 380454
rect 54986 379898 55222 380134
rect 54986 344218 55222 344454
rect 54986 343898 55222 344134
rect 54986 308218 55222 308454
rect 54986 307898 55222 308134
rect 54986 272218 55222 272454
rect 54986 271898 55222 272134
rect 54986 236218 55222 236454
rect 54986 235898 55222 236134
rect 54986 200218 55222 200454
rect 54986 199898 55222 200134
rect 54986 164218 55222 164454
rect 54986 163898 55222 164134
rect 54986 128218 55222 128454
rect 54986 127898 55222 128134
rect 54986 92218 55222 92454
rect 54986 91898 55222 92134
rect 54986 56218 55222 56454
rect 54986 55898 55222 56134
rect 54986 20218 55222 20454
rect 54986 19898 55222 20134
rect 54986 -1502 55222 -1266
rect 54986 -1822 55222 -1586
rect 58586 671818 58822 672054
rect 58586 671498 58822 671734
rect 58586 635818 58822 636054
rect 58586 635498 58822 635734
rect 58586 599818 58822 600054
rect 58586 599498 58822 599734
rect 58586 563818 58822 564054
rect 58586 563498 58822 563734
rect 58586 527818 58822 528054
rect 58586 527498 58822 527734
rect 58586 491818 58822 492054
rect 58586 491498 58822 491734
rect 58586 455818 58822 456054
rect 58586 455498 58822 455734
rect 58586 419818 58822 420054
rect 58586 419498 58822 419734
rect 58586 383818 58822 384054
rect 58586 383498 58822 383734
rect 58586 347818 58822 348054
rect 58586 347498 58822 347734
rect 58586 311818 58822 312054
rect 58586 311498 58822 311734
rect 58586 275818 58822 276054
rect 58586 275498 58822 275734
rect 58586 239818 58822 240054
rect 58586 239498 58822 239734
rect 58586 203818 58822 204054
rect 58586 203498 58822 203734
rect 58586 167818 58822 168054
rect 58586 167498 58822 167734
rect 58586 131818 58822 132054
rect 58586 131498 58822 131734
rect 58586 95818 58822 96054
rect 58586 95498 58822 95734
rect 58586 59818 58822 60054
rect 58586 59498 58822 59734
rect 58586 23818 58822 24054
rect 58586 23498 58822 23734
rect 58586 -3342 58822 -3106
rect 58586 -3662 58822 -3426
rect 62186 675418 62422 675654
rect 62186 675098 62422 675334
rect 62186 639418 62422 639654
rect 62186 639098 62422 639334
rect 62186 603418 62422 603654
rect 62186 603098 62422 603334
rect 62186 567418 62422 567654
rect 62186 567098 62422 567334
rect 62186 531418 62422 531654
rect 62186 531098 62422 531334
rect 62186 495418 62422 495654
rect 62186 495098 62422 495334
rect 62186 459418 62422 459654
rect 62186 459098 62422 459334
rect 62186 423418 62422 423654
rect 62186 423098 62422 423334
rect 62186 387418 62422 387654
rect 62186 387098 62422 387334
rect 62186 351418 62422 351654
rect 62186 351098 62422 351334
rect 62186 315418 62422 315654
rect 62186 315098 62422 315334
rect 62186 279418 62422 279654
rect 62186 279098 62422 279334
rect 62186 243418 62422 243654
rect 62186 243098 62422 243334
rect 62186 207418 62422 207654
rect 62186 207098 62422 207334
rect 62186 171418 62422 171654
rect 62186 171098 62422 171334
rect 62186 135418 62422 135654
rect 62186 135098 62422 135334
rect 62186 99418 62422 99654
rect 62186 99098 62422 99334
rect 62186 63418 62422 63654
rect 62186 63098 62422 63334
rect 62186 27418 62422 27654
rect 62186 27098 62422 27334
rect 62186 -5182 62422 -4946
rect 62186 -5502 62422 -5266
rect 83786 710122 84022 710358
rect 83786 709802 84022 710038
rect 80186 708282 80422 708518
rect 80186 707962 80422 708198
rect 76586 706442 76822 706678
rect 76586 706122 76822 706358
rect 65786 679018 66022 679254
rect 65786 678698 66022 678934
rect 65786 643018 66022 643254
rect 65786 642698 66022 642934
rect 65786 607018 66022 607254
rect 65786 606698 66022 606934
rect 65786 571018 66022 571254
rect 65786 570698 66022 570934
rect 65786 535018 66022 535254
rect 65786 534698 66022 534934
rect 65786 499018 66022 499254
rect 65786 498698 66022 498934
rect 65786 463018 66022 463254
rect 65786 462698 66022 462934
rect 65786 427018 66022 427254
rect 65786 426698 66022 426934
rect 65786 391018 66022 391254
rect 65786 390698 66022 390934
rect 65786 355018 66022 355254
rect 65786 354698 66022 354934
rect 65786 319018 66022 319254
rect 65786 318698 66022 318934
rect 65786 283018 66022 283254
rect 65786 282698 66022 282934
rect 65786 247018 66022 247254
rect 65786 246698 66022 246934
rect 65786 211018 66022 211254
rect 65786 210698 66022 210934
rect 65786 175018 66022 175254
rect 65786 174698 66022 174934
rect 65786 139018 66022 139254
rect 65786 138698 66022 138934
rect 65786 103018 66022 103254
rect 65786 102698 66022 102934
rect 65786 67018 66022 67254
rect 65786 66698 66022 66934
rect 65786 31018 66022 31254
rect 65786 30698 66022 30934
rect 47786 -6102 48022 -5866
rect 47786 -6422 48022 -6186
rect 72986 704602 73222 704838
rect 72986 704282 73222 704518
rect 72986 686218 73222 686454
rect 72986 685898 73222 686134
rect 72986 650218 73222 650454
rect 72986 649898 73222 650134
rect 72986 614218 73222 614454
rect 72986 613898 73222 614134
rect 72986 578218 73222 578454
rect 72986 577898 73222 578134
rect 72986 542218 73222 542454
rect 72986 541898 73222 542134
rect 72986 506218 73222 506454
rect 72986 505898 73222 506134
rect 72986 470218 73222 470454
rect 72986 469898 73222 470134
rect 72986 434218 73222 434454
rect 72986 433898 73222 434134
rect 72986 398218 73222 398454
rect 72986 397898 73222 398134
rect 72986 362218 73222 362454
rect 72986 361898 73222 362134
rect 72986 326218 73222 326454
rect 72986 325898 73222 326134
rect 72986 290218 73222 290454
rect 72986 289898 73222 290134
rect 72986 254218 73222 254454
rect 72986 253898 73222 254134
rect 72986 218218 73222 218454
rect 72986 217898 73222 218134
rect 72986 182218 73222 182454
rect 72986 181898 73222 182134
rect 72986 146218 73222 146454
rect 72986 145898 73222 146134
rect 72986 110218 73222 110454
rect 72986 109898 73222 110134
rect 72986 74218 73222 74454
rect 72986 73898 73222 74134
rect 72986 38218 73222 38454
rect 72986 37898 73222 38134
rect 72986 2218 73222 2454
rect 72986 1898 73222 2134
rect 72986 -582 73222 -346
rect 72986 -902 73222 -666
rect 76586 689818 76822 690054
rect 76586 689498 76822 689734
rect 76586 653818 76822 654054
rect 76586 653498 76822 653734
rect 76586 617818 76822 618054
rect 76586 617498 76822 617734
rect 76586 581818 76822 582054
rect 76586 581498 76822 581734
rect 76586 545818 76822 546054
rect 76586 545498 76822 545734
rect 76586 509818 76822 510054
rect 76586 509498 76822 509734
rect 76586 473818 76822 474054
rect 76586 473498 76822 473734
rect 76586 437818 76822 438054
rect 76586 437498 76822 437734
rect 76586 401818 76822 402054
rect 76586 401498 76822 401734
rect 76586 365818 76822 366054
rect 76586 365498 76822 365734
rect 76586 329818 76822 330054
rect 76586 329498 76822 329734
rect 76586 293818 76822 294054
rect 76586 293498 76822 293734
rect 76586 257818 76822 258054
rect 76586 257498 76822 257734
rect 76586 221818 76822 222054
rect 76586 221498 76822 221734
rect 76586 185818 76822 186054
rect 76586 185498 76822 185734
rect 76586 149818 76822 150054
rect 76586 149498 76822 149734
rect 76586 113818 76822 114054
rect 76586 113498 76822 113734
rect 76586 77818 76822 78054
rect 76586 77498 76822 77734
rect 76586 41818 76822 42054
rect 76586 41498 76822 41734
rect 76586 5818 76822 6054
rect 76586 5498 76822 5734
rect 76586 -2422 76822 -2186
rect 76586 -2742 76822 -2506
rect 80186 693418 80422 693654
rect 80186 693098 80422 693334
rect 80186 657418 80422 657654
rect 80186 657098 80422 657334
rect 80186 621418 80422 621654
rect 80186 621098 80422 621334
rect 80186 585418 80422 585654
rect 80186 585098 80422 585334
rect 80186 549418 80422 549654
rect 80186 549098 80422 549334
rect 80186 513418 80422 513654
rect 80186 513098 80422 513334
rect 80186 477418 80422 477654
rect 80186 477098 80422 477334
rect 80186 441418 80422 441654
rect 80186 441098 80422 441334
rect 80186 405418 80422 405654
rect 80186 405098 80422 405334
rect 80186 369418 80422 369654
rect 80186 369098 80422 369334
rect 80186 333418 80422 333654
rect 80186 333098 80422 333334
rect 80186 297418 80422 297654
rect 80186 297098 80422 297334
rect 80186 261418 80422 261654
rect 80186 261098 80422 261334
rect 80186 225418 80422 225654
rect 80186 225098 80422 225334
rect 80186 189418 80422 189654
rect 80186 189098 80422 189334
rect 80186 153418 80422 153654
rect 80186 153098 80422 153334
rect 80186 117418 80422 117654
rect 80186 117098 80422 117334
rect 80186 81418 80422 81654
rect 80186 81098 80422 81334
rect 80186 45418 80422 45654
rect 80186 45098 80422 45334
rect 80186 9418 80422 9654
rect 80186 9098 80422 9334
rect 80186 -4262 80422 -4026
rect 80186 -4582 80422 -4346
rect 101786 711042 102022 711278
rect 101786 710722 102022 710958
rect 98186 709202 98422 709438
rect 98186 708882 98422 709118
rect 94586 707362 94822 707598
rect 94586 707042 94822 707278
rect 83786 697018 84022 697254
rect 83786 696698 84022 696934
rect 83786 661018 84022 661254
rect 83786 660698 84022 660934
rect 83786 625018 84022 625254
rect 83786 624698 84022 624934
rect 83786 589018 84022 589254
rect 83786 588698 84022 588934
rect 83786 553018 84022 553254
rect 83786 552698 84022 552934
rect 83786 517018 84022 517254
rect 83786 516698 84022 516934
rect 83786 481018 84022 481254
rect 83786 480698 84022 480934
rect 83786 445018 84022 445254
rect 83786 444698 84022 444934
rect 83786 409018 84022 409254
rect 83786 408698 84022 408934
rect 83786 373018 84022 373254
rect 83786 372698 84022 372934
rect 83786 337018 84022 337254
rect 83786 336698 84022 336934
rect 83786 301018 84022 301254
rect 83786 300698 84022 300934
rect 83786 265018 84022 265254
rect 83786 264698 84022 264934
rect 83786 229018 84022 229254
rect 83786 228698 84022 228934
rect 83786 193018 84022 193254
rect 83786 192698 84022 192934
rect 83786 157018 84022 157254
rect 83786 156698 84022 156934
rect 83786 121018 84022 121254
rect 83786 120698 84022 120934
rect 83786 85018 84022 85254
rect 83786 84698 84022 84934
rect 83786 49018 84022 49254
rect 83786 48698 84022 48934
rect 83786 13018 84022 13254
rect 83786 12698 84022 12934
rect 65786 -7022 66022 -6786
rect 65786 -7342 66022 -7106
rect 90986 705522 91222 705758
rect 90986 705202 91222 705438
rect 90986 668218 91222 668454
rect 90986 667898 91222 668134
rect 90986 632218 91222 632454
rect 90986 631898 91222 632134
rect 90986 596218 91222 596454
rect 90986 595898 91222 596134
rect 90986 560218 91222 560454
rect 90986 559898 91222 560134
rect 90986 524218 91222 524454
rect 90986 523898 91222 524134
rect 90986 488218 91222 488454
rect 90986 487898 91222 488134
rect 90986 452218 91222 452454
rect 90986 451898 91222 452134
rect 90986 416218 91222 416454
rect 90986 415898 91222 416134
rect 90986 380218 91222 380454
rect 90986 379898 91222 380134
rect 90986 344218 91222 344454
rect 90986 343898 91222 344134
rect 90986 308218 91222 308454
rect 90986 307898 91222 308134
rect 90986 272218 91222 272454
rect 90986 271898 91222 272134
rect 90986 236218 91222 236454
rect 90986 235898 91222 236134
rect 90986 200218 91222 200454
rect 90986 199898 91222 200134
rect 90986 164218 91222 164454
rect 90986 163898 91222 164134
rect 90986 128218 91222 128454
rect 90986 127898 91222 128134
rect 90986 92218 91222 92454
rect 90986 91898 91222 92134
rect 90986 56218 91222 56454
rect 90986 55898 91222 56134
rect 90986 20218 91222 20454
rect 90986 19898 91222 20134
rect 90986 -1502 91222 -1266
rect 90986 -1822 91222 -1586
rect 94586 671818 94822 672054
rect 94586 671498 94822 671734
rect 94586 635818 94822 636054
rect 94586 635498 94822 635734
rect 94586 599818 94822 600054
rect 94586 599498 94822 599734
rect 94586 563818 94822 564054
rect 94586 563498 94822 563734
rect 94586 527818 94822 528054
rect 94586 527498 94822 527734
rect 94586 491818 94822 492054
rect 94586 491498 94822 491734
rect 94586 455818 94822 456054
rect 94586 455498 94822 455734
rect 94586 419818 94822 420054
rect 94586 419498 94822 419734
rect 94586 383818 94822 384054
rect 94586 383498 94822 383734
rect 94586 347818 94822 348054
rect 94586 347498 94822 347734
rect 94586 311818 94822 312054
rect 94586 311498 94822 311734
rect 94586 275818 94822 276054
rect 94586 275498 94822 275734
rect 94586 239818 94822 240054
rect 94586 239498 94822 239734
rect 94586 203818 94822 204054
rect 94586 203498 94822 203734
rect 94586 167818 94822 168054
rect 94586 167498 94822 167734
rect 94586 131818 94822 132054
rect 94586 131498 94822 131734
rect 94586 95818 94822 96054
rect 94586 95498 94822 95734
rect 94586 59818 94822 60054
rect 94586 59498 94822 59734
rect 94586 23818 94822 24054
rect 94586 23498 94822 23734
rect 94586 -3342 94822 -3106
rect 94586 -3662 94822 -3426
rect 98186 675418 98422 675654
rect 98186 675098 98422 675334
rect 98186 639418 98422 639654
rect 98186 639098 98422 639334
rect 98186 603418 98422 603654
rect 98186 603098 98422 603334
rect 98186 567418 98422 567654
rect 98186 567098 98422 567334
rect 98186 531418 98422 531654
rect 98186 531098 98422 531334
rect 98186 495418 98422 495654
rect 98186 495098 98422 495334
rect 98186 459418 98422 459654
rect 98186 459098 98422 459334
rect 98186 423418 98422 423654
rect 98186 423098 98422 423334
rect 98186 387418 98422 387654
rect 98186 387098 98422 387334
rect 98186 351418 98422 351654
rect 98186 351098 98422 351334
rect 98186 315418 98422 315654
rect 98186 315098 98422 315334
rect 98186 279418 98422 279654
rect 98186 279098 98422 279334
rect 98186 243418 98422 243654
rect 98186 243098 98422 243334
rect 98186 207418 98422 207654
rect 98186 207098 98422 207334
rect 98186 171418 98422 171654
rect 98186 171098 98422 171334
rect 98186 135418 98422 135654
rect 98186 135098 98422 135334
rect 98186 99418 98422 99654
rect 98186 99098 98422 99334
rect 98186 63418 98422 63654
rect 98186 63098 98422 63334
rect 98186 27418 98422 27654
rect 98186 27098 98422 27334
rect 98186 -5182 98422 -4946
rect 98186 -5502 98422 -5266
rect 119786 710122 120022 710358
rect 119786 709802 120022 710038
rect 116186 708282 116422 708518
rect 116186 707962 116422 708198
rect 112586 706442 112822 706678
rect 112586 706122 112822 706358
rect 101786 679018 102022 679254
rect 101786 678698 102022 678934
rect 101786 643018 102022 643254
rect 101786 642698 102022 642934
rect 101786 607018 102022 607254
rect 101786 606698 102022 606934
rect 101786 571018 102022 571254
rect 101786 570698 102022 570934
rect 101786 535018 102022 535254
rect 101786 534698 102022 534934
rect 101786 499018 102022 499254
rect 101786 498698 102022 498934
rect 101786 463018 102022 463254
rect 101786 462698 102022 462934
rect 101786 427018 102022 427254
rect 101786 426698 102022 426934
rect 101786 391018 102022 391254
rect 101786 390698 102022 390934
rect 101786 355018 102022 355254
rect 101786 354698 102022 354934
rect 101786 319018 102022 319254
rect 101786 318698 102022 318934
rect 101786 283018 102022 283254
rect 101786 282698 102022 282934
rect 101786 247018 102022 247254
rect 101786 246698 102022 246934
rect 101786 211018 102022 211254
rect 101786 210698 102022 210934
rect 101786 175018 102022 175254
rect 101786 174698 102022 174934
rect 101786 139018 102022 139254
rect 101786 138698 102022 138934
rect 101786 103018 102022 103254
rect 101786 102698 102022 102934
rect 101786 67018 102022 67254
rect 101786 66698 102022 66934
rect 101786 31018 102022 31254
rect 101786 30698 102022 30934
rect 83786 -6102 84022 -5866
rect 83786 -6422 84022 -6186
rect 108986 704602 109222 704838
rect 108986 704282 109222 704518
rect 108986 686218 109222 686454
rect 108986 685898 109222 686134
rect 108986 650218 109222 650454
rect 108986 649898 109222 650134
rect 108986 614218 109222 614454
rect 108986 613898 109222 614134
rect 108986 578218 109222 578454
rect 108986 577898 109222 578134
rect 108986 542218 109222 542454
rect 108986 541898 109222 542134
rect 108986 506218 109222 506454
rect 108986 505898 109222 506134
rect 108986 470218 109222 470454
rect 108986 469898 109222 470134
rect 108986 434218 109222 434454
rect 108986 433898 109222 434134
rect 108986 398218 109222 398454
rect 108986 397898 109222 398134
rect 108986 362218 109222 362454
rect 108986 361898 109222 362134
rect 108986 326218 109222 326454
rect 108986 325898 109222 326134
rect 108986 290218 109222 290454
rect 108986 289898 109222 290134
rect 108986 254218 109222 254454
rect 108986 253898 109222 254134
rect 108986 218218 109222 218454
rect 108986 217898 109222 218134
rect 108986 182218 109222 182454
rect 108986 181898 109222 182134
rect 108986 146218 109222 146454
rect 108986 145898 109222 146134
rect 108986 110218 109222 110454
rect 108986 109898 109222 110134
rect 108986 74218 109222 74454
rect 108986 73898 109222 74134
rect 108986 38218 109222 38454
rect 108986 37898 109222 38134
rect 108986 2218 109222 2454
rect 108986 1898 109222 2134
rect 108986 -582 109222 -346
rect 108986 -902 109222 -666
rect 112586 689818 112822 690054
rect 112586 689498 112822 689734
rect 112586 653818 112822 654054
rect 112586 653498 112822 653734
rect 112586 617818 112822 618054
rect 112586 617498 112822 617734
rect 112586 581818 112822 582054
rect 112586 581498 112822 581734
rect 112586 545818 112822 546054
rect 112586 545498 112822 545734
rect 112586 509818 112822 510054
rect 112586 509498 112822 509734
rect 112586 473818 112822 474054
rect 112586 473498 112822 473734
rect 112586 437818 112822 438054
rect 112586 437498 112822 437734
rect 112586 401818 112822 402054
rect 112586 401498 112822 401734
rect 112586 365818 112822 366054
rect 112586 365498 112822 365734
rect 112586 329818 112822 330054
rect 112586 329498 112822 329734
rect 112586 293818 112822 294054
rect 112586 293498 112822 293734
rect 112586 257818 112822 258054
rect 112586 257498 112822 257734
rect 112586 221818 112822 222054
rect 112586 221498 112822 221734
rect 112586 185818 112822 186054
rect 112586 185498 112822 185734
rect 112586 149818 112822 150054
rect 112586 149498 112822 149734
rect 112586 113818 112822 114054
rect 112586 113498 112822 113734
rect 112586 77818 112822 78054
rect 112586 77498 112822 77734
rect 112586 41818 112822 42054
rect 112586 41498 112822 41734
rect 112586 5818 112822 6054
rect 112586 5498 112822 5734
rect 112586 -2422 112822 -2186
rect 112586 -2742 112822 -2506
rect 116186 693418 116422 693654
rect 116186 693098 116422 693334
rect 116186 657418 116422 657654
rect 116186 657098 116422 657334
rect 116186 621418 116422 621654
rect 116186 621098 116422 621334
rect 116186 585418 116422 585654
rect 116186 585098 116422 585334
rect 116186 549418 116422 549654
rect 116186 549098 116422 549334
rect 116186 513418 116422 513654
rect 116186 513098 116422 513334
rect 116186 477418 116422 477654
rect 116186 477098 116422 477334
rect 116186 441418 116422 441654
rect 116186 441098 116422 441334
rect 116186 405418 116422 405654
rect 116186 405098 116422 405334
rect 116186 369418 116422 369654
rect 116186 369098 116422 369334
rect 116186 333418 116422 333654
rect 116186 333098 116422 333334
rect 116186 297418 116422 297654
rect 116186 297098 116422 297334
rect 116186 261418 116422 261654
rect 116186 261098 116422 261334
rect 116186 225418 116422 225654
rect 116186 225098 116422 225334
rect 116186 189418 116422 189654
rect 116186 189098 116422 189334
rect 116186 153418 116422 153654
rect 116186 153098 116422 153334
rect 116186 117418 116422 117654
rect 116186 117098 116422 117334
rect 116186 81418 116422 81654
rect 116186 81098 116422 81334
rect 116186 45418 116422 45654
rect 116186 45098 116422 45334
rect 116186 9418 116422 9654
rect 116186 9098 116422 9334
rect 116186 -4262 116422 -4026
rect 116186 -4582 116422 -4346
rect 137786 711042 138022 711278
rect 137786 710722 138022 710958
rect 134186 709202 134422 709438
rect 134186 708882 134422 709118
rect 130586 707362 130822 707598
rect 130586 707042 130822 707278
rect 119786 697018 120022 697254
rect 119786 696698 120022 696934
rect 119786 661018 120022 661254
rect 119786 660698 120022 660934
rect 119786 625018 120022 625254
rect 119786 624698 120022 624934
rect 119786 589018 120022 589254
rect 119786 588698 120022 588934
rect 119786 553018 120022 553254
rect 119786 552698 120022 552934
rect 119786 517018 120022 517254
rect 119786 516698 120022 516934
rect 119786 481018 120022 481254
rect 119786 480698 120022 480934
rect 119786 445018 120022 445254
rect 119786 444698 120022 444934
rect 119786 409018 120022 409254
rect 119786 408698 120022 408934
rect 119786 373018 120022 373254
rect 119786 372698 120022 372934
rect 119786 337018 120022 337254
rect 119786 336698 120022 336934
rect 119786 301018 120022 301254
rect 119786 300698 120022 300934
rect 119786 265018 120022 265254
rect 119786 264698 120022 264934
rect 119786 229018 120022 229254
rect 119786 228698 120022 228934
rect 119786 193018 120022 193254
rect 119786 192698 120022 192934
rect 119786 157018 120022 157254
rect 119786 156698 120022 156934
rect 119786 121018 120022 121254
rect 119786 120698 120022 120934
rect 119786 85018 120022 85254
rect 119786 84698 120022 84934
rect 119786 49018 120022 49254
rect 119786 48698 120022 48934
rect 119786 13018 120022 13254
rect 119786 12698 120022 12934
rect 101786 -7022 102022 -6786
rect 101786 -7342 102022 -7106
rect 126986 705522 127222 705758
rect 126986 705202 127222 705438
rect 126986 668218 127222 668454
rect 126986 667898 127222 668134
rect 126986 632218 127222 632454
rect 126986 631898 127222 632134
rect 126986 596218 127222 596454
rect 126986 595898 127222 596134
rect 126986 560218 127222 560454
rect 126986 559898 127222 560134
rect 126986 524218 127222 524454
rect 126986 523898 127222 524134
rect 126986 488218 127222 488454
rect 126986 487898 127222 488134
rect 126986 452218 127222 452454
rect 126986 451898 127222 452134
rect 126986 416218 127222 416454
rect 126986 415898 127222 416134
rect 126986 380218 127222 380454
rect 126986 379898 127222 380134
rect 126986 344218 127222 344454
rect 126986 343898 127222 344134
rect 126986 308218 127222 308454
rect 126986 307898 127222 308134
rect 126986 272218 127222 272454
rect 126986 271898 127222 272134
rect 126986 236218 127222 236454
rect 126986 235898 127222 236134
rect 126986 200218 127222 200454
rect 126986 199898 127222 200134
rect 126986 164218 127222 164454
rect 126986 163898 127222 164134
rect 126986 128218 127222 128454
rect 126986 127898 127222 128134
rect 126986 92218 127222 92454
rect 126986 91898 127222 92134
rect 126986 56218 127222 56454
rect 126986 55898 127222 56134
rect 126986 20218 127222 20454
rect 126986 19898 127222 20134
rect 126986 -1502 127222 -1266
rect 126986 -1822 127222 -1586
rect 130586 671818 130822 672054
rect 130586 671498 130822 671734
rect 130586 635818 130822 636054
rect 130586 635498 130822 635734
rect 130586 599818 130822 600054
rect 130586 599498 130822 599734
rect 130586 563818 130822 564054
rect 130586 563498 130822 563734
rect 130586 527818 130822 528054
rect 130586 527498 130822 527734
rect 130586 491818 130822 492054
rect 130586 491498 130822 491734
rect 130586 455818 130822 456054
rect 130586 455498 130822 455734
rect 130586 419818 130822 420054
rect 130586 419498 130822 419734
rect 130586 383818 130822 384054
rect 130586 383498 130822 383734
rect 130586 347818 130822 348054
rect 130586 347498 130822 347734
rect 130586 311818 130822 312054
rect 130586 311498 130822 311734
rect 130586 275818 130822 276054
rect 130586 275498 130822 275734
rect 130586 239818 130822 240054
rect 130586 239498 130822 239734
rect 130586 203818 130822 204054
rect 130586 203498 130822 203734
rect 130586 167818 130822 168054
rect 130586 167498 130822 167734
rect 130586 131818 130822 132054
rect 130586 131498 130822 131734
rect 130586 95818 130822 96054
rect 130586 95498 130822 95734
rect 130586 59818 130822 60054
rect 130586 59498 130822 59734
rect 130586 23818 130822 24054
rect 130586 23498 130822 23734
rect 130586 -3342 130822 -3106
rect 130586 -3662 130822 -3426
rect 134186 675418 134422 675654
rect 134186 675098 134422 675334
rect 134186 639418 134422 639654
rect 134186 639098 134422 639334
rect 134186 603418 134422 603654
rect 134186 603098 134422 603334
rect 134186 567418 134422 567654
rect 134186 567098 134422 567334
rect 134186 531418 134422 531654
rect 134186 531098 134422 531334
rect 134186 495418 134422 495654
rect 134186 495098 134422 495334
rect 134186 459418 134422 459654
rect 134186 459098 134422 459334
rect 134186 423418 134422 423654
rect 134186 423098 134422 423334
rect 134186 387418 134422 387654
rect 134186 387098 134422 387334
rect 134186 351418 134422 351654
rect 134186 351098 134422 351334
rect 134186 315418 134422 315654
rect 134186 315098 134422 315334
rect 134186 279418 134422 279654
rect 134186 279098 134422 279334
rect 134186 243418 134422 243654
rect 134186 243098 134422 243334
rect 134186 207418 134422 207654
rect 134186 207098 134422 207334
rect 134186 171418 134422 171654
rect 134186 171098 134422 171334
rect 134186 135418 134422 135654
rect 134186 135098 134422 135334
rect 134186 99418 134422 99654
rect 134186 99098 134422 99334
rect 134186 63418 134422 63654
rect 134186 63098 134422 63334
rect 134186 27418 134422 27654
rect 134186 27098 134422 27334
rect 134186 -5182 134422 -4946
rect 134186 -5502 134422 -5266
rect 155786 710122 156022 710358
rect 155786 709802 156022 710038
rect 152186 708282 152422 708518
rect 152186 707962 152422 708198
rect 148586 706442 148822 706678
rect 148586 706122 148822 706358
rect 137786 679018 138022 679254
rect 137786 678698 138022 678934
rect 137786 643018 138022 643254
rect 137786 642698 138022 642934
rect 137786 607018 138022 607254
rect 137786 606698 138022 606934
rect 137786 571018 138022 571254
rect 137786 570698 138022 570934
rect 137786 535018 138022 535254
rect 137786 534698 138022 534934
rect 137786 499018 138022 499254
rect 137786 498698 138022 498934
rect 137786 463018 138022 463254
rect 137786 462698 138022 462934
rect 137786 427018 138022 427254
rect 137786 426698 138022 426934
rect 137786 391018 138022 391254
rect 137786 390698 138022 390934
rect 137786 355018 138022 355254
rect 137786 354698 138022 354934
rect 137786 319018 138022 319254
rect 137786 318698 138022 318934
rect 137786 283018 138022 283254
rect 137786 282698 138022 282934
rect 137786 247018 138022 247254
rect 137786 246698 138022 246934
rect 137786 211018 138022 211254
rect 137786 210698 138022 210934
rect 137786 175018 138022 175254
rect 137786 174698 138022 174934
rect 137786 139018 138022 139254
rect 137786 138698 138022 138934
rect 137786 103018 138022 103254
rect 137786 102698 138022 102934
rect 137786 67018 138022 67254
rect 137786 66698 138022 66934
rect 137786 31018 138022 31254
rect 137786 30698 138022 30934
rect 119786 -6102 120022 -5866
rect 119786 -6422 120022 -6186
rect 144986 704602 145222 704838
rect 144986 704282 145222 704518
rect 144986 686218 145222 686454
rect 144986 685898 145222 686134
rect 144986 650218 145222 650454
rect 144986 649898 145222 650134
rect 144986 614218 145222 614454
rect 144986 613898 145222 614134
rect 144986 578218 145222 578454
rect 144986 577898 145222 578134
rect 144986 542218 145222 542454
rect 144986 541898 145222 542134
rect 144986 506218 145222 506454
rect 144986 505898 145222 506134
rect 144986 470218 145222 470454
rect 144986 469898 145222 470134
rect 144986 434218 145222 434454
rect 144986 433898 145222 434134
rect 144986 398218 145222 398454
rect 144986 397898 145222 398134
rect 144986 362218 145222 362454
rect 144986 361898 145222 362134
rect 144986 326218 145222 326454
rect 144986 325898 145222 326134
rect 144986 290218 145222 290454
rect 144986 289898 145222 290134
rect 144986 254218 145222 254454
rect 144986 253898 145222 254134
rect 144986 218218 145222 218454
rect 144986 217898 145222 218134
rect 144986 182218 145222 182454
rect 144986 181898 145222 182134
rect 144986 146218 145222 146454
rect 144986 145898 145222 146134
rect 144986 110218 145222 110454
rect 144986 109898 145222 110134
rect 144986 74218 145222 74454
rect 144986 73898 145222 74134
rect 144986 38218 145222 38454
rect 144986 37898 145222 38134
rect 144986 2218 145222 2454
rect 144986 1898 145222 2134
rect 144986 -582 145222 -346
rect 144986 -902 145222 -666
rect 148586 689818 148822 690054
rect 148586 689498 148822 689734
rect 148586 653818 148822 654054
rect 148586 653498 148822 653734
rect 148586 617818 148822 618054
rect 148586 617498 148822 617734
rect 148586 581818 148822 582054
rect 148586 581498 148822 581734
rect 148586 545818 148822 546054
rect 148586 545498 148822 545734
rect 148586 509818 148822 510054
rect 148586 509498 148822 509734
rect 148586 473818 148822 474054
rect 148586 473498 148822 473734
rect 148586 437818 148822 438054
rect 148586 437498 148822 437734
rect 148586 401818 148822 402054
rect 148586 401498 148822 401734
rect 148586 365818 148822 366054
rect 148586 365498 148822 365734
rect 148586 329818 148822 330054
rect 148586 329498 148822 329734
rect 148586 293818 148822 294054
rect 148586 293498 148822 293734
rect 148586 257818 148822 258054
rect 148586 257498 148822 257734
rect 148586 221818 148822 222054
rect 148586 221498 148822 221734
rect 148586 185818 148822 186054
rect 148586 185498 148822 185734
rect 148586 149818 148822 150054
rect 148586 149498 148822 149734
rect 148586 113818 148822 114054
rect 148586 113498 148822 113734
rect 148586 77818 148822 78054
rect 148586 77498 148822 77734
rect 148586 41818 148822 42054
rect 148586 41498 148822 41734
rect 148586 5818 148822 6054
rect 148586 5498 148822 5734
rect 148586 -2422 148822 -2186
rect 148586 -2742 148822 -2506
rect 152186 693418 152422 693654
rect 152186 693098 152422 693334
rect 152186 657418 152422 657654
rect 152186 657098 152422 657334
rect 152186 621418 152422 621654
rect 152186 621098 152422 621334
rect 152186 585418 152422 585654
rect 152186 585098 152422 585334
rect 152186 549418 152422 549654
rect 152186 549098 152422 549334
rect 152186 513418 152422 513654
rect 152186 513098 152422 513334
rect 152186 477418 152422 477654
rect 152186 477098 152422 477334
rect 152186 441418 152422 441654
rect 152186 441098 152422 441334
rect 152186 405418 152422 405654
rect 152186 405098 152422 405334
rect 152186 369418 152422 369654
rect 152186 369098 152422 369334
rect 152186 333418 152422 333654
rect 152186 333098 152422 333334
rect 152186 297418 152422 297654
rect 152186 297098 152422 297334
rect 152186 261418 152422 261654
rect 152186 261098 152422 261334
rect 152186 225418 152422 225654
rect 152186 225098 152422 225334
rect 152186 189418 152422 189654
rect 152186 189098 152422 189334
rect 152186 153418 152422 153654
rect 152186 153098 152422 153334
rect 152186 117418 152422 117654
rect 152186 117098 152422 117334
rect 152186 81418 152422 81654
rect 152186 81098 152422 81334
rect 152186 45418 152422 45654
rect 152186 45098 152422 45334
rect 152186 9418 152422 9654
rect 152186 9098 152422 9334
rect 152186 -4262 152422 -4026
rect 152186 -4582 152422 -4346
rect 173786 711042 174022 711278
rect 173786 710722 174022 710958
rect 170186 709202 170422 709438
rect 170186 708882 170422 709118
rect 166586 707362 166822 707598
rect 166586 707042 166822 707278
rect 155786 697018 156022 697254
rect 155786 696698 156022 696934
rect 155786 661018 156022 661254
rect 155786 660698 156022 660934
rect 155786 625018 156022 625254
rect 155786 624698 156022 624934
rect 155786 589018 156022 589254
rect 155786 588698 156022 588934
rect 155786 553018 156022 553254
rect 155786 552698 156022 552934
rect 155786 517018 156022 517254
rect 155786 516698 156022 516934
rect 155786 481018 156022 481254
rect 155786 480698 156022 480934
rect 155786 445018 156022 445254
rect 155786 444698 156022 444934
rect 155786 409018 156022 409254
rect 155786 408698 156022 408934
rect 155786 373018 156022 373254
rect 155786 372698 156022 372934
rect 155786 337018 156022 337254
rect 155786 336698 156022 336934
rect 155786 301018 156022 301254
rect 155786 300698 156022 300934
rect 155786 265018 156022 265254
rect 155786 264698 156022 264934
rect 155786 229018 156022 229254
rect 155786 228698 156022 228934
rect 155786 193018 156022 193254
rect 155786 192698 156022 192934
rect 155786 157018 156022 157254
rect 155786 156698 156022 156934
rect 155786 121018 156022 121254
rect 155786 120698 156022 120934
rect 155786 85018 156022 85254
rect 155786 84698 156022 84934
rect 155786 49018 156022 49254
rect 155786 48698 156022 48934
rect 155786 13018 156022 13254
rect 155786 12698 156022 12934
rect 137786 -7022 138022 -6786
rect 137786 -7342 138022 -7106
rect 162986 705522 163222 705758
rect 162986 705202 163222 705438
rect 162986 668218 163222 668454
rect 162986 667898 163222 668134
rect 162986 632218 163222 632454
rect 162986 631898 163222 632134
rect 162986 596218 163222 596454
rect 162986 595898 163222 596134
rect 162986 560218 163222 560454
rect 162986 559898 163222 560134
rect 162986 524218 163222 524454
rect 162986 523898 163222 524134
rect 162986 488218 163222 488454
rect 162986 487898 163222 488134
rect 162986 452218 163222 452454
rect 162986 451898 163222 452134
rect 162986 416218 163222 416454
rect 162986 415898 163222 416134
rect 162986 380218 163222 380454
rect 162986 379898 163222 380134
rect 162986 344218 163222 344454
rect 162986 343898 163222 344134
rect 162986 308218 163222 308454
rect 162986 307898 163222 308134
rect 162986 272218 163222 272454
rect 162986 271898 163222 272134
rect 162986 236218 163222 236454
rect 162986 235898 163222 236134
rect 162986 200218 163222 200454
rect 162986 199898 163222 200134
rect 162986 164218 163222 164454
rect 162986 163898 163222 164134
rect 162986 128218 163222 128454
rect 162986 127898 163222 128134
rect 162986 92218 163222 92454
rect 162986 91898 163222 92134
rect 162986 56218 163222 56454
rect 162986 55898 163222 56134
rect 162986 20218 163222 20454
rect 162986 19898 163222 20134
rect 162986 -1502 163222 -1266
rect 162986 -1822 163222 -1586
rect 166586 671818 166822 672054
rect 166586 671498 166822 671734
rect 166586 635818 166822 636054
rect 166586 635498 166822 635734
rect 166586 599818 166822 600054
rect 166586 599498 166822 599734
rect 166586 563818 166822 564054
rect 166586 563498 166822 563734
rect 166586 527818 166822 528054
rect 166586 527498 166822 527734
rect 166586 491818 166822 492054
rect 166586 491498 166822 491734
rect 166586 455818 166822 456054
rect 166586 455498 166822 455734
rect 166586 419818 166822 420054
rect 166586 419498 166822 419734
rect 166586 383818 166822 384054
rect 166586 383498 166822 383734
rect 166586 347818 166822 348054
rect 166586 347498 166822 347734
rect 166586 311818 166822 312054
rect 166586 311498 166822 311734
rect 166586 275818 166822 276054
rect 166586 275498 166822 275734
rect 166586 239818 166822 240054
rect 166586 239498 166822 239734
rect 166586 203818 166822 204054
rect 166586 203498 166822 203734
rect 166586 167818 166822 168054
rect 166586 167498 166822 167734
rect 166586 131818 166822 132054
rect 166586 131498 166822 131734
rect 166586 95818 166822 96054
rect 166586 95498 166822 95734
rect 166586 59818 166822 60054
rect 166586 59498 166822 59734
rect 166586 23818 166822 24054
rect 166586 23498 166822 23734
rect 166586 -3342 166822 -3106
rect 166586 -3662 166822 -3426
rect 170186 675418 170422 675654
rect 170186 675098 170422 675334
rect 170186 639418 170422 639654
rect 170186 639098 170422 639334
rect 170186 603418 170422 603654
rect 170186 603098 170422 603334
rect 170186 567418 170422 567654
rect 170186 567098 170422 567334
rect 170186 531418 170422 531654
rect 170186 531098 170422 531334
rect 170186 495418 170422 495654
rect 170186 495098 170422 495334
rect 170186 459418 170422 459654
rect 170186 459098 170422 459334
rect 170186 423418 170422 423654
rect 170186 423098 170422 423334
rect 170186 387418 170422 387654
rect 170186 387098 170422 387334
rect 170186 351418 170422 351654
rect 170186 351098 170422 351334
rect 170186 315418 170422 315654
rect 170186 315098 170422 315334
rect 170186 279418 170422 279654
rect 170186 279098 170422 279334
rect 170186 243418 170422 243654
rect 170186 243098 170422 243334
rect 170186 207418 170422 207654
rect 170186 207098 170422 207334
rect 170186 171418 170422 171654
rect 170186 171098 170422 171334
rect 170186 135418 170422 135654
rect 170186 135098 170422 135334
rect 170186 99418 170422 99654
rect 170186 99098 170422 99334
rect 170186 63418 170422 63654
rect 170186 63098 170422 63334
rect 170186 27418 170422 27654
rect 170186 27098 170422 27334
rect 170186 -5182 170422 -4946
rect 170186 -5502 170422 -5266
rect 191786 710122 192022 710358
rect 191786 709802 192022 710038
rect 188186 708282 188422 708518
rect 188186 707962 188422 708198
rect 184586 706442 184822 706678
rect 184586 706122 184822 706358
rect 173786 679018 174022 679254
rect 173786 678698 174022 678934
rect 173786 643018 174022 643254
rect 173786 642698 174022 642934
rect 173786 607018 174022 607254
rect 173786 606698 174022 606934
rect 173786 571018 174022 571254
rect 173786 570698 174022 570934
rect 173786 535018 174022 535254
rect 173786 534698 174022 534934
rect 173786 499018 174022 499254
rect 173786 498698 174022 498934
rect 173786 463018 174022 463254
rect 173786 462698 174022 462934
rect 173786 427018 174022 427254
rect 173786 426698 174022 426934
rect 173786 391018 174022 391254
rect 173786 390698 174022 390934
rect 173786 355018 174022 355254
rect 173786 354698 174022 354934
rect 173786 319018 174022 319254
rect 173786 318698 174022 318934
rect 173786 283018 174022 283254
rect 173786 282698 174022 282934
rect 173786 247018 174022 247254
rect 173786 246698 174022 246934
rect 173786 211018 174022 211254
rect 173786 210698 174022 210934
rect 173786 175018 174022 175254
rect 173786 174698 174022 174934
rect 173786 139018 174022 139254
rect 173786 138698 174022 138934
rect 173786 103018 174022 103254
rect 173786 102698 174022 102934
rect 173786 67018 174022 67254
rect 173786 66698 174022 66934
rect 173786 31018 174022 31254
rect 173786 30698 174022 30934
rect 155786 -6102 156022 -5866
rect 155786 -6422 156022 -6186
rect 180986 704602 181222 704838
rect 180986 704282 181222 704518
rect 180986 686218 181222 686454
rect 180986 685898 181222 686134
rect 180986 650218 181222 650454
rect 180986 649898 181222 650134
rect 180986 614218 181222 614454
rect 180986 613898 181222 614134
rect 180986 578218 181222 578454
rect 180986 577898 181222 578134
rect 180986 542218 181222 542454
rect 180986 541898 181222 542134
rect 180986 506218 181222 506454
rect 180986 505898 181222 506134
rect 180986 470218 181222 470454
rect 180986 469898 181222 470134
rect 180986 434218 181222 434454
rect 180986 433898 181222 434134
rect 180986 398218 181222 398454
rect 180986 397898 181222 398134
rect 180986 362218 181222 362454
rect 180986 361898 181222 362134
rect 180986 326218 181222 326454
rect 180986 325898 181222 326134
rect 180986 290218 181222 290454
rect 180986 289898 181222 290134
rect 180986 254218 181222 254454
rect 180986 253898 181222 254134
rect 180986 218218 181222 218454
rect 180986 217898 181222 218134
rect 180986 182218 181222 182454
rect 180986 181898 181222 182134
rect 180986 146218 181222 146454
rect 180986 145898 181222 146134
rect 180986 110218 181222 110454
rect 180986 109898 181222 110134
rect 180986 74218 181222 74454
rect 180986 73898 181222 74134
rect 180986 38218 181222 38454
rect 180986 37898 181222 38134
rect 180986 2218 181222 2454
rect 180986 1898 181222 2134
rect 180986 -582 181222 -346
rect 180986 -902 181222 -666
rect 184586 689818 184822 690054
rect 184586 689498 184822 689734
rect 184586 653818 184822 654054
rect 184586 653498 184822 653734
rect 184586 617818 184822 618054
rect 184586 617498 184822 617734
rect 184586 581818 184822 582054
rect 184586 581498 184822 581734
rect 184586 545818 184822 546054
rect 184586 545498 184822 545734
rect 184586 509818 184822 510054
rect 184586 509498 184822 509734
rect 184586 473818 184822 474054
rect 184586 473498 184822 473734
rect 184586 437818 184822 438054
rect 184586 437498 184822 437734
rect 184586 401818 184822 402054
rect 184586 401498 184822 401734
rect 184586 365818 184822 366054
rect 184586 365498 184822 365734
rect 184586 329818 184822 330054
rect 184586 329498 184822 329734
rect 184586 293818 184822 294054
rect 184586 293498 184822 293734
rect 184586 257818 184822 258054
rect 184586 257498 184822 257734
rect 184586 221818 184822 222054
rect 184586 221498 184822 221734
rect 184586 185818 184822 186054
rect 184586 185498 184822 185734
rect 184586 149818 184822 150054
rect 184586 149498 184822 149734
rect 184586 113818 184822 114054
rect 184586 113498 184822 113734
rect 184586 77818 184822 78054
rect 184586 77498 184822 77734
rect 184586 41818 184822 42054
rect 184586 41498 184822 41734
rect 184586 5818 184822 6054
rect 184586 5498 184822 5734
rect 184586 -2422 184822 -2186
rect 184586 -2742 184822 -2506
rect 188186 693418 188422 693654
rect 188186 693098 188422 693334
rect 188186 657418 188422 657654
rect 188186 657098 188422 657334
rect 188186 621418 188422 621654
rect 188186 621098 188422 621334
rect 188186 585418 188422 585654
rect 188186 585098 188422 585334
rect 188186 549418 188422 549654
rect 188186 549098 188422 549334
rect 188186 513418 188422 513654
rect 188186 513098 188422 513334
rect 188186 477418 188422 477654
rect 188186 477098 188422 477334
rect 188186 441418 188422 441654
rect 188186 441098 188422 441334
rect 188186 405418 188422 405654
rect 188186 405098 188422 405334
rect 188186 369418 188422 369654
rect 188186 369098 188422 369334
rect 188186 333418 188422 333654
rect 188186 333098 188422 333334
rect 188186 297418 188422 297654
rect 188186 297098 188422 297334
rect 188186 261418 188422 261654
rect 188186 261098 188422 261334
rect 188186 225418 188422 225654
rect 188186 225098 188422 225334
rect 188186 189418 188422 189654
rect 188186 189098 188422 189334
rect 188186 153418 188422 153654
rect 188186 153098 188422 153334
rect 188186 117418 188422 117654
rect 188186 117098 188422 117334
rect 188186 81418 188422 81654
rect 188186 81098 188422 81334
rect 188186 45418 188422 45654
rect 188186 45098 188422 45334
rect 188186 9418 188422 9654
rect 188186 9098 188422 9334
rect 188186 -4262 188422 -4026
rect 188186 -4582 188422 -4346
rect 209786 711042 210022 711278
rect 209786 710722 210022 710958
rect 206186 709202 206422 709438
rect 206186 708882 206422 709118
rect 202586 707362 202822 707598
rect 202586 707042 202822 707278
rect 191786 697018 192022 697254
rect 191786 696698 192022 696934
rect 191786 661018 192022 661254
rect 191786 660698 192022 660934
rect 191786 625018 192022 625254
rect 191786 624698 192022 624934
rect 191786 589018 192022 589254
rect 191786 588698 192022 588934
rect 191786 553018 192022 553254
rect 191786 552698 192022 552934
rect 191786 517018 192022 517254
rect 191786 516698 192022 516934
rect 191786 481018 192022 481254
rect 191786 480698 192022 480934
rect 191786 445018 192022 445254
rect 191786 444698 192022 444934
rect 191786 409018 192022 409254
rect 191786 408698 192022 408934
rect 191786 373018 192022 373254
rect 191786 372698 192022 372934
rect 191786 337018 192022 337254
rect 191786 336698 192022 336934
rect 191786 301018 192022 301254
rect 191786 300698 192022 300934
rect 191786 265018 192022 265254
rect 191786 264698 192022 264934
rect 191786 229018 192022 229254
rect 191786 228698 192022 228934
rect 191786 193018 192022 193254
rect 191786 192698 192022 192934
rect 191786 157018 192022 157254
rect 191786 156698 192022 156934
rect 191786 121018 192022 121254
rect 191786 120698 192022 120934
rect 191786 85018 192022 85254
rect 191786 84698 192022 84934
rect 191786 49018 192022 49254
rect 191786 48698 192022 48934
rect 191786 13018 192022 13254
rect 191786 12698 192022 12934
rect 173786 -7022 174022 -6786
rect 173786 -7342 174022 -7106
rect 198986 705522 199222 705758
rect 198986 705202 199222 705438
rect 198986 668218 199222 668454
rect 198986 667898 199222 668134
rect 198986 632218 199222 632454
rect 198986 631898 199222 632134
rect 198986 596218 199222 596454
rect 198986 595898 199222 596134
rect 198986 560218 199222 560454
rect 198986 559898 199222 560134
rect 198986 524218 199222 524454
rect 198986 523898 199222 524134
rect 198986 488218 199222 488454
rect 198986 487898 199222 488134
rect 198986 452218 199222 452454
rect 198986 451898 199222 452134
rect 198986 416218 199222 416454
rect 198986 415898 199222 416134
rect 198986 380218 199222 380454
rect 198986 379898 199222 380134
rect 198986 344218 199222 344454
rect 198986 343898 199222 344134
rect 198986 308218 199222 308454
rect 198986 307898 199222 308134
rect 198986 272218 199222 272454
rect 198986 271898 199222 272134
rect 198986 236218 199222 236454
rect 198986 235898 199222 236134
rect 198986 200218 199222 200454
rect 198986 199898 199222 200134
rect 198986 164218 199222 164454
rect 198986 163898 199222 164134
rect 198986 128218 199222 128454
rect 198986 127898 199222 128134
rect 198986 92218 199222 92454
rect 198986 91898 199222 92134
rect 198986 56218 199222 56454
rect 198986 55898 199222 56134
rect 198986 20218 199222 20454
rect 198986 19898 199222 20134
rect 198986 -1502 199222 -1266
rect 198986 -1822 199222 -1586
rect 202586 671818 202822 672054
rect 202586 671498 202822 671734
rect 202586 635818 202822 636054
rect 202586 635498 202822 635734
rect 202586 599818 202822 600054
rect 202586 599498 202822 599734
rect 202586 563818 202822 564054
rect 202586 563498 202822 563734
rect 202586 527818 202822 528054
rect 202586 527498 202822 527734
rect 202586 491818 202822 492054
rect 202586 491498 202822 491734
rect 202586 455818 202822 456054
rect 202586 455498 202822 455734
rect 202586 419818 202822 420054
rect 202586 419498 202822 419734
rect 202586 383818 202822 384054
rect 202586 383498 202822 383734
rect 202586 347818 202822 348054
rect 202586 347498 202822 347734
rect 202586 311818 202822 312054
rect 202586 311498 202822 311734
rect 202586 275818 202822 276054
rect 202586 275498 202822 275734
rect 202586 239818 202822 240054
rect 202586 239498 202822 239734
rect 202586 203818 202822 204054
rect 202586 203498 202822 203734
rect 202586 167818 202822 168054
rect 202586 167498 202822 167734
rect 202586 131818 202822 132054
rect 202586 131498 202822 131734
rect 202586 95818 202822 96054
rect 202586 95498 202822 95734
rect 202586 59818 202822 60054
rect 202586 59498 202822 59734
rect 202586 23818 202822 24054
rect 202586 23498 202822 23734
rect 202586 -3342 202822 -3106
rect 202586 -3662 202822 -3426
rect 206186 675418 206422 675654
rect 206186 675098 206422 675334
rect 206186 639418 206422 639654
rect 206186 639098 206422 639334
rect 206186 603418 206422 603654
rect 206186 603098 206422 603334
rect 206186 567418 206422 567654
rect 206186 567098 206422 567334
rect 206186 531418 206422 531654
rect 206186 531098 206422 531334
rect 206186 495418 206422 495654
rect 206186 495098 206422 495334
rect 206186 459418 206422 459654
rect 206186 459098 206422 459334
rect 206186 423418 206422 423654
rect 206186 423098 206422 423334
rect 206186 387418 206422 387654
rect 206186 387098 206422 387334
rect 206186 351418 206422 351654
rect 206186 351098 206422 351334
rect 206186 315418 206422 315654
rect 206186 315098 206422 315334
rect 206186 279418 206422 279654
rect 206186 279098 206422 279334
rect 206186 243418 206422 243654
rect 206186 243098 206422 243334
rect 206186 207418 206422 207654
rect 206186 207098 206422 207334
rect 206186 171418 206422 171654
rect 206186 171098 206422 171334
rect 206186 135418 206422 135654
rect 206186 135098 206422 135334
rect 206186 99418 206422 99654
rect 206186 99098 206422 99334
rect 206186 63418 206422 63654
rect 206186 63098 206422 63334
rect 206186 27418 206422 27654
rect 206186 27098 206422 27334
rect 206186 -5182 206422 -4946
rect 206186 -5502 206422 -5266
rect 227786 710122 228022 710358
rect 227786 709802 228022 710038
rect 224186 708282 224422 708518
rect 224186 707962 224422 708198
rect 220586 706442 220822 706678
rect 220586 706122 220822 706358
rect 209786 679018 210022 679254
rect 209786 678698 210022 678934
rect 209786 643018 210022 643254
rect 209786 642698 210022 642934
rect 209786 607018 210022 607254
rect 209786 606698 210022 606934
rect 209786 571018 210022 571254
rect 209786 570698 210022 570934
rect 209786 535018 210022 535254
rect 209786 534698 210022 534934
rect 209786 499018 210022 499254
rect 209786 498698 210022 498934
rect 209786 463018 210022 463254
rect 209786 462698 210022 462934
rect 209786 427018 210022 427254
rect 209786 426698 210022 426934
rect 209786 391018 210022 391254
rect 209786 390698 210022 390934
rect 209786 355018 210022 355254
rect 209786 354698 210022 354934
rect 209786 319018 210022 319254
rect 209786 318698 210022 318934
rect 209786 283018 210022 283254
rect 209786 282698 210022 282934
rect 209786 247018 210022 247254
rect 209786 246698 210022 246934
rect 209786 211018 210022 211254
rect 209786 210698 210022 210934
rect 209786 175018 210022 175254
rect 209786 174698 210022 174934
rect 209786 139018 210022 139254
rect 209786 138698 210022 138934
rect 209786 103018 210022 103254
rect 209786 102698 210022 102934
rect 209786 67018 210022 67254
rect 209786 66698 210022 66934
rect 209786 31018 210022 31254
rect 209786 30698 210022 30934
rect 191786 -6102 192022 -5866
rect 191786 -6422 192022 -6186
rect 216986 704602 217222 704838
rect 216986 704282 217222 704518
rect 216986 686218 217222 686454
rect 216986 685898 217222 686134
rect 216986 650218 217222 650454
rect 216986 649898 217222 650134
rect 216986 614218 217222 614454
rect 216986 613898 217222 614134
rect 216986 578218 217222 578454
rect 216986 577898 217222 578134
rect 216986 542218 217222 542454
rect 216986 541898 217222 542134
rect 216986 506218 217222 506454
rect 216986 505898 217222 506134
rect 216986 470218 217222 470454
rect 216986 469898 217222 470134
rect 216986 434218 217222 434454
rect 216986 433898 217222 434134
rect 216986 398218 217222 398454
rect 216986 397898 217222 398134
rect 216986 362218 217222 362454
rect 216986 361898 217222 362134
rect 216986 326218 217222 326454
rect 216986 325898 217222 326134
rect 216986 290218 217222 290454
rect 216986 289898 217222 290134
rect 216986 254218 217222 254454
rect 216986 253898 217222 254134
rect 216986 218218 217222 218454
rect 216986 217898 217222 218134
rect 216986 182218 217222 182454
rect 216986 181898 217222 182134
rect 216986 146218 217222 146454
rect 216986 145898 217222 146134
rect 216986 110218 217222 110454
rect 216986 109898 217222 110134
rect 216986 74218 217222 74454
rect 216986 73898 217222 74134
rect 216986 38218 217222 38454
rect 216986 37898 217222 38134
rect 216986 2218 217222 2454
rect 216986 1898 217222 2134
rect 216986 -582 217222 -346
rect 216986 -902 217222 -666
rect 220586 689818 220822 690054
rect 220586 689498 220822 689734
rect 220586 653818 220822 654054
rect 220586 653498 220822 653734
rect 220586 617818 220822 618054
rect 220586 617498 220822 617734
rect 220586 581818 220822 582054
rect 220586 581498 220822 581734
rect 220586 545818 220822 546054
rect 220586 545498 220822 545734
rect 220586 509818 220822 510054
rect 220586 509498 220822 509734
rect 220586 473818 220822 474054
rect 220586 473498 220822 473734
rect 220586 437818 220822 438054
rect 220586 437498 220822 437734
rect 220586 401818 220822 402054
rect 220586 401498 220822 401734
rect 220586 365818 220822 366054
rect 220586 365498 220822 365734
rect 220586 329818 220822 330054
rect 220586 329498 220822 329734
rect 220586 293818 220822 294054
rect 220586 293498 220822 293734
rect 220586 257818 220822 258054
rect 220586 257498 220822 257734
rect 220586 221818 220822 222054
rect 220586 221498 220822 221734
rect 220586 185818 220822 186054
rect 220586 185498 220822 185734
rect 220586 149818 220822 150054
rect 220586 149498 220822 149734
rect 220586 113818 220822 114054
rect 220586 113498 220822 113734
rect 220586 77818 220822 78054
rect 220586 77498 220822 77734
rect 220586 41818 220822 42054
rect 220586 41498 220822 41734
rect 220586 5818 220822 6054
rect 220586 5498 220822 5734
rect 220586 -2422 220822 -2186
rect 220586 -2742 220822 -2506
rect 224186 693418 224422 693654
rect 224186 693098 224422 693334
rect 224186 657418 224422 657654
rect 224186 657098 224422 657334
rect 224186 621418 224422 621654
rect 224186 621098 224422 621334
rect 224186 585418 224422 585654
rect 224186 585098 224422 585334
rect 224186 549418 224422 549654
rect 224186 549098 224422 549334
rect 224186 513418 224422 513654
rect 224186 513098 224422 513334
rect 224186 477418 224422 477654
rect 224186 477098 224422 477334
rect 224186 441418 224422 441654
rect 224186 441098 224422 441334
rect 224186 405418 224422 405654
rect 224186 405098 224422 405334
rect 224186 369418 224422 369654
rect 224186 369098 224422 369334
rect 224186 333418 224422 333654
rect 224186 333098 224422 333334
rect 224186 297418 224422 297654
rect 224186 297098 224422 297334
rect 224186 261418 224422 261654
rect 224186 261098 224422 261334
rect 224186 225418 224422 225654
rect 224186 225098 224422 225334
rect 224186 189418 224422 189654
rect 224186 189098 224422 189334
rect 224186 153418 224422 153654
rect 224186 153098 224422 153334
rect 224186 117418 224422 117654
rect 224186 117098 224422 117334
rect 224186 81418 224422 81654
rect 224186 81098 224422 81334
rect 224186 45418 224422 45654
rect 224186 45098 224422 45334
rect 224186 9418 224422 9654
rect 224186 9098 224422 9334
rect 224186 -4262 224422 -4026
rect 224186 -4582 224422 -4346
rect 245786 711042 246022 711278
rect 245786 710722 246022 710958
rect 242186 709202 242422 709438
rect 242186 708882 242422 709118
rect 238586 707362 238822 707598
rect 238586 707042 238822 707278
rect 227786 697018 228022 697254
rect 227786 696698 228022 696934
rect 227786 661018 228022 661254
rect 227786 660698 228022 660934
rect 227786 625018 228022 625254
rect 227786 624698 228022 624934
rect 227786 589018 228022 589254
rect 227786 588698 228022 588934
rect 227786 553018 228022 553254
rect 227786 552698 228022 552934
rect 227786 517018 228022 517254
rect 227786 516698 228022 516934
rect 227786 481018 228022 481254
rect 227786 480698 228022 480934
rect 227786 445018 228022 445254
rect 227786 444698 228022 444934
rect 227786 409018 228022 409254
rect 227786 408698 228022 408934
rect 234986 705522 235222 705758
rect 234986 705202 235222 705438
rect 234986 668218 235222 668454
rect 234986 667898 235222 668134
rect 234986 632218 235222 632454
rect 234986 631898 235222 632134
rect 234986 596218 235222 596454
rect 234986 595898 235222 596134
rect 234986 560218 235222 560454
rect 234986 559898 235222 560134
rect 234986 524218 235222 524454
rect 234986 523898 235222 524134
rect 234986 488218 235222 488454
rect 234986 487898 235222 488134
rect 234986 452218 235222 452454
rect 234986 451898 235222 452134
rect 234986 416218 235222 416454
rect 234986 415898 235222 416134
rect 227786 373018 228022 373254
rect 227786 372698 228022 372934
rect 227786 337018 228022 337254
rect 227786 336698 228022 336934
rect 227786 301018 228022 301254
rect 227786 300698 228022 300934
rect 227786 265018 228022 265254
rect 227786 264698 228022 264934
rect 227786 229018 228022 229254
rect 227786 228698 228022 228934
rect 227786 193018 228022 193254
rect 227786 192698 228022 192934
rect 227786 157018 228022 157254
rect 227786 156698 228022 156934
rect 227786 121018 228022 121254
rect 227786 120698 228022 120934
rect 227786 85018 228022 85254
rect 227786 84698 228022 84934
rect 227786 49018 228022 49254
rect 227786 48698 228022 48934
rect 238586 671818 238822 672054
rect 238586 671498 238822 671734
rect 238586 635818 238822 636054
rect 238586 635498 238822 635734
rect 238586 599818 238822 600054
rect 238586 599498 238822 599734
rect 238586 563818 238822 564054
rect 238586 563498 238822 563734
rect 238586 527818 238822 528054
rect 238586 527498 238822 527734
rect 238586 491818 238822 492054
rect 238586 491498 238822 491734
rect 238586 455818 238822 456054
rect 238586 455498 238822 455734
rect 238586 419818 238822 420054
rect 238586 419498 238822 419734
rect 234986 380218 235222 380454
rect 234986 379898 235222 380134
rect 234986 344218 235222 344454
rect 234986 343898 235222 344134
rect 234986 308218 235222 308454
rect 234986 307898 235222 308134
rect 234986 272218 235222 272454
rect 234986 271898 235222 272134
rect 234986 236218 235222 236454
rect 234986 235898 235222 236134
rect 238586 383818 238822 384054
rect 238586 383498 238822 383734
rect 238586 347818 238822 348054
rect 238586 347498 238822 347734
rect 238586 311818 238822 312054
rect 238586 311498 238822 311734
rect 238586 275818 238822 276054
rect 238586 275498 238822 275734
rect 238586 239818 238822 240054
rect 238586 239498 238822 239734
rect 234986 200218 235222 200454
rect 234986 199898 235222 200134
rect 234986 164218 235222 164454
rect 234986 163898 235222 164134
rect 234986 128218 235222 128454
rect 234986 127898 235222 128134
rect 234986 92218 235222 92454
rect 234986 91898 235222 92134
rect 234986 56218 235222 56454
rect 234986 55898 235222 56134
rect 227786 13018 228022 13254
rect 227786 12698 228022 12934
rect 209786 -7022 210022 -6786
rect 209786 -7342 210022 -7106
rect 234986 20218 235222 20454
rect 234986 19898 235222 20134
rect 234986 -1502 235222 -1266
rect 234986 -1822 235222 -1586
rect 238586 203818 238822 204054
rect 238586 203498 238822 203734
rect 238586 167818 238822 168054
rect 238586 167498 238822 167734
rect 238586 131818 238822 132054
rect 238586 131498 238822 131734
rect 238586 95818 238822 96054
rect 238586 95498 238822 95734
rect 238586 59818 238822 60054
rect 238586 59498 238822 59734
rect 238586 23818 238822 24054
rect 238586 23498 238822 23734
rect 238586 -3342 238822 -3106
rect 238586 -3662 238822 -3426
rect 242186 675418 242422 675654
rect 242186 675098 242422 675334
rect 242186 639418 242422 639654
rect 242186 639098 242422 639334
rect 242186 603418 242422 603654
rect 242186 603098 242422 603334
rect 242186 567418 242422 567654
rect 242186 567098 242422 567334
rect 242186 531418 242422 531654
rect 242186 531098 242422 531334
rect 242186 495418 242422 495654
rect 242186 495098 242422 495334
rect 242186 459418 242422 459654
rect 242186 459098 242422 459334
rect 242186 423418 242422 423654
rect 242186 423098 242422 423334
rect 263786 710122 264022 710358
rect 263786 709802 264022 710038
rect 260186 708282 260422 708518
rect 260186 707962 260422 708198
rect 256586 706442 256822 706678
rect 256586 706122 256822 706358
rect 245786 679018 246022 679254
rect 245786 678698 246022 678934
rect 245786 643018 246022 643254
rect 245786 642698 246022 642934
rect 245786 607018 246022 607254
rect 245786 606698 246022 606934
rect 245786 571018 246022 571254
rect 245786 570698 246022 570934
rect 245786 535018 246022 535254
rect 245786 534698 246022 534934
rect 245786 499018 246022 499254
rect 245786 498698 246022 498934
rect 245786 463018 246022 463254
rect 245786 462698 246022 462934
rect 245786 427018 246022 427254
rect 245786 426698 246022 426934
rect 242186 387418 242422 387654
rect 242186 387098 242422 387334
rect 242186 351418 242422 351654
rect 242186 351098 242422 351334
rect 242186 315418 242422 315654
rect 242186 315098 242422 315334
rect 242186 279418 242422 279654
rect 242186 279098 242422 279334
rect 242186 243418 242422 243654
rect 242186 243098 242422 243334
rect 242186 207418 242422 207654
rect 242186 207098 242422 207334
rect 242186 171418 242422 171654
rect 242186 171098 242422 171334
rect 242186 135418 242422 135654
rect 242186 135098 242422 135334
rect 242186 99418 242422 99654
rect 242186 99098 242422 99334
rect 242186 63418 242422 63654
rect 242186 63098 242422 63334
rect 242186 27418 242422 27654
rect 242186 27098 242422 27334
rect 242186 -5182 242422 -4946
rect 242186 -5502 242422 -5266
rect 245786 391018 246022 391254
rect 245786 390698 246022 390934
rect 245786 355018 246022 355254
rect 245786 354698 246022 354934
rect 245786 319018 246022 319254
rect 245786 318698 246022 318934
rect 245786 283018 246022 283254
rect 245786 282698 246022 282934
rect 245786 247018 246022 247254
rect 245786 246698 246022 246934
rect 245786 211018 246022 211254
rect 245786 210698 246022 210934
rect 245786 175018 246022 175254
rect 245786 174698 246022 174934
rect 245786 139018 246022 139254
rect 245786 138698 246022 138934
rect 245786 103018 246022 103254
rect 245786 102698 246022 102934
rect 245786 67018 246022 67254
rect 245786 66698 246022 66934
rect 245786 31018 246022 31254
rect 245786 30698 246022 30934
rect 227786 -6102 228022 -5866
rect 227786 -6422 228022 -6186
rect 252986 704602 253222 704838
rect 252986 704282 253222 704518
rect 252986 686218 253222 686454
rect 252986 685898 253222 686134
rect 252986 650218 253222 650454
rect 252986 649898 253222 650134
rect 252986 614218 253222 614454
rect 252986 613898 253222 614134
rect 252986 578218 253222 578454
rect 252986 577898 253222 578134
rect 252986 542218 253222 542454
rect 252986 541898 253222 542134
rect 252986 506218 253222 506454
rect 252986 505898 253222 506134
rect 252986 470218 253222 470454
rect 252986 469898 253222 470134
rect 252986 434218 253222 434454
rect 252986 433898 253222 434134
rect 252986 398218 253222 398454
rect 252986 397898 253222 398134
rect 252986 362218 253222 362454
rect 252986 361898 253222 362134
rect 252986 326218 253222 326454
rect 252986 325898 253222 326134
rect 256586 689818 256822 690054
rect 256586 689498 256822 689734
rect 256586 653818 256822 654054
rect 256586 653498 256822 653734
rect 256586 617818 256822 618054
rect 256586 617498 256822 617734
rect 256586 581818 256822 582054
rect 256586 581498 256822 581734
rect 256586 545818 256822 546054
rect 256586 545498 256822 545734
rect 256586 509818 256822 510054
rect 256586 509498 256822 509734
rect 256586 473818 256822 474054
rect 256586 473498 256822 473734
rect 256586 437818 256822 438054
rect 256586 437498 256822 437734
rect 256586 401818 256822 402054
rect 256586 401498 256822 401734
rect 256586 365818 256822 366054
rect 256586 365498 256822 365734
rect 256586 329818 256822 330054
rect 256586 329498 256822 329734
rect 252986 290218 253222 290454
rect 252986 289898 253222 290134
rect 256586 293818 256822 294054
rect 256586 293498 256822 293734
rect 252986 254218 253222 254454
rect 252986 253898 253222 254134
rect 252986 218218 253222 218454
rect 252986 217898 253222 218134
rect 252986 182218 253222 182454
rect 252986 181898 253222 182134
rect 252986 146218 253222 146454
rect 252986 145898 253222 146134
rect 252986 110218 253222 110454
rect 252986 109898 253222 110134
rect 252986 74218 253222 74454
rect 252986 73898 253222 74134
rect 252986 38218 253222 38454
rect 252986 37898 253222 38134
rect 252986 2218 253222 2454
rect 252986 1898 253222 2134
rect 252986 -582 253222 -346
rect 252986 -902 253222 -666
rect 256586 257818 256822 258054
rect 256586 257498 256822 257734
rect 256586 221818 256822 222054
rect 256586 221498 256822 221734
rect 256586 185818 256822 186054
rect 256586 185498 256822 185734
rect 256586 149818 256822 150054
rect 256586 149498 256822 149734
rect 256586 113818 256822 114054
rect 256586 113498 256822 113734
rect 256586 77818 256822 78054
rect 256586 77498 256822 77734
rect 256586 41818 256822 42054
rect 256586 41498 256822 41734
rect 256586 5818 256822 6054
rect 256586 5498 256822 5734
rect 256586 -2422 256822 -2186
rect 256586 -2742 256822 -2506
rect 260186 693418 260422 693654
rect 260186 693098 260422 693334
rect 260186 657418 260422 657654
rect 260186 657098 260422 657334
rect 260186 621418 260422 621654
rect 260186 621098 260422 621334
rect 260186 585418 260422 585654
rect 260186 585098 260422 585334
rect 260186 549418 260422 549654
rect 260186 549098 260422 549334
rect 260186 513418 260422 513654
rect 260186 513098 260422 513334
rect 260186 477418 260422 477654
rect 260186 477098 260422 477334
rect 260186 441418 260422 441654
rect 260186 441098 260422 441334
rect 260186 405418 260422 405654
rect 260186 405098 260422 405334
rect 260186 369418 260422 369654
rect 260186 369098 260422 369334
rect 260186 333418 260422 333654
rect 260186 333098 260422 333334
rect 260186 297418 260422 297654
rect 260186 297098 260422 297334
rect 260186 261418 260422 261654
rect 260186 261098 260422 261334
rect 260186 225418 260422 225654
rect 260186 225098 260422 225334
rect 260186 189418 260422 189654
rect 260186 189098 260422 189334
rect 260186 153418 260422 153654
rect 260186 153098 260422 153334
rect 260186 117418 260422 117654
rect 260186 117098 260422 117334
rect 260186 81418 260422 81654
rect 260186 81098 260422 81334
rect 260186 45418 260422 45654
rect 260186 45098 260422 45334
rect 260186 9418 260422 9654
rect 260186 9098 260422 9334
rect 260186 -4262 260422 -4026
rect 260186 -4582 260422 -4346
rect 281786 711042 282022 711278
rect 281786 710722 282022 710958
rect 278186 709202 278422 709438
rect 278186 708882 278422 709118
rect 274586 707362 274822 707598
rect 274586 707042 274822 707278
rect 263786 697018 264022 697254
rect 263786 696698 264022 696934
rect 263786 661018 264022 661254
rect 263786 660698 264022 660934
rect 263786 625018 264022 625254
rect 263786 624698 264022 624934
rect 263786 589018 264022 589254
rect 263786 588698 264022 588934
rect 263786 553018 264022 553254
rect 263786 552698 264022 552934
rect 263786 517018 264022 517254
rect 263786 516698 264022 516934
rect 263786 481018 264022 481254
rect 263786 480698 264022 480934
rect 263786 445018 264022 445254
rect 263786 444698 264022 444934
rect 263786 409018 264022 409254
rect 263786 408698 264022 408934
rect 263786 373018 264022 373254
rect 263786 372698 264022 372934
rect 263786 337018 264022 337254
rect 263786 336698 264022 336934
rect 263786 301018 264022 301254
rect 263786 300698 264022 300934
rect 263786 265018 264022 265254
rect 263786 264698 264022 264934
rect 263786 229018 264022 229254
rect 263786 228698 264022 228934
rect 263786 193018 264022 193254
rect 263786 192698 264022 192934
rect 263786 157018 264022 157254
rect 263786 156698 264022 156934
rect 263786 121018 264022 121254
rect 263786 120698 264022 120934
rect 263786 85018 264022 85254
rect 263786 84698 264022 84934
rect 263786 49018 264022 49254
rect 263786 48698 264022 48934
rect 263786 13018 264022 13254
rect 263786 12698 264022 12934
rect 245786 -7022 246022 -6786
rect 245786 -7342 246022 -7106
rect 270986 705522 271222 705758
rect 270986 705202 271222 705438
rect 270986 668218 271222 668454
rect 270986 667898 271222 668134
rect 270986 632218 271222 632454
rect 270986 631898 271222 632134
rect 270986 596218 271222 596454
rect 270986 595898 271222 596134
rect 270986 560218 271222 560454
rect 270986 559898 271222 560134
rect 270986 524218 271222 524454
rect 270986 523898 271222 524134
rect 270986 488218 271222 488454
rect 270986 487898 271222 488134
rect 270986 452218 271222 452454
rect 270986 451898 271222 452134
rect 270986 416218 271222 416454
rect 270986 415898 271222 416134
rect 270986 380218 271222 380454
rect 270986 379898 271222 380134
rect 270986 344218 271222 344454
rect 270986 343898 271222 344134
rect 270986 308218 271222 308454
rect 270986 307898 271222 308134
rect 270986 272218 271222 272454
rect 270986 271898 271222 272134
rect 270986 236218 271222 236454
rect 270986 235898 271222 236134
rect 270986 200218 271222 200454
rect 270986 199898 271222 200134
rect 270986 164218 271222 164454
rect 270986 163898 271222 164134
rect 270986 128218 271222 128454
rect 270986 127898 271222 128134
rect 270986 92218 271222 92454
rect 270986 91898 271222 92134
rect 270986 56218 271222 56454
rect 270986 55898 271222 56134
rect 270986 20218 271222 20454
rect 270986 19898 271222 20134
rect 270986 -1502 271222 -1266
rect 270986 -1822 271222 -1586
rect 274586 671818 274822 672054
rect 274586 671498 274822 671734
rect 274586 635818 274822 636054
rect 274586 635498 274822 635734
rect 274586 599818 274822 600054
rect 274586 599498 274822 599734
rect 274586 563818 274822 564054
rect 274586 563498 274822 563734
rect 274586 527818 274822 528054
rect 274586 527498 274822 527734
rect 274586 491818 274822 492054
rect 274586 491498 274822 491734
rect 274586 455818 274822 456054
rect 274586 455498 274822 455734
rect 274586 419818 274822 420054
rect 274586 419498 274822 419734
rect 278186 675418 278422 675654
rect 278186 675098 278422 675334
rect 278186 639418 278422 639654
rect 278186 639098 278422 639334
rect 278186 603418 278422 603654
rect 278186 603098 278422 603334
rect 278186 567418 278422 567654
rect 278186 567098 278422 567334
rect 278186 531418 278422 531654
rect 278186 531098 278422 531334
rect 278186 495418 278422 495654
rect 278186 495098 278422 495334
rect 278186 459418 278422 459654
rect 278186 459098 278422 459334
rect 278186 423418 278422 423654
rect 278186 423098 278422 423334
rect 274586 383818 274822 384054
rect 274586 383498 274822 383734
rect 274586 347818 274822 348054
rect 274586 347498 274822 347734
rect 274586 311818 274822 312054
rect 274586 311498 274822 311734
rect 274586 275818 274822 276054
rect 274586 275498 274822 275734
rect 274586 239818 274822 240054
rect 274586 239498 274822 239734
rect 274586 203818 274822 204054
rect 274586 203498 274822 203734
rect 274586 167818 274822 168054
rect 274586 167498 274822 167734
rect 274586 131818 274822 132054
rect 274586 131498 274822 131734
rect 274586 95818 274822 96054
rect 274586 95498 274822 95734
rect 274586 59818 274822 60054
rect 274586 59498 274822 59734
rect 274586 23818 274822 24054
rect 274586 23498 274822 23734
rect 274586 -3342 274822 -3106
rect 274586 -3662 274822 -3426
rect 278186 387418 278422 387654
rect 278186 387098 278422 387334
rect 278186 351418 278422 351654
rect 278186 351098 278422 351334
rect 278186 315418 278422 315654
rect 278186 315098 278422 315334
rect 278186 279418 278422 279654
rect 278186 279098 278422 279334
rect 278186 243418 278422 243654
rect 278186 243098 278422 243334
rect 278186 207418 278422 207654
rect 278186 207098 278422 207334
rect 278186 171418 278422 171654
rect 278186 171098 278422 171334
rect 278186 135418 278422 135654
rect 278186 135098 278422 135334
rect 278186 99418 278422 99654
rect 278186 99098 278422 99334
rect 278186 63418 278422 63654
rect 278186 63098 278422 63334
rect 278186 27418 278422 27654
rect 278186 27098 278422 27334
rect 278186 -5182 278422 -4946
rect 278186 -5502 278422 -5266
rect 299786 710122 300022 710358
rect 299786 709802 300022 710038
rect 296186 708282 296422 708518
rect 296186 707962 296422 708198
rect 292586 706442 292822 706678
rect 292586 706122 292822 706358
rect 281786 679018 282022 679254
rect 281786 678698 282022 678934
rect 281786 643018 282022 643254
rect 281786 642698 282022 642934
rect 281786 607018 282022 607254
rect 281786 606698 282022 606934
rect 281786 571018 282022 571254
rect 281786 570698 282022 570934
rect 281786 535018 282022 535254
rect 281786 534698 282022 534934
rect 281786 499018 282022 499254
rect 281786 498698 282022 498934
rect 281786 463018 282022 463254
rect 281786 462698 282022 462934
rect 281786 427018 282022 427254
rect 281786 426698 282022 426934
rect 288986 704602 289222 704838
rect 288986 704282 289222 704518
rect 288986 686218 289222 686454
rect 288986 685898 289222 686134
rect 288986 650218 289222 650454
rect 288986 649898 289222 650134
rect 288986 614218 289222 614454
rect 288986 613898 289222 614134
rect 288986 578218 289222 578454
rect 288986 577898 289222 578134
rect 288986 542218 289222 542454
rect 288986 541898 289222 542134
rect 288986 506218 289222 506454
rect 288986 505898 289222 506134
rect 288986 470218 289222 470454
rect 288986 469898 289222 470134
rect 288986 434218 289222 434454
rect 288986 433898 289222 434134
rect 281786 391018 282022 391254
rect 281786 390698 282022 390934
rect 281786 355018 282022 355254
rect 281786 354698 282022 354934
rect 281786 319018 282022 319254
rect 281786 318698 282022 318934
rect 281786 283018 282022 283254
rect 281786 282698 282022 282934
rect 281786 247018 282022 247254
rect 281786 246698 282022 246934
rect 281786 211018 282022 211254
rect 281786 210698 282022 210934
rect 281786 175018 282022 175254
rect 281786 174698 282022 174934
rect 281786 139018 282022 139254
rect 281786 138698 282022 138934
rect 288986 398218 289222 398454
rect 288986 397898 289222 398134
rect 288986 362218 289222 362454
rect 288986 361898 289222 362134
rect 288986 326218 289222 326454
rect 288986 325898 289222 326134
rect 288986 290218 289222 290454
rect 288986 289898 289222 290134
rect 288986 254218 289222 254454
rect 288986 253898 289222 254134
rect 288986 218218 289222 218454
rect 288986 217898 289222 218134
rect 288986 182218 289222 182454
rect 288986 181898 289222 182134
rect 288986 146218 289222 146454
rect 288986 145898 289222 146134
rect 288986 110218 289222 110454
rect 288986 109898 289222 110134
rect 281786 103018 282022 103254
rect 281786 102698 282022 102934
rect 281786 67018 282022 67254
rect 281786 66698 282022 66934
rect 281786 31018 282022 31254
rect 281786 30698 282022 30934
rect 263786 -6102 264022 -5866
rect 263786 -6422 264022 -6186
rect 288986 74218 289222 74454
rect 288986 73898 289222 74134
rect 288986 38218 289222 38454
rect 288986 37898 289222 38134
rect 288986 2218 289222 2454
rect 288986 1898 289222 2134
rect 288986 -582 289222 -346
rect 288986 -902 289222 -666
rect 292586 689818 292822 690054
rect 292586 689498 292822 689734
rect 292586 653818 292822 654054
rect 292586 653498 292822 653734
rect 292586 617818 292822 618054
rect 292586 617498 292822 617734
rect 292586 581818 292822 582054
rect 292586 581498 292822 581734
rect 292586 545818 292822 546054
rect 292586 545498 292822 545734
rect 292586 509818 292822 510054
rect 292586 509498 292822 509734
rect 292586 473818 292822 474054
rect 292586 473498 292822 473734
rect 292586 437818 292822 438054
rect 292586 437498 292822 437734
rect 292586 401818 292822 402054
rect 292586 401498 292822 401734
rect 292586 365818 292822 366054
rect 292586 365498 292822 365734
rect 292586 329818 292822 330054
rect 292586 329498 292822 329734
rect 292586 293818 292822 294054
rect 292586 293498 292822 293734
rect 292586 257818 292822 258054
rect 292586 257498 292822 257734
rect 292586 221818 292822 222054
rect 292586 221498 292822 221734
rect 292586 185818 292822 186054
rect 292586 185498 292822 185734
rect 292586 149818 292822 150054
rect 292586 149498 292822 149734
rect 292586 113818 292822 114054
rect 292586 113498 292822 113734
rect 292586 77818 292822 78054
rect 292586 77498 292822 77734
rect 292586 41818 292822 42054
rect 292586 41498 292822 41734
rect 292586 5818 292822 6054
rect 292586 5498 292822 5734
rect 292586 -2422 292822 -2186
rect 292586 -2742 292822 -2506
rect 296186 693418 296422 693654
rect 296186 693098 296422 693334
rect 296186 657418 296422 657654
rect 296186 657098 296422 657334
rect 296186 621418 296422 621654
rect 296186 621098 296422 621334
rect 296186 585418 296422 585654
rect 296186 585098 296422 585334
rect 296186 549418 296422 549654
rect 296186 549098 296422 549334
rect 296186 513418 296422 513654
rect 296186 513098 296422 513334
rect 296186 477418 296422 477654
rect 296186 477098 296422 477334
rect 296186 441418 296422 441654
rect 296186 441098 296422 441334
rect 296186 405418 296422 405654
rect 296186 405098 296422 405334
rect 296186 369418 296422 369654
rect 296186 369098 296422 369334
rect 296186 333418 296422 333654
rect 296186 333098 296422 333334
rect 296186 297418 296422 297654
rect 296186 297098 296422 297334
rect 296186 261418 296422 261654
rect 296186 261098 296422 261334
rect 296186 225418 296422 225654
rect 296186 225098 296422 225334
rect 296186 189418 296422 189654
rect 296186 189098 296422 189334
rect 296186 153418 296422 153654
rect 296186 153098 296422 153334
rect 296186 117418 296422 117654
rect 296186 117098 296422 117334
rect 296186 81418 296422 81654
rect 296186 81098 296422 81334
rect 296186 45418 296422 45654
rect 296186 45098 296422 45334
rect 296186 9418 296422 9654
rect 296186 9098 296422 9334
rect 296186 -4262 296422 -4026
rect 296186 -4582 296422 -4346
rect 317786 711042 318022 711278
rect 317786 710722 318022 710958
rect 314186 709202 314422 709438
rect 314186 708882 314422 709118
rect 310586 707362 310822 707598
rect 310586 707042 310822 707278
rect 299786 697018 300022 697254
rect 299786 696698 300022 696934
rect 299786 661018 300022 661254
rect 299786 660698 300022 660934
rect 299786 625018 300022 625254
rect 299786 624698 300022 624934
rect 299786 589018 300022 589254
rect 299786 588698 300022 588934
rect 299786 553018 300022 553254
rect 299786 552698 300022 552934
rect 299786 517018 300022 517254
rect 299786 516698 300022 516934
rect 299786 481018 300022 481254
rect 299786 480698 300022 480934
rect 299786 445018 300022 445254
rect 299786 444698 300022 444934
rect 299786 409018 300022 409254
rect 299786 408698 300022 408934
rect 299786 373018 300022 373254
rect 299786 372698 300022 372934
rect 299786 337018 300022 337254
rect 299786 336698 300022 336934
rect 299786 301018 300022 301254
rect 299786 300698 300022 300934
rect 299786 265018 300022 265254
rect 299786 264698 300022 264934
rect 299786 229018 300022 229254
rect 299786 228698 300022 228934
rect 299786 193018 300022 193254
rect 299786 192698 300022 192934
rect 299786 157018 300022 157254
rect 299786 156698 300022 156934
rect 299786 121018 300022 121254
rect 299786 120698 300022 120934
rect 299786 85018 300022 85254
rect 299786 84698 300022 84934
rect 299786 49018 300022 49254
rect 299786 48698 300022 48934
rect 299786 13018 300022 13254
rect 299786 12698 300022 12934
rect 281786 -7022 282022 -6786
rect 281786 -7342 282022 -7106
rect 306986 705522 307222 705758
rect 306986 705202 307222 705438
rect 306986 668218 307222 668454
rect 306986 667898 307222 668134
rect 306986 632218 307222 632454
rect 306986 631898 307222 632134
rect 306986 596218 307222 596454
rect 306986 595898 307222 596134
rect 306986 560218 307222 560454
rect 306986 559898 307222 560134
rect 306986 524218 307222 524454
rect 306986 523898 307222 524134
rect 306986 488218 307222 488454
rect 306986 487898 307222 488134
rect 306986 452218 307222 452454
rect 306986 451898 307222 452134
rect 306986 416218 307222 416454
rect 306986 415898 307222 416134
rect 306986 380218 307222 380454
rect 306986 379898 307222 380134
rect 306986 344218 307222 344454
rect 306986 343898 307222 344134
rect 306986 308218 307222 308454
rect 306986 307898 307222 308134
rect 306986 272218 307222 272454
rect 306986 271898 307222 272134
rect 306986 236218 307222 236454
rect 306986 235898 307222 236134
rect 306986 200218 307222 200454
rect 306986 199898 307222 200134
rect 306986 164218 307222 164454
rect 306986 163898 307222 164134
rect 306986 128218 307222 128454
rect 306986 127898 307222 128134
rect 306986 92218 307222 92454
rect 306986 91898 307222 92134
rect 306986 56218 307222 56454
rect 306986 55898 307222 56134
rect 306986 20218 307222 20454
rect 306986 19898 307222 20134
rect 306986 -1502 307222 -1266
rect 306986 -1822 307222 -1586
rect 310586 671818 310822 672054
rect 310586 671498 310822 671734
rect 310586 635818 310822 636054
rect 310586 635498 310822 635734
rect 310586 599818 310822 600054
rect 310586 599498 310822 599734
rect 310586 563818 310822 564054
rect 310586 563498 310822 563734
rect 310586 527818 310822 528054
rect 310586 527498 310822 527734
rect 310586 491818 310822 492054
rect 310586 491498 310822 491734
rect 310586 455818 310822 456054
rect 310586 455498 310822 455734
rect 310586 419818 310822 420054
rect 310586 419498 310822 419734
rect 310586 383818 310822 384054
rect 310586 383498 310822 383734
rect 310586 347818 310822 348054
rect 310586 347498 310822 347734
rect 310586 311818 310822 312054
rect 310586 311498 310822 311734
rect 310586 275818 310822 276054
rect 310586 275498 310822 275734
rect 310586 239818 310822 240054
rect 310586 239498 310822 239734
rect 310586 203818 310822 204054
rect 310586 203498 310822 203734
rect 310586 167818 310822 168054
rect 310586 167498 310822 167734
rect 310586 131818 310822 132054
rect 310586 131498 310822 131734
rect 310586 95818 310822 96054
rect 310586 95498 310822 95734
rect 310586 59818 310822 60054
rect 310586 59498 310822 59734
rect 310586 23818 310822 24054
rect 310586 23498 310822 23734
rect 310586 -3342 310822 -3106
rect 310586 -3662 310822 -3426
rect 314186 675418 314422 675654
rect 314186 675098 314422 675334
rect 314186 639418 314422 639654
rect 314186 639098 314422 639334
rect 314186 603418 314422 603654
rect 314186 603098 314422 603334
rect 314186 567418 314422 567654
rect 314186 567098 314422 567334
rect 314186 531418 314422 531654
rect 314186 531098 314422 531334
rect 314186 495418 314422 495654
rect 314186 495098 314422 495334
rect 314186 459418 314422 459654
rect 314186 459098 314422 459334
rect 314186 423418 314422 423654
rect 314186 423098 314422 423334
rect 314186 387418 314422 387654
rect 314186 387098 314422 387334
rect 314186 351418 314422 351654
rect 314186 351098 314422 351334
rect 314186 315418 314422 315654
rect 314186 315098 314422 315334
rect 314186 279418 314422 279654
rect 314186 279098 314422 279334
rect 314186 243418 314422 243654
rect 314186 243098 314422 243334
rect 314186 207418 314422 207654
rect 314186 207098 314422 207334
rect 314186 171418 314422 171654
rect 314186 171098 314422 171334
rect 314186 135418 314422 135654
rect 314186 135098 314422 135334
rect 314186 99418 314422 99654
rect 314186 99098 314422 99334
rect 314186 63418 314422 63654
rect 314186 63098 314422 63334
rect 314186 27418 314422 27654
rect 314186 27098 314422 27334
rect 314186 -5182 314422 -4946
rect 314186 -5502 314422 -5266
rect 335786 710122 336022 710358
rect 335786 709802 336022 710038
rect 332186 708282 332422 708518
rect 332186 707962 332422 708198
rect 328586 706442 328822 706678
rect 328586 706122 328822 706358
rect 317786 679018 318022 679254
rect 317786 678698 318022 678934
rect 317786 643018 318022 643254
rect 317786 642698 318022 642934
rect 317786 607018 318022 607254
rect 317786 606698 318022 606934
rect 317786 571018 318022 571254
rect 317786 570698 318022 570934
rect 317786 535018 318022 535254
rect 317786 534698 318022 534934
rect 317786 499018 318022 499254
rect 317786 498698 318022 498934
rect 317786 463018 318022 463254
rect 317786 462698 318022 462934
rect 317786 427018 318022 427254
rect 317786 426698 318022 426934
rect 317786 391018 318022 391254
rect 317786 390698 318022 390934
rect 317786 355018 318022 355254
rect 317786 354698 318022 354934
rect 317786 319018 318022 319254
rect 317786 318698 318022 318934
rect 317786 283018 318022 283254
rect 317786 282698 318022 282934
rect 317786 247018 318022 247254
rect 317786 246698 318022 246934
rect 324986 704602 325222 704838
rect 324986 704282 325222 704518
rect 324986 686218 325222 686454
rect 324986 685898 325222 686134
rect 324986 650218 325222 650454
rect 324986 649898 325222 650134
rect 324986 614218 325222 614454
rect 324986 613898 325222 614134
rect 324986 578218 325222 578454
rect 324986 577898 325222 578134
rect 324986 542218 325222 542454
rect 324986 541898 325222 542134
rect 324986 506218 325222 506454
rect 324986 505898 325222 506134
rect 324986 470218 325222 470454
rect 324986 469898 325222 470134
rect 324986 434218 325222 434454
rect 324986 433898 325222 434134
rect 324986 398218 325222 398454
rect 324986 397898 325222 398134
rect 324986 362218 325222 362454
rect 324986 361898 325222 362134
rect 324986 326218 325222 326454
rect 324986 325898 325222 326134
rect 324986 290218 325222 290454
rect 324986 289898 325222 290134
rect 324986 254218 325222 254454
rect 324986 253898 325222 254134
rect 317786 211018 318022 211254
rect 317786 210698 318022 210934
rect 317786 175018 318022 175254
rect 317786 174698 318022 174934
rect 317786 139018 318022 139254
rect 317786 138698 318022 138934
rect 317786 103018 318022 103254
rect 317786 102698 318022 102934
rect 324986 218218 325222 218454
rect 324986 217898 325222 218134
rect 324986 182218 325222 182454
rect 324986 181898 325222 182134
rect 324986 146218 325222 146454
rect 324986 145898 325222 146134
rect 324986 110218 325222 110454
rect 324986 109898 325222 110134
rect 317786 67018 318022 67254
rect 317786 66698 318022 66934
rect 317786 31018 318022 31254
rect 317786 30698 318022 30934
rect 299786 -6102 300022 -5866
rect 299786 -6422 300022 -6186
rect 324986 74218 325222 74454
rect 324986 73898 325222 74134
rect 324986 38218 325222 38454
rect 324986 37898 325222 38134
rect 324986 2218 325222 2454
rect 324986 1898 325222 2134
rect 324986 -582 325222 -346
rect 324986 -902 325222 -666
rect 328586 689818 328822 690054
rect 328586 689498 328822 689734
rect 328586 653818 328822 654054
rect 328586 653498 328822 653734
rect 328586 617818 328822 618054
rect 328586 617498 328822 617734
rect 328586 581818 328822 582054
rect 328586 581498 328822 581734
rect 328586 545818 328822 546054
rect 328586 545498 328822 545734
rect 328586 509818 328822 510054
rect 328586 509498 328822 509734
rect 328586 473818 328822 474054
rect 328586 473498 328822 473734
rect 328586 437818 328822 438054
rect 328586 437498 328822 437734
rect 328586 401818 328822 402054
rect 328586 401498 328822 401734
rect 328586 365818 328822 366054
rect 328586 365498 328822 365734
rect 328586 329818 328822 330054
rect 328586 329498 328822 329734
rect 328586 293818 328822 294054
rect 328586 293498 328822 293734
rect 328586 257818 328822 258054
rect 328586 257498 328822 257734
rect 328586 221818 328822 222054
rect 328586 221498 328822 221734
rect 328586 185818 328822 186054
rect 328586 185498 328822 185734
rect 328586 149818 328822 150054
rect 328586 149498 328822 149734
rect 328586 113818 328822 114054
rect 328586 113498 328822 113734
rect 328586 77818 328822 78054
rect 328586 77498 328822 77734
rect 328586 41818 328822 42054
rect 328586 41498 328822 41734
rect 328586 5818 328822 6054
rect 328586 5498 328822 5734
rect 328586 -2422 328822 -2186
rect 328586 -2742 328822 -2506
rect 332186 693418 332422 693654
rect 332186 693098 332422 693334
rect 332186 657418 332422 657654
rect 332186 657098 332422 657334
rect 332186 621418 332422 621654
rect 332186 621098 332422 621334
rect 332186 585418 332422 585654
rect 332186 585098 332422 585334
rect 332186 549418 332422 549654
rect 332186 549098 332422 549334
rect 332186 513418 332422 513654
rect 332186 513098 332422 513334
rect 332186 477418 332422 477654
rect 332186 477098 332422 477334
rect 332186 441418 332422 441654
rect 332186 441098 332422 441334
rect 332186 405418 332422 405654
rect 332186 405098 332422 405334
rect 332186 369418 332422 369654
rect 332186 369098 332422 369334
rect 332186 333418 332422 333654
rect 332186 333098 332422 333334
rect 332186 297418 332422 297654
rect 332186 297098 332422 297334
rect 332186 261418 332422 261654
rect 332186 261098 332422 261334
rect 332186 225418 332422 225654
rect 332186 225098 332422 225334
rect 332186 189418 332422 189654
rect 332186 189098 332422 189334
rect 332186 153418 332422 153654
rect 332186 153098 332422 153334
rect 332186 117418 332422 117654
rect 332186 117098 332422 117334
rect 332186 81418 332422 81654
rect 332186 81098 332422 81334
rect 332186 45418 332422 45654
rect 332186 45098 332422 45334
rect 332186 9418 332422 9654
rect 332186 9098 332422 9334
rect 332186 -4262 332422 -4026
rect 332186 -4582 332422 -4346
rect 353786 711042 354022 711278
rect 353786 710722 354022 710958
rect 350186 709202 350422 709438
rect 350186 708882 350422 709118
rect 346586 707362 346822 707598
rect 346586 707042 346822 707278
rect 335786 697018 336022 697254
rect 335786 696698 336022 696934
rect 335786 661018 336022 661254
rect 335786 660698 336022 660934
rect 335786 625018 336022 625254
rect 335786 624698 336022 624934
rect 335786 589018 336022 589254
rect 335786 588698 336022 588934
rect 335786 553018 336022 553254
rect 335786 552698 336022 552934
rect 335786 517018 336022 517254
rect 335786 516698 336022 516934
rect 335786 481018 336022 481254
rect 335786 480698 336022 480934
rect 335786 445018 336022 445254
rect 335786 444698 336022 444934
rect 335786 409018 336022 409254
rect 335786 408698 336022 408934
rect 335786 373018 336022 373254
rect 335786 372698 336022 372934
rect 335786 337018 336022 337254
rect 335786 336698 336022 336934
rect 335786 301018 336022 301254
rect 335786 300698 336022 300934
rect 335786 265018 336022 265254
rect 335786 264698 336022 264934
rect 335786 229018 336022 229254
rect 335786 228698 336022 228934
rect 342986 705522 343222 705758
rect 342986 705202 343222 705438
rect 342986 668218 343222 668454
rect 342986 667898 343222 668134
rect 342986 632218 343222 632454
rect 342986 631898 343222 632134
rect 342986 596218 343222 596454
rect 342986 595898 343222 596134
rect 342986 560218 343222 560454
rect 342986 559898 343222 560134
rect 342986 524218 343222 524454
rect 342986 523898 343222 524134
rect 342986 488218 343222 488454
rect 342986 487898 343222 488134
rect 342986 452218 343222 452454
rect 342986 451898 343222 452134
rect 342986 416218 343222 416454
rect 342986 415898 343222 416134
rect 342986 380218 343222 380454
rect 342986 379898 343222 380134
rect 342986 344218 343222 344454
rect 342986 343898 343222 344134
rect 342986 308218 343222 308454
rect 342986 307898 343222 308134
rect 342986 272218 343222 272454
rect 342986 271898 343222 272134
rect 342986 236218 343222 236454
rect 342986 235898 343222 236134
rect 335786 193018 336022 193254
rect 335786 192698 336022 192934
rect 335786 157018 336022 157254
rect 335786 156698 336022 156934
rect 335786 121018 336022 121254
rect 335786 120698 336022 120934
rect 335786 85018 336022 85254
rect 335786 84698 336022 84934
rect 342986 200218 343222 200454
rect 342986 199898 343222 200134
rect 342986 164218 343222 164454
rect 342986 163898 343222 164134
rect 342986 128218 343222 128454
rect 342986 127898 343222 128134
rect 342986 92218 343222 92454
rect 342986 91898 343222 92134
rect 335786 49018 336022 49254
rect 335786 48698 336022 48934
rect 335786 13018 336022 13254
rect 335786 12698 336022 12934
rect 317786 -7022 318022 -6786
rect 317786 -7342 318022 -7106
rect 342986 56218 343222 56454
rect 342986 55898 343222 56134
rect 342986 20218 343222 20454
rect 342986 19898 343222 20134
rect 342986 -1502 343222 -1266
rect 342986 -1822 343222 -1586
rect 346586 671818 346822 672054
rect 346586 671498 346822 671734
rect 346586 635818 346822 636054
rect 346586 635498 346822 635734
rect 346586 599818 346822 600054
rect 346586 599498 346822 599734
rect 346586 563818 346822 564054
rect 346586 563498 346822 563734
rect 346586 527818 346822 528054
rect 346586 527498 346822 527734
rect 346586 491818 346822 492054
rect 346586 491498 346822 491734
rect 346586 455818 346822 456054
rect 346586 455498 346822 455734
rect 346586 419818 346822 420054
rect 346586 419498 346822 419734
rect 346586 383818 346822 384054
rect 346586 383498 346822 383734
rect 346586 347818 346822 348054
rect 346586 347498 346822 347734
rect 346586 311818 346822 312054
rect 346586 311498 346822 311734
rect 346586 275818 346822 276054
rect 346586 275498 346822 275734
rect 346586 239818 346822 240054
rect 346586 239498 346822 239734
rect 346586 203818 346822 204054
rect 346586 203498 346822 203734
rect 346586 167818 346822 168054
rect 346586 167498 346822 167734
rect 346586 131818 346822 132054
rect 346586 131498 346822 131734
rect 346586 95818 346822 96054
rect 346586 95498 346822 95734
rect 346586 59818 346822 60054
rect 346586 59498 346822 59734
rect 346586 23818 346822 24054
rect 346586 23498 346822 23734
rect 346586 -3342 346822 -3106
rect 346586 -3662 346822 -3426
rect 350186 675418 350422 675654
rect 350186 675098 350422 675334
rect 350186 639418 350422 639654
rect 350186 639098 350422 639334
rect 350186 603418 350422 603654
rect 350186 603098 350422 603334
rect 350186 567418 350422 567654
rect 350186 567098 350422 567334
rect 350186 531418 350422 531654
rect 350186 531098 350422 531334
rect 350186 495418 350422 495654
rect 350186 495098 350422 495334
rect 350186 459418 350422 459654
rect 350186 459098 350422 459334
rect 350186 423418 350422 423654
rect 350186 423098 350422 423334
rect 350186 387418 350422 387654
rect 350186 387098 350422 387334
rect 350186 351418 350422 351654
rect 350186 351098 350422 351334
rect 350186 315418 350422 315654
rect 350186 315098 350422 315334
rect 350186 279418 350422 279654
rect 350186 279098 350422 279334
rect 350186 243418 350422 243654
rect 350186 243098 350422 243334
rect 350186 207418 350422 207654
rect 350186 207098 350422 207334
rect 350186 171418 350422 171654
rect 350186 171098 350422 171334
rect 350186 135418 350422 135654
rect 350186 135098 350422 135334
rect 350186 99418 350422 99654
rect 350186 99098 350422 99334
rect 350186 63418 350422 63654
rect 350186 63098 350422 63334
rect 350186 27418 350422 27654
rect 350186 27098 350422 27334
rect 350186 -5182 350422 -4946
rect 350186 -5502 350422 -5266
rect 371786 710122 372022 710358
rect 371786 709802 372022 710038
rect 368186 708282 368422 708518
rect 368186 707962 368422 708198
rect 364586 706442 364822 706678
rect 364586 706122 364822 706358
rect 353786 679018 354022 679254
rect 353786 678698 354022 678934
rect 353786 643018 354022 643254
rect 353786 642698 354022 642934
rect 353786 607018 354022 607254
rect 353786 606698 354022 606934
rect 353786 571018 354022 571254
rect 353786 570698 354022 570934
rect 353786 535018 354022 535254
rect 353786 534698 354022 534934
rect 353786 499018 354022 499254
rect 353786 498698 354022 498934
rect 353786 463018 354022 463254
rect 353786 462698 354022 462934
rect 353786 427018 354022 427254
rect 353786 426698 354022 426934
rect 353786 391018 354022 391254
rect 353786 390698 354022 390934
rect 353786 355018 354022 355254
rect 353786 354698 354022 354934
rect 353786 319018 354022 319254
rect 353786 318698 354022 318934
rect 353786 283018 354022 283254
rect 353786 282698 354022 282934
rect 353786 247018 354022 247254
rect 353786 246698 354022 246934
rect 353786 211018 354022 211254
rect 353786 210698 354022 210934
rect 353786 175018 354022 175254
rect 353786 174698 354022 174934
rect 353786 139018 354022 139254
rect 353786 138698 354022 138934
rect 353786 103018 354022 103254
rect 353786 102698 354022 102934
rect 353786 67018 354022 67254
rect 353786 66698 354022 66934
rect 353786 31018 354022 31254
rect 353786 30698 354022 30934
rect 335786 -6102 336022 -5866
rect 335786 -6422 336022 -6186
rect 360986 704602 361222 704838
rect 360986 704282 361222 704518
rect 360986 686218 361222 686454
rect 360986 685898 361222 686134
rect 360986 650218 361222 650454
rect 360986 649898 361222 650134
rect 360986 614218 361222 614454
rect 360986 613898 361222 614134
rect 360986 578218 361222 578454
rect 360986 577898 361222 578134
rect 360986 542218 361222 542454
rect 360986 541898 361222 542134
rect 360986 506218 361222 506454
rect 360986 505898 361222 506134
rect 360986 470218 361222 470454
rect 360986 469898 361222 470134
rect 360986 434218 361222 434454
rect 360986 433898 361222 434134
rect 360986 398218 361222 398454
rect 360986 397898 361222 398134
rect 360986 362218 361222 362454
rect 360986 361898 361222 362134
rect 360986 326218 361222 326454
rect 360986 325898 361222 326134
rect 360986 290218 361222 290454
rect 360986 289898 361222 290134
rect 360986 254218 361222 254454
rect 360986 253898 361222 254134
rect 360986 218218 361222 218454
rect 360986 217898 361222 218134
rect 360986 182218 361222 182454
rect 360986 181898 361222 182134
rect 360986 146218 361222 146454
rect 360986 145898 361222 146134
rect 360986 110218 361222 110454
rect 360986 109898 361222 110134
rect 360986 74218 361222 74454
rect 360986 73898 361222 74134
rect 360986 38218 361222 38454
rect 360986 37898 361222 38134
rect 360986 2218 361222 2454
rect 360986 1898 361222 2134
rect 360986 -582 361222 -346
rect 360986 -902 361222 -666
rect 364586 689818 364822 690054
rect 364586 689498 364822 689734
rect 364586 653818 364822 654054
rect 364586 653498 364822 653734
rect 364586 617818 364822 618054
rect 364586 617498 364822 617734
rect 364586 581818 364822 582054
rect 364586 581498 364822 581734
rect 364586 545818 364822 546054
rect 364586 545498 364822 545734
rect 364586 509818 364822 510054
rect 364586 509498 364822 509734
rect 364586 473818 364822 474054
rect 364586 473498 364822 473734
rect 364586 437818 364822 438054
rect 364586 437498 364822 437734
rect 364586 401818 364822 402054
rect 364586 401498 364822 401734
rect 364586 365818 364822 366054
rect 364586 365498 364822 365734
rect 364586 329818 364822 330054
rect 364586 329498 364822 329734
rect 364586 293818 364822 294054
rect 364586 293498 364822 293734
rect 364586 257818 364822 258054
rect 364586 257498 364822 257734
rect 364586 221818 364822 222054
rect 364586 221498 364822 221734
rect 364586 185818 364822 186054
rect 364586 185498 364822 185734
rect 364586 149818 364822 150054
rect 364586 149498 364822 149734
rect 364586 113818 364822 114054
rect 364586 113498 364822 113734
rect 364586 77818 364822 78054
rect 364586 77498 364822 77734
rect 364586 41818 364822 42054
rect 364586 41498 364822 41734
rect 364586 5818 364822 6054
rect 364586 5498 364822 5734
rect 364586 -2422 364822 -2186
rect 364586 -2742 364822 -2506
rect 368186 693418 368422 693654
rect 368186 693098 368422 693334
rect 368186 657418 368422 657654
rect 368186 657098 368422 657334
rect 368186 621418 368422 621654
rect 368186 621098 368422 621334
rect 368186 585418 368422 585654
rect 368186 585098 368422 585334
rect 368186 549418 368422 549654
rect 368186 549098 368422 549334
rect 368186 513418 368422 513654
rect 368186 513098 368422 513334
rect 368186 477418 368422 477654
rect 368186 477098 368422 477334
rect 368186 441418 368422 441654
rect 368186 441098 368422 441334
rect 368186 405418 368422 405654
rect 368186 405098 368422 405334
rect 368186 369418 368422 369654
rect 368186 369098 368422 369334
rect 368186 333418 368422 333654
rect 368186 333098 368422 333334
rect 368186 297418 368422 297654
rect 368186 297098 368422 297334
rect 368186 261418 368422 261654
rect 368186 261098 368422 261334
rect 368186 225418 368422 225654
rect 368186 225098 368422 225334
rect 368186 189418 368422 189654
rect 368186 189098 368422 189334
rect 368186 153418 368422 153654
rect 368186 153098 368422 153334
rect 368186 117418 368422 117654
rect 368186 117098 368422 117334
rect 368186 81418 368422 81654
rect 368186 81098 368422 81334
rect 368186 45418 368422 45654
rect 368186 45098 368422 45334
rect 368186 9418 368422 9654
rect 368186 9098 368422 9334
rect 368186 -4262 368422 -4026
rect 368186 -4582 368422 -4346
rect 389786 711042 390022 711278
rect 389786 710722 390022 710958
rect 386186 709202 386422 709438
rect 386186 708882 386422 709118
rect 382586 707362 382822 707598
rect 382586 707042 382822 707278
rect 371786 697018 372022 697254
rect 371786 696698 372022 696934
rect 371786 661018 372022 661254
rect 371786 660698 372022 660934
rect 371786 625018 372022 625254
rect 371786 624698 372022 624934
rect 371786 589018 372022 589254
rect 371786 588698 372022 588934
rect 371786 553018 372022 553254
rect 371786 552698 372022 552934
rect 371786 517018 372022 517254
rect 371786 516698 372022 516934
rect 371786 481018 372022 481254
rect 371786 480698 372022 480934
rect 371786 445018 372022 445254
rect 371786 444698 372022 444934
rect 371786 409018 372022 409254
rect 371786 408698 372022 408934
rect 371786 373018 372022 373254
rect 371786 372698 372022 372934
rect 371786 337018 372022 337254
rect 371786 336698 372022 336934
rect 371786 301018 372022 301254
rect 371786 300698 372022 300934
rect 371786 265018 372022 265254
rect 371786 264698 372022 264934
rect 371786 229018 372022 229254
rect 371786 228698 372022 228934
rect 371786 193018 372022 193254
rect 371786 192698 372022 192934
rect 371786 157018 372022 157254
rect 371786 156698 372022 156934
rect 371786 121018 372022 121254
rect 371786 120698 372022 120934
rect 371786 85018 372022 85254
rect 371786 84698 372022 84934
rect 371786 49018 372022 49254
rect 371786 48698 372022 48934
rect 371786 13018 372022 13254
rect 371786 12698 372022 12934
rect 353786 -7022 354022 -6786
rect 353786 -7342 354022 -7106
rect 378986 705522 379222 705758
rect 378986 705202 379222 705438
rect 378986 668218 379222 668454
rect 378986 667898 379222 668134
rect 378986 632218 379222 632454
rect 378986 631898 379222 632134
rect 378986 596218 379222 596454
rect 378986 595898 379222 596134
rect 378986 560218 379222 560454
rect 378986 559898 379222 560134
rect 378986 524218 379222 524454
rect 378986 523898 379222 524134
rect 378986 488218 379222 488454
rect 378986 487898 379222 488134
rect 378986 452218 379222 452454
rect 378986 451898 379222 452134
rect 378986 416218 379222 416454
rect 378986 415898 379222 416134
rect 378986 380218 379222 380454
rect 378986 379898 379222 380134
rect 378986 344218 379222 344454
rect 378986 343898 379222 344134
rect 378986 308218 379222 308454
rect 378986 307898 379222 308134
rect 378986 272218 379222 272454
rect 378986 271898 379222 272134
rect 378986 236218 379222 236454
rect 378986 235898 379222 236134
rect 378986 200218 379222 200454
rect 378986 199898 379222 200134
rect 378986 164218 379222 164454
rect 378986 163898 379222 164134
rect 378986 128218 379222 128454
rect 378986 127898 379222 128134
rect 378986 92218 379222 92454
rect 378986 91898 379222 92134
rect 378986 56218 379222 56454
rect 378986 55898 379222 56134
rect 378986 20218 379222 20454
rect 378986 19898 379222 20134
rect 378986 -1502 379222 -1266
rect 378986 -1822 379222 -1586
rect 382586 671818 382822 672054
rect 382586 671498 382822 671734
rect 382586 635818 382822 636054
rect 382586 635498 382822 635734
rect 382586 599818 382822 600054
rect 382586 599498 382822 599734
rect 382586 563818 382822 564054
rect 382586 563498 382822 563734
rect 382586 527818 382822 528054
rect 382586 527498 382822 527734
rect 382586 491818 382822 492054
rect 382586 491498 382822 491734
rect 382586 455818 382822 456054
rect 382586 455498 382822 455734
rect 382586 419818 382822 420054
rect 382586 419498 382822 419734
rect 382586 383818 382822 384054
rect 382586 383498 382822 383734
rect 382586 347818 382822 348054
rect 382586 347498 382822 347734
rect 382586 311818 382822 312054
rect 382586 311498 382822 311734
rect 382586 275818 382822 276054
rect 382586 275498 382822 275734
rect 382586 239818 382822 240054
rect 382586 239498 382822 239734
rect 382586 203818 382822 204054
rect 382586 203498 382822 203734
rect 382586 167818 382822 168054
rect 382586 167498 382822 167734
rect 382586 131818 382822 132054
rect 382586 131498 382822 131734
rect 382586 95818 382822 96054
rect 382586 95498 382822 95734
rect 382586 59818 382822 60054
rect 382586 59498 382822 59734
rect 382586 23818 382822 24054
rect 382586 23498 382822 23734
rect 382586 -3342 382822 -3106
rect 382586 -3662 382822 -3426
rect 386186 675418 386422 675654
rect 386186 675098 386422 675334
rect 386186 639418 386422 639654
rect 386186 639098 386422 639334
rect 386186 603418 386422 603654
rect 386186 603098 386422 603334
rect 386186 567418 386422 567654
rect 386186 567098 386422 567334
rect 386186 531418 386422 531654
rect 386186 531098 386422 531334
rect 386186 495418 386422 495654
rect 386186 495098 386422 495334
rect 386186 459418 386422 459654
rect 386186 459098 386422 459334
rect 386186 423418 386422 423654
rect 386186 423098 386422 423334
rect 386186 387418 386422 387654
rect 386186 387098 386422 387334
rect 386186 351418 386422 351654
rect 386186 351098 386422 351334
rect 386186 315418 386422 315654
rect 386186 315098 386422 315334
rect 386186 279418 386422 279654
rect 386186 279098 386422 279334
rect 386186 243418 386422 243654
rect 386186 243098 386422 243334
rect 386186 207418 386422 207654
rect 386186 207098 386422 207334
rect 386186 171418 386422 171654
rect 386186 171098 386422 171334
rect 386186 135418 386422 135654
rect 386186 135098 386422 135334
rect 386186 99418 386422 99654
rect 386186 99098 386422 99334
rect 386186 63418 386422 63654
rect 386186 63098 386422 63334
rect 386186 27418 386422 27654
rect 386186 27098 386422 27334
rect 386186 -5182 386422 -4946
rect 386186 -5502 386422 -5266
rect 407786 710122 408022 710358
rect 407786 709802 408022 710038
rect 404186 708282 404422 708518
rect 404186 707962 404422 708198
rect 400586 706442 400822 706678
rect 400586 706122 400822 706358
rect 389786 679018 390022 679254
rect 389786 678698 390022 678934
rect 389786 643018 390022 643254
rect 389786 642698 390022 642934
rect 389786 607018 390022 607254
rect 389786 606698 390022 606934
rect 389786 571018 390022 571254
rect 389786 570698 390022 570934
rect 389786 535018 390022 535254
rect 389786 534698 390022 534934
rect 389786 499018 390022 499254
rect 389786 498698 390022 498934
rect 389786 463018 390022 463254
rect 389786 462698 390022 462934
rect 389786 427018 390022 427254
rect 389786 426698 390022 426934
rect 389786 391018 390022 391254
rect 389786 390698 390022 390934
rect 389786 355018 390022 355254
rect 389786 354698 390022 354934
rect 389786 319018 390022 319254
rect 389786 318698 390022 318934
rect 389786 283018 390022 283254
rect 389786 282698 390022 282934
rect 389786 247018 390022 247254
rect 389786 246698 390022 246934
rect 389786 211018 390022 211254
rect 389786 210698 390022 210934
rect 389786 175018 390022 175254
rect 389786 174698 390022 174934
rect 389786 139018 390022 139254
rect 389786 138698 390022 138934
rect 389786 103018 390022 103254
rect 389786 102698 390022 102934
rect 389786 67018 390022 67254
rect 389786 66698 390022 66934
rect 389786 31018 390022 31254
rect 389786 30698 390022 30934
rect 371786 -6102 372022 -5866
rect 371786 -6422 372022 -6186
rect 396986 704602 397222 704838
rect 396986 704282 397222 704518
rect 396986 686218 397222 686454
rect 396986 685898 397222 686134
rect 396986 650218 397222 650454
rect 396986 649898 397222 650134
rect 396986 614218 397222 614454
rect 396986 613898 397222 614134
rect 396986 578218 397222 578454
rect 396986 577898 397222 578134
rect 396986 542218 397222 542454
rect 396986 541898 397222 542134
rect 396986 506218 397222 506454
rect 396986 505898 397222 506134
rect 396986 470218 397222 470454
rect 396986 469898 397222 470134
rect 396986 434218 397222 434454
rect 396986 433898 397222 434134
rect 396986 398218 397222 398454
rect 396986 397898 397222 398134
rect 396986 362218 397222 362454
rect 396986 361898 397222 362134
rect 396986 326218 397222 326454
rect 396986 325898 397222 326134
rect 396986 290218 397222 290454
rect 396986 289898 397222 290134
rect 396986 254218 397222 254454
rect 396986 253898 397222 254134
rect 396986 218218 397222 218454
rect 396986 217898 397222 218134
rect 396986 182218 397222 182454
rect 396986 181898 397222 182134
rect 396986 146218 397222 146454
rect 396986 145898 397222 146134
rect 396986 110218 397222 110454
rect 396986 109898 397222 110134
rect 396986 74218 397222 74454
rect 396986 73898 397222 74134
rect 396986 38218 397222 38454
rect 396986 37898 397222 38134
rect 396986 2218 397222 2454
rect 396986 1898 397222 2134
rect 396986 -582 397222 -346
rect 396986 -902 397222 -666
rect 400586 689818 400822 690054
rect 400586 689498 400822 689734
rect 400586 653818 400822 654054
rect 400586 653498 400822 653734
rect 400586 617818 400822 618054
rect 400586 617498 400822 617734
rect 400586 581818 400822 582054
rect 400586 581498 400822 581734
rect 400586 545818 400822 546054
rect 400586 545498 400822 545734
rect 400586 509818 400822 510054
rect 400586 509498 400822 509734
rect 400586 473818 400822 474054
rect 400586 473498 400822 473734
rect 400586 437818 400822 438054
rect 400586 437498 400822 437734
rect 400586 401818 400822 402054
rect 400586 401498 400822 401734
rect 400586 365818 400822 366054
rect 400586 365498 400822 365734
rect 400586 329818 400822 330054
rect 400586 329498 400822 329734
rect 400586 293818 400822 294054
rect 400586 293498 400822 293734
rect 400586 257818 400822 258054
rect 400586 257498 400822 257734
rect 400586 221818 400822 222054
rect 400586 221498 400822 221734
rect 400586 185818 400822 186054
rect 400586 185498 400822 185734
rect 400586 149818 400822 150054
rect 400586 149498 400822 149734
rect 400586 113818 400822 114054
rect 400586 113498 400822 113734
rect 400586 77818 400822 78054
rect 400586 77498 400822 77734
rect 400586 41818 400822 42054
rect 400586 41498 400822 41734
rect 400586 5818 400822 6054
rect 400586 5498 400822 5734
rect 400586 -2422 400822 -2186
rect 400586 -2742 400822 -2506
rect 404186 693418 404422 693654
rect 404186 693098 404422 693334
rect 404186 657418 404422 657654
rect 404186 657098 404422 657334
rect 404186 621418 404422 621654
rect 404186 621098 404422 621334
rect 404186 585418 404422 585654
rect 404186 585098 404422 585334
rect 404186 549418 404422 549654
rect 404186 549098 404422 549334
rect 404186 513418 404422 513654
rect 404186 513098 404422 513334
rect 404186 477418 404422 477654
rect 404186 477098 404422 477334
rect 404186 441418 404422 441654
rect 404186 441098 404422 441334
rect 404186 405418 404422 405654
rect 404186 405098 404422 405334
rect 404186 369418 404422 369654
rect 404186 369098 404422 369334
rect 404186 333418 404422 333654
rect 404186 333098 404422 333334
rect 404186 297418 404422 297654
rect 404186 297098 404422 297334
rect 404186 261418 404422 261654
rect 404186 261098 404422 261334
rect 404186 225418 404422 225654
rect 404186 225098 404422 225334
rect 404186 189418 404422 189654
rect 404186 189098 404422 189334
rect 404186 153418 404422 153654
rect 404186 153098 404422 153334
rect 404186 117418 404422 117654
rect 404186 117098 404422 117334
rect 404186 81418 404422 81654
rect 404186 81098 404422 81334
rect 404186 45418 404422 45654
rect 404186 45098 404422 45334
rect 404186 9418 404422 9654
rect 404186 9098 404422 9334
rect 404186 -4262 404422 -4026
rect 404186 -4582 404422 -4346
rect 425786 711042 426022 711278
rect 425786 710722 426022 710958
rect 422186 709202 422422 709438
rect 422186 708882 422422 709118
rect 418586 707362 418822 707598
rect 418586 707042 418822 707278
rect 407786 697018 408022 697254
rect 407786 696698 408022 696934
rect 407786 661018 408022 661254
rect 407786 660698 408022 660934
rect 407786 625018 408022 625254
rect 407786 624698 408022 624934
rect 407786 589018 408022 589254
rect 407786 588698 408022 588934
rect 407786 553018 408022 553254
rect 407786 552698 408022 552934
rect 407786 517018 408022 517254
rect 407786 516698 408022 516934
rect 407786 481018 408022 481254
rect 407786 480698 408022 480934
rect 407786 445018 408022 445254
rect 407786 444698 408022 444934
rect 407786 409018 408022 409254
rect 407786 408698 408022 408934
rect 407786 373018 408022 373254
rect 407786 372698 408022 372934
rect 407786 337018 408022 337254
rect 407786 336698 408022 336934
rect 407786 301018 408022 301254
rect 407786 300698 408022 300934
rect 407786 265018 408022 265254
rect 407786 264698 408022 264934
rect 407786 229018 408022 229254
rect 407786 228698 408022 228934
rect 407786 193018 408022 193254
rect 407786 192698 408022 192934
rect 407786 157018 408022 157254
rect 407786 156698 408022 156934
rect 407786 121018 408022 121254
rect 407786 120698 408022 120934
rect 407786 85018 408022 85254
rect 407786 84698 408022 84934
rect 407786 49018 408022 49254
rect 407786 48698 408022 48934
rect 407786 13018 408022 13254
rect 407786 12698 408022 12934
rect 389786 -7022 390022 -6786
rect 389786 -7342 390022 -7106
rect 414986 705522 415222 705758
rect 414986 705202 415222 705438
rect 414986 668218 415222 668454
rect 414986 667898 415222 668134
rect 414986 632218 415222 632454
rect 414986 631898 415222 632134
rect 414986 596218 415222 596454
rect 414986 595898 415222 596134
rect 414986 560218 415222 560454
rect 414986 559898 415222 560134
rect 414986 524218 415222 524454
rect 414986 523898 415222 524134
rect 414986 488218 415222 488454
rect 414986 487898 415222 488134
rect 414986 452218 415222 452454
rect 414986 451898 415222 452134
rect 414986 416218 415222 416454
rect 414986 415898 415222 416134
rect 414986 380218 415222 380454
rect 414986 379898 415222 380134
rect 414986 344218 415222 344454
rect 414986 343898 415222 344134
rect 414986 308218 415222 308454
rect 414986 307898 415222 308134
rect 414986 272218 415222 272454
rect 414986 271898 415222 272134
rect 414986 236218 415222 236454
rect 414986 235898 415222 236134
rect 414986 200218 415222 200454
rect 414986 199898 415222 200134
rect 414986 164218 415222 164454
rect 414986 163898 415222 164134
rect 414986 128218 415222 128454
rect 414986 127898 415222 128134
rect 414986 92218 415222 92454
rect 414986 91898 415222 92134
rect 414986 56218 415222 56454
rect 414986 55898 415222 56134
rect 414986 20218 415222 20454
rect 414986 19898 415222 20134
rect 414986 -1502 415222 -1266
rect 414986 -1822 415222 -1586
rect 418586 671818 418822 672054
rect 418586 671498 418822 671734
rect 418586 635818 418822 636054
rect 418586 635498 418822 635734
rect 418586 599818 418822 600054
rect 418586 599498 418822 599734
rect 418586 563818 418822 564054
rect 418586 563498 418822 563734
rect 418586 527818 418822 528054
rect 418586 527498 418822 527734
rect 418586 491818 418822 492054
rect 418586 491498 418822 491734
rect 418586 455818 418822 456054
rect 418586 455498 418822 455734
rect 418586 419818 418822 420054
rect 418586 419498 418822 419734
rect 418586 383818 418822 384054
rect 418586 383498 418822 383734
rect 418586 347818 418822 348054
rect 418586 347498 418822 347734
rect 418586 311818 418822 312054
rect 418586 311498 418822 311734
rect 418586 275818 418822 276054
rect 418586 275498 418822 275734
rect 418586 239818 418822 240054
rect 418586 239498 418822 239734
rect 418586 203818 418822 204054
rect 418586 203498 418822 203734
rect 418586 167818 418822 168054
rect 418586 167498 418822 167734
rect 418586 131818 418822 132054
rect 418586 131498 418822 131734
rect 418586 95818 418822 96054
rect 418586 95498 418822 95734
rect 418586 59818 418822 60054
rect 418586 59498 418822 59734
rect 418586 23818 418822 24054
rect 418586 23498 418822 23734
rect 418586 -3342 418822 -3106
rect 418586 -3662 418822 -3426
rect 422186 675418 422422 675654
rect 422186 675098 422422 675334
rect 422186 639418 422422 639654
rect 422186 639098 422422 639334
rect 422186 603418 422422 603654
rect 422186 603098 422422 603334
rect 422186 567418 422422 567654
rect 422186 567098 422422 567334
rect 422186 531418 422422 531654
rect 422186 531098 422422 531334
rect 422186 495418 422422 495654
rect 422186 495098 422422 495334
rect 422186 459418 422422 459654
rect 422186 459098 422422 459334
rect 422186 423418 422422 423654
rect 422186 423098 422422 423334
rect 422186 387418 422422 387654
rect 422186 387098 422422 387334
rect 422186 351418 422422 351654
rect 422186 351098 422422 351334
rect 422186 315418 422422 315654
rect 422186 315098 422422 315334
rect 422186 279418 422422 279654
rect 422186 279098 422422 279334
rect 422186 243418 422422 243654
rect 422186 243098 422422 243334
rect 422186 207418 422422 207654
rect 422186 207098 422422 207334
rect 422186 171418 422422 171654
rect 422186 171098 422422 171334
rect 422186 135418 422422 135654
rect 422186 135098 422422 135334
rect 422186 99418 422422 99654
rect 422186 99098 422422 99334
rect 422186 63418 422422 63654
rect 422186 63098 422422 63334
rect 422186 27418 422422 27654
rect 422186 27098 422422 27334
rect 422186 -5182 422422 -4946
rect 422186 -5502 422422 -5266
rect 443786 710122 444022 710358
rect 443786 709802 444022 710038
rect 440186 708282 440422 708518
rect 440186 707962 440422 708198
rect 436586 706442 436822 706678
rect 436586 706122 436822 706358
rect 425786 679018 426022 679254
rect 425786 678698 426022 678934
rect 425786 643018 426022 643254
rect 425786 642698 426022 642934
rect 425786 607018 426022 607254
rect 425786 606698 426022 606934
rect 425786 571018 426022 571254
rect 425786 570698 426022 570934
rect 425786 535018 426022 535254
rect 425786 534698 426022 534934
rect 425786 499018 426022 499254
rect 425786 498698 426022 498934
rect 425786 463018 426022 463254
rect 425786 462698 426022 462934
rect 425786 427018 426022 427254
rect 425786 426698 426022 426934
rect 425786 391018 426022 391254
rect 425786 390698 426022 390934
rect 425786 355018 426022 355254
rect 425786 354698 426022 354934
rect 425786 319018 426022 319254
rect 425786 318698 426022 318934
rect 425786 283018 426022 283254
rect 425786 282698 426022 282934
rect 425786 247018 426022 247254
rect 425786 246698 426022 246934
rect 425786 211018 426022 211254
rect 425786 210698 426022 210934
rect 425786 175018 426022 175254
rect 425786 174698 426022 174934
rect 425786 139018 426022 139254
rect 425786 138698 426022 138934
rect 425786 103018 426022 103254
rect 425786 102698 426022 102934
rect 425786 67018 426022 67254
rect 425786 66698 426022 66934
rect 425786 31018 426022 31254
rect 425786 30698 426022 30934
rect 407786 -6102 408022 -5866
rect 407786 -6422 408022 -6186
rect 432986 704602 433222 704838
rect 432986 704282 433222 704518
rect 432986 686218 433222 686454
rect 432986 685898 433222 686134
rect 432986 650218 433222 650454
rect 432986 649898 433222 650134
rect 432986 614218 433222 614454
rect 432986 613898 433222 614134
rect 432986 578218 433222 578454
rect 432986 577898 433222 578134
rect 432986 542218 433222 542454
rect 432986 541898 433222 542134
rect 432986 506218 433222 506454
rect 432986 505898 433222 506134
rect 432986 470218 433222 470454
rect 432986 469898 433222 470134
rect 432986 434218 433222 434454
rect 432986 433898 433222 434134
rect 432986 398218 433222 398454
rect 432986 397898 433222 398134
rect 432986 362218 433222 362454
rect 432986 361898 433222 362134
rect 432986 326218 433222 326454
rect 432986 325898 433222 326134
rect 432986 290218 433222 290454
rect 432986 289898 433222 290134
rect 432986 254218 433222 254454
rect 432986 253898 433222 254134
rect 432986 218218 433222 218454
rect 432986 217898 433222 218134
rect 432986 182218 433222 182454
rect 432986 181898 433222 182134
rect 432986 146218 433222 146454
rect 432986 145898 433222 146134
rect 432986 110218 433222 110454
rect 432986 109898 433222 110134
rect 432986 74218 433222 74454
rect 432986 73898 433222 74134
rect 432986 38218 433222 38454
rect 432986 37898 433222 38134
rect 432986 2218 433222 2454
rect 432986 1898 433222 2134
rect 432986 -582 433222 -346
rect 432986 -902 433222 -666
rect 436586 689818 436822 690054
rect 436586 689498 436822 689734
rect 436586 653818 436822 654054
rect 436586 653498 436822 653734
rect 436586 617818 436822 618054
rect 436586 617498 436822 617734
rect 436586 581818 436822 582054
rect 436586 581498 436822 581734
rect 436586 545818 436822 546054
rect 436586 545498 436822 545734
rect 436586 509818 436822 510054
rect 436586 509498 436822 509734
rect 436586 473818 436822 474054
rect 436586 473498 436822 473734
rect 436586 437818 436822 438054
rect 436586 437498 436822 437734
rect 436586 401818 436822 402054
rect 436586 401498 436822 401734
rect 436586 365818 436822 366054
rect 436586 365498 436822 365734
rect 436586 329818 436822 330054
rect 436586 329498 436822 329734
rect 436586 293818 436822 294054
rect 436586 293498 436822 293734
rect 436586 257818 436822 258054
rect 436586 257498 436822 257734
rect 436586 221818 436822 222054
rect 436586 221498 436822 221734
rect 436586 185818 436822 186054
rect 436586 185498 436822 185734
rect 436586 149818 436822 150054
rect 436586 149498 436822 149734
rect 436586 113818 436822 114054
rect 436586 113498 436822 113734
rect 436586 77818 436822 78054
rect 436586 77498 436822 77734
rect 436586 41818 436822 42054
rect 436586 41498 436822 41734
rect 436586 5818 436822 6054
rect 436586 5498 436822 5734
rect 436586 -2422 436822 -2186
rect 436586 -2742 436822 -2506
rect 440186 693418 440422 693654
rect 440186 693098 440422 693334
rect 440186 657418 440422 657654
rect 440186 657098 440422 657334
rect 440186 621418 440422 621654
rect 440186 621098 440422 621334
rect 440186 585418 440422 585654
rect 440186 585098 440422 585334
rect 440186 549418 440422 549654
rect 440186 549098 440422 549334
rect 440186 513418 440422 513654
rect 440186 513098 440422 513334
rect 440186 477418 440422 477654
rect 440186 477098 440422 477334
rect 440186 441418 440422 441654
rect 440186 441098 440422 441334
rect 440186 405418 440422 405654
rect 440186 405098 440422 405334
rect 440186 369418 440422 369654
rect 440186 369098 440422 369334
rect 440186 333418 440422 333654
rect 440186 333098 440422 333334
rect 440186 297418 440422 297654
rect 440186 297098 440422 297334
rect 440186 261418 440422 261654
rect 440186 261098 440422 261334
rect 440186 225418 440422 225654
rect 440186 225098 440422 225334
rect 440186 189418 440422 189654
rect 440186 189098 440422 189334
rect 440186 153418 440422 153654
rect 440186 153098 440422 153334
rect 440186 117418 440422 117654
rect 440186 117098 440422 117334
rect 440186 81418 440422 81654
rect 440186 81098 440422 81334
rect 440186 45418 440422 45654
rect 440186 45098 440422 45334
rect 440186 9418 440422 9654
rect 440186 9098 440422 9334
rect 440186 -4262 440422 -4026
rect 440186 -4582 440422 -4346
rect 461786 711042 462022 711278
rect 461786 710722 462022 710958
rect 458186 709202 458422 709438
rect 458186 708882 458422 709118
rect 454586 707362 454822 707598
rect 454586 707042 454822 707278
rect 443786 697018 444022 697254
rect 443786 696698 444022 696934
rect 443786 661018 444022 661254
rect 443786 660698 444022 660934
rect 443786 625018 444022 625254
rect 443786 624698 444022 624934
rect 443786 589018 444022 589254
rect 443786 588698 444022 588934
rect 443786 553018 444022 553254
rect 443786 552698 444022 552934
rect 443786 517018 444022 517254
rect 443786 516698 444022 516934
rect 443786 481018 444022 481254
rect 443786 480698 444022 480934
rect 443786 445018 444022 445254
rect 443786 444698 444022 444934
rect 443786 409018 444022 409254
rect 443786 408698 444022 408934
rect 443786 373018 444022 373254
rect 443786 372698 444022 372934
rect 443786 337018 444022 337254
rect 443786 336698 444022 336934
rect 443786 301018 444022 301254
rect 443786 300698 444022 300934
rect 443786 265018 444022 265254
rect 443786 264698 444022 264934
rect 443786 229018 444022 229254
rect 443786 228698 444022 228934
rect 443786 193018 444022 193254
rect 443786 192698 444022 192934
rect 443786 157018 444022 157254
rect 443786 156698 444022 156934
rect 443786 121018 444022 121254
rect 443786 120698 444022 120934
rect 443786 85018 444022 85254
rect 443786 84698 444022 84934
rect 443786 49018 444022 49254
rect 443786 48698 444022 48934
rect 443786 13018 444022 13254
rect 443786 12698 444022 12934
rect 425786 -7022 426022 -6786
rect 425786 -7342 426022 -7106
rect 450986 705522 451222 705758
rect 450986 705202 451222 705438
rect 450986 668218 451222 668454
rect 450986 667898 451222 668134
rect 450986 632218 451222 632454
rect 450986 631898 451222 632134
rect 450986 596218 451222 596454
rect 450986 595898 451222 596134
rect 450986 560218 451222 560454
rect 450986 559898 451222 560134
rect 450986 524218 451222 524454
rect 450986 523898 451222 524134
rect 450986 488218 451222 488454
rect 450986 487898 451222 488134
rect 450986 452218 451222 452454
rect 450986 451898 451222 452134
rect 450986 416218 451222 416454
rect 450986 415898 451222 416134
rect 450986 380218 451222 380454
rect 450986 379898 451222 380134
rect 450986 344218 451222 344454
rect 450986 343898 451222 344134
rect 450986 308218 451222 308454
rect 450986 307898 451222 308134
rect 450986 272218 451222 272454
rect 450986 271898 451222 272134
rect 450986 236218 451222 236454
rect 450986 235898 451222 236134
rect 450986 200218 451222 200454
rect 450986 199898 451222 200134
rect 450986 164218 451222 164454
rect 450986 163898 451222 164134
rect 450986 128218 451222 128454
rect 450986 127898 451222 128134
rect 450986 92218 451222 92454
rect 450986 91898 451222 92134
rect 450986 56218 451222 56454
rect 450986 55898 451222 56134
rect 450986 20218 451222 20454
rect 450986 19898 451222 20134
rect 450986 -1502 451222 -1266
rect 450986 -1822 451222 -1586
rect 454586 671818 454822 672054
rect 454586 671498 454822 671734
rect 454586 635818 454822 636054
rect 454586 635498 454822 635734
rect 454586 599818 454822 600054
rect 454586 599498 454822 599734
rect 454586 563818 454822 564054
rect 454586 563498 454822 563734
rect 454586 527818 454822 528054
rect 454586 527498 454822 527734
rect 454586 491818 454822 492054
rect 454586 491498 454822 491734
rect 454586 455818 454822 456054
rect 454586 455498 454822 455734
rect 454586 419818 454822 420054
rect 454586 419498 454822 419734
rect 454586 383818 454822 384054
rect 454586 383498 454822 383734
rect 454586 347818 454822 348054
rect 454586 347498 454822 347734
rect 454586 311818 454822 312054
rect 454586 311498 454822 311734
rect 454586 275818 454822 276054
rect 454586 275498 454822 275734
rect 454586 239818 454822 240054
rect 454586 239498 454822 239734
rect 454586 203818 454822 204054
rect 454586 203498 454822 203734
rect 454586 167818 454822 168054
rect 454586 167498 454822 167734
rect 454586 131818 454822 132054
rect 454586 131498 454822 131734
rect 454586 95818 454822 96054
rect 454586 95498 454822 95734
rect 454586 59818 454822 60054
rect 454586 59498 454822 59734
rect 454586 23818 454822 24054
rect 454586 23498 454822 23734
rect 454586 -3342 454822 -3106
rect 454586 -3662 454822 -3426
rect 458186 675418 458422 675654
rect 458186 675098 458422 675334
rect 458186 639418 458422 639654
rect 458186 639098 458422 639334
rect 458186 603418 458422 603654
rect 458186 603098 458422 603334
rect 458186 567418 458422 567654
rect 458186 567098 458422 567334
rect 458186 531418 458422 531654
rect 458186 531098 458422 531334
rect 458186 495418 458422 495654
rect 458186 495098 458422 495334
rect 458186 459418 458422 459654
rect 458186 459098 458422 459334
rect 458186 423418 458422 423654
rect 458186 423098 458422 423334
rect 458186 387418 458422 387654
rect 458186 387098 458422 387334
rect 458186 351418 458422 351654
rect 458186 351098 458422 351334
rect 458186 315418 458422 315654
rect 458186 315098 458422 315334
rect 458186 279418 458422 279654
rect 458186 279098 458422 279334
rect 458186 243418 458422 243654
rect 458186 243098 458422 243334
rect 458186 207418 458422 207654
rect 458186 207098 458422 207334
rect 458186 171418 458422 171654
rect 458186 171098 458422 171334
rect 458186 135418 458422 135654
rect 458186 135098 458422 135334
rect 458186 99418 458422 99654
rect 458186 99098 458422 99334
rect 458186 63418 458422 63654
rect 458186 63098 458422 63334
rect 458186 27418 458422 27654
rect 458186 27098 458422 27334
rect 458186 -5182 458422 -4946
rect 458186 -5502 458422 -5266
rect 479786 710122 480022 710358
rect 479786 709802 480022 710038
rect 476186 708282 476422 708518
rect 476186 707962 476422 708198
rect 472586 706442 472822 706678
rect 472586 706122 472822 706358
rect 461786 679018 462022 679254
rect 461786 678698 462022 678934
rect 461786 643018 462022 643254
rect 461786 642698 462022 642934
rect 461786 607018 462022 607254
rect 461786 606698 462022 606934
rect 461786 571018 462022 571254
rect 461786 570698 462022 570934
rect 461786 535018 462022 535254
rect 461786 534698 462022 534934
rect 461786 499018 462022 499254
rect 461786 498698 462022 498934
rect 461786 463018 462022 463254
rect 461786 462698 462022 462934
rect 461786 427018 462022 427254
rect 461786 426698 462022 426934
rect 461786 391018 462022 391254
rect 461786 390698 462022 390934
rect 461786 355018 462022 355254
rect 461786 354698 462022 354934
rect 461786 319018 462022 319254
rect 461786 318698 462022 318934
rect 461786 283018 462022 283254
rect 461786 282698 462022 282934
rect 461786 247018 462022 247254
rect 461786 246698 462022 246934
rect 461786 211018 462022 211254
rect 461786 210698 462022 210934
rect 461786 175018 462022 175254
rect 461786 174698 462022 174934
rect 461786 139018 462022 139254
rect 461786 138698 462022 138934
rect 461786 103018 462022 103254
rect 461786 102698 462022 102934
rect 461786 67018 462022 67254
rect 461786 66698 462022 66934
rect 461786 31018 462022 31254
rect 461786 30698 462022 30934
rect 443786 -6102 444022 -5866
rect 443786 -6422 444022 -6186
rect 468986 704602 469222 704838
rect 468986 704282 469222 704518
rect 468986 686218 469222 686454
rect 468986 685898 469222 686134
rect 468986 650218 469222 650454
rect 468986 649898 469222 650134
rect 468986 614218 469222 614454
rect 468986 613898 469222 614134
rect 468986 578218 469222 578454
rect 468986 577898 469222 578134
rect 468986 542218 469222 542454
rect 468986 541898 469222 542134
rect 468986 506218 469222 506454
rect 468986 505898 469222 506134
rect 468986 470218 469222 470454
rect 468986 469898 469222 470134
rect 468986 434218 469222 434454
rect 468986 433898 469222 434134
rect 468986 398218 469222 398454
rect 468986 397898 469222 398134
rect 468986 362218 469222 362454
rect 468986 361898 469222 362134
rect 468986 326218 469222 326454
rect 468986 325898 469222 326134
rect 468986 290218 469222 290454
rect 468986 289898 469222 290134
rect 468986 254218 469222 254454
rect 468986 253898 469222 254134
rect 468986 218218 469222 218454
rect 468986 217898 469222 218134
rect 468986 182218 469222 182454
rect 468986 181898 469222 182134
rect 468986 146218 469222 146454
rect 468986 145898 469222 146134
rect 468986 110218 469222 110454
rect 468986 109898 469222 110134
rect 468986 74218 469222 74454
rect 468986 73898 469222 74134
rect 468986 38218 469222 38454
rect 468986 37898 469222 38134
rect 468986 2218 469222 2454
rect 468986 1898 469222 2134
rect 468986 -582 469222 -346
rect 468986 -902 469222 -666
rect 472586 689818 472822 690054
rect 472586 689498 472822 689734
rect 472586 653818 472822 654054
rect 472586 653498 472822 653734
rect 472586 617818 472822 618054
rect 472586 617498 472822 617734
rect 472586 581818 472822 582054
rect 472586 581498 472822 581734
rect 472586 545818 472822 546054
rect 472586 545498 472822 545734
rect 472586 509818 472822 510054
rect 472586 509498 472822 509734
rect 472586 473818 472822 474054
rect 472586 473498 472822 473734
rect 472586 437818 472822 438054
rect 472586 437498 472822 437734
rect 472586 401818 472822 402054
rect 472586 401498 472822 401734
rect 472586 365818 472822 366054
rect 472586 365498 472822 365734
rect 472586 329818 472822 330054
rect 472586 329498 472822 329734
rect 472586 293818 472822 294054
rect 472586 293498 472822 293734
rect 472586 257818 472822 258054
rect 472586 257498 472822 257734
rect 472586 221818 472822 222054
rect 472586 221498 472822 221734
rect 472586 185818 472822 186054
rect 472586 185498 472822 185734
rect 472586 149818 472822 150054
rect 472586 149498 472822 149734
rect 472586 113818 472822 114054
rect 472586 113498 472822 113734
rect 472586 77818 472822 78054
rect 472586 77498 472822 77734
rect 472586 41818 472822 42054
rect 472586 41498 472822 41734
rect 472586 5818 472822 6054
rect 472586 5498 472822 5734
rect 472586 -2422 472822 -2186
rect 472586 -2742 472822 -2506
rect 476186 693418 476422 693654
rect 476186 693098 476422 693334
rect 476186 657418 476422 657654
rect 476186 657098 476422 657334
rect 476186 621418 476422 621654
rect 476186 621098 476422 621334
rect 476186 585418 476422 585654
rect 476186 585098 476422 585334
rect 476186 549418 476422 549654
rect 476186 549098 476422 549334
rect 476186 513418 476422 513654
rect 476186 513098 476422 513334
rect 476186 477418 476422 477654
rect 476186 477098 476422 477334
rect 476186 441418 476422 441654
rect 476186 441098 476422 441334
rect 476186 405418 476422 405654
rect 476186 405098 476422 405334
rect 476186 369418 476422 369654
rect 476186 369098 476422 369334
rect 476186 333418 476422 333654
rect 476186 333098 476422 333334
rect 476186 297418 476422 297654
rect 476186 297098 476422 297334
rect 476186 261418 476422 261654
rect 476186 261098 476422 261334
rect 476186 225418 476422 225654
rect 476186 225098 476422 225334
rect 476186 189418 476422 189654
rect 476186 189098 476422 189334
rect 476186 153418 476422 153654
rect 476186 153098 476422 153334
rect 476186 117418 476422 117654
rect 476186 117098 476422 117334
rect 476186 81418 476422 81654
rect 476186 81098 476422 81334
rect 476186 45418 476422 45654
rect 476186 45098 476422 45334
rect 476186 9418 476422 9654
rect 476186 9098 476422 9334
rect 476186 -4262 476422 -4026
rect 476186 -4582 476422 -4346
rect 497786 711042 498022 711278
rect 497786 710722 498022 710958
rect 494186 709202 494422 709438
rect 494186 708882 494422 709118
rect 490586 707362 490822 707598
rect 490586 707042 490822 707278
rect 479786 697018 480022 697254
rect 479786 696698 480022 696934
rect 479786 661018 480022 661254
rect 479786 660698 480022 660934
rect 479786 625018 480022 625254
rect 479786 624698 480022 624934
rect 479786 589018 480022 589254
rect 479786 588698 480022 588934
rect 479786 553018 480022 553254
rect 479786 552698 480022 552934
rect 479786 517018 480022 517254
rect 479786 516698 480022 516934
rect 479786 481018 480022 481254
rect 479786 480698 480022 480934
rect 479786 445018 480022 445254
rect 479786 444698 480022 444934
rect 479786 409018 480022 409254
rect 479786 408698 480022 408934
rect 479786 373018 480022 373254
rect 479786 372698 480022 372934
rect 479786 337018 480022 337254
rect 479786 336698 480022 336934
rect 479786 301018 480022 301254
rect 479786 300698 480022 300934
rect 479786 265018 480022 265254
rect 479786 264698 480022 264934
rect 479786 229018 480022 229254
rect 479786 228698 480022 228934
rect 479786 193018 480022 193254
rect 479786 192698 480022 192934
rect 479786 157018 480022 157254
rect 479786 156698 480022 156934
rect 479786 121018 480022 121254
rect 479786 120698 480022 120934
rect 479786 85018 480022 85254
rect 479786 84698 480022 84934
rect 479786 49018 480022 49254
rect 479786 48698 480022 48934
rect 479786 13018 480022 13254
rect 479786 12698 480022 12934
rect 461786 -7022 462022 -6786
rect 461786 -7342 462022 -7106
rect 486986 705522 487222 705758
rect 486986 705202 487222 705438
rect 486986 668218 487222 668454
rect 486986 667898 487222 668134
rect 486986 632218 487222 632454
rect 486986 631898 487222 632134
rect 486986 596218 487222 596454
rect 486986 595898 487222 596134
rect 486986 560218 487222 560454
rect 486986 559898 487222 560134
rect 486986 524218 487222 524454
rect 486986 523898 487222 524134
rect 486986 488218 487222 488454
rect 486986 487898 487222 488134
rect 486986 452218 487222 452454
rect 486986 451898 487222 452134
rect 486986 416218 487222 416454
rect 486986 415898 487222 416134
rect 486986 380218 487222 380454
rect 486986 379898 487222 380134
rect 486986 344218 487222 344454
rect 486986 343898 487222 344134
rect 486986 308218 487222 308454
rect 486986 307898 487222 308134
rect 486986 272218 487222 272454
rect 486986 271898 487222 272134
rect 486986 236218 487222 236454
rect 486986 235898 487222 236134
rect 486986 200218 487222 200454
rect 486986 199898 487222 200134
rect 486986 164218 487222 164454
rect 486986 163898 487222 164134
rect 486986 128218 487222 128454
rect 486986 127898 487222 128134
rect 486986 92218 487222 92454
rect 486986 91898 487222 92134
rect 486986 56218 487222 56454
rect 486986 55898 487222 56134
rect 486986 20218 487222 20454
rect 486986 19898 487222 20134
rect 486986 -1502 487222 -1266
rect 486986 -1822 487222 -1586
rect 490586 671818 490822 672054
rect 490586 671498 490822 671734
rect 490586 635818 490822 636054
rect 490586 635498 490822 635734
rect 490586 599818 490822 600054
rect 490586 599498 490822 599734
rect 490586 563818 490822 564054
rect 490586 563498 490822 563734
rect 490586 527818 490822 528054
rect 490586 527498 490822 527734
rect 490586 491818 490822 492054
rect 490586 491498 490822 491734
rect 490586 455818 490822 456054
rect 490586 455498 490822 455734
rect 490586 419818 490822 420054
rect 490586 419498 490822 419734
rect 490586 383818 490822 384054
rect 490586 383498 490822 383734
rect 490586 347818 490822 348054
rect 490586 347498 490822 347734
rect 490586 311818 490822 312054
rect 490586 311498 490822 311734
rect 490586 275818 490822 276054
rect 490586 275498 490822 275734
rect 490586 239818 490822 240054
rect 490586 239498 490822 239734
rect 490586 203818 490822 204054
rect 490586 203498 490822 203734
rect 490586 167818 490822 168054
rect 490586 167498 490822 167734
rect 490586 131818 490822 132054
rect 490586 131498 490822 131734
rect 490586 95818 490822 96054
rect 490586 95498 490822 95734
rect 494186 675418 494422 675654
rect 494186 675098 494422 675334
rect 494186 639418 494422 639654
rect 494186 639098 494422 639334
rect 494186 603418 494422 603654
rect 494186 603098 494422 603334
rect 494186 567418 494422 567654
rect 494186 567098 494422 567334
rect 494186 531418 494422 531654
rect 494186 531098 494422 531334
rect 494186 495418 494422 495654
rect 494186 495098 494422 495334
rect 494186 459418 494422 459654
rect 494186 459098 494422 459334
rect 494186 423418 494422 423654
rect 494186 423098 494422 423334
rect 494186 387418 494422 387654
rect 494186 387098 494422 387334
rect 494186 351418 494422 351654
rect 494186 351098 494422 351334
rect 494186 315418 494422 315654
rect 494186 315098 494422 315334
rect 494186 279418 494422 279654
rect 494186 279098 494422 279334
rect 494186 243418 494422 243654
rect 494186 243098 494422 243334
rect 494186 207418 494422 207654
rect 494186 207098 494422 207334
rect 494186 171418 494422 171654
rect 494186 171098 494422 171334
rect 494186 135418 494422 135654
rect 494186 135098 494422 135334
rect 494186 99418 494422 99654
rect 494186 99098 494422 99334
rect 490586 59818 490822 60054
rect 490586 59498 490822 59734
rect 490586 23818 490822 24054
rect 490586 23498 490822 23734
rect 490586 -3342 490822 -3106
rect 490586 -3662 490822 -3426
rect 494186 63418 494422 63654
rect 494186 63098 494422 63334
rect 494186 27418 494422 27654
rect 494186 27098 494422 27334
rect 494186 -5182 494422 -4946
rect 494186 -5502 494422 -5266
rect 515786 710122 516022 710358
rect 515786 709802 516022 710038
rect 512186 708282 512422 708518
rect 512186 707962 512422 708198
rect 508586 706442 508822 706678
rect 508586 706122 508822 706358
rect 497786 679018 498022 679254
rect 497786 678698 498022 678934
rect 497786 643018 498022 643254
rect 497786 642698 498022 642934
rect 497786 607018 498022 607254
rect 497786 606698 498022 606934
rect 497786 571018 498022 571254
rect 497786 570698 498022 570934
rect 497786 535018 498022 535254
rect 497786 534698 498022 534934
rect 497786 499018 498022 499254
rect 497786 498698 498022 498934
rect 497786 463018 498022 463254
rect 497786 462698 498022 462934
rect 497786 427018 498022 427254
rect 497786 426698 498022 426934
rect 497786 391018 498022 391254
rect 497786 390698 498022 390934
rect 497786 355018 498022 355254
rect 497786 354698 498022 354934
rect 497786 319018 498022 319254
rect 497786 318698 498022 318934
rect 497786 283018 498022 283254
rect 497786 282698 498022 282934
rect 497786 247018 498022 247254
rect 497786 246698 498022 246934
rect 497786 211018 498022 211254
rect 497786 210698 498022 210934
rect 497786 175018 498022 175254
rect 497786 174698 498022 174934
rect 497786 139018 498022 139254
rect 497786 138698 498022 138934
rect 497786 103018 498022 103254
rect 497786 102698 498022 102934
rect 497786 67018 498022 67254
rect 497786 66698 498022 66934
rect 497786 31018 498022 31254
rect 497786 30698 498022 30934
rect 479786 -6102 480022 -5866
rect 479786 -6422 480022 -6186
rect 504986 704602 505222 704838
rect 504986 704282 505222 704518
rect 504986 686218 505222 686454
rect 504986 685898 505222 686134
rect 504986 650218 505222 650454
rect 504986 649898 505222 650134
rect 504986 614218 505222 614454
rect 504986 613898 505222 614134
rect 504986 578218 505222 578454
rect 504986 577898 505222 578134
rect 504986 542218 505222 542454
rect 504986 541898 505222 542134
rect 504986 506218 505222 506454
rect 504986 505898 505222 506134
rect 504986 470218 505222 470454
rect 504986 469898 505222 470134
rect 504986 434218 505222 434454
rect 504986 433898 505222 434134
rect 504986 398218 505222 398454
rect 504986 397898 505222 398134
rect 504986 362218 505222 362454
rect 504986 361898 505222 362134
rect 504986 326218 505222 326454
rect 504986 325898 505222 326134
rect 504986 290218 505222 290454
rect 504986 289898 505222 290134
rect 504986 254218 505222 254454
rect 504986 253898 505222 254134
rect 504986 218218 505222 218454
rect 504986 217898 505222 218134
rect 504986 182218 505222 182454
rect 504986 181898 505222 182134
rect 504986 146218 505222 146454
rect 504986 145898 505222 146134
rect 504986 110218 505222 110454
rect 504986 109898 505222 110134
rect 504986 74218 505222 74454
rect 504986 73898 505222 74134
rect 504986 38218 505222 38454
rect 504986 37898 505222 38134
rect 504986 2218 505222 2454
rect 504986 1898 505222 2134
rect 504986 -582 505222 -346
rect 504986 -902 505222 -666
rect 508586 689818 508822 690054
rect 508586 689498 508822 689734
rect 508586 653818 508822 654054
rect 508586 653498 508822 653734
rect 508586 617818 508822 618054
rect 508586 617498 508822 617734
rect 508586 581818 508822 582054
rect 508586 581498 508822 581734
rect 508586 545818 508822 546054
rect 508586 545498 508822 545734
rect 508586 509818 508822 510054
rect 508586 509498 508822 509734
rect 508586 473818 508822 474054
rect 508586 473498 508822 473734
rect 508586 437818 508822 438054
rect 508586 437498 508822 437734
rect 508586 401818 508822 402054
rect 508586 401498 508822 401734
rect 508586 365818 508822 366054
rect 508586 365498 508822 365734
rect 508586 329818 508822 330054
rect 508586 329498 508822 329734
rect 508586 293818 508822 294054
rect 508586 293498 508822 293734
rect 508586 257818 508822 258054
rect 508586 257498 508822 257734
rect 508586 221818 508822 222054
rect 508586 221498 508822 221734
rect 508586 185818 508822 186054
rect 508586 185498 508822 185734
rect 508586 149818 508822 150054
rect 508586 149498 508822 149734
rect 508586 113818 508822 114054
rect 508586 113498 508822 113734
rect 508586 77818 508822 78054
rect 508586 77498 508822 77734
rect 508586 41818 508822 42054
rect 508586 41498 508822 41734
rect 508586 5818 508822 6054
rect 508586 5498 508822 5734
rect 508586 -2422 508822 -2186
rect 508586 -2742 508822 -2506
rect 512186 693418 512422 693654
rect 512186 693098 512422 693334
rect 512186 657418 512422 657654
rect 512186 657098 512422 657334
rect 512186 621418 512422 621654
rect 512186 621098 512422 621334
rect 512186 585418 512422 585654
rect 512186 585098 512422 585334
rect 512186 549418 512422 549654
rect 512186 549098 512422 549334
rect 512186 513418 512422 513654
rect 512186 513098 512422 513334
rect 512186 477418 512422 477654
rect 512186 477098 512422 477334
rect 512186 441418 512422 441654
rect 512186 441098 512422 441334
rect 512186 405418 512422 405654
rect 512186 405098 512422 405334
rect 512186 369418 512422 369654
rect 512186 369098 512422 369334
rect 512186 333418 512422 333654
rect 512186 333098 512422 333334
rect 512186 297418 512422 297654
rect 512186 297098 512422 297334
rect 512186 261418 512422 261654
rect 512186 261098 512422 261334
rect 512186 225418 512422 225654
rect 512186 225098 512422 225334
rect 512186 189418 512422 189654
rect 512186 189098 512422 189334
rect 512186 153418 512422 153654
rect 512186 153098 512422 153334
rect 512186 117418 512422 117654
rect 512186 117098 512422 117334
rect 512186 81418 512422 81654
rect 512186 81098 512422 81334
rect 512186 45418 512422 45654
rect 512186 45098 512422 45334
rect 512186 9418 512422 9654
rect 512186 9098 512422 9334
rect 512186 -4262 512422 -4026
rect 512186 -4582 512422 -4346
rect 533786 711042 534022 711278
rect 533786 710722 534022 710958
rect 530186 709202 530422 709438
rect 530186 708882 530422 709118
rect 526586 707362 526822 707598
rect 526586 707042 526822 707278
rect 515786 697018 516022 697254
rect 515786 696698 516022 696934
rect 515786 661018 516022 661254
rect 515786 660698 516022 660934
rect 515786 625018 516022 625254
rect 515786 624698 516022 624934
rect 515786 589018 516022 589254
rect 515786 588698 516022 588934
rect 515786 553018 516022 553254
rect 515786 552698 516022 552934
rect 515786 517018 516022 517254
rect 515786 516698 516022 516934
rect 515786 481018 516022 481254
rect 515786 480698 516022 480934
rect 515786 445018 516022 445254
rect 515786 444698 516022 444934
rect 515786 409018 516022 409254
rect 515786 408698 516022 408934
rect 515786 373018 516022 373254
rect 515786 372698 516022 372934
rect 515786 337018 516022 337254
rect 515786 336698 516022 336934
rect 515786 301018 516022 301254
rect 515786 300698 516022 300934
rect 515786 265018 516022 265254
rect 515786 264698 516022 264934
rect 515786 229018 516022 229254
rect 515786 228698 516022 228934
rect 515786 193018 516022 193254
rect 515786 192698 516022 192934
rect 515786 157018 516022 157254
rect 515786 156698 516022 156934
rect 515786 121018 516022 121254
rect 515786 120698 516022 120934
rect 515786 85018 516022 85254
rect 515786 84698 516022 84934
rect 515786 49018 516022 49254
rect 515786 48698 516022 48934
rect 515786 13018 516022 13254
rect 515786 12698 516022 12934
rect 497786 -7022 498022 -6786
rect 497786 -7342 498022 -7106
rect 522986 705522 523222 705758
rect 522986 705202 523222 705438
rect 522986 668218 523222 668454
rect 522986 667898 523222 668134
rect 522986 632218 523222 632454
rect 522986 631898 523222 632134
rect 522986 596218 523222 596454
rect 522986 595898 523222 596134
rect 522986 560218 523222 560454
rect 522986 559898 523222 560134
rect 522986 524218 523222 524454
rect 522986 523898 523222 524134
rect 522986 488218 523222 488454
rect 522986 487898 523222 488134
rect 522986 452218 523222 452454
rect 522986 451898 523222 452134
rect 522986 416218 523222 416454
rect 522986 415898 523222 416134
rect 522986 380218 523222 380454
rect 522986 379898 523222 380134
rect 522986 344218 523222 344454
rect 522986 343898 523222 344134
rect 522986 308218 523222 308454
rect 522986 307898 523222 308134
rect 522986 272218 523222 272454
rect 522986 271898 523222 272134
rect 522986 236218 523222 236454
rect 522986 235898 523222 236134
rect 522986 200218 523222 200454
rect 522986 199898 523222 200134
rect 522986 164218 523222 164454
rect 522986 163898 523222 164134
rect 522986 128218 523222 128454
rect 522986 127898 523222 128134
rect 522986 92218 523222 92454
rect 522986 91898 523222 92134
rect 522986 56218 523222 56454
rect 522986 55898 523222 56134
rect 522986 20218 523222 20454
rect 522986 19898 523222 20134
rect 522986 -1502 523222 -1266
rect 522986 -1822 523222 -1586
rect 526586 671818 526822 672054
rect 526586 671498 526822 671734
rect 526586 635818 526822 636054
rect 526586 635498 526822 635734
rect 526586 599818 526822 600054
rect 526586 599498 526822 599734
rect 526586 563818 526822 564054
rect 526586 563498 526822 563734
rect 526586 527818 526822 528054
rect 526586 527498 526822 527734
rect 526586 491818 526822 492054
rect 526586 491498 526822 491734
rect 526586 455818 526822 456054
rect 526586 455498 526822 455734
rect 526586 419818 526822 420054
rect 526586 419498 526822 419734
rect 526586 383818 526822 384054
rect 526586 383498 526822 383734
rect 526586 347818 526822 348054
rect 526586 347498 526822 347734
rect 526586 311818 526822 312054
rect 526586 311498 526822 311734
rect 526586 275818 526822 276054
rect 526586 275498 526822 275734
rect 526586 239818 526822 240054
rect 526586 239498 526822 239734
rect 526586 203818 526822 204054
rect 526586 203498 526822 203734
rect 526586 167818 526822 168054
rect 526586 167498 526822 167734
rect 526586 131818 526822 132054
rect 526586 131498 526822 131734
rect 526586 95818 526822 96054
rect 526586 95498 526822 95734
rect 526586 59818 526822 60054
rect 526586 59498 526822 59734
rect 526586 23818 526822 24054
rect 526586 23498 526822 23734
rect 526586 -3342 526822 -3106
rect 526586 -3662 526822 -3426
rect 530186 675418 530422 675654
rect 530186 675098 530422 675334
rect 530186 639418 530422 639654
rect 530186 639098 530422 639334
rect 530186 603418 530422 603654
rect 530186 603098 530422 603334
rect 530186 567418 530422 567654
rect 530186 567098 530422 567334
rect 530186 531418 530422 531654
rect 530186 531098 530422 531334
rect 530186 495418 530422 495654
rect 530186 495098 530422 495334
rect 530186 459418 530422 459654
rect 530186 459098 530422 459334
rect 530186 423418 530422 423654
rect 530186 423098 530422 423334
rect 530186 387418 530422 387654
rect 530186 387098 530422 387334
rect 530186 351418 530422 351654
rect 530186 351098 530422 351334
rect 530186 315418 530422 315654
rect 530186 315098 530422 315334
rect 530186 279418 530422 279654
rect 530186 279098 530422 279334
rect 530186 243418 530422 243654
rect 530186 243098 530422 243334
rect 530186 207418 530422 207654
rect 530186 207098 530422 207334
rect 530186 171418 530422 171654
rect 530186 171098 530422 171334
rect 530186 135418 530422 135654
rect 530186 135098 530422 135334
rect 530186 99418 530422 99654
rect 530186 99098 530422 99334
rect 530186 63418 530422 63654
rect 530186 63098 530422 63334
rect 530186 27418 530422 27654
rect 530186 27098 530422 27334
rect 530186 -5182 530422 -4946
rect 530186 -5502 530422 -5266
rect 551786 710122 552022 710358
rect 551786 709802 552022 710038
rect 548186 708282 548422 708518
rect 548186 707962 548422 708198
rect 544586 706442 544822 706678
rect 544586 706122 544822 706358
rect 533786 679018 534022 679254
rect 533786 678698 534022 678934
rect 533786 643018 534022 643254
rect 533786 642698 534022 642934
rect 533786 607018 534022 607254
rect 533786 606698 534022 606934
rect 533786 571018 534022 571254
rect 533786 570698 534022 570934
rect 533786 535018 534022 535254
rect 533786 534698 534022 534934
rect 533786 499018 534022 499254
rect 533786 498698 534022 498934
rect 533786 463018 534022 463254
rect 533786 462698 534022 462934
rect 533786 427018 534022 427254
rect 533786 426698 534022 426934
rect 533786 391018 534022 391254
rect 533786 390698 534022 390934
rect 533786 355018 534022 355254
rect 533786 354698 534022 354934
rect 533786 319018 534022 319254
rect 533786 318698 534022 318934
rect 533786 283018 534022 283254
rect 533786 282698 534022 282934
rect 533786 247018 534022 247254
rect 533786 246698 534022 246934
rect 533786 211018 534022 211254
rect 533786 210698 534022 210934
rect 533786 175018 534022 175254
rect 533786 174698 534022 174934
rect 533786 139018 534022 139254
rect 533786 138698 534022 138934
rect 533786 103018 534022 103254
rect 533786 102698 534022 102934
rect 533786 67018 534022 67254
rect 533786 66698 534022 66934
rect 533786 31018 534022 31254
rect 533786 30698 534022 30934
rect 515786 -6102 516022 -5866
rect 515786 -6422 516022 -6186
rect 540986 704602 541222 704838
rect 540986 704282 541222 704518
rect 540986 686218 541222 686454
rect 540986 685898 541222 686134
rect 540986 650218 541222 650454
rect 540986 649898 541222 650134
rect 540986 614218 541222 614454
rect 540986 613898 541222 614134
rect 540986 578218 541222 578454
rect 540986 577898 541222 578134
rect 540986 542218 541222 542454
rect 540986 541898 541222 542134
rect 540986 506218 541222 506454
rect 540986 505898 541222 506134
rect 540986 470218 541222 470454
rect 540986 469898 541222 470134
rect 540986 434218 541222 434454
rect 540986 433898 541222 434134
rect 540986 398218 541222 398454
rect 540986 397898 541222 398134
rect 540986 362218 541222 362454
rect 540986 361898 541222 362134
rect 540986 326218 541222 326454
rect 540986 325898 541222 326134
rect 540986 290218 541222 290454
rect 540986 289898 541222 290134
rect 540986 254218 541222 254454
rect 540986 253898 541222 254134
rect 540986 218218 541222 218454
rect 540986 217898 541222 218134
rect 540986 182218 541222 182454
rect 540986 181898 541222 182134
rect 540986 146218 541222 146454
rect 540986 145898 541222 146134
rect 540986 110218 541222 110454
rect 540986 109898 541222 110134
rect 540986 74218 541222 74454
rect 540986 73898 541222 74134
rect 540986 38218 541222 38454
rect 540986 37898 541222 38134
rect 540986 2218 541222 2454
rect 540986 1898 541222 2134
rect 540986 -582 541222 -346
rect 540986 -902 541222 -666
rect 544586 689818 544822 690054
rect 544586 689498 544822 689734
rect 544586 653818 544822 654054
rect 544586 653498 544822 653734
rect 544586 617818 544822 618054
rect 544586 617498 544822 617734
rect 544586 581818 544822 582054
rect 544586 581498 544822 581734
rect 544586 545818 544822 546054
rect 544586 545498 544822 545734
rect 544586 509818 544822 510054
rect 544586 509498 544822 509734
rect 544586 473818 544822 474054
rect 544586 473498 544822 473734
rect 544586 437818 544822 438054
rect 544586 437498 544822 437734
rect 544586 401818 544822 402054
rect 544586 401498 544822 401734
rect 544586 365818 544822 366054
rect 544586 365498 544822 365734
rect 544586 329818 544822 330054
rect 544586 329498 544822 329734
rect 544586 293818 544822 294054
rect 544586 293498 544822 293734
rect 544586 257818 544822 258054
rect 544586 257498 544822 257734
rect 544586 221818 544822 222054
rect 544586 221498 544822 221734
rect 544586 185818 544822 186054
rect 544586 185498 544822 185734
rect 544586 149818 544822 150054
rect 544586 149498 544822 149734
rect 544586 113818 544822 114054
rect 544586 113498 544822 113734
rect 544586 77818 544822 78054
rect 544586 77498 544822 77734
rect 544586 41818 544822 42054
rect 544586 41498 544822 41734
rect 544586 5818 544822 6054
rect 544586 5498 544822 5734
rect 544586 -2422 544822 -2186
rect 544586 -2742 544822 -2506
rect 548186 693418 548422 693654
rect 548186 693098 548422 693334
rect 548186 657418 548422 657654
rect 548186 657098 548422 657334
rect 548186 621418 548422 621654
rect 548186 621098 548422 621334
rect 548186 585418 548422 585654
rect 548186 585098 548422 585334
rect 548186 549418 548422 549654
rect 548186 549098 548422 549334
rect 548186 513418 548422 513654
rect 548186 513098 548422 513334
rect 548186 477418 548422 477654
rect 548186 477098 548422 477334
rect 548186 441418 548422 441654
rect 548186 441098 548422 441334
rect 548186 405418 548422 405654
rect 548186 405098 548422 405334
rect 548186 369418 548422 369654
rect 548186 369098 548422 369334
rect 548186 333418 548422 333654
rect 548186 333098 548422 333334
rect 548186 297418 548422 297654
rect 548186 297098 548422 297334
rect 548186 261418 548422 261654
rect 548186 261098 548422 261334
rect 548186 225418 548422 225654
rect 548186 225098 548422 225334
rect 548186 189418 548422 189654
rect 548186 189098 548422 189334
rect 548186 153418 548422 153654
rect 548186 153098 548422 153334
rect 548186 117418 548422 117654
rect 548186 117098 548422 117334
rect 548186 81418 548422 81654
rect 548186 81098 548422 81334
rect 548186 45418 548422 45654
rect 548186 45098 548422 45334
rect 548186 9418 548422 9654
rect 548186 9098 548422 9334
rect 548186 -4262 548422 -4026
rect 548186 -4582 548422 -4346
rect 569786 711042 570022 711278
rect 569786 710722 570022 710958
rect 566186 709202 566422 709438
rect 566186 708882 566422 709118
rect 562586 707362 562822 707598
rect 562586 707042 562822 707278
rect 551786 697018 552022 697254
rect 551786 696698 552022 696934
rect 551786 661018 552022 661254
rect 551786 660698 552022 660934
rect 551786 625018 552022 625254
rect 551786 624698 552022 624934
rect 551786 589018 552022 589254
rect 551786 588698 552022 588934
rect 551786 553018 552022 553254
rect 551786 552698 552022 552934
rect 551786 517018 552022 517254
rect 551786 516698 552022 516934
rect 551786 481018 552022 481254
rect 551786 480698 552022 480934
rect 551786 445018 552022 445254
rect 551786 444698 552022 444934
rect 551786 409018 552022 409254
rect 551786 408698 552022 408934
rect 551786 373018 552022 373254
rect 551786 372698 552022 372934
rect 551786 337018 552022 337254
rect 551786 336698 552022 336934
rect 551786 301018 552022 301254
rect 551786 300698 552022 300934
rect 551786 265018 552022 265254
rect 551786 264698 552022 264934
rect 551786 229018 552022 229254
rect 551786 228698 552022 228934
rect 551786 193018 552022 193254
rect 551786 192698 552022 192934
rect 551786 157018 552022 157254
rect 551786 156698 552022 156934
rect 551786 121018 552022 121254
rect 551786 120698 552022 120934
rect 551786 85018 552022 85254
rect 551786 84698 552022 84934
rect 551786 49018 552022 49254
rect 551786 48698 552022 48934
rect 551786 13018 552022 13254
rect 551786 12698 552022 12934
rect 533786 -7022 534022 -6786
rect 533786 -7342 534022 -7106
rect 558986 705522 559222 705758
rect 558986 705202 559222 705438
rect 558986 668218 559222 668454
rect 558986 667898 559222 668134
rect 558986 632218 559222 632454
rect 558986 631898 559222 632134
rect 558986 596218 559222 596454
rect 558986 595898 559222 596134
rect 558986 560218 559222 560454
rect 558986 559898 559222 560134
rect 558986 524218 559222 524454
rect 558986 523898 559222 524134
rect 558986 488218 559222 488454
rect 558986 487898 559222 488134
rect 558986 452218 559222 452454
rect 558986 451898 559222 452134
rect 558986 416218 559222 416454
rect 558986 415898 559222 416134
rect 558986 380218 559222 380454
rect 558986 379898 559222 380134
rect 558986 344218 559222 344454
rect 558986 343898 559222 344134
rect 558986 308218 559222 308454
rect 558986 307898 559222 308134
rect 558986 272218 559222 272454
rect 558986 271898 559222 272134
rect 558986 236218 559222 236454
rect 558986 235898 559222 236134
rect 558986 200218 559222 200454
rect 558986 199898 559222 200134
rect 558986 164218 559222 164454
rect 558986 163898 559222 164134
rect 558986 128218 559222 128454
rect 558986 127898 559222 128134
rect 558986 92218 559222 92454
rect 558986 91898 559222 92134
rect 558986 56218 559222 56454
rect 558986 55898 559222 56134
rect 558986 20218 559222 20454
rect 558986 19898 559222 20134
rect 558986 -1502 559222 -1266
rect 558986 -1822 559222 -1586
rect 562586 671818 562822 672054
rect 562586 671498 562822 671734
rect 562586 635818 562822 636054
rect 562586 635498 562822 635734
rect 562586 599818 562822 600054
rect 562586 599498 562822 599734
rect 562586 563818 562822 564054
rect 562586 563498 562822 563734
rect 562586 527818 562822 528054
rect 562586 527498 562822 527734
rect 562586 491818 562822 492054
rect 562586 491498 562822 491734
rect 562586 455818 562822 456054
rect 562586 455498 562822 455734
rect 562586 419818 562822 420054
rect 562586 419498 562822 419734
rect 562586 383818 562822 384054
rect 562586 383498 562822 383734
rect 562586 347818 562822 348054
rect 562586 347498 562822 347734
rect 562586 311818 562822 312054
rect 562586 311498 562822 311734
rect 562586 275818 562822 276054
rect 562586 275498 562822 275734
rect 562586 239818 562822 240054
rect 562586 239498 562822 239734
rect 562586 203818 562822 204054
rect 562586 203498 562822 203734
rect 562586 167818 562822 168054
rect 562586 167498 562822 167734
rect 562586 131818 562822 132054
rect 562586 131498 562822 131734
rect 562586 95818 562822 96054
rect 562586 95498 562822 95734
rect 562586 59818 562822 60054
rect 562586 59498 562822 59734
rect 562586 23818 562822 24054
rect 562586 23498 562822 23734
rect 562586 -3342 562822 -3106
rect 562586 -3662 562822 -3426
rect 566186 675418 566422 675654
rect 566186 675098 566422 675334
rect 566186 639418 566422 639654
rect 566186 639098 566422 639334
rect 566186 603418 566422 603654
rect 566186 603098 566422 603334
rect 566186 567418 566422 567654
rect 566186 567098 566422 567334
rect 566186 531418 566422 531654
rect 566186 531098 566422 531334
rect 566186 495418 566422 495654
rect 566186 495098 566422 495334
rect 566186 459418 566422 459654
rect 566186 459098 566422 459334
rect 566186 423418 566422 423654
rect 566186 423098 566422 423334
rect 566186 387418 566422 387654
rect 566186 387098 566422 387334
rect 566186 351418 566422 351654
rect 566186 351098 566422 351334
rect 566186 315418 566422 315654
rect 566186 315098 566422 315334
rect 566186 279418 566422 279654
rect 566186 279098 566422 279334
rect 566186 243418 566422 243654
rect 566186 243098 566422 243334
rect 566186 207418 566422 207654
rect 566186 207098 566422 207334
rect 566186 171418 566422 171654
rect 566186 171098 566422 171334
rect 566186 135418 566422 135654
rect 566186 135098 566422 135334
rect 566186 99418 566422 99654
rect 566186 99098 566422 99334
rect 566186 63418 566422 63654
rect 566186 63098 566422 63334
rect 566186 27418 566422 27654
rect 566186 27098 566422 27334
rect 566186 -5182 566422 -4946
rect 566186 -5502 566422 -5266
rect 591942 711042 592178 711278
rect 591942 710722 592178 710958
rect 591022 710122 591258 710358
rect 591022 709802 591258 710038
rect 590102 709202 590338 709438
rect 590102 708882 590338 709118
rect 589182 708282 589418 708518
rect 589182 707962 589418 708198
rect 588262 707362 588498 707598
rect 588262 707042 588498 707278
rect 580586 706442 580822 706678
rect 580586 706122 580822 706358
rect 569786 679018 570022 679254
rect 569786 678698 570022 678934
rect 569786 643018 570022 643254
rect 569786 642698 570022 642934
rect 569786 607018 570022 607254
rect 569786 606698 570022 606934
rect 569786 571018 570022 571254
rect 569786 570698 570022 570934
rect 569786 535018 570022 535254
rect 569786 534698 570022 534934
rect 569786 499018 570022 499254
rect 569786 498698 570022 498934
rect 569786 463018 570022 463254
rect 569786 462698 570022 462934
rect 569786 427018 570022 427254
rect 569786 426698 570022 426934
rect 569786 391018 570022 391254
rect 569786 390698 570022 390934
rect 569786 355018 570022 355254
rect 569786 354698 570022 354934
rect 569786 319018 570022 319254
rect 569786 318698 570022 318934
rect 569786 283018 570022 283254
rect 569786 282698 570022 282934
rect 569786 247018 570022 247254
rect 569786 246698 570022 246934
rect 569786 211018 570022 211254
rect 569786 210698 570022 210934
rect 569786 175018 570022 175254
rect 569786 174698 570022 174934
rect 569786 139018 570022 139254
rect 569786 138698 570022 138934
rect 569786 103018 570022 103254
rect 569786 102698 570022 102934
rect 569786 67018 570022 67254
rect 569786 66698 570022 66934
rect 569786 31018 570022 31254
rect 569786 30698 570022 30934
rect 551786 -6102 552022 -5866
rect 551786 -6422 552022 -6186
rect 576986 704602 577222 704838
rect 576986 704282 577222 704518
rect 576986 686218 577222 686454
rect 576986 685898 577222 686134
rect 576986 650218 577222 650454
rect 576986 649898 577222 650134
rect 576986 614218 577222 614454
rect 576986 613898 577222 614134
rect 576986 578218 577222 578454
rect 576986 577898 577222 578134
rect 576986 542218 577222 542454
rect 576986 541898 577222 542134
rect 576986 506218 577222 506454
rect 576986 505898 577222 506134
rect 576986 470218 577222 470454
rect 576986 469898 577222 470134
rect 576986 434218 577222 434454
rect 576986 433898 577222 434134
rect 576986 398218 577222 398454
rect 576986 397898 577222 398134
rect 576986 362218 577222 362454
rect 576986 361898 577222 362134
rect 576986 326218 577222 326454
rect 576986 325898 577222 326134
rect 576986 290218 577222 290454
rect 576986 289898 577222 290134
rect 576986 254218 577222 254454
rect 576986 253898 577222 254134
rect 576986 218218 577222 218454
rect 576986 217898 577222 218134
rect 576986 182218 577222 182454
rect 576986 181898 577222 182134
rect 576986 146218 577222 146454
rect 576986 145898 577222 146134
rect 576986 110218 577222 110454
rect 576986 109898 577222 110134
rect 576986 74218 577222 74454
rect 576986 73898 577222 74134
rect 576986 38218 577222 38454
rect 576986 37898 577222 38134
rect 576986 2218 577222 2454
rect 576986 1898 577222 2134
rect 576986 -582 577222 -346
rect 576986 -902 577222 -666
rect 587342 706442 587578 706678
rect 587342 706122 587578 706358
rect 586422 705522 586658 705758
rect 586422 705202 586658 705438
rect 580586 689818 580822 690054
rect 580586 689498 580822 689734
rect 580586 653818 580822 654054
rect 580586 653498 580822 653734
rect 580586 617818 580822 618054
rect 580586 617498 580822 617734
rect 580586 581818 580822 582054
rect 580586 581498 580822 581734
rect 580586 545818 580822 546054
rect 580586 545498 580822 545734
rect 580586 509818 580822 510054
rect 580586 509498 580822 509734
rect 580586 473818 580822 474054
rect 580586 473498 580822 473734
rect 580586 437818 580822 438054
rect 580586 437498 580822 437734
rect 580586 401818 580822 402054
rect 580586 401498 580822 401734
rect 580586 365818 580822 366054
rect 580586 365498 580822 365734
rect 580586 329818 580822 330054
rect 580586 329498 580822 329734
rect 580586 293818 580822 294054
rect 580586 293498 580822 293734
rect 580586 257818 580822 258054
rect 580586 257498 580822 257734
rect 580586 221818 580822 222054
rect 580586 221498 580822 221734
rect 580586 185818 580822 186054
rect 580586 185498 580822 185734
rect 580586 149818 580822 150054
rect 580586 149498 580822 149734
rect 580586 113818 580822 114054
rect 580586 113498 580822 113734
rect 580586 77818 580822 78054
rect 580586 77498 580822 77734
rect 580586 41818 580822 42054
rect 580586 41498 580822 41734
rect 580586 5818 580822 6054
rect 580586 5498 580822 5734
rect 585502 704602 585738 704838
rect 585502 704282 585738 704518
rect 585502 686218 585738 686454
rect 585502 685898 585738 686134
rect 585502 650218 585738 650454
rect 585502 649898 585738 650134
rect 585502 614218 585738 614454
rect 585502 613898 585738 614134
rect 585502 578218 585738 578454
rect 585502 577898 585738 578134
rect 585502 542218 585738 542454
rect 585502 541898 585738 542134
rect 585502 506218 585738 506454
rect 585502 505898 585738 506134
rect 585502 470218 585738 470454
rect 585502 469898 585738 470134
rect 585502 434218 585738 434454
rect 585502 433898 585738 434134
rect 585502 398218 585738 398454
rect 585502 397898 585738 398134
rect 585502 362218 585738 362454
rect 585502 361898 585738 362134
rect 585502 326218 585738 326454
rect 585502 325898 585738 326134
rect 585502 290218 585738 290454
rect 585502 289898 585738 290134
rect 585502 254218 585738 254454
rect 585502 253898 585738 254134
rect 585502 218218 585738 218454
rect 585502 217898 585738 218134
rect 585502 182218 585738 182454
rect 585502 181898 585738 182134
rect 585502 146218 585738 146454
rect 585502 145898 585738 146134
rect 585502 110218 585738 110454
rect 585502 109898 585738 110134
rect 585502 74218 585738 74454
rect 585502 73898 585738 74134
rect 585502 38218 585738 38454
rect 585502 37898 585738 38134
rect 585502 2218 585738 2454
rect 585502 1898 585738 2134
rect 585502 -582 585738 -346
rect 585502 -902 585738 -666
rect 586422 668218 586658 668454
rect 586422 667898 586658 668134
rect 586422 632218 586658 632454
rect 586422 631898 586658 632134
rect 586422 596218 586658 596454
rect 586422 595898 586658 596134
rect 586422 560218 586658 560454
rect 586422 559898 586658 560134
rect 586422 524218 586658 524454
rect 586422 523898 586658 524134
rect 586422 488218 586658 488454
rect 586422 487898 586658 488134
rect 586422 452218 586658 452454
rect 586422 451898 586658 452134
rect 586422 416218 586658 416454
rect 586422 415898 586658 416134
rect 586422 380218 586658 380454
rect 586422 379898 586658 380134
rect 586422 344218 586658 344454
rect 586422 343898 586658 344134
rect 586422 308218 586658 308454
rect 586422 307898 586658 308134
rect 586422 272218 586658 272454
rect 586422 271898 586658 272134
rect 586422 236218 586658 236454
rect 586422 235898 586658 236134
rect 586422 200218 586658 200454
rect 586422 199898 586658 200134
rect 586422 164218 586658 164454
rect 586422 163898 586658 164134
rect 586422 128218 586658 128454
rect 586422 127898 586658 128134
rect 586422 92218 586658 92454
rect 586422 91898 586658 92134
rect 586422 56218 586658 56454
rect 586422 55898 586658 56134
rect 586422 20218 586658 20454
rect 586422 19898 586658 20134
rect 586422 -1502 586658 -1266
rect 586422 -1822 586658 -1586
rect 587342 689818 587578 690054
rect 587342 689498 587578 689734
rect 587342 653818 587578 654054
rect 587342 653498 587578 653734
rect 587342 617818 587578 618054
rect 587342 617498 587578 617734
rect 587342 581818 587578 582054
rect 587342 581498 587578 581734
rect 587342 545818 587578 546054
rect 587342 545498 587578 545734
rect 587342 509818 587578 510054
rect 587342 509498 587578 509734
rect 587342 473818 587578 474054
rect 587342 473498 587578 473734
rect 587342 437818 587578 438054
rect 587342 437498 587578 437734
rect 587342 401818 587578 402054
rect 587342 401498 587578 401734
rect 587342 365818 587578 366054
rect 587342 365498 587578 365734
rect 587342 329818 587578 330054
rect 587342 329498 587578 329734
rect 587342 293818 587578 294054
rect 587342 293498 587578 293734
rect 587342 257818 587578 258054
rect 587342 257498 587578 257734
rect 587342 221818 587578 222054
rect 587342 221498 587578 221734
rect 587342 185818 587578 186054
rect 587342 185498 587578 185734
rect 587342 149818 587578 150054
rect 587342 149498 587578 149734
rect 587342 113818 587578 114054
rect 587342 113498 587578 113734
rect 587342 77818 587578 78054
rect 587342 77498 587578 77734
rect 587342 41818 587578 42054
rect 587342 41498 587578 41734
rect 587342 5818 587578 6054
rect 587342 5498 587578 5734
rect 580586 -2422 580822 -2186
rect 580586 -2742 580822 -2506
rect 587342 -2422 587578 -2186
rect 587342 -2742 587578 -2506
rect 588262 671818 588498 672054
rect 588262 671498 588498 671734
rect 588262 635818 588498 636054
rect 588262 635498 588498 635734
rect 588262 599818 588498 600054
rect 588262 599498 588498 599734
rect 588262 563818 588498 564054
rect 588262 563498 588498 563734
rect 588262 527818 588498 528054
rect 588262 527498 588498 527734
rect 588262 491818 588498 492054
rect 588262 491498 588498 491734
rect 588262 455818 588498 456054
rect 588262 455498 588498 455734
rect 588262 419818 588498 420054
rect 588262 419498 588498 419734
rect 588262 383818 588498 384054
rect 588262 383498 588498 383734
rect 588262 347818 588498 348054
rect 588262 347498 588498 347734
rect 588262 311818 588498 312054
rect 588262 311498 588498 311734
rect 588262 275818 588498 276054
rect 588262 275498 588498 275734
rect 588262 239818 588498 240054
rect 588262 239498 588498 239734
rect 588262 203818 588498 204054
rect 588262 203498 588498 203734
rect 588262 167818 588498 168054
rect 588262 167498 588498 167734
rect 588262 131818 588498 132054
rect 588262 131498 588498 131734
rect 588262 95818 588498 96054
rect 588262 95498 588498 95734
rect 588262 59818 588498 60054
rect 588262 59498 588498 59734
rect 588262 23818 588498 24054
rect 588262 23498 588498 23734
rect 588262 -3342 588498 -3106
rect 588262 -3662 588498 -3426
rect 589182 693418 589418 693654
rect 589182 693098 589418 693334
rect 589182 657418 589418 657654
rect 589182 657098 589418 657334
rect 589182 621418 589418 621654
rect 589182 621098 589418 621334
rect 589182 585418 589418 585654
rect 589182 585098 589418 585334
rect 589182 549418 589418 549654
rect 589182 549098 589418 549334
rect 589182 513418 589418 513654
rect 589182 513098 589418 513334
rect 589182 477418 589418 477654
rect 589182 477098 589418 477334
rect 589182 441418 589418 441654
rect 589182 441098 589418 441334
rect 589182 405418 589418 405654
rect 589182 405098 589418 405334
rect 589182 369418 589418 369654
rect 589182 369098 589418 369334
rect 589182 333418 589418 333654
rect 589182 333098 589418 333334
rect 589182 297418 589418 297654
rect 589182 297098 589418 297334
rect 589182 261418 589418 261654
rect 589182 261098 589418 261334
rect 589182 225418 589418 225654
rect 589182 225098 589418 225334
rect 589182 189418 589418 189654
rect 589182 189098 589418 189334
rect 589182 153418 589418 153654
rect 589182 153098 589418 153334
rect 589182 117418 589418 117654
rect 589182 117098 589418 117334
rect 589182 81418 589418 81654
rect 589182 81098 589418 81334
rect 589182 45418 589418 45654
rect 589182 45098 589418 45334
rect 589182 9418 589418 9654
rect 589182 9098 589418 9334
rect 589182 -4262 589418 -4026
rect 589182 -4582 589418 -4346
rect 590102 675418 590338 675654
rect 590102 675098 590338 675334
rect 590102 639418 590338 639654
rect 590102 639098 590338 639334
rect 590102 603418 590338 603654
rect 590102 603098 590338 603334
rect 590102 567418 590338 567654
rect 590102 567098 590338 567334
rect 590102 531418 590338 531654
rect 590102 531098 590338 531334
rect 590102 495418 590338 495654
rect 590102 495098 590338 495334
rect 590102 459418 590338 459654
rect 590102 459098 590338 459334
rect 590102 423418 590338 423654
rect 590102 423098 590338 423334
rect 590102 387418 590338 387654
rect 590102 387098 590338 387334
rect 590102 351418 590338 351654
rect 590102 351098 590338 351334
rect 590102 315418 590338 315654
rect 590102 315098 590338 315334
rect 590102 279418 590338 279654
rect 590102 279098 590338 279334
rect 590102 243418 590338 243654
rect 590102 243098 590338 243334
rect 590102 207418 590338 207654
rect 590102 207098 590338 207334
rect 590102 171418 590338 171654
rect 590102 171098 590338 171334
rect 590102 135418 590338 135654
rect 590102 135098 590338 135334
rect 590102 99418 590338 99654
rect 590102 99098 590338 99334
rect 590102 63418 590338 63654
rect 590102 63098 590338 63334
rect 590102 27418 590338 27654
rect 590102 27098 590338 27334
rect 590102 -5182 590338 -4946
rect 590102 -5502 590338 -5266
rect 591022 697018 591258 697254
rect 591022 696698 591258 696934
rect 591022 661018 591258 661254
rect 591022 660698 591258 660934
rect 591022 625018 591258 625254
rect 591022 624698 591258 624934
rect 591022 589018 591258 589254
rect 591022 588698 591258 588934
rect 591022 553018 591258 553254
rect 591022 552698 591258 552934
rect 591022 517018 591258 517254
rect 591022 516698 591258 516934
rect 591022 481018 591258 481254
rect 591022 480698 591258 480934
rect 591022 445018 591258 445254
rect 591022 444698 591258 444934
rect 591022 409018 591258 409254
rect 591022 408698 591258 408934
rect 591022 373018 591258 373254
rect 591022 372698 591258 372934
rect 591022 337018 591258 337254
rect 591022 336698 591258 336934
rect 591022 301018 591258 301254
rect 591022 300698 591258 300934
rect 591022 265018 591258 265254
rect 591022 264698 591258 264934
rect 591022 229018 591258 229254
rect 591022 228698 591258 228934
rect 591022 193018 591258 193254
rect 591022 192698 591258 192934
rect 591022 157018 591258 157254
rect 591022 156698 591258 156934
rect 591022 121018 591258 121254
rect 591022 120698 591258 120934
rect 591022 85018 591258 85254
rect 591022 84698 591258 84934
rect 591022 49018 591258 49254
rect 591022 48698 591258 48934
rect 591022 13018 591258 13254
rect 591022 12698 591258 12934
rect 591022 -6102 591258 -5866
rect 591022 -6422 591258 -6186
rect 591942 679018 592178 679254
rect 591942 678698 592178 678934
rect 591942 643018 592178 643254
rect 591942 642698 592178 642934
rect 591942 607018 592178 607254
rect 591942 606698 592178 606934
rect 591942 571018 592178 571254
rect 591942 570698 592178 570934
rect 591942 535018 592178 535254
rect 591942 534698 592178 534934
rect 591942 499018 592178 499254
rect 591942 498698 592178 498934
rect 591942 463018 592178 463254
rect 591942 462698 592178 462934
rect 591942 427018 592178 427254
rect 591942 426698 592178 426934
rect 591942 391018 592178 391254
rect 591942 390698 592178 390934
rect 591942 355018 592178 355254
rect 591942 354698 592178 354934
rect 591942 319018 592178 319254
rect 591942 318698 592178 318934
rect 591942 283018 592178 283254
rect 591942 282698 592178 282934
rect 591942 247018 592178 247254
rect 591942 246698 592178 246934
rect 591942 211018 592178 211254
rect 591942 210698 592178 210934
rect 591942 175018 592178 175254
rect 591942 174698 592178 174934
rect 591942 139018 592178 139254
rect 591942 138698 592178 138934
rect 591942 103018 592178 103254
rect 591942 102698 592178 102934
rect 591942 67018 592178 67254
rect 591942 66698 592178 66934
rect 591942 31018 592178 31254
rect 591942 30698 592178 30934
rect 569786 -7022 570022 -6786
rect 569786 -7342 570022 -7106
rect 591942 -7022 592178 -6786
rect 591942 -7342 592178 -7106
<< metal5 >>
rect -8436 711300 -7836 711302
rect 29604 711300 30204 711302
rect 65604 711300 66204 711302
rect 101604 711300 102204 711302
rect 137604 711300 138204 711302
rect 173604 711300 174204 711302
rect 209604 711300 210204 711302
rect 245604 711300 246204 711302
rect 281604 711300 282204 711302
rect 317604 711300 318204 711302
rect 353604 711300 354204 711302
rect 389604 711300 390204 711302
rect 425604 711300 426204 711302
rect 461604 711300 462204 711302
rect 497604 711300 498204 711302
rect 533604 711300 534204 711302
rect 569604 711300 570204 711302
rect 591760 711300 592360 711302
rect -8436 711278 592360 711300
rect -8436 711042 -8254 711278
rect -8018 711042 29786 711278
rect 30022 711042 65786 711278
rect 66022 711042 101786 711278
rect 102022 711042 137786 711278
rect 138022 711042 173786 711278
rect 174022 711042 209786 711278
rect 210022 711042 245786 711278
rect 246022 711042 281786 711278
rect 282022 711042 317786 711278
rect 318022 711042 353786 711278
rect 354022 711042 389786 711278
rect 390022 711042 425786 711278
rect 426022 711042 461786 711278
rect 462022 711042 497786 711278
rect 498022 711042 533786 711278
rect 534022 711042 569786 711278
rect 570022 711042 591942 711278
rect 592178 711042 592360 711278
rect -8436 710958 592360 711042
rect -8436 710722 -8254 710958
rect -8018 710722 29786 710958
rect 30022 710722 65786 710958
rect 66022 710722 101786 710958
rect 102022 710722 137786 710958
rect 138022 710722 173786 710958
rect 174022 710722 209786 710958
rect 210022 710722 245786 710958
rect 246022 710722 281786 710958
rect 282022 710722 317786 710958
rect 318022 710722 353786 710958
rect 354022 710722 389786 710958
rect 390022 710722 425786 710958
rect 426022 710722 461786 710958
rect 462022 710722 497786 710958
rect 498022 710722 533786 710958
rect 534022 710722 569786 710958
rect 570022 710722 591942 710958
rect 592178 710722 592360 710958
rect -8436 710700 592360 710722
rect -8436 710698 -7836 710700
rect 29604 710698 30204 710700
rect 65604 710698 66204 710700
rect 101604 710698 102204 710700
rect 137604 710698 138204 710700
rect 173604 710698 174204 710700
rect 209604 710698 210204 710700
rect 245604 710698 246204 710700
rect 281604 710698 282204 710700
rect 317604 710698 318204 710700
rect 353604 710698 354204 710700
rect 389604 710698 390204 710700
rect 425604 710698 426204 710700
rect 461604 710698 462204 710700
rect 497604 710698 498204 710700
rect 533604 710698 534204 710700
rect 569604 710698 570204 710700
rect 591760 710698 592360 710700
rect -7516 710380 -6916 710382
rect 11604 710380 12204 710382
rect 47604 710380 48204 710382
rect 83604 710380 84204 710382
rect 119604 710380 120204 710382
rect 155604 710380 156204 710382
rect 191604 710380 192204 710382
rect 227604 710380 228204 710382
rect 263604 710380 264204 710382
rect 299604 710380 300204 710382
rect 335604 710380 336204 710382
rect 371604 710380 372204 710382
rect 407604 710380 408204 710382
rect 443604 710380 444204 710382
rect 479604 710380 480204 710382
rect 515604 710380 516204 710382
rect 551604 710380 552204 710382
rect 590840 710380 591440 710382
rect -7516 710358 591440 710380
rect -7516 710122 -7334 710358
rect -7098 710122 11786 710358
rect 12022 710122 47786 710358
rect 48022 710122 83786 710358
rect 84022 710122 119786 710358
rect 120022 710122 155786 710358
rect 156022 710122 191786 710358
rect 192022 710122 227786 710358
rect 228022 710122 263786 710358
rect 264022 710122 299786 710358
rect 300022 710122 335786 710358
rect 336022 710122 371786 710358
rect 372022 710122 407786 710358
rect 408022 710122 443786 710358
rect 444022 710122 479786 710358
rect 480022 710122 515786 710358
rect 516022 710122 551786 710358
rect 552022 710122 591022 710358
rect 591258 710122 591440 710358
rect -7516 710038 591440 710122
rect -7516 709802 -7334 710038
rect -7098 709802 11786 710038
rect 12022 709802 47786 710038
rect 48022 709802 83786 710038
rect 84022 709802 119786 710038
rect 120022 709802 155786 710038
rect 156022 709802 191786 710038
rect 192022 709802 227786 710038
rect 228022 709802 263786 710038
rect 264022 709802 299786 710038
rect 300022 709802 335786 710038
rect 336022 709802 371786 710038
rect 372022 709802 407786 710038
rect 408022 709802 443786 710038
rect 444022 709802 479786 710038
rect 480022 709802 515786 710038
rect 516022 709802 551786 710038
rect 552022 709802 591022 710038
rect 591258 709802 591440 710038
rect -7516 709780 591440 709802
rect -7516 709778 -6916 709780
rect 11604 709778 12204 709780
rect 47604 709778 48204 709780
rect 83604 709778 84204 709780
rect 119604 709778 120204 709780
rect 155604 709778 156204 709780
rect 191604 709778 192204 709780
rect 227604 709778 228204 709780
rect 263604 709778 264204 709780
rect 299604 709778 300204 709780
rect 335604 709778 336204 709780
rect 371604 709778 372204 709780
rect 407604 709778 408204 709780
rect 443604 709778 444204 709780
rect 479604 709778 480204 709780
rect 515604 709778 516204 709780
rect 551604 709778 552204 709780
rect 590840 709778 591440 709780
rect -6596 709460 -5996 709462
rect 26004 709460 26604 709462
rect 62004 709460 62604 709462
rect 98004 709460 98604 709462
rect 134004 709460 134604 709462
rect 170004 709460 170604 709462
rect 206004 709460 206604 709462
rect 242004 709460 242604 709462
rect 278004 709460 278604 709462
rect 314004 709460 314604 709462
rect 350004 709460 350604 709462
rect 386004 709460 386604 709462
rect 422004 709460 422604 709462
rect 458004 709460 458604 709462
rect 494004 709460 494604 709462
rect 530004 709460 530604 709462
rect 566004 709460 566604 709462
rect 589920 709460 590520 709462
rect -6596 709438 590520 709460
rect -6596 709202 -6414 709438
rect -6178 709202 26186 709438
rect 26422 709202 62186 709438
rect 62422 709202 98186 709438
rect 98422 709202 134186 709438
rect 134422 709202 170186 709438
rect 170422 709202 206186 709438
rect 206422 709202 242186 709438
rect 242422 709202 278186 709438
rect 278422 709202 314186 709438
rect 314422 709202 350186 709438
rect 350422 709202 386186 709438
rect 386422 709202 422186 709438
rect 422422 709202 458186 709438
rect 458422 709202 494186 709438
rect 494422 709202 530186 709438
rect 530422 709202 566186 709438
rect 566422 709202 590102 709438
rect 590338 709202 590520 709438
rect -6596 709118 590520 709202
rect -6596 708882 -6414 709118
rect -6178 708882 26186 709118
rect 26422 708882 62186 709118
rect 62422 708882 98186 709118
rect 98422 708882 134186 709118
rect 134422 708882 170186 709118
rect 170422 708882 206186 709118
rect 206422 708882 242186 709118
rect 242422 708882 278186 709118
rect 278422 708882 314186 709118
rect 314422 708882 350186 709118
rect 350422 708882 386186 709118
rect 386422 708882 422186 709118
rect 422422 708882 458186 709118
rect 458422 708882 494186 709118
rect 494422 708882 530186 709118
rect 530422 708882 566186 709118
rect 566422 708882 590102 709118
rect 590338 708882 590520 709118
rect -6596 708860 590520 708882
rect -6596 708858 -5996 708860
rect 26004 708858 26604 708860
rect 62004 708858 62604 708860
rect 98004 708858 98604 708860
rect 134004 708858 134604 708860
rect 170004 708858 170604 708860
rect 206004 708858 206604 708860
rect 242004 708858 242604 708860
rect 278004 708858 278604 708860
rect 314004 708858 314604 708860
rect 350004 708858 350604 708860
rect 386004 708858 386604 708860
rect 422004 708858 422604 708860
rect 458004 708858 458604 708860
rect 494004 708858 494604 708860
rect 530004 708858 530604 708860
rect 566004 708858 566604 708860
rect 589920 708858 590520 708860
rect -5676 708540 -5076 708542
rect 8004 708540 8604 708542
rect 44004 708540 44604 708542
rect 80004 708540 80604 708542
rect 116004 708540 116604 708542
rect 152004 708540 152604 708542
rect 188004 708540 188604 708542
rect 224004 708540 224604 708542
rect 260004 708540 260604 708542
rect 296004 708540 296604 708542
rect 332004 708540 332604 708542
rect 368004 708540 368604 708542
rect 404004 708540 404604 708542
rect 440004 708540 440604 708542
rect 476004 708540 476604 708542
rect 512004 708540 512604 708542
rect 548004 708540 548604 708542
rect 589000 708540 589600 708542
rect -5676 708518 589600 708540
rect -5676 708282 -5494 708518
rect -5258 708282 8186 708518
rect 8422 708282 44186 708518
rect 44422 708282 80186 708518
rect 80422 708282 116186 708518
rect 116422 708282 152186 708518
rect 152422 708282 188186 708518
rect 188422 708282 224186 708518
rect 224422 708282 260186 708518
rect 260422 708282 296186 708518
rect 296422 708282 332186 708518
rect 332422 708282 368186 708518
rect 368422 708282 404186 708518
rect 404422 708282 440186 708518
rect 440422 708282 476186 708518
rect 476422 708282 512186 708518
rect 512422 708282 548186 708518
rect 548422 708282 589182 708518
rect 589418 708282 589600 708518
rect -5676 708198 589600 708282
rect -5676 707962 -5494 708198
rect -5258 707962 8186 708198
rect 8422 707962 44186 708198
rect 44422 707962 80186 708198
rect 80422 707962 116186 708198
rect 116422 707962 152186 708198
rect 152422 707962 188186 708198
rect 188422 707962 224186 708198
rect 224422 707962 260186 708198
rect 260422 707962 296186 708198
rect 296422 707962 332186 708198
rect 332422 707962 368186 708198
rect 368422 707962 404186 708198
rect 404422 707962 440186 708198
rect 440422 707962 476186 708198
rect 476422 707962 512186 708198
rect 512422 707962 548186 708198
rect 548422 707962 589182 708198
rect 589418 707962 589600 708198
rect -5676 707940 589600 707962
rect -5676 707938 -5076 707940
rect 8004 707938 8604 707940
rect 44004 707938 44604 707940
rect 80004 707938 80604 707940
rect 116004 707938 116604 707940
rect 152004 707938 152604 707940
rect 188004 707938 188604 707940
rect 224004 707938 224604 707940
rect 260004 707938 260604 707940
rect 296004 707938 296604 707940
rect 332004 707938 332604 707940
rect 368004 707938 368604 707940
rect 404004 707938 404604 707940
rect 440004 707938 440604 707940
rect 476004 707938 476604 707940
rect 512004 707938 512604 707940
rect 548004 707938 548604 707940
rect 589000 707938 589600 707940
rect -4756 707620 -4156 707622
rect 22404 707620 23004 707622
rect 58404 707620 59004 707622
rect 94404 707620 95004 707622
rect 130404 707620 131004 707622
rect 166404 707620 167004 707622
rect 202404 707620 203004 707622
rect 238404 707620 239004 707622
rect 274404 707620 275004 707622
rect 310404 707620 311004 707622
rect 346404 707620 347004 707622
rect 382404 707620 383004 707622
rect 418404 707620 419004 707622
rect 454404 707620 455004 707622
rect 490404 707620 491004 707622
rect 526404 707620 527004 707622
rect 562404 707620 563004 707622
rect 588080 707620 588680 707622
rect -4756 707598 588680 707620
rect -4756 707362 -4574 707598
rect -4338 707362 22586 707598
rect 22822 707362 58586 707598
rect 58822 707362 94586 707598
rect 94822 707362 130586 707598
rect 130822 707362 166586 707598
rect 166822 707362 202586 707598
rect 202822 707362 238586 707598
rect 238822 707362 274586 707598
rect 274822 707362 310586 707598
rect 310822 707362 346586 707598
rect 346822 707362 382586 707598
rect 382822 707362 418586 707598
rect 418822 707362 454586 707598
rect 454822 707362 490586 707598
rect 490822 707362 526586 707598
rect 526822 707362 562586 707598
rect 562822 707362 588262 707598
rect 588498 707362 588680 707598
rect -4756 707278 588680 707362
rect -4756 707042 -4574 707278
rect -4338 707042 22586 707278
rect 22822 707042 58586 707278
rect 58822 707042 94586 707278
rect 94822 707042 130586 707278
rect 130822 707042 166586 707278
rect 166822 707042 202586 707278
rect 202822 707042 238586 707278
rect 238822 707042 274586 707278
rect 274822 707042 310586 707278
rect 310822 707042 346586 707278
rect 346822 707042 382586 707278
rect 382822 707042 418586 707278
rect 418822 707042 454586 707278
rect 454822 707042 490586 707278
rect 490822 707042 526586 707278
rect 526822 707042 562586 707278
rect 562822 707042 588262 707278
rect 588498 707042 588680 707278
rect -4756 707020 588680 707042
rect -4756 707018 -4156 707020
rect 22404 707018 23004 707020
rect 58404 707018 59004 707020
rect 94404 707018 95004 707020
rect 130404 707018 131004 707020
rect 166404 707018 167004 707020
rect 202404 707018 203004 707020
rect 238404 707018 239004 707020
rect 274404 707018 275004 707020
rect 310404 707018 311004 707020
rect 346404 707018 347004 707020
rect 382404 707018 383004 707020
rect 418404 707018 419004 707020
rect 454404 707018 455004 707020
rect 490404 707018 491004 707020
rect 526404 707018 527004 707020
rect 562404 707018 563004 707020
rect 588080 707018 588680 707020
rect -3836 706700 -3236 706702
rect 4404 706700 5004 706702
rect 40404 706700 41004 706702
rect 76404 706700 77004 706702
rect 112404 706700 113004 706702
rect 148404 706700 149004 706702
rect 184404 706700 185004 706702
rect 220404 706700 221004 706702
rect 256404 706700 257004 706702
rect 292404 706700 293004 706702
rect 328404 706700 329004 706702
rect 364404 706700 365004 706702
rect 400404 706700 401004 706702
rect 436404 706700 437004 706702
rect 472404 706700 473004 706702
rect 508404 706700 509004 706702
rect 544404 706700 545004 706702
rect 580404 706700 581004 706702
rect 587160 706700 587760 706702
rect -3836 706678 587760 706700
rect -3836 706442 -3654 706678
rect -3418 706442 4586 706678
rect 4822 706442 40586 706678
rect 40822 706442 76586 706678
rect 76822 706442 112586 706678
rect 112822 706442 148586 706678
rect 148822 706442 184586 706678
rect 184822 706442 220586 706678
rect 220822 706442 256586 706678
rect 256822 706442 292586 706678
rect 292822 706442 328586 706678
rect 328822 706442 364586 706678
rect 364822 706442 400586 706678
rect 400822 706442 436586 706678
rect 436822 706442 472586 706678
rect 472822 706442 508586 706678
rect 508822 706442 544586 706678
rect 544822 706442 580586 706678
rect 580822 706442 587342 706678
rect 587578 706442 587760 706678
rect -3836 706358 587760 706442
rect -3836 706122 -3654 706358
rect -3418 706122 4586 706358
rect 4822 706122 40586 706358
rect 40822 706122 76586 706358
rect 76822 706122 112586 706358
rect 112822 706122 148586 706358
rect 148822 706122 184586 706358
rect 184822 706122 220586 706358
rect 220822 706122 256586 706358
rect 256822 706122 292586 706358
rect 292822 706122 328586 706358
rect 328822 706122 364586 706358
rect 364822 706122 400586 706358
rect 400822 706122 436586 706358
rect 436822 706122 472586 706358
rect 472822 706122 508586 706358
rect 508822 706122 544586 706358
rect 544822 706122 580586 706358
rect 580822 706122 587342 706358
rect 587578 706122 587760 706358
rect -3836 706100 587760 706122
rect -3836 706098 -3236 706100
rect 4404 706098 5004 706100
rect 40404 706098 41004 706100
rect 76404 706098 77004 706100
rect 112404 706098 113004 706100
rect 148404 706098 149004 706100
rect 184404 706098 185004 706100
rect 220404 706098 221004 706100
rect 256404 706098 257004 706100
rect 292404 706098 293004 706100
rect 328404 706098 329004 706100
rect 364404 706098 365004 706100
rect 400404 706098 401004 706100
rect 436404 706098 437004 706100
rect 472404 706098 473004 706100
rect 508404 706098 509004 706100
rect 544404 706098 545004 706100
rect 580404 706098 581004 706100
rect 587160 706098 587760 706100
rect -2916 705780 -2316 705782
rect 18804 705780 19404 705782
rect 54804 705780 55404 705782
rect 90804 705780 91404 705782
rect 126804 705780 127404 705782
rect 162804 705780 163404 705782
rect 198804 705780 199404 705782
rect 234804 705780 235404 705782
rect 270804 705780 271404 705782
rect 306804 705780 307404 705782
rect 342804 705780 343404 705782
rect 378804 705780 379404 705782
rect 414804 705780 415404 705782
rect 450804 705780 451404 705782
rect 486804 705780 487404 705782
rect 522804 705780 523404 705782
rect 558804 705780 559404 705782
rect 586240 705780 586840 705782
rect -2916 705758 586840 705780
rect -2916 705522 -2734 705758
rect -2498 705522 18986 705758
rect 19222 705522 54986 705758
rect 55222 705522 90986 705758
rect 91222 705522 126986 705758
rect 127222 705522 162986 705758
rect 163222 705522 198986 705758
rect 199222 705522 234986 705758
rect 235222 705522 270986 705758
rect 271222 705522 306986 705758
rect 307222 705522 342986 705758
rect 343222 705522 378986 705758
rect 379222 705522 414986 705758
rect 415222 705522 450986 705758
rect 451222 705522 486986 705758
rect 487222 705522 522986 705758
rect 523222 705522 558986 705758
rect 559222 705522 586422 705758
rect 586658 705522 586840 705758
rect -2916 705438 586840 705522
rect -2916 705202 -2734 705438
rect -2498 705202 18986 705438
rect 19222 705202 54986 705438
rect 55222 705202 90986 705438
rect 91222 705202 126986 705438
rect 127222 705202 162986 705438
rect 163222 705202 198986 705438
rect 199222 705202 234986 705438
rect 235222 705202 270986 705438
rect 271222 705202 306986 705438
rect 307222 705202 342986 705438
rect 343222 705202 378986 705438
rect 379222 705202 414986 705438
rect 415222 705202 450986 705438
rect 451222 705202 486986 705438
rect 487222 705202 522986 705438
rect 523222 705202 558986 705438
rect 559222 705202 586422 705438
rect 586658 705202 586840 705438
rect -2916 705180 586840 705202
rect -2916 705178 -2316 705180
rect 18804 705178 19404 705180
rect 54804 705178 55404 705180
rect 90804 705178 91404 705180
rect 126804 705178 127404 705180
rect 162804 705178 163404 705180
rect 198804 705178 199404 705180
rect 234804 705178 235404 705180
rect 270804 705178 271404 705180
rect 306804 705178 307404 705180
rect 342804 705178 343404 705180
rect 378804 705178 379404 705180
rect 414804 705178 415404 705180
rect 450804 705178 451404 705180
rect 486804 705178 487404 705180
rect 522804 705178 523404 705180
rect 558804 705178 559404 705180
rect 586240 705178 586840 705180
rect -1996 704860 -1396 704862
rect 804 704860 1404 704862
rect 36804 704860 37404 704862
rect 72804 704860 73404 704862
rect 108804 704860 109404 704862
rect 144804 704860 145404 704862
rect 180804 704860 181404 704862
rect 216804 704860 217404 704862
rect 252804 704860 253404 704862
rect 288804 704860 289404 704862
rect 324804 704860 325404 704862
rect 360804 704860 361404 704862
rect 396804 704860 397404 704862
rect 432804 704860 433404 704862
rect 468804 704860 469404 704862
rect 504804 704860 505404 704862
rect 540804 704860 541404 704862
rect 576804 704860 577404 704862
rect 585320 704860 585920 704862
rect -1996 704838 585920 704860
rect -1996 704602 -1814 704838
rect -1578 704602 986 704838
rect 1222 704602 36986 704838
rect 37222 704602 72986 704838
rect 73222 704602 108986 704838
rect 109222 704602 144986 704838
rect 145222 704602 180986 704838
rect 181222 704602 216986 704838
rect 217222 704602 252986 704838
rect 253222 704602 288986 704838
rect 289222 704602 324986 704838
rect 325222 704602 360986 704838
rect 361222 704602 396986 704838
rect 397222 704602 432986 704838
rect 433222 704602 468986 704838
rect 469222 704602 504986 704838
rect 505222 704602 540986 704838
rect 541222 704602 576986 704838
rect 577222 704602 585502 704838
rect 585738 704602 585920 704838
rect -1996 704518 585920 704602
rect -1996 704282 -1814 704518
rect -1578 704282 986 704518
rect 1222 704282 36986 704518
rect 37222 704282 72986 704518
rect 73222 704282 108986 704518
rect 109222 704282 144986 704518
rect 145222 704282 180986 704518
rect 181222 704282 216986 704518
rect 217222 704282 252986 704518
rect 253222 704282 288986 704518
rect 289222 704282 324986 704518
rect 325222 704282 360986 704518
rect 361222 704282 396986 704518
rect 397222 704282 432986 704518
rect 433222 704282 468986 704518
rect 469222 704282 504986 704518
rect 505222 704282 540986 704518
rect 541222 704282 576986 704518
rect 577222 704282 585502 704518
rect 585738 704282 585920 704518
rect -1996 704260 585920 704282
rect -1996 704258 -1396 704260
rect 804 704258 1404 704260
rect 36804 704258 37404 704260
rect 72804 704258 73404 704260
rect 108804 704258 109404 704260
rect 144804 704258 145404 704260
rect 180804 704258 181404 704260
rect 216804 704258 217404 704260
rect 252804 704258 253404 704260
rect 288804 704258 289404 704260
rect 324804 704258 325404 704260
rect 360804 704258 361404 704260
rect 396804 704258 397404 704260
rect 432804 704258 433404 704260
rect 468804 704258 469404 704260
rect 504804 704258 505404 704260
rect 540804 704258 541404 704260
rect 576804 704258 577404 704260
rect 585320 704258 585920 704260
rect -7516 697276 -6916 697278
rect 11604 697276 12204 697278
rect 47604 697276 48204 697278
rect 83604 697276 84204 697278
rect 119604 697276 120204 697278
rect 155604 697276 156204 697278
rect 191604 697276 192204 697278
rect 227604 697276 228204 697278
rect 263604 697276 264204 697278
rect 299604 697276 300204 697278
rect 335604 697276 336204 697278
rect 371604 697276 372204 697278
rect 407604 697276 408204 697278
rect 443604 697276 444204 697278
rect 479604 697276 480204 697278
rect 515604 697276 516204 697278
rect 551604 697276 552204 697278
rect 590840 697276 591440 697278
rect -8436 697254 592360 697276
rect -8436 697018 -7334 697254
rect -7098 697018 11786 697254
rect 12022 697018 47786 697254
rect 48022 697018 83786 697254
rect 84022 697018 119786 697254
rect 120022 697018 155786 697254
rect 156022 697018 191786 697254
rect 192022 697018 227786 697254
rect 228022 697018 263786 697254
rect 264022 697018 299786 697254
rect 300022 697018 335786 697254
rect 336022 697018 371786 697254
rect 372022 697018 407786 697254
rect 408022 697018 443786 697254
rect 444022 697018 479786 697254
rect 480022 697018 515786 697254
rect 516022 697018 551786 697254
rect 552022 697018 591022 697254
rect 591258 697018 592360 697254
rect -8436 696934 592360 697018
rect -8436 696698 -7334 696934
rect -7098 696698 11786 696934
rect 12022 696698 47786 696934
rect 48022 696698 83786 696934
rect 84022 696698 119786 696934
rect 120022 696698 155786 696934
rect 156022 696698 191786 696934
rect 192022 696698 227786 696934
rect 228022 696698 263786 696934
rect 264022 696698 299786 696934
rect 300022 696698 335786 696934
rect 336022 696698 371786 696934
rect 372022 696698 407786 696934
rect 408022 696698 443786 696934
rect 444022 696698 479786 696934
rect 480022 696698 515786 696934
rect 516022 696698 551786 696934
rect 552022 696698 591022 696934
rect 591258 696698 592360 696934
rect -8436 696676 592360 696698
rect -7516 696674 -6916 696676
rect 11604 696674 12204 696676
rect 47604 696674 48204 696676
rect 83604 696674 84204 696676
rect 119604 696674 120204 696676
rect 155604 696674 156204 696676
rect 191604 696674 192204 696676
rect 227604 696674 228204 696676
rect 263604 696674 264204 696676
rect 299604 696674 300204 696676
rect 335604 696674 336204 696676
rect 371604 696674 372204 696676
rect 407604 696674 408204 696676
rect 443604 696674 444204 696676
rect 479604 696674 480204 696676
rect 515604 696674 516204 696676
rect 551604 696674 552204 696676
rect 590840 696674 591440 696676
rect -5676 693676 -5076 693678
rect 8004 693676 8604 693678
rect 44004 693676 44604 693678
rect 80004 693676 80604 693678
rect 116004 693676 116604 693678
rect 152004 693676 152604 693678
rect 188004 693676 188604 693678
rect 224004 693676 224604 693678
rect 260004 693676 260604 693678
rect 296004 693676 296604 693678
rect 332004 693676 332604 693678
rect 368004 693676 368604 693678
rect 404004 693676 404604 693678
rect 440004 693676 440604 693678
rect 476004 693676 476604 693678
rect 512004 693676 512604 693678
rect 548004 693676 548604 693678
rect 589000 693676 589600 693678
rect -6596 693654 590520 693676
rect -6596 693418 -5494 693654
rect -5258 693418 8186 693654
rect 8422 693418 44186 693654
rect 44422 693418 80186 693654
rect 80422 693418 116186 693654
rect 116422 693418 152186 693654
rect 152422 693418 188186 693654
rect 188422 693418 224186 693654
rect 224422 693418 260186 693654
rect 260422 693418 296186 693654
rect 296422 693418 332186 693654
rect 332422 693418 368186 693654
rect 368422 693418 404186 693654
rect 404422 693418 440186 693654
rect 440422 693418 476186 693654
rect 476422 693418 512186 693654
rect 512422 693418 548186 693654
rect 548422 693418 589182 693654
rect 589418 693418 590520 693654
rect -6596 693334 590520 693418
rect -6596 693098 -5494 693334
rect -5258 693098 8186 693334
rect 8422 693098 44186 693334
rect 44422 693098 80186 693334
rect 80422 693098 116186 693334
rect 116422 693098 152186 693334
rect 152422 693098 188186 693334
rect 188422 693098 224186 693334
rect 224422 693098 260186 693334
rect 260422 693098 296186 693334
rect 296422 693098 332186 693334
rect 332422 693098 368186 693334
rect 368422 693098 404186 693334
rect 404422 693098 440186 693334
rect 440422 693098 476186 693334
rect 476422 693098 512186 693334
rect 512422 693098 548186 693334
rect 548422 693098 589182 693334
rect 589418 693098 590520 693334
rect -6596 693076 590520 693098
rect -5676 693074 -5076 693076
rect 8004 693074 8604 693076
rect 44004 693074 44604 693076
rect 80004 693074 80604 693076
rect 116004 693074 116604 693076
rect 152004 693074 152604 693076
rect 188004 693074 188604 693076
rect 224004 693074 224604 693076
rect 260004 693074 260604 693076
rect 296004 693074 296604 693076
rect 332004 693074 332604 693076
rect 368004 693074 368604 693076
rect 404004 693074 404604 693076
rect 440004 693074 440604 693076
rect 476004 693074 476604 693076
rect 512004 693074 512604 693076
rect 548004 693074 548604 693076
rect 589000 693074 589600 693076
rect -3836 690076 -3236 690078
rect 4404 690076 5004 690078
rect 40404 690076 41004 690078
rect 76404 690076 77004 690078
rect 112404 690076 113004 690078
rect 148404 690076 149004 690078
rect 184404 690076 185004 690078
rect 220404 690076 221004 690078
rect 256404 690076 257004 690078
rect 292404 690076 293004 690078
rect 328404 690076 329004 690078
rect 364404 690076 365004 690078
rect 400404 690076 401004 690078
rect 436404 690076 437004 690078
rect 472404 690076 473004 690078
rect 508404 690076 509004 690078
rect 544404 690076 545004 690078
rect 580404 690076 581004 690078
rect 587160 690076 587760 690078
rect -4756 690054 588680 690076
rect -4756 689818 -3654 690054
rect -3418 689818 4586 690054
rect 4822 689818 40586 690054
rect 40822 689818 76586 690054
rect 76822 689818 112586 690054
rect 112822 689818 148586 690054
rect 148822 689818 184586 690054
rect 184822 689818 220586 690054
rect 220822 689818 256586 690054
rect 256822 689818 292586 690054
rect 292822 689818 328586 690054
rect 328822 689818 364586 690054
rect 364822 689818 400586 690054
rect 400822 689818 436586 690054
rect 436822 689818 472586 690054
rect 472822 689818 508586 690054
rect 508822 689818 544586 690054
rect 544822 689818 580586 690054
rect 580822 689818 587342 690054
rect 587578 689818 588680 690054
rect -4756 689734 588680 689818
rect -4756 689498 -3654 689734
rect -3418 689498 4586 689734
rect 4822 689498 40586 689734
rect 40822 689498 76586 689734
rect 76822 689498 112586 689734
rect 112822 689498 148586 689734
rect 148822 689498 184586 689734
rect 184822 689498 220586 689734
rect 220822 689498 256586 689734
rect 256822 689498 292586 689734
rect 292822 689498 328586 689734
rect 328822 689498 364586 689734
rect 364822 689498 400586 689734
rect 400822 689498 436586 689734
rect 436822 689498 472586 689734
rect 472822 689498 508586 689734
rect 508822 689498 544586 689734
rect 544822 689498 580586 689734
rect 580822 689498 587342 689734
rect 587578 689498 588680 689734
rect -4756 689476 588680 689498
rect -3836 689474 -3236 689476
rect 4404 689474 5004 689476
rect 40404 689474 41004 689476
rect 76404 689474 77004 689476
rect 112404 689474 113004 689476
rect 148404 689474 149004 689476
rect 184404 689474 185004 689476
rect 220404 689474 221004 689476
rect 256404 689474 257004 689476
rect 292404 689474 293004 689476
rect 328404 689474 329004 689476
rect 364404 689474 365004 689476
rect 400404 689474 401004 689476
rect 436404 689474 437004 689476
rect 472404 689474 473004 689476
rect 508404 689474 509004 689476
rect 544404 689474 545004 689476
rect 580404 689474 581004 689476
rect 587160 689474 587760 689476
rect -1996 686476 -1396 686478
rect 804 686476 1404 686478
rect 36804 686476 37404 686478
rect 72804 686476 73404 686478
rect 108804 686476 109404 686478
rect 144804 686476 145404 686478
rect 180804 686476 181404 686478
rect 216804 686476 217404 686478
rect 252804 686476 253404 686478
rect 288804 686476 289404 686478
rect 324804 686476 325404 686478
rect 360804 686476 361404 686478
rect 396804 686476 397404 686478
rect 432804 686476 433404 686478
rect 468804 686476 469404 686478
rect 504804 686476 505404 686478
rect 540804 686476 541404 686478
rect 576804 686476 577404 686478
rect 585320 686476 585920 686478
rect -2916 686454 586840 686476
rect -2916 686218 -1814 686454
rect -1578 686218 986 686454
rect 1222 686218 36986 686454
rect 37222 686218 72986 686454
rect 73222 686218 108986 686454
rect 109222 686218 144986 686454
rect 145222 686218 180986 686454
rect 181222 686218 216986 686454
rect 217222 686218 252986 686454
rect 253222 686218 288986 686454
rect 289222 686218 324986 686454
rect 325222 686218 360986 686454
rect 361222 686218 396986 686454
rect 397222 686218 432986 686454
rect 433222 686218 468986 686454
rect 469222 686218 504986 686454
rect 505222 686218 540986 686454
rect 541222 686218 576986 686454
rect 577222 686218 585502 686454
rect 585738 686218 586840 686454
rect -2916 686134 586840 686218
rect -2916 685898 -1814 686134
rect -1578 685898 986 686134
rect 1222 685898 36986 686134
rect 37222 685898 72986 686134
rect 73222 685898 108986 686134
rect 109222 685898 144986 686134
rect 145222 685898 180986 686134
rect 181222 685898 216986 686134
rect 217222 685898 252986 686134
rect 253222 685898 288986 686134
rect 289222 685898 324986 686134
rect 325222 685898 360986 686134
rect 361222 685898 396986 686134
rect 397222 685898 432986 686134
rect 433222 685898 468986 686134
rect 469222 685898 504986 686134
rect 505222 685898 540986 686134
rect 541222 685898 576986 686134
rect 577222 685898 585502 686134
rect 585738 685898 586840 686134
rect -2916 685876 586840 685898
rect -1996 685874 -1396 685876
rect 804 685874 1404 685876
rect 36804 685874 37404 685876
rect 72804 685874 73404 685876
rect 108804 685874 109404 685876
rect 144804 685874 145404 685876
rect 180804 685874 181404 685876
rect 216804 685874 217404 685876
rect 252804 685874 253404 685876
rect 288804 685874 289404 685876
rect 324804 685874 325404 685876
rect 360804 685874 361404 685876
rect 396804 685874 397404 685876
rect 432804 685874 433404 685876
rect 468804 685874 469404 685876
rect 504804 685874 505404 685876
rect 540804 685874 541404 685876
rect 576804 685874 577404 685876
rect 585320 685874 585920 685876
rect -8436 679276 -7836 679278
rect 29604 679276 30204 679278
rect 65604 679276 66204 679278
rect 101604 679276 102204 679278
rect 137604 679276 138204 679278
rect 173604 679276 174204 679278
rect 209604 679276 210204 679278
rect 245604 679276 246204 679278
rect 281604 679276 282204 679278
rect 317604 679276 318204 679278
rect 353604 679276 354204 679278
rect 389604 679276 390204 679278
rect 425604 679276 426204 679278
rect 461604 679276 462204 679278
rect 497604 679276 498204 679278
rect 533604 679276 534204 679278
rect 569604 679276 570204 679278
rect 591760 679276 592360 679278
rect -8436 679254 592360 679276
rect -8436 679018 -8254 679254
rect -8018 679018 29786 679254
rect 30022 679018 65786 679254
rect 66022 679018 101786 679254
rect 102022 679018 137786 679254
rect 138022 679018 173786 679254
rect 174022 679018 209786 679254
rect 210022 679018 245786 679254
rect 246022 679018 281786 679254
rect 282022 679018 317786 679254
rect 318022 679018 353786 679254
rect 354022 679018 389786 679254
rect 390022 679018 425786 679254
rect 426022 679018 461786 679254
rect 462022 679018 497786 679254
rect 498022 679018 533786 679254
rect 534022 679018 569786 679254
rect 570022 679018 591942 679254
rect 592178 679018 592360 679254
rect -8436 678934 592360 679018
rect -8436 678698 -8254 678934
rect -8018 678698 29786 678934
rect 30022 678698 65786 678934
rect 66022 678698 101786 678934
rect 102022 678698 137786 678934
rect 138022 678698 173786 678934
rect 174022 678698 209786 678934
rect 210022 678698 245786 678934
rect 246022 678698 281786 678934
rect 282022 678698 317786 678934
rect 318022 678698 353786 678934
rect 354022 678698 389786 678934
rect 390022 678698 425786 678934
rect 426022 678698 461786 678934
rect 462022 678698 497786 678934
rect 498022 678698 533786 678934
rect 534022 678698 569786 678934
rect 570022 678698 591942 678934
rect 592178 678698 592360 678934
rect -8436 678676 592360 678698
rect -8436 678674 -7836 678676
rect 29604 678674 30204 678676
rect 65604 678674 66204 678676
rect 101604 678674 102204 678676
rect 137604 678674 138204 678676
rect 173604 678674 174204 678676
rect 209604 678674 210204 678676
rect 245604 678674 246204 678676
rect 281604 678674 282204 678676
rect 317604 678674 318204 678676
rect 353604 678674 354204 678676
rect 389604 678674 390204 678676
rect 425604 678674 426204 678676
rect 461604 678674 462204 678676
rect 497604 678674 498204 678676
rect 533604 678674 534204 678676
rect 569604 678674 570204 678676
rect 591760 678674 592360 678676
rect -6596 675676 -5996 675678
rect 26004 675676 26604 675678
rect 62004 675676 62604 675678
rect 98004 675676 98604 675678
rect 134004 675676 134604 675678
rect 170004 675676 170604 675678
rect 206004 675676 206604 675678
rect 242004 675676 242604 675678
rect 278004 675676 278604 675678
rect 314004 675676 314604 675678
rect 350004 675676 350604 675678
rect 386004 675676 386604 675678
rect 422004 675676 422604 675678
rect 458004 675676 458604 675678
rect 494004 675676 494604 675678
rect 530004 675676 530604 675678
rect 566004 675676 566604 675678
rect 589920 675676 590520 675678
rect -6596 675654 590520 675676
rect -6596 675418 -6414 675654
rect -6178 675418 26186 675654
rect 26422 675418 62186 675654
rect 62422 675418 98186 675654
rect 98422 675418 134186 675654
rect 134422 675418 170186 675654
rect 170422 675418 206186 675654
rect 206422 675418 242186 675654
rect 242422 675418 278186 675654
rect 278422 675418 314186 675654
rect 314422 675418 350186 675654
rect 350422 675418 386186 675654
rect 386422 675418 422186 675654
rect 422422 675418 458186 675654
rect 458422 675418 494186 675654
rect 494422 675418 530186 675654
rect 530422 675418 566186 675654
rect 566422 675418 590102 675654
rect 590338 675418 590520 675654
rect -6596 675334 590520 675418
rect -6596 675098 -6414 675334
rect -6178 675098 26186 675334
rect 26422 675098 62186 675334
rect 62422 675098 98186 675334
rect 98422 675098 134186 675334
rect 134422 675098 170186 675334
rect 170422 675098 206186 675334
rect 206422 675098 242186 675334
rect 242422 675098 278186 675334
rect 278422 675098 314186 675334
rect 314422 675098 350186 675334
rect 350422 675098 386186 675334
rect 386422 675098 422186 675334
rect 422422 675098 458186 675334
rect 458422 675098 494186 675334
rect 494422 675098 530186 675334
rect 530422 675098 566186 675334
rect 566422 675098 590102 675334
rect 590338 675098 590520 675334
rect -6596 675076 590520 675098
rect -6596 675074 -5996 675076
rect 26004 675074 26604 675076
rect 62004 675074 62604 675076
rect 98004 675074 98604 675076
rect 134004 675074 134604 675076
rect 170004 675074 170604 675076
rect 206004 675074 206604 675076
rect 242004 675074 242604 675076
rect 278004 675074 278604 675076
rect 314004 675074 314604 675076
rect 350004 675074 350604 675076
rect 386004 675074 386604 675076
rect 422004 675074 422604 675076
rect 458004 675074 458604 675076
rect 494004 675074 494604 675076
rect 530004 675074 530604 675076
rect 566004 675074 566604 675076
rect 589920 675074 590520 675076
rect -4756 672076 -4156 672078
rect 22404 672076 23004 672078
rect 58404 672076 59004 672078
rect 94404 672076 95004 672078
rect 130404 672076 131004 672078
rect 166404 672076 167004 672078
rect 202404 672076 203004 672078
rect 238404 672076 239004 672078
rect 274404 672076 275004 672078
rect 310404 672076 311004 672078
rect 346404 672076 347004 672078
rect 382404 672076 383004 672078
rect 418404 672076 419004 672078
rect 454404 672076 455004 672078
rect 490404 672076 491004 672078
rect 526404 672076 527004 672078
rect 562404 672076 563004 672078
rect 588080 672076 588680 672078
rect -4756 672054 588680 672076
rect -4756 671818 -4574 672054
rect -4338 671818 22586 672054
rect 22822 671818 58586 672054
rect 58822 671818 94586 672054
rect 94822 671818 130586 672054
rect 130822 671818 166586 672054
rect 166822 671818 202586 672054
rect 202822 671818 238586 672054
rect 238822 671818 274586 672054
rect 274822 671818 310586 672054
rect 310822 671818 346586 672054
rect 346822 671818 382586 672054
rect 382822 671818 418586 672054
rect 418822 671818 454586 672054
rect 454822 671818 490586 672054
rect 490822 671818 526586 672054
rect 526822 671818 562586 672054
rect 562822 671818 588262 672054
rect 588498 671818 588680 672054
rect -4756 671734 588680 671818
rect -4756 671498 -4574 671734
rect -4338 671498 22586 671734
rect 22822 671498 58586 671734
rect 58822 671498 94586 671734
rect 94822 671498 130586 671734
rect 130822 671498 166586 671734
rect 166822 671498 202586 671734
rect 202822 671498 238586 671734
rect 238822 671498 274586 671734
rect 274822 671498 310586 671734
rect 310822 671498 346586 671734
rect 346822 671498 382586 671734
rect 382822 671498 418586 671734
rect 418822 671498 454586 671734
rect 454822 671498 490586 671734
rect 490822 671498 526586 671734
rect 526822 671498 562586 671734
rect 562822 671498 588262 671734
rect 588498 671498 588680 671734
rect -4756 671476 588680 671498
rect -4756 671474 -4156 671476
rect 22404 671474 23004 671476
rect 58404 671474 59004 671476
rect 94404 671474 95004 671476
rect 130404 671474 131004 671476
rect 166404 671474 167004 671476
rect 202404 671474 203004 671476
rect 238404 671474 239004 671476
rect 274404 671474 275004 671476
rect 310404 671474 311004 671476
rect 346404 671474 347004 671476
rect 382404 671474 383004 671476
rect 418404 671474 419004 671476
rect 454404 671474 455004 671476
rect 490404 671474 491004 671476
rect 526404 671474 527004 671476
rect 562404 671474 563004 671476
rect 588080 671474 588680 671476
rect -2916 668476 -2316 668478
rect 18804 668476 19404 668478
rect 54804 668476 55404 668478
rect 90804 668476 91404 668478
rect 126804 668476 127404 668478
rect 162804 668476 163404 668478
rect 198804 668476 199404 668478
rect 234804 668476 235404 668478
rect 270804 668476 271404 668478
rect 306804 668476 307404 668478
rect 342804 668476 343404 668478
rect 378804 668476 379404 668478
rect 414804 668476 415404 668478
rect 450804 668476 451404 668478
rect 486804 668476 487404 668478
rect 522804 668476 523404 668478
rect 558804 668476 559404 668478
rect 586240 668476 586840 668478
rect -2916 668454 586840 668476
rect -2916 668218 -2734 668454
rect -2498 668218 18986 668454
rect 19222 668218 54986 668454
rect 55222 668218 90986 668454
rect 91222 668218 126986 668454
rect 127222 668218 162986 668454
rect 163222 668218 198986 668454
rect 199222 668218 234986 668454
rect 235222 668218 270986 668454
rect 271222 668218 306986 668454
rect 307222 668218 342986 668454
rect 343222 668218 378986 668454
rect 379222 668218 414986 668454
rect 415222 668218 450986 668454
rect 451222 668218 486986 668454
rect 487222 668218 522986 668454
rect 523222 668218 558986 668454
rect 559222 668218 586422 668454
rect 586658 668218 586840 668454
rect -2916 668134 586840 668218
rect -2916 667898 -2734 668134
rect -2498 667898 18986 668134
rect 19222 667898 54986 668134
rect 55222 667898 90986 668134
rect 91222 667898 126986 668134
rect 127222 667898 162986 668134
rect 163222 667898 198986 668134
rect 199222 667898 234986 668134
rect 235222 667898 270986 668134
rect 271222 667898 306986 668134
rect 307222 667898 342986 668134
rect 343222 667898 378986 668134
rect 379222 667898 414986 668134
rect 415222 667898 450986 668134
rect 451222 667898 486986 668134
rect 487222 667898 522986 668134
rect 523222 667898 558986 668134
rect 559222 667898 586422 668134
rect 586658 667898 586840 668134
rect -2916 667876 586840 667898
rect -2916 667874 -2316 667876
rect 18804 667874 19404 667876
rect 54804 667874 55404 667876
rect 90804 667874 91404 667876
rect 126804 667874 127404 667876
rect 162804 667874 163404 667876
rect 198804 667874 199404 667876
rect 234804 667874 235404 667876
rect 270804 667874 271404 667876
rect 306804 667874 307404 667876
rect 342804 667874 343404 667876
rect 378804 667874 379404 667876
rect 414804 667874 415404 667876
rect 450804 667874 451404 667876
rect 486804 667874 487404 667876
rect 522804 667874 523404 667876
rect 558804 667874 559404 667876
rect 586240 667874 586840 667876
rect -7516 661276 -6916 661278
rect 11604 661276 12204 661278
rect 47604 661276 48204 661278
rect 83604 661276 84204 661278
rect 119604 661276 120204 661278
rect 155604 661276 156204 661278
rect 191604 661276 192204 661278
rect 227604 661276 228204 661278
rect 263604 661276 264204 661278
rect 299604 661276 300204 661278
rect 335604 661276 336204 661278
rect 371604 661276 372204 661278
rect 407604 661276 408204 661278
rect 443604 661276 444204 661278
rect 479604 661276 480204 661278
rect 515604 661276 516204 661278
rect 551604 661276 552204 661278
rect 590840 661276 591440 661278
rect -8436 661254 592360 661276
rect -8436 661018 -7334 661254
rect -7098 661018 11786 661254
rect 12022 661018 47786 661254
rect 48022 661018 83786 661254
rect 84022 661018 119786 661254
rect 120022 661018 155786 661254
rect 156022 661018 191786 661254
rect 192022 661018 227786 661254
rect 228022 661018 263786 661254
rect 264022 661018 299786 661254
rect 300022 661018 335786 661254
rect 336022 661018 371786 661254
rect 372022 661018 407786 661254
rect 408022 661018 443786 661254
rect 444022 661018 479786 661254
rect 480022 661018 515786 661254
rect 516022 661018 551786 661254
rect 552022 661018 591022 661254
rect 591258 661018 592360 661254
rect -8436 660934 592360 661018
rect -8436 660698 -7334 660934
rect -7098 660698 11786 660934
rect 12022 660698 47786 660934
rect 48022 660698 83786 660934
rect 84022 660698 119786 660934
rect 120022 660698 155786 660934
rect 156022 660698 191786 660934
rect 192022 660698 227786 660934
rect 228022 660698 263786 660934
rect 264022 660698 299786 660934
rect 300022 660698 335786 660934
rect 336022 660698 371786 660934
rect 372022 660698 407786 660934
rect 408022 660698 443786 660934
rect 444022 660698 479786 660934
rect 480022 660698 515786 660934
rect 516022 660698 551786 660934
rect 552022 660698 591022 660934
rect 591258 660698 592360 660934
rect -8436 660676 592360 660698
rect -7516 660674 -6916 660676
rect 11604 660674 12204 660676
rect 47604 660674 48204 660676
rect 83604 660674 84204 660676
rect 119604 660674 120204 660676
rect 155604 660674 156204 660676
rect 191604 660674 192204 660676
rect 227604 660674 228204 660676
rect 263604 660674 264204 660676
rect 299604 660674 300204 660676
rect 335604 660674 336204 660676
rect 371604 660674 372204 660676
rect 407604 660674 408204 660676
rect 443604 660674 444204 660676
rect 479604 660674 480204 660676
rect 515604 660674 516204 660676
rect 551604 660674 552204 660676
rect 590840 660674 591440 660676
rect -5676 657676 -5076 657678
rect 8004 657676 8604 657678
rect 44004 657676 44604 657678
rect 80004 657676 80604 657678
rect 116004 657676 116604 657678
rect 152004 657676 152604 657678
rect 188004 657676 188604 657678
rect 224004 657676 224604 657678
rect 260004 657676 260604 657678
rect 296004 657676 296604 657678
rect 332004 657676 332604 657678
rect 368004 657676 368604 657678
rect 404004 657676 404604 657678
rect 440004 657676 440604 657678
rect 476004 657676 476604 657678
rect 512004 657676 512604 657678
rect 548004 657676 548604 657678
rect 589000 657676 589600 657678
rect -6596 657654 590520 657676
rect -6596 657418 -5494 657654
rect -5258 657418 8186 657654
rect 8422 657418 44186 657654
rect 44422 657418 80186 657654
rect 80422 657418 116186 657654
rect 116422 657418 152186 657654
rect 152422 657418 188186 657654
rect 188422 657418 224186 657654
rect 224422 657418 260186 657654
rect 260422 657418 296186 657654
rect 296422 657418 332186 657654
rect 332422 657418 368186 657654
rect 368422 657418 404186 657654
rect 404422 657418 440186 657654
rect 440422 657418 476186 657654
rect 476422 657418 512186 657654
rect 512422 657418 548186 657654
rect 548422 657418 589182 657654
rect 589418 657418 590520 657654
rect -6596 657334 590520 657418
rect -6596 657098 -5494 657334
rect -5258 657098 8186 657334
rect 8422 657098 44186 657334
rect 44422 657098 80186 657334
rect 80422 657098 116186 657334
rect 116422 657098 152186 657334
rect 152422 657098 188186 657334
rect 188422 657098 224186 657334
rect 224422 657098 260186 657334
rect 260422 657098 296186 657334
rect 296422 657098 332186 657334
rect 332422 657098 368186 657334
rect 368422 657098 404186 657334
rect 404422 657098 440186 657334
rect 440422 657098 476186 657334
rect 476422 657098 512186 657334
rect 512422 657098 548186 657334
rect 548422 657098 589182 657334
rect 589418 657098 590520 657334
rect -6596 657076 590520 657098
rect -5676 657074 -5076 657076
rect 8004 657074 8604 657076
rect 44004 657074 44604 657076
rect 80004 657074 80604 657076
rect 116004 657074 116604 657076
rect 152004 657074 152604 657076
rect 188004 657074 188604 657076
rect 224004 657074 224604 657076
rect 260004 657074 260604 657076
rect 296004 657074 296604 657076
rect 332004 657074 332604 657076
rect 368004 657074 368604 657076
rect 404004 657074 404604 657076
rect 440004 657074 440604 657076
rect 476004 657074 476604 657076
rect 512004 657074 512604 657076
rect 548004 657074 548604 657076
rect 589000 657074 589600 657076
rect -3836 654076 -3236 654078
rect 4404 654076 5004 654078
rect 40404 654076 41004 654078
rect 76404 654076 77004 654078
rect 112404 654076 113004 654078
rect 148404 654076 149004 654078
rect 184404 654076 185004 654078
rect 220404 654076 221004 654078
rect 256404 654076 257004 654078
rect 292404 654076 293004 654078
rect 328404 654076 329004 654078
rect 364404 654076 365004 654078
rect 400404 654076 401004 654078
rect 436404 654076 437004 654078
rect 472404 654076 473004 654078
rect 508404 654076 509004 654078
rect 544404 654076 545004 654078
rect 580404 654076 581004 654078
rect 587160 654076 587760 654078
rect -4756 654054 588680 654076
rect -4756 653818 -3654 654054
rect -3418 653818 4586 654054
rect 4822 653818 40586 654054
rect 40822 653818 76586 654054
rect 76822 653818 112586 654054
rect 112822 653818 148586 654054
rect 148822 653818 184586 654054
rect 184822 653818 220586 654054
rect 220822 653818 256586 654054
rect 256822 653818 292586 654054
rect 292822 653818 328586 654054
rect 328822 653818 364586 654054
rect 364822 653818 400586 654054
rect 400822 653818 436586 654054
rect 436822 653818 472586 654054
rect 472822 653818 508586 654054
rect 508822 653818 544586 654054
rect 544822 653818 580586 654054
rect 580822 653818 587342 654054
rect 587578 653818 588680 654054
rect -4756 653734 588680 653818
rect -4756 653498 -3654 653734
rect -3418 653498 4586 653734
rect 4822 653498 40586 653734
rect 40822 653498 76586 653734
rect 76822 653498 112586 653734
rect 112822 653498 148586 653734
rect 148822 653498 184586 653734
rect 184822 653498 220586 653734
rect 220822 653498 256586 653734
rect 256822 653498 292586 653734
rect 292822 653498 328586 653734
rect 328822 653498 364586 653734
rect 364822 653498 400586 653734
rect 400822 653498 436586 653734
rect 436822 653498 472586 653734
rect 472822 653498 508586 653734
rect 508822 653498 544586 653734
rect 544822 653498 580586 653734
rect 580822 653498 587342 653734
rect 587578 653498 588680 653734
rect -4756 653476 588680 653498
rect -3836 653474 -3236 653476
rect 4404 653474 5004 653476
rect 40404 653474 41004 653476
rect 76404 653474 77004 653476
rect 112404 653474 113004 653476
rect 148404 653474 149004 653476
rect 184404 653474 185004 653476
rect 220404 653474 221004 653476
rect 256404 653474 257004 653476
rect 292404 653474 293004 653476
rect 328404 653474 329004 653476
rect 364404 653474 365004 653476
rect 400404 653474 401004 653476
rect 436404 653474 437004 653476
rect 472404 653474 473004 653476
rect 508404 653474 509004 653476
rect 544404 653474 545004 653476
rect 580404 653474 581004 653476
rect 587160 653474 587760 653476
rect -1996 650476 -1396 650478
rect 804 650476 1404 650478
rect 36804 650476 37404 650478
rect 72804 650476 73404 650478
rect 108804 650476 109404 650478
rect 144804 650476 145404 650478
rect 180804 650476 181404 650478
rect 216804 650476 217404 650478
rect 252804 650476 253404 650478
rect 288804 650476 289404 650478
rect 324804 650476 325404 650478
rect 360804 650476 361404 650478
rect 396804 650476 397404 650478
rect 432804 650476 433404 650478
rect 468804 650476 469404 650478
rect 504804 650476 505404 650478
rect 540804 650476 541404 650478
rect 576804 650476 577404 650478
rect 585320 650476 585920 650478
rect -2916 650454 586840 650476
rect -2916 650218 -1814 650454
rect -1578 650218 986 650454
rect 1222 650218 36986 650454
rect 37222 650218 72986 650454
rect 73222 650218 108986 650454
rect 109222 650218 144986 650454
rect 145222 650218 180986 650454
rect 181222 650218 216986 650454
rect 217222 650218 252986 650454
rect 253222 650218 288986 650454
rect 289222 650218 324986 650454
rect 325222 650218 360986 650454
rect 361222 650218 396986 650454
rect 397222 650218 432986 650454
rect 433222 650218 468986 650454
rect 469222 650218 504986 650454
rect 505222 650218 540986 650454
rect 541222 650218 576986 650454
rect 577222 650218 585502 650454
rect 585738 650218 586840 650454
rect -2916 650134 586840 650218
rect -2916 649898 -1814 650134
rect -1578 649898 986 650134
rect 1222 649898 36986 650134
rect 37222 649898 72986 650134
rect 73222 649898 108986 650134
rect 109222 649898 144986 650134
rect 145222 649898 180986 650134
rect 181222 649898 216986 650134
rect 217222 649898 252986 650134
rect 253222 649898 288986 650134
rect 289222 649898 324986 650134
rect 325222 649898 360986 650134
rect 361222 649898 396986 650134
rect 397222 649898 432986 650134
rect 433222 649898 468986 650134
rect 469222 649898 504986 650134
rect 505222 649898 540986 650134
rect 541222 649898 576986 650134
rect 577222 649898 585502 650134
rect 585738 649898 586840 650134
rect -2916 649876 586840 649898
rect -1996 649874 -1396 649876
rect 804 649874 1404 649876
rect 36804 649874 37404 649876
rect 72804 649874 73404 649876
rect 108804 649874 109404 649876
rect 144804 649874 145404 649876
rect 180804 649874 181404 649876
rect 216804 649874 217404 649876
rect 252804 649874 253404 649876
rect 288804 649874 289404 649876
rect 324804 649874 325404 649876
rect 360804 649874 361404 649876
rect 396804 649874 397404 649876
rect 432804 649874 433404 649876
rect 468804 649874 469404 649876
rect 504804 649874 505404 649876
rect 540804 649874 541404 649876
rect 576804 649874 577404 649876
rect 585320 649874 585920 649876
rect -8436 643276 -7836 643278
rect 29604 643276 30204 643278
rect 65604 643276 66204 643278
rect 101604 643276 102204 643278
rect 137604 643276 138204 643278
rect 173604 643276 174204 643278
rect 209604 643276 210204 643278
rect 245604 643276 246204 643278
rect 281604 643276 282204 643278
rect 317604 643276 318204 643278
rect 353604 643276 354204 643278
rect 389604 643276 390204 643278
rect 425604 643276 426204 643278
rect 461604 643276 462204 643278
rect 497604 643276 498204 643278
rect 533604 643276 534204 643278
rect 569604 643276 570204 643278
rect 591760 643276 592360 643278
rect -8436 643254 592360 643276
rect -8436 643018 -8254 643254
rect -8018 643018 29786 643254
rect 30022 643018 65786 643254
rect 66022 643018 101786 643254
rect 102022 643018 137786 643254
rect 138022 643018 173786 643254
rect 174022 643018 209786 643254
rect 210022 643018 245786 643254
rect 246022 643018 281786 643254
rect 282022 643018 317786 643254
rect 318022 643018 353786 643254
rect 354022 643018 389786 643254
rect 390022 643018 425786 643254
rect 426022 643018 461786 643254
rect 462022 643018 497786 643254
rect 498022 643018 533786 643254
rect 534022 643018 569786 643254
rect 570022 643018 591942 643254
rect 592178 643018 592360 643254
rect -8436 642934 592360 643018
rect -8436 642698 -8254 642934
rect -8018 642698 29786 642934
rect 30022 642698 65786 642934
rect 66022 642698 101786 642934
rect 102022 642698 137786 642934
rect 138022 642698 173786 642934
rect 174022 642698 209786 642934
rect 210022 642698 245786 642934
rect 246022 642698 281786 642934
rect 282022 642698 317786 642934
rect 318022 642698 353786 642934
rect 354022 642698 389786 642934
rect 390022 642698 425786 642934
rect 426022 642698 461786 642934
rect 462022 642698 497786 642934
rect 498022 642698 533786 642934
rect 534022 642698 569786 642934
rect 570022 642698 591942 642934
rect 592178 642698 592360 642934
rect -8436 642676 592360 642698
rect -8436 642674 -7836 642676
rect 29604 642674 30204 642676
rect 65604 642674 66204 642676
rect 101604 642674 102204 642676
rect 137604 642674 138204 642676
rect 173604 642674 174204 642676
rect 209604 642674 210204 642676
rect 245604 642674 246204 642676
rect 281604 642674 282204 642676
rect 317604 642674 318204 642676
rect 353604 642674 354204 642676
rect 389604 642674 390204 642676
rect 425604 642674 426204 642676
rect 461604 642674 462204 642676
rect 497604 642674 498204 642676
rect 533604 642674 534204 642676
rect 569604 642674 570204 642676
rect 591760 642674 592360 642676
rect -6596 639676 -5996 639678
rect 26004 639676 26604 639678
rect 62004 639676 62604 639678
rect 98004 639676 98604 639678
rect 134004 639676 134604 639678
rect 170004 639676 170604 639678
rect 206004 639676 206604 639678
rect 242004 639676 242604 639678
rect 278004 639676 278604 639678
rect 314004 639676 314604 639678
rect 350004 639676 350604 639678
rect 386004 639676 386604 639678
rect 422004 639676 422604 639678
rect 458004 639676 458604 639678
rect 494004 639676 494604 639678
rect 530004 639676 530604 639678
rect 566004 639676 566604 639678
rect 589920 639676 590520 639678
rect -6596 639654 590520 639676
rect -6596 639418 -6414 639654
rect -6178 639418 26186 639654
rect 26422 639418 62186 639654
rect 62422 639418 98186 639654
rect 98422 639418 134186 639654
rect 134422 639418 170186 639654
rect 170422 639418 206186 639654
rect 206422 639418 242186 639654
rect 242422 639418 278186 639654
rect 278422 639418 314186 639654
rect 314422 639418 350186 639654
rect 350422 639418 386186 639654
rect 386422 639418 422186 639654
rect 422422 639418 458186 639654
rect 458422 639418 494186 639654
rect 494422 639418 530186 639654
rect 530422 639418 566186 639654
rect 566422 639418 590102 639654
rect 590338 639418 590520 639654
rect -6596 639334 590520 639418
rect -6596 639098 -6414 639334
rect -6178 639098 26186 639334
rect 26422 639098 62186 639334
rect 62422 639098 98186 639334
rect 98422 639098 134186 639334
rect 134422 639098 170186 639334
rect 170422 639098 206186 639334
rect 206422 639098 242186 639334
rect 242422 639098 278186 639334
rect 278422 639098 314186 639334
rect 314422 639098 350186 639334
rect 350422 639098 386186 639334
rect 386422 639098 422186 639334
rect 422422 639098 458186 639334
rect 458422 639098 494186 639334
rect 494422 639098 530186 639334
rect 530422 639098 566186 639334
rect 566422 639098 590102 639334
rect 590338 639098 590520 639334
rect -6596 639076 590520 639098
rect -6596 639074 -5996 639076
rect 26004 639074 26604 639076
rect 62004 639074 62604 639076
rect 98004 639074 98604 639076
rect 134004 639074 134604 639076
rect 170004 639074 170604 639076
rect 206004 639074 206604 639076
rect 242004 639074 242604 639076
rect 278004 639074 278604 639076
rect 314004 639074 314604 639076
rect 350004 639074 350604 639076
rect 386004 639074 386604 639076
rect 422004 639074 422604 639076
rect 458004 639074 458604 639076
rect 494004 639074 494604 639076
rect 530004 639074 530604 639076
rect 566004 639074 566604 639076
rect 589920 639074 590520 639076
rect -4756 636076 -4156 636078
rect 22404 636076 23004 636078
rect 58404 636076 59004 636078
rect 94404 636076 95004 636078
rect 130404 636076 131004 636078
rect 166404 636076 167004 636078
rect 202404 636076 203004 636078
rect 238404 636076 239004 636078
rect 274404 636076 275004 636078
rect 310404 636076 311004 636078
rect 346404 636076 347004 636078
rect 382404 636076 383004 636078
rect 418404 636076 419004 636078
rect 454404 636076 455004 636078
rect 490404 636076 491004 636078
rect 526404 636076 527004 636078
rect 562404 636076 563004 636078
rect 588080 636076 588680 636078
rect -4756 636054 588680 636076
rect -4756 635818 -4574 636054
rect -4338 635818 22586 636054
rect 22822 635818 58586 636054
rect 58822 635818 94586 636054
rect 94822 635818 130586 636054
rect 130822 635818 166586 636054
rect 166822 635818 202586 636054
rect 202822 635818 238586 636054
rect 238822 635818 274586 636054
rect 274822 635818 310586 636054
rect 310822 635818 346586 636054
rect 346822 635818 382586 636054
rect 382822 635818 418586 636054
rect 418822 635818 454586 636054
rect 454822 635818 490586 636054
rect 490822 635818 526586 636054
rect 526822 635818 562586 636054
rect 562822 635818 588262 636054
rect 588498 635818 588680 636054
rect -4756 635734 588680 635818
rect -4756 635498 -4574 635734
rect -4338 635498 22586 635734
rect 22822 635498 58586 635734
rect 58822 635498 94586 635734
rect 94822 635498 130586 635734
rect 130822 635498 166586 635734
rect 166822 635498 202586 635734
rect 202822 635498 238586 635734
rect 238822 635498 274586 635734
rect 274822 635498 310586 635734
rect 310822 635498 346586 635734
rect 346822 635498 382586 635734
rect 382822 635498 418586 635734
rect 418822 635498 454586 635734
rect 454822 635498 490586 635734
rect 490822 635498 526586 635734
rect 526822 635498 562586 635734
rect 562822 635498 588262 635734
rect 588498 635498 588680 635734
rect -4756 635476 588680 635498
rect -4756 635474 -4156 635476
rect 22404 635474 23004 635476
rect 58404 635474 59004 635476
rect 94404 635474 95004 635476
rect 130404 635474 131004 635476
rect 166404 635474 167004 635476
rect 202404 635474 203004 635476
rect 238404 635474 239004 635476
rect 274404 635474 275004 635476
rect 310404 635474 311004 635476
rect 346404 635474 347004 635476
rect 382404 635474 383004 635476
rect 418404 635474 419004 635476
rect 454404 635474 455004 635476
rect 490404 635474 491004 635476
rect 526404 635474 527004 635476
rect 562404 635474 563004 635476
rect 588080 635474 588680 635476
rect -2916 632476 -2316 632478
rect 18804 632476 19404 632478
rect 54804 632476 55404 632478
rect 90804 632476 91404 632478
rect 126804 632476 127404 632478
rect 162804 632476 163404 632478
rect 198804 632476 199404 632478
rect 234804 632476 235404 632478
rect 270804 632476 271404 632478
rect 306804 632476 307404 632478
rect 342804 632476 343404 632478
rect 378804 632476 379404 632478
rect 414804 632476 415404 632478
rect 450804 632476 451404 632478
rect 486804 632476 487404 632478
rect 522804 632476 523404 632478
rect 558804 632476 559404 632478
rect 586240 632476 586840 632478
rect -2916 632454 586840 632476
rect -2916 632218 -2734 632454
rect -2498 632218 18986 632454
rect 19222 632218 54986 632454
rect 55222 632218 90986 632454
rect 91222 632218 126986 632454
rect 127222 632218 162986 632454
rect 163222 632218 198986 632454
rect 199222 632218 234986 632454
rect 235222 632218 270986 632454
rect 271222 632218 306986 632454
rect 307222 632218 342986 632454
rect 343222 632218 378986 632454
rect 379222 632218 414986 632454
rect 415222 632218 450986 632454
rect 451222 632218 486986 632454
rect 487222 632218 522986 632454
rect 523222 632218 558986 632454
rect 559222 632218 586422 632454
rect 586658 632218 586840 632454
rect -2916 632134 586840 632218
rect -2916 631898 -2734 632134
rect -2498 631898 18986 632134
rect 19222 631898 54986 632134
rect 55222 631898 90986 632134
rect 91222 631898 126986 632134
rect 127222 631898 162986 632134
rect 163222 631898 198986 632134
rect 199222 631898 234986 632134
rect 235222 631898 270986 632134
rect 271222 631898 306986 632134
rect 307222 631898 342986 632134
rect 343222 631898 378986 632134
rect 379222 631898 414986 632134
rect 415222 631898 450986 632134
rect 451222 631898 486986 632134
rect 487222 631898 522986 632134
rect 523222 631898 558986 632134
rect 559222 631898 586422 632134
rect 586658 631898 586840 632134
rect -2916 631876 586840 631898
rect -2916 631874 -2316 631876
rect 18804 631874 19404 631876
rect 54804 631874 55404 631876
rect 90804 631874 91404 631876
rect 126804 631874 127404 631876
rect 162804 631874 163404 631876
rect 198804 631874 199404 631876
rect 234804 631874 235404 631876
rect 270804 631874 271404 631876
rect 306804 631874 307404 631876
rect 342804 631874 343404 631876
rect 378804 631874 379404 631876
rect 414804 631874 415404 631876
rect 450804 631874 451404 631876
rect 486804 631874 487404 631876
rect 522804 631874 523404 631876
rect 558804 631874 559404 631876
rect 586240 631874 586840 631876
rect -7516 625276 -6916 625278
rect 11604 625276 12204 625278
rect 47604 625276 48204 625278
rect 83604 625276 84204 625278
rect 119604 625276 120204 625278
rect 155604 625276 156204 625278
rect 191604 625276 192204 625278
rect 227604 625276 228204 625278
rect 263604 625276 264204 625278
rect 299604 625276 300204 625278
rect 335604 625276 336204 625278
rect 371604 625276 372204 625278
rect 407604 625276 408204 625278
rect 443604 625276 444204 625278
rect 479604 625276 480204 625278
rect 515604 625276 516204 625278
rect 551604 625276 552204 625278
rect 590840 625276 591440 625278
rect -8436 625254 592360 625276
rect -8436 625018 -7334 625254
rect -7098 625018 11786 625254
rect 12022 625018 47786 625254
rect 48022 625018 83786 625254
rect 84022 625018 119786 625254
rect 120022 625018 155786 625254
rect 156022 625018 191786 625254
rect 192022 625018 227786 625254
rect 228022 625018 263786 625254
rect 264022 625018 299786 625254
rect 300022 625018 335786 625254
rect 336022 625018 371786 625254
rect 372022 625018 407786 625254
rect 408022 625018 443786 625254
rect 444022 625018 479786 625254
rect 480022 625018 515786 625254
rect 516022 625018 551786 625254
rect 552022 625018 591022 625254
rect 591258 625018 592360 625254
rect -8436 624934 592360 625018
rect -8436 624698 -7334 624934
rect -7098 624698 11786 624934
rect 12022 624698 47786 624934
rect 48022 624698 83786 624934
rect 84022 624698 119786 624934
rect 120022 624698 155786 624934
rect 156022 624698 191786 624934
rect 192022 624698 227786 624934
rect 228022 624698 263786 624934
rect 264022 624698 299786 624934
rect 300022 624698 335786 624934
rect 336022 624698 371786 624934
rect 372022 624698 407786 624934
rect 408022 624698 443786 624934
rect 444022 624698 479786 624934
rect 480022 624698 515786 624934
rect 516022 624698 551786 624934
rect 552022 624698 591022 624934
rect 591258 624698 592360 624934
rect -8436 624676 592360 624698
rect -7516 624674 -6916 624676
rect 11604 624674 12204 624676
rect 47604 624674 48204 624676
rect 83604 624674 84204 624676
rect 119604 624674 120204 624676
rect 155604 624674 156204 624676
rect 191604 624674 192204 624676
rect 227604 624674 228204 624676
rect 263604 624674 264204 624676
rect 299604 624674 300204 624676
rect 335604 624674 336204 624676
rect 371604 624674 372204 624676
rect 407604 624674 408204 624676
rect 443604 624674 444204 624676
rect 479604 624674 480204 624676
rect 515604 624674 516204 624676
rect 551604 624674 552204 624676
rect 590840 624674 591440 624676
rect -5676 621676 -5076 621678
rect 8004 621676 8604 621678
rect 44004 621676 44604 621678
rect 80004 621676 80604 621678
rect 116004 621676 116604 621678
rect 152004 621676 152604 621678
rect 188004 621676 188604 621678
rect 224004 621676 224604 621678
rect 260004 621676 260604 621678
rect 296004 621676 296604 621678
rect 332004 621676 332604 621678
rect 368004 621676 368604 621678
rect 404004 621676 404604 621678
rect 440004 621676 440604 621678
rect 476004 621676 476604 621678
rect 512004 621676 512604 621678
rect 548004 621676 548604 621678
rect 589000 621676 589600 621678
rect -6596 621654 590520 621676
rect -6596 621418 -5494 621654
rect -5258 621418 8186 621654
rect 8422 621418 44186 621654
rect 44422 621418 80186 621654
rect 80422 621418 116186 621654
rect 116422 621418 152186 621654
rect 152422 621418 188186 621654
rect 188422 621418 224186 621654
rect 224422 621418 260186 621654
rect 260422 621418 296186 621654
rect 296422 621418 332186 621654
rect 332422 621418 368186 621654
rect 368422 621418 404186 621654
rect 404422 621418 440186 621654
rect 440422 621418 476186 621654
rect 476422 621418 512186 621654
rect 512422 621418 548186 621654
rect 548422 621418 589182 621654
rect 589418 621418 590520 621654
rect -6596 621334 590520 621418
rect -6596 621098 -5494 621334
rect -5258 621098 8186 621334
rect 8422 621098 44186 621334
rect 44422 621098 80186 621334
rect 80422 621098 116186 621334
rect 116422 621098 152186 621334
rect 152422 621098 188186 621334
rect 188422 621098 224186 621334
rect 224422 621098 260186 621334
rect 260422 621098 296186 621334
rect 296422 621098 332186 621334
rect 332422 621098 368186 621334
rect 368422 621098 404186 621334
rect 404422 621098 440186 621334
rect 440422 621098 476186 621334
rect 476422 621098 512186 621334
rect 512422 621098 548186 621334
rect 548422 621098 589182 621334
rect 589418 621098 590520 621334
rect -6596 621076 590520 621098
rect -5676 621074 -5076 621076
rect 8004 621074 8604 621076
rect 44004 621074 44604 621076
rect 80004 621074 80604 621076
rect 116004 621074 116604 621076
rect 152004 621074 152604 621076
rect 188004 621074 188604 621076
rect 224004 621074 224604 621076
rect 260004 621074 260604 621076
rect 296004 621074 296604 621076
rect 332004 621074 332604 621076
rect 368004 621074 368604 621076
rect 404004 621074 404604 621076
rect 440004 621074 440604 621076
rect 476004 621074 476604 621076
rect 512004 621074 512604 621076
rect 548004 621074 548604 621076
rect 589000 621074 589600 621076
rect -3836 618076 -3236 618078
rect 4404 618076 5004 618078
rect 40404 618076 41004 618078
rect 76404 618076 77004 618078
rect 112404 618076 113004 618078
rect 148404 618076 149004 618078
rect 184404 618076 185004 618078
rect 220404 618076 221004 618078
rect 256404 618076 257004 618078
rect 292404 618076 293004 618078
rect 328404 618076 329004 618078
rect 364404 618076 365004 618078
rect 400404 618076 401004 618078
rect 436404 618076 437004 618078
rect 472404 618076 473004 618078
rect 508404 618076 509004 618078
rect 544404 618076 545004 618078
rect 580404 618076 581004 618078
rect 587160 618076 587760 618078
rect -4756 618054 588680 618076
rect -4756 617818 -3654 618054
rect -3418 617818 4586 618054
rect 4822 617818 40586 618054
rect 40822 617818 76586 618054
rect 76822 617818 112586 618054
rect 112822 617818 148586 618054
rect 148822 617818 184586 618054
rect 184822 617818 220586 618054
rect 220822 617818 256586 618054
rect 256822 617818 292586 618054
rect 292822 617818 328586 618054
rect 328822 617818 364586 618054
rect 364822 617818 400586 618054
rect 400822 617818 436586 618054
rect 436822 617818 472586 618054
rect 472822 617818 508586 618054
rect 508822 617818 544586 618054
rect 544822 617818 580586 618054
rect 580822 617818 587342 618054
rect 587578 617818 588680 618054
rect -4756 617734 588680 617818
rect -4756 617498 -3654 617734
rect -3418 617498 4586 617734
rect 4822 617498 40586 617734
rect 40822 617498 76586 617734
rect 76822 617498 112586 617734
rect 112822 617498 148586 617734
rect 148822 617498 184586 617734
rect 184822 617498 220586 617734
rect 220822 617498 256586 617734
rect 256822 617498 292586 617734
rect 292822 617498 328586 617734
rect 328822 617498 364586 617734
rect 364822 617498 400586 617734
rect 400822 617498 436586 617734
rect 436822 617498 472586 617734
rect 472822 617498 508586 617734
rect 508822 617498 544586 617734
rect 544822 617498 580586 617734
rect 580822 617498 587342 617734
rect 587578 617498 588680 617734
rect -4756 617476 588680 617498
rect -3836 617474 -3236 617476
rect 4404 617474 5004 617476
rect 40404 617474 41004 617476
rect 76404 617474 77004 617476
rect 112404 617474 113004 617476
rect 148404 617474 149004 617476
rect 184404 617474 185004 617476
rect 220404 617474 221004 617476
rect 256404 617474 257004 617476
rect 292404 617474 293004 617476
rect 328404 617474 329004 617476
rect 364404 617474 365004 617476
rect 400404 617474 401004 617476
rect 436404 617474 437004 617476
rect 472404 617474 473004 617476
rect 508404 617474 509004 617476
rect 544404 617474 545004 617476
rect 580404 617474 581004 617476
rect 587160 617474 587760 617476
rect -1996 614476 -1396 614478
rect 804 614476 1404 614478
rect 36804 614476 37404 614478
rect 72804 614476 73404 614478
rect 108804 614476 109404 614478
rect 144804 614476 145404 614478
rect 180804 614476 181404 614478
rect 216804 614476 217404 614478
rect 252804 614476 253404 614478
rect 288804 614476 289404 614478
rect 324804 614476 325404 614478
rect 360804 614476 361404 614478
rect 396804 614476 397404 614478
rect 432804 614476 433404 614478
rect 468804 614476 469404 614478
rect 504804 614476 505404 614478
rect 540804 614476 541404 614478
rect 576804 614476 577404 614478
rect 585320 614476 585920 614478
rect -2916 614454 586840 614476
rect -2916 614218 -1814 614454
rect -1578 614218 986 614454
rect 1222 614218 36986 614454
rect 37222 614218 72986 614454
rect 73222 614218 108986 614454
rect 109222 614218 144986 614454
rect 145222 614218 180986 614454
rect 181222 614218 216986 614454
rect 217222 614218 252986 614454
rect 253222 614218 288986 614454
rect 289222 614218 324986 614454
rect 325222 614218 360986 614454
rect 361222 614218 396986 614454
rect 397222 614218 432986 614454
rect 433222 614218 468986 614454
rect 469222 614218 504986 614454
rect 505222 614218 540986 614454
rect 541222 614218 576986 614454
rect 577222 614218 585502 614454
rect 585738 614218 586840 614454
rect -2916 614134 586840 614218
rect -2916 613898 -1814 614134
rect -1578 613898 986 614134
rect 1222 613898 36986 614134
rect 37222 613898 72986 614134
rect 73222 613898 108986 614134
rect 109222 613898 144986 614134
rect 145222 613898 180986 614134
rect 181222 613898 216986 614134
rect 217222 613898 252986 614134
rect 253222 613898 288986 614134
rect 289222 613898 324986 614134
rect 325222 613898 360986 614134
rect 361222 613898 396986 614134
rect 397222 613898 432986 614134
rect 433222 613898 468986 614134
rect 469222 613898 504986 614134
rect 505222 613898 540986 614134
rect 541222 613898 576986 614134
rect 577222 613898 585502 614134
rect 585738 613898 586840 614134
rect -2916 613876 586840 613898
rect -1996 613874 -1396 613876
rect 804 613874 1404 613876
rect 36804 613874 37404 613876
rect 72804 613874 73404 613876
rect 108804 613874 109404 613876
rect 144804 613874 145404 613876
rect 180804 613874 181404 613876
rect 216804 613874 217404 613876
rect 252804 613874 253404 613876
rect 288804 613874 289404 613876
rect 324804 613874 325404 613876
rect 360804 613874 361404 613876
rect 396804 613874 397404 613876
rect 432804 613874 433404 613876
rect 468804 613874 469404 613876
rect 504804 613874 505404 613876
rect 540804 613874 541404 613876
rect 576804 613874 577404 613876
rect 585320 613874 585920 613876
rect -8436 607276 -7836 607278
rect 29604 607276 30204 607278
rect 65604 607276 66204 607278
rect 101604 607276 102204 607278
rect 137604 607276 138204 607278
rect 173604 607276 174204 607278
rect 209604 607276 210204 607278
rect 245604 607276 246204 607278
rect 281604 607276 282204 607278
rect 317604 607276 318204 607278
rect 353604 607276 354204 607278
rect 389604 607276 390204 607278
rect 425604 607276 426204 607278
rect 461604 607276 462204 607278
rect 497604 607276 498204 607278
rect 533604 607276 534204 607278
rect 569604 607276 570204 607278
rect 591760 607276 592360 607278
rect -8436 607254 592360 607276
rect -8436 607018 -8254 607254
rect -8018 607018 29786 607254
rect 30022 607018 65786 607254
rect 66022 607018 101786 607254
rect 102022 607018 137786 607254
rect 138022 607018 173786 607254
rect 174022 607018 209786 607254
rect 210022 607018 245786 607254
rect 246022 607018 281786 607254
rect 282022 607018 317786 607254
rect 318022 607018 353786 607254
rect 354022 607018 389786 607254
rect 390022 607018 425786 607254
rect 426022 607018 461786 607254
rect 462022 607018 497786 607254
rect 498022 607018 533786 607254
rect 534022 607018 569786 607254
rect 570022 607018 591942 607254
rect 592178 607018 592360 607254
rect -8436 606934 592360 607018
rect -8436 606698 -8254 606934
rect -8018 606698 29786 606934
rect 30022 606698 65786 606934
rect 66022 606698 101786 606934
rect 102022 606698 137786 606934
rect 138022 606698 173786 606934
rect 174022 606698 209786 606934
rect 210022 606698 245786 606934
rect 246022 606698 281786 606934
rect 282022 606698 317786 606934
rect 318022 606698 353786 606934
rect 354022 606698 389786 606934
rect 390022 606698 425786 606934
rect 426022 606698 461786 606934
rect 462022 606698 497786 606934
rect 498022 606698 533786 606934
rect 534022 606698 569786 606934
rect 570022 606698 591942 606934
rect 592178 606698 592360 606934
rect -8436 606676 592360 606698
rect -8436 606674 -7836 606676
rect 29604 606674 30204 606676
rect 65604 606674 66204 606676
rect 101604 606674 102204 606676
rect 137604 606674 138204 606676
rect 173604 606674 174204 606676
rect 209604 606674 210204 606676
rect 245604 606674 246204 606676
rect 281604 606674 282204 606676
rect 317604 606674 318204 606676
rect 353604 606674 354204 606676
rect 389604 606674 390204 606676
rect 425604 606674 426204 606676
rect 461604 606674 462204 606676
rect 497604 606674 498204 606676
rect 533604 606674 534204 606676
rect 569604 606674 570204 606676
rect 591760 606674 592360 606676
rect -6596 603676 -5996 603678
rect 26004 603676 26604 603678
rect 62004 603676 62604 603678
rect 98004 603676 98604 603678
rect 134004 603676 134604 603678
rect 170004 603676 170604 603678
rect 206004 603676 206604 603678
rect 242004 603676 242604 603678
rect 278004 603676 278604 603678
rect 314004 603676 314604 603678
rect 350004 603676 350604 603678
rect 386004 603676 386604 603678
rect 422004 603676 422604 603678
rect 458004 603676 458604 603678
rect 494004 603676 494604 603678
rect 530004 603676 530604 603678
rect 566004 603676 566604 603678
rect 589920 603676 590520 603678
rect -6596 603654 590520 603676
rect -6596 603418 -6414 603654
rect -6178 603418 26186 603654
rect 26422 603418 62186 603654
rect 62422 603418 98186 603654
rect 98422 603418 134186 603654
rect 134422 603418 170186 603654
rect 170422 603418 206186 603654
rect 206422 603418 242186 603654
rect 242422 603418 278186 603654
rect 278422 603418 314186 603654
rect 314422 603418 350186 603654
rect 350422 603418 386186 603654
rect 386422 603418 422186 603654
rect 422422 603418 458186 603654
rect 458422 603418 494186 603654
rect 494422 603418 530186 603654
rect 530422 603418 566186 603654
rect 566422 603418 590102 603654
rect 590338 603418 590520 603654
rect -6596 603334 590520 603418
rect -6596 603098 -6414 603334
rect -6178 603098 26186 603334
rect 26422 603098 62186 603334
rect 62422 603098 98186 603334
rect 98422 603098 134186 603334
rect 134422 603098 170186 603334
rect 170422 603098 206186 603334
rect 206422 603098 242186 603334
rect 242422 603098 278186 603334
rect 278422 603098 314186 603334
rect 314422 603098 350186 603334
rect 350422 603098 386186 603334
rect 386422 603098 422186 603334
rect 422422 603098 458186 603334
rect 458422 603098 494186 603334
rect 494422 603098 530186 603334
rect 530422 603098 566186 603334
rect 566422 603098 590102 603334
rect 590338 603098 590520 603334
rect -6596 603076 590520 603098
rect -6596 603074 -5996 603076
rect 26004 603074 26604 603076
rect 62004 603074 62604 603076
rect 98004 603074 98604 603076
rect 134004 603074 134604 603076
rect 170004 603074 170604 603076
rect 206004 603074 206604 603076
rect 242004 603074 242604 603076
rect 278004 603074 278604 603076
rect 314004 603074 314604 603076
rect 350004 603074 350604 603076
rect 386004 603074 386604 603076
rect 422004 603074 422604 603076
rect 458004 603074 458604 603076
rect 494004 603074 494604 603076
rect 530004 603074 530604 603076
rect 566004 603074 566604 603076
rect 589920 603074 590520 603076
rect -4756 600076 -4156 600078
rect 22404 600076 23004 600078
rect 58404 600076 59004 600078
rect 94404 600076 95004 600078
rect 130404 600076 131004 600078
rect 166404 600076 167004 600078
rect 202404 600076 203004 600078
rect 238404 600076 239004 600078
rect 274404 600076 275004 600078
rect 310404 600076 311004 600078
rect 346404 600076 347004 600078
rect 382404 600076 383004 600078
rect 418404 600076 419004 600078
rect 454404 600076 455004 600078
rect 490404 600076 491004 600078
rect 526404 600076 527004 600078
rect 562404 600076 563004 600078
rect 588080 600076 588680 600078
rect -4756 600054 588680 600076
rect -4756 599818 -4574 600054
rect -4338 599818 22586 600054
rect 22822 599818 58586 600054
rect 58822 599818 94586 600054
rect 94822 599818 130586 600054
rect 130822 599818 166586 600054
rect 166822 599818 202586 600054
rect 202822 599818 238586 600054
rect 238822 599818 274586 600054
rect 274822 599818 310586 600054
rect 310822 599818 346586 600054
rect 346822 599818 382586 600054
rect 382822 599818 418586 600054
rect 418822 599818 454586 600054
rect 454822 599818 490586 600054
rect 490822 599818 526586 600054
rect 526822 599818 562586 600054
rect 562822 599818 588262 600054
rect 588498 599818 588680 600054
rect -4756 599734 588680 599818
rect -4756 599498 -4574 599734
rect -4338 599498 22586 599734
rect 22822 599498 58586 599734
rect 58822 599498 94586 599734
rect 94822 599498 130586 599734
rect 130822 599498 166586 599734
rect 166822 599498 202586 599734
rect 202822 599498 238586 599734
rect 238822 599498 274586 599734
rect 274822 599498 310586 599734
rect 310822 599498 346586 599734
rect 346822 599498 382586 599734
rect 382822 599498 418586 599734
rect 418822 599498 454586 599734
rect 454822 599498 490586 599734
rect 490822 599498 526586 599734
rect 526822 599498 562586 599734
rect 562822 599498 588262 599734
rect 588498 599498 588680 599734
rect -4756 599476 588680 599498
rect -4756 599474 -4156 599476
rect 22404 599474 23004 599476
rect 58404 599474 59004 599476
rect 94404 599474 95004 599476
rect 130404 599474 131004 599476
rect 166404 599474 167004 599476
rect 202404 599474 203004 599476
rect 238404 599474 239004 599476
rect 274404 599474 275004 599476
rect 310404 599474 311004 599476
rect 346404 599474 347004 599476
rect 382404 599474 383004 599476
rect 418404 599474 419004 599476
rect 454404 599474 455004 599476
rect 490404 599474 491004 599476
rect 526404 599474 527004 599476
rect 562404 599474 563004 599476
rect 588080 599474 588680 599476
rect -2916 596476 -2316 596478
rect 18804 596476 19404 596478
rect 54804 596476 55404 596478
rect 90804 596476 91404 596478
rect 126804 596476 127404 596478
rect 162804 596476 163404 596478
rect 198804 596476 199404 596478
rect 234804 596476 235404 596478
rect 270804 596476 271404 596478
rect 306804 596476 307404 596478
rect 342804 596476 343404 596478
rect 378804 596476 379404 596478
rect 414804 596476 415404 596478
rect 450804 596476 451404 596478
rect 486804 596476 487404 596478
rect 522804 596476 523404 596478
rect 558804 596476 559404 596478
rect 586240 596476 586840 596478
rect -2916 596454 586840 596476
rect -2916 596218 -2734 596454
rect -2498 596218 18986 596454
rect 19222 596218 54986 596454
rect 55222 596218 90986 596454
rect 91222 596218 126986 596454
rect 127222 596218 162986 596454
rect 163222 596218 198986 596454
rect 199222 596218 234986 596454
rect 235222 596218 270986 596454
rect 271222 596218 306986 596454
rect 307222 596218 342986 596454
rect 343222 596218 378986 596454
rect 379222 596218 414986 596454
rect 415222 596218 450986 596454
rect 451222 596218 486986 596454
rect 487222 596218 522986 596454
rect 523222 596218 558986 596454
rect 559222 596218 586422 596454
rect 586658 596218 586840 596454
rect -2916 596134 586840 596218
rect -2916 595898 -2734 596134
rect -2498 595898 18986 596134
rect 19222 595898 54986 596134
rect 55222 595898 90986 596134
rect 91222 595898 126986 596134
rect 127222 595898 162986 596134
rect 163222 595898 198986 596134
rect 199222 595898 234986 596134
rect 235222 595898 270986 596134
rect 271222 595898 306986 596134
rect 307222 595898 342986 596134
rect 343222 595898 378986 596134
rect 379222 595898 414986 596134
rect 415222 595898 450986 596134
rect 451222 595898 486986 596134
rect 487222 595898 522986 596134
rect 523222 595898 558986 596134
rect 559222 595898 586422 596134
rect 586658 595898 586840 596134
rect -2916 595876 586840 595898
rect -2916 595874 -2316 595876
rect 18804 595874 19404 595876
rect 54804 595874 55404 595876
rect 90804 595874 91404 595876
rect 126804 595874 127404 595876
rect 162804 595874 163404 595876
rect 198804 595874 199404 595876
rect 234804 595874 235404 595876
rect 270804 595874 271404 595876
rect 306804 595874 307404 595876
rect 342804 595874 343404 595876
rect 378804 595874 379404 595876
rect 414804 595874 415404 595876
rect 450804 595874 451404 595876
rect 486804 595874 487404 595876
rect 522804 595874 523404 595876
rect 558804 595874 559404 595876
rect 586240 595874 586840 595876
rect -7516 589276 -6916 589278
rect 11604 589276 12204 589278
rect 47604 589276 48204 589278
rect 83604 589276 84204 589278
rect 119604 589276 120204 589278
rect 155604 589276 156204 589278
rect 191604 589276 192204 589278
rect 227604 589276 228204 589278
rect 263604 589276 264204 589278
rect 299604 589276 300204 589278
rect 335604 589276 336204 589278
rect 371604 589276 372204 589278
rect 407604 589276 408204 589278
rect 443604 589276 444204 589278
rect 479604 589276 480204 589278
rect 515604 589276 516204 589278
rect 551604 589276 552204 589278
rect 590840 589276 591440 589278
rect -8436 589254 592360 589276
rect -8436 589018 -7334 589254
rect -7098 589018 11786 589254
rect 12022 589018 47786 589254
rect 48022 589018 83786 589254
rect 84022 589018 119786 589254
rect 120022 589018 155786 589254
rect 156022 589018 191786 589254
rect 192022 589018 227786 589254
rect 228022 589018 263786 589254
rect 264022 589018 299786 589254
rect 300022 589018 335786 589254
rect 336022 589018 371786 589254
rect 372022 589018 407786 589254
rect 408022 589018 443786 589254
rect 444022 589018 479786 589254
rect 480022 589018 515786 589254
rect 516022 589018 551786 589254
rect 552022 589018 591022 589254
rect 591258 589018 592360 589254
rect -8436 588934 592360 589018
rect -8436 588698 -7334 588934
rect -7098 588698 11786 588934
rect 12022 588698 47786 588934
rect 48022 588698 83786 588934
rect 84022 588698 119786 588934
rect 120022 588698 155786 588934
rect 156022 588698 191786 588934
rect 192022 588698 227786 588934
rect 228022 588698 263786 588934
rect 264022 588698 299786 588934
rect 300022 588698 335786 588934
rect 336022 588698 371786 588934
rect 372022 588698 407786 588934
rect 408022 588698 443786 588934
rect 444022 588698 479786 588934
rect 480022 588698 515786 588934
rect 516022 588698 551786 588934
rect 552022 588698 591022 588934
rect 591258 588698 592360 588934
rect -8436 588676 592360 588698
rect -7516 588674 -6916 588676
rect 11604 588674 12204 588676
rect 47604 588674 48204 588676
rect 83604 588674 84204 588676
rect 119604 588674 120204 588676
rect 155604 588674 156204 588676
rect 191604 588674 192204 588676
rect 227604 588674 228204 588676
rect 263604 588674 264204 588676
rect 299604 588674 300204 588676
rect 335604 588674 336204 588676
rect 371604 588674 372204 588676
rect 407604 588674 408204 588676
rect 443604 588674 444204 588676
rect 479604 588674 480204 588676
rect 515604 588674 516204 588676
rect 551604 588674 552204 588676
rect 590840 588674 591440 588676
rect -5676 585676 -5076 585678
rect 8004 585676 8604 585678
rect 44004 585676 44604 585678
rect 80004 585676 80604 585678
rect 116004 585676 116604 585678
rect 152004 585676 152604 585678
rect 188004 585676 188604 585678
rect 224004 585676 224604 585678
rect 260004 585676 260604 585678
rect 296004 585676 296604 585678
rect 332004 585676 332604 585678
rect 368004 585676 368604 585678
rect 404004 585676 404604 585678
rect 440004 585676 440604 585678
rect 476004 585676 476604 585678
rect 512004 585676 512604 585678
rect 548004 585676 548604 585678
rect 589000 585676 589600 585678
rect -6596 585654 590520 585676
rect -6596 585418 -5494 585654
rect -5258 585418 8186 585654
rect 8422 585418 44186 585654
rect 44422 585418 80186 585654
rect 80422 585418 116186 585654
rect 116422 585418 152186 585654
rect 152422 585418 188186 585654
rect 188422 585418 224186 585654
rect 224422 585418 260186 585654
rect 260422 585418 296186 585654
rect 296422 585418 332186 585654
rect 332422 585418 368186 585654
rect 368422 585418 404186 585654
rect 404422 585418 440186 585654
rect 440422 585418 476186 585654
rect 476422 585418 512186 585654
rect 512422 585418 548186 585654
rect 548422 585418 589182 585654
rect 589418 585418 590520 585654
rect -6596 585334 590520 585418
rect -6596 585098 -5494 585334
rect -5258 585098 8186 585334
rect 8422 585098 44186 585334
rect 44422 585098 80186 585334
rect 80422 585098 116186 585334
rect 116422 585098 152186 585334
rect 152422 585098 188186 585334
rect 188422 585098 224186 585334
rect 224422 585098 260186 585334
rect 260422 585098 296186 585334
rect 296422 585098 332186 585334
rect 332422 585098 368186 585334
rect 368422 585098 404186 585334
rect 404422 585098 440186 585334
rect 440422 585098 476186 585334
rect 476422 585098 512186 585334
rect 512422 585098 548186 585334
rect 548422 585098 589182 585334
rect 589418 585098 590520 585334
rect -6596 585076 590520 585098
rect -5676 585074 -5076 585076
rect 8004 585074 8604 585076
rect 44004 585074 44604 585076
rect 80004 585074 80604 585076
rect 116004 585074 116604 585076
rect 152004 585074 152604 585076
rect 188004 585074 188604 585076
rect 224004 585074 224604 585076
rect 260004 585074 260604 585076
rect 296004 585074 296604 585076
rect 332004 585074 332604 585076
rect 368004 585074 368604 585076
rect 404004 585074 404604 585076
rect 440004 585074 440604 585076
rect 476004 585074 476604 585076
rect 512004 585074 512604 585076
rect 548004 585074 548604 585076
rect 589000 585074 589600 585076
rect -3836 582076 -3236 582078
rect 4404 582076 5004 582078
rect 40404 582076 41004 582078
rect 76404 582076 77004 582078
rect 112404 582076 113004 582078
rect 148404 582076 149004 582078
rect 184404 582076 185004 582078
rect 220404 582076 221004 582078
rect 256404 582076 257004 582078
rect 292404 582076 293004 582078
rect 328404 582076 329004 582078
rect 364404 582076 365004 582078
rect 400404 582076 401004 582078
rect 436404 582076 437004 582078
rect 472404 582076 473004 582078
rect 508404 582076 509004 582078
rect 544404 582076 545004 582078
rect 580404 582076 581004 582078
rect 587160 582076 587760 582078
rect -4756 582054 588680 582076
rect -4756 581818 -3654 582054
rect -3418 581818 4586 582054
rect 4822 581818 40586 582054
rect 40822 581818 76586 582054
rect 76822 581818 112586 582054
rect 112822 581818 148586 582054
rect 148822 581818 184586 582054
rect 184822 581818 220586 582054
rect 220822 581818 256586 582054
rect 256822 581818 292586 582054
rect 292822 581818 328586 582054
rect 328822 581818 364586 582054
rect 364822 581818 400586 582054
rect 400822 581818 436586 582054
rect 436822 581818 472586 582054
rect 472822 581818 508586 582054
rect 508822 581818 544586 582054
rect 544822 581818 580586 582054
rect 580822 581818 587342 582054
rect 587578 581818 588680 582054
rect -4756 581734 588680 581818
rect -4756 581498 -3654 581734
rect -3418 581498 4586 581734
rect 4822 581498 40586 581734
rect 40822 581498 76586 581734
rect 76822 581498 112586 581734
rect 112822 581498 148586 581734
rect 148822 581498 184586 581734
rect 184822 581498 220586 581734
rect 220822 581498 256586 581734
rect 256822 581498 292586 581734
rect 292822 581498 328586 581734
rect 328822 581498 364586 581734
rect 364822 581498 400586 581734
rect 400822 581498 436586 581734
rect 436822 581498 472586 581734
rect 472822 581498 508586 581734
rect 508822 581498 544586 581734
rect 544822 581498 580586 581734
rect 580822 581498 587342 581734
rect 587578 581498 588680 581734
rect -4756 581476 588680 581498
rect -3836 581474 -3236 581476
rect 4404 581474 5004 581476
rect 40404 581474 41004 581476
rect 76404 581474 77004 581476
rect 112404 581474 113004 581476
rect 148404 581474 149004 581476
rect 184404 581474 185004 581476
rect 220404 581474 221004 581476
rect 256404 581474 257004 581476
rect 292404 581474 293004 581476
rect 328404 581474 329004 581476
rect 364404 581474 365004 581476
rect 400404 581474 401004 581476
rect 436404 581474 437004 581476
rect 472404 581474 473004 581476
rect 508404 581474 509004 581476
rect 544404 581474 545004 581476
rect 580404 581474 581004 581476
rect 587160 581474 587760 581476
rect -1996 578476 -1396 578478
rect 804 578476 1404 578478
rect 36804 578476 37404 578478
rect 72804 578476 73404 578478
rect 108804 578476 109404 578478
rect 144804 578476 145404 578478
rect 180804 578476 181404 578478
rect 216804 578476 217404 578478
rect 252804 578476 253404 578478
rect 288804 578476 289404 578478
rect 324804 578476 325404 578478
rect 360804 578476 361404 578478
rect 396804 578476 397404 578478
rect 432804 578476 433404 578478
rect 468804 578476 469404 578478
rect 504804 578476 505404 578478
rect 540804 578476 541404 578478
rect 576804 578476 577404 578478
rect 585320 578476 585920 578478
rect -2916 578454 586840 578476
rect -2916 578218 -1814 578454
rect -1578 578218 986 578454
rect 1222 578218 36986 578454
rect 37222 578218 72986 578454
rect 73222 578218 108986 578454
rect 109222 578218 144986 578454
rect 145222 578218 180986 578454
rect 181222 578218 216986 578454
rect 217222 578218 252986 578454
rect 253222 578218 288986 578454
rect 289222 578218 324986 578454
rect 325222 578218 360986 578454
rect 361222 578218 396986 578454
rect 397222 578218 432986 578454
rect 433222 578218 468986 578454
rect 469222 578218 504986 578454
rect 505222 578218 540986 578454
rect 541222 578218 576986 578454
rect 577222 578218 585502 578454
rect 585738 578218 586840 578454
rect -2916 578134 586840 578218
rect -2916 577898 -1814 578134
rect -1578 577898 986 578134
rect 1222 577898 36986 578134
rect 37222 577898 72986 578134
rect 73222 577898 108986 578134
rect 109222 577898 144986 578134
rect 145222 577898 180986 578134
rect 181222 577898 216986 578134
rect 217222 577898 252986 578134
rect 253222 577898 288986 578134
rect 289222 577898 324986 578134
rect 325222 577898 360986 578134
rect 361222 577898 396986 578134
rect 397222 577898 432986 578134
rect 433222 577898 468986 578134
rect 469222 577898 504986 578134
rect 505222 577898 540986 578134
rect 541222 577898 576986 578134
rect 577222 577898 585502 578134
rect 585738 577898 586840 578134
rect -2916 577876 586840 577898
rect -1996 577874 -1396 577876
rect 804 577874 1404 577876
rect 36804 577874 37404 577876
rect 72804 577874 73404 577876
rect 108804 577874 109404 577876
rect 144804 577874 145404 577876
rect 180804 577874 181404 577876
rect 216804 577874 217404 577876
rect 252804 577874 253404 577876
rect 288804 577874 289404 577876
rect 324804 577874 325404 577876
rect 360804 577874 361404 577876
rect 396804 577874 397404 577876
rect 432804 577874 433404 577876
rect 468804 577874 469404 577876
rect 504804 577874 505404 577876
rect 540804 577874 541404 577876
rect 576804 577874 577404 577876
rect 585320 577874 585920 577876
rect -8436 571276 -7836 571278
rect 29604 571276 30204 571278
rect 65604 571276 66204 571278
rect 101604 571276 102204 571278
rect 137604 571276 138204 571278
rect 173604 571276 174204 571278
rect 209604 571276 210204 571278
rect 245604 571276 246204 571278
rect 281604 571276 282204 571278
rect 317604 571276 318204 571278
rect 353604 571276 354204 571278
rect 389604 571276 390204 571278
rect 425604 571276 426204 571278
rect 461604 571276 462204 571278
rect 497604 571276 498204 571278
rect 533604 571276 534204 571278
rect 569604 571276 570204 571278
rect 591760 571276 592360 571278
rect -8436 571254 592360 571276
rect -8436 571018 -8254 571254
rect -8018 571018 29786 571254
rect 30022 571018 65786 571254
rect 66022 571018 101786 571254
rect 102022 571018 137786 571254
rect 138022 571018 173786 571254
rect 174022 571018 209786 571254
rect 210022 571018 245786 571254
rect 246022 571018 281786 571254
rect 282022 571018 317786 571254
rect 318022 571018 353786 571254
rect 354022 571018 389786 571254
rect 390022 571018 425786 571254
rect 426022 571018 461786 571254
rect 462022 571018 497786 571254
rect 498022 571018 533786 571254
rect 534022 571018 569786 571254
rect 570022 571018 591942 571254
rect 592178 571018 592360 571254
rect -8436 570934 592360 571018
rect -8436 570698 -8254 570934
rect -8018 570698 29786 570934
rect 30022 570698 65786 570934
rect 66022 570698 101786 570934
rect 102022 570698 137786 570934
rect 138022 570698 173786 570934
rect 174022 570698 209786 570934
rect 210022 570698 245786 570934
rect 246022 570698 281786 570934
rect 282022 570698 317786 570934
rect 318022 570698 353786 570934
rect 354022 570698 389786 570934
rect 390022 570698 425786 570934
rect 426022 570698 461786 570934
rect 462022 570698 497786 570934
rect 498022 570698 533786 570934
rect 534022 570698 569786 570934
rect 570022 570698 591942 570934
rect 592178 570698 592360 570934
rect -8436 570676 592360 570698
rect -8436 570674 -7836 570676
rect 29604 570674 30204 570676
rect 65604 570674 66204 570676
rect 101604 570674 102204 570676
rect 137604 570674 138204 570676
rect 173604 570674 174204 570676
rect 209604 570674 210204 570676
rect 245604 570674 246204 570676
rect 281604 570674 282204 570676
rect 317604 570674 318204 570676
rect 353604 570674 354204 570676
rect 389604 570674 390204 570676
rect 425604 570674 426204 570676
rect 461604 570674 462204 570676
rect 497604 570674 498204 570676
rect 533604 570674 534204 570676
rect 569604 570674 570204 570676
rect 591760 570674 592360 570676
rect -6596 567676 -5996 567678
rect 26004 567676 26604 567678
rect 62004 567676 62604 567678
rect 98004 567676 98604 567678
rect 134004 567676 134604 567678
rect 170004 567676 170604 567678
rect 206004 567676 206604 567678
rect 242004 567676 242604 567678
rect 278004 567676 278604 567678
rect 314004 567676 314604 567678
rect 350004 567676 350604 567678
rect 386004 567676 386604 567678
rect 422004 567676 422604 567678
rect 458004 567676 458604 567678
rect 494004 567676 494604 567678
rect 530004 567676 530604 567678
rect 566004 567676 566604 567678
rect 589920 567676 590520 567678
rect -6596 567654 590520 567676
rect -6596 567418 -6414 567654
rect -6178 567418 26186 567654
rect 26422 567418 62186 567654
rect 62422 567418 98186 567654
rect 98422 567418 134186 567654
rect 134422 567418 170186 567654
rect 170422 567418 206186 567654
rect 206422 567418 242186 567654
rect 242422 567418 278186 567654
rect 278422 567418 314186 567654
rect 314422 567418 350186 567654
rect 350422 567418 386186 567654
rect 386422 567418 422186 567654
rect 422422 567418 458186 567654
rect 458422 567418 494186 567654
rect 494422 567418 530186 567654
rect 530422 567418 566186 567654
rect 566422 567418 590102 567654
rect 590338 567418 590520 567654
rect -6596 567334 590520 567418
rect -6596 567098 -6414 567334
rect -6178 567098 26186 567334
rect 26422 567098 62186 567334
rect 62422 567098 98186 567334
rect 98422 567098 134186 567334
rect 134422 567098 170186 567334
rect 170422 567098 206186 567334
rect 206422 567098 242186 567334
rect 242422 567098 278186 567334
rect 278422 567098 314186 567334
rect 314422 567098 350186 567334
rect 350422 567098 386186 567334
rect 386422 567098 422186 567334
rect 422422 567098 458186 567334
rect 458422 567098 494186 567334
rect 494422 567098 530186 567334
rect 530422 567098 566186 567334
rect 566422 567098 590102 567334
rect 590338 567098 590520 567334
rect -6596 567076 590520 567098
rect -6596 567074 -5996 567076
rect 26004 567074 26604 567076
rect 62004 567074 62604 567076
rect 98004 567074 98604 567076
rect 134004 567074 134604 567076
rect 170004 567074 170604 567076
rect 206004 567074 206604 567076
rect 242004 567074 242604 567076
rect 278004 567074 278604 567076
rect 314004 567074 314604 567076
rect 350004 567074 350604 567076
rect 386004 567074 386604 567076
rect 422004 567074 422604 567076
rect 458004 567074 458604 567076
rect 494004 567074 494604 567076
rect 530004 567074 530604 567076
rect 566004 567074 566604 567076
rect 589920 567074 590520 567076
rect -4756 564076 -4156 564078
rect 22404 564076 23004 564078
rect 58404 564076 59004 564078
rect 94404 564076 95004 564078
rect 130404 564076 131004 564078
rect 166404 564076 167004 564078
rect 202404 564076 203004 564078
rect 238404 564076 239004 564078
rect 274404 564076 275004 564078
rect 310404 564076 311004 564078
rect 346404 564076 347004 564078
rect 382404 564076 383004 564078
rect 418404 564076 419004 564078
rect 454404 564076 455004 564078
rect 490404 564076 491004 564078
rect 526404 564076 527004 564078
rect 562404 564076 563004 564078
rect 588080 564076 588680 564078
rect -4756 564054 588680 564076
rect -4756 563818 -4574 564054
rect -4338 563818 22586 564054
rect 22822 563818 58586 564054
rect 58822 563818 94586 564054
rect 94822 563818 130586 564054
rect 130822 563818 166586 564054
rect 166822 563818 202586 564054
rect 202822 563818 238586 564054
rect 238822 563818 274586 564054
rect 274822 563818 310586 564054
rect 310822 563818 346586 564054
rect 346822 563818 382586 564054
rect 382822 563818 418586 564054
rect 418822 563818 454586 564054
rect 454822 563818 490586 564054
rect 490822 563818 526586 564054
rect 526822 563818 562586 564054
rect 562822 563818 588262 564054
rect 588498 563818 588680 564054
rect -4756 563734 588680 563818
rect -4756 563498 -4574 563734
rect -4338 563498 22586 563734
rect 22822 563498 58586 563734
rect 58822 563498 94586 563734
rect 94822 563498 130586 563734
rect 130822 563498 166586 563734
rect 166822 563498 202586 563734
rect 202822 563498 238586 563734
rect 238822 563498 274586 563734
rect 274822 563498 310586 563734
rect 310822 563498 346586 563734
rect 346822 563498 382586 563734
rect 382822 563498 418586 563734
rect 418822 563498 454586 563734
rect 454822 563498 490586 563734
rect 490822 563498 526586 563734
rect 526822 563498 562586 563734
rect 562822 563498 588262 563734
rect 588498 563498 588680 563734
rect -4756 563476 588680 563498
rect -4756 563474 -4156 563476
rect 22404 563474 23004 563476
rect 58404 563474 59004 563476
rect 94404 563474 95004 563476
rect 130404 563474 131004 563476
rect 166404 563474 167004 563476
rect 202404 563474 203004 563476
rect 238404 563474 239004 563476
rect 274404 563474 275004 563476
rect 310404 563474 311004 563476
rect 346404 563474 347004 563476
rect 382404 563474 383004 563476
rect 418404 563474 419004 563476
rect 454404 563474 455004 563476
rect 490404 563474 491004 563476
rect 526404 563474 527004 563476
rect 562404 563474 563004 563476
rect 588080 563474 588680 563476
rect -2916 560476 -2316 560478
rect 18804 560476 19404 560478
rect 54804 560476 55404 560478
rect 90804 560476 91404 560478
rect 126804 560476 127404 560478
rect 162804 560476 163404 560478
rect 198804 560476 199404 560478
rect 234804 560476 235404 560478
rect 270804 560476 271404 560478
rect 306804 560476 307404 560478
rect 342804 560476 343404 560478
rect 378804 560476 379404 560478
rect 414804 560476 415404 560478
rect 450804 560476 451404 560478
rect 486804 560476 487404 560478
rect 522804 560476 523404 560478
rect 558804 560476 559404 560478
rect 586240 560476 586840 560478
rect -2916 560454 586840 560476
rect -2916 560218 -2734 560454
rect -2498 560218 18986 560454
rect 19222 560218 54986 560454
rect 55222 560218 90986 560454
rect 91222 560218 126986 560454
rect 127222 560218 162986 560454
rect 163222 560218 198986 560454
rect 199222 560218 234986 560454
rect 235222 560218 270986 560454
rect 271222 560218 306986 560454
rect 307222 560218 342986 560454
rect 343222 560218 378986 560454
rect 379222 560218 414986 560454
rect 415222 560218 450986 560454
rect 451222 560218 486986 560454
rect 487222 560218 522986 560454
rect 523222 560218 558986 560454
rect 559222 560218 586422 560454
rect 586658 560218 586840 560454
rect -2916 560134 586840 560218
rect -2916 559898 -2734 560134
rect -2498 559898 18986 560134
rect 19222 559898 54986 560134
rect 55222 559898 90986 560134
rect 91222 559898 126986 560134
rect 127222 559898 162986 560134
rect 163222 559898 198986 560134
rect 199222 559898 234986 560134
rect 235222 559898 270986 560134
rect 271222 559898 306986 560134
rect 307222 559898 342986 560134
rect 343222 559898 378986 560134
rect 379222 559898 414986 560134
rect 415222 559898 450986 560134
rect 451222 559898 486986 560134
rect 487222 559898 522986 560134
rect 523222 559898 558986 560134
rect 559222 559898 586422 560134
rect 586658 559898 586840 560134
rect -2916 559876 586840 559898
rect -2916 559874 -2316 559876
rect 18804 559874 19404 559876
rect 54804 559874 55404 559876
rect 90804 559874 91404 559876
rect 126804 559874 127404 559876
rect 162804 559874 163404 559876
rect 198804 559874 199404 559876
rect 234804 559874 235404 559876
rect 270804 559874 271404 559876
rect 306804 559874 307404 559876
rect 342804 559874 343404 559876
rect 378804 559874 379404 559876
rect 414804 559874 415404 559876
rect 450804 559874 451404 559876
rect 486804 559874 487404 559876
rect 522804 559874 523404 559876
rect 558804 559874 559404 559876
rect 586240 559874 586840 559876
rect -7516 553276 -6916 553278
rect 11604 553276 12204 553278
rect 47604 553276 48204 553278
rect 83604 553276 84204 553278
rect 119604 553276 120204 553278
rect 155604 553276 156204 553278
rect 191604 553276 192204 553278
rect 227604 553276 228204 553278
rect 263604 553276 264204 553278
rect 299604 553276 300204 553278
rect 335604 553276 336204 553278
rect 371604 553276 372204 553278
rect 407604 553276 408204 553278
rect 443604 553276 444204 553278
rect 479604 553276 480204 553278
rect 515604 553276 516204 553278
rect 551604 553276 552204 553278
rect 590840 553276 591440 553278
rect -8436 553254 592360 553276
rect -8436 553018 -7334 553254
rect -7098 553018 11786 553254
rect 12022 553018 47786 553254
rect 48022 553018 83786 553254
rect 84022 553018 119786 553254
rect 120022 553018 155786 553254
rect 156022 553018 191786 553254
rect 192022 553018 227786 553254
rect 228022 553018 263786 553254
rect 264022 553018 299786 553254
rect 300022 553018 335786 553254
rect 336022 553018 371786 553254
rect 372022 553018 407786 553254
rect 408022 553018 443786 553254
rect 444022 553018 479786 553254
rect 480022 553018 515786 553254
rect 516022 553018 551786 553254
rect 552022 553018 591022 553254
rect 591258 553018 592360 553254
rect -8436 552934 592360 553018
rect -8436 552698 -7334 552934
rect -7098 552698 11786 552934
rect 12022 552698 47786 552934
rect 48022 552698 83786 552934
rect 84022 552698 119786 552934
rect 120022 552698 155786 552934
rect 156022 552698 191786 552934
rect 192022 552698 227786 552934
rect 228022 552698 263786 552934
rect 264022 552698 299786 552934
rect 300022 552698 335786 552934
rect 336022 552698 371786 552934
rect 372022 552698 407786 552934
rect 408022 552698 443786 552934
rect 444022 552698 479786 552934
rect 480022 552698 515786 552934
rect 516022 552698 551786 552934
rect 552022 552698 591022 552934
rect 591258 552698 592360 552934
rect -8436 552676 592360 552698
rect -7516 552674 -6916 552676
rect 11604 552674 12204 552676
rect 47604 552674 48204 552676
rect 83604 552674 84204 552676
rect 119604 552674 120204 552676
rect 155604 552674 156204 552676
rect 191604 552674 192204 552676
rect 227604 552674 228204 552676
rect 263604 552674 264204 552676
rect 299604 552674 300204 552676
rect 335604 552674 336204 552676
rect 371604 552674 372204 552676
rect 407604 552674 408204 552676
rect 443604 552674 444204 552676
rect 479604 552674 480204 552676
rect 515604 552674 516204 552676
rect 551604 552674 552204 552676
rect 590840 552674 591440 552676
rect -5676 549676 -5076 549678
rect 8004 549676 8604 549678
rect 44004 549676 44604 549678
rect 80004 549676 80604 549678
rect 116004 549676 116604 549678
rect 152004 549676 152604 549678
rect 188004 549676 188604 549678
rect 224004 549676 224604 549678
rect 260004 549676 260604 549678
rect 296004 549676 296604 549678
rect 332004 549676 332604 549678
rect 368004 549676 368604 549678
rect 404004 549676 404604 549678
rect 440004 549676 440604 549678
rect 476004 549676 476604 549678
rect 512004 549676 512604 549678
rect 548004 549676 548604 549678
rect 589000 549676 589600 549678
rect -6596 549654 590520 549676
rect -6596 549418 -5494 549654
rect -5258 549418 8186 549654
rect 8422 549418 44186 549654
rect 44422 549418 80186 549654
rect 80422 549418 116186 549654
rect 116422 549418 152186 549654
rect 152422 549418 188186 549654
rect 188422 549418 224186 549654
rect 224422 549418 260186 549654
rect 260422 549418 296186 549654
rect 296422 549418 332186 549654
rect 332422 549418 368186 549654
rect 368422 549418 404186 549654
rect 404422 549418 440186 549654
rect 440422 549418 476186 549654
rect 476422 549418 512186 549654
rect 512422 549418 548186 549654
rect 548422 549418 589182 549654
rect 589418 549418 590520 549654
rect -6596 549334 590520 549418
rect -6596 549098 -5494 549334
rect -5258 549098 8186 549334
rect 8422 549098 44186 549334
rect 44422 549098 80186 549334
rect 80422 549098 116186 549334
rect 116422 549098 152186 549334
rect 152422 549098 188186 549334
rect 188422 549098 224186 549334
rect 224422 549098 260186 549334
rect 260422 549098 296186 549334
rect 296422 549098 332186 549334
rect 332422 549098 368186 549334
rect 368422 549098 404186 549334
rect 404422 549098 440186 549334
rect 440422 549098 476186 549334
rect 476422 549098 512186 549334
rect 512422 549098 548186 549334
rect 548422 549098 589182 549334
rect 589418 549098 590520 549334
rect -6596 549076 590520 549098
rect -5676 549074 -5076 549076
rect 8004 549074 8604 549076
rect 44004 549074 44604 549076
rect 80004 549074 80604 549076
rect 116004 549074 116604 549076
rect 152004 549074 152604 549076
rect 188004 549074 188604 549076
rect 224004 549074 224604 549076
rect 260004 549074 260604 549076
rect 296004 549074 296604 549076
rect 332004 549074 332604 549076
rect 368004 549074 368604 549076
rect 404004 549074 404604 549076
rect 440004 549074 440604 549076
rect 476004 549074 476604 549076
rect 512004 549074 512604 549076
rect 548004 549074 548604 549076
rect 589000 549074 589600 549076
rect -3836 546076 -3236 546078
rect 4404 546076 5004 546078
rect 40404 546076 41004 546078
rect 76404 546076 77004 546078
rect 112404 546076 113004 546078
rect 148404 546076 149004 546078
rect 184404 546076 185004 546078
rect 220404 546076 221004 546078
rect 256404 546076 257004 546078
rect 292404 546076 293004 546078
rect 328404 546076 329004 546078
rect 364404 546076 365004 546078
rect 400404 546076 401004 546078
rect 436404 546076 437004 546078
rect 472404 546076 473004 546078
rect 508404 546076 509004 546078
rect 544404 546076 545004 546078
rect 580404 546076 581004 546078
rect 587160 546076 587760 546078
rect -4756 546054 588680 546076
rect -4756 545818 -3654 546054
rect -3418 545818 4586 546054
rect 4822 545818 40586 546054
rect 40822 545818 76586 546054
rect 76822 545818 112586 546054
rect 112822 545818 148586 546054
rect 148822 545818 184586 546054
rect 184822 545818 220586 546054
rect 220822 545818 256586 546054
rect 256822 545818 292586 546054
rect 292822 545818 328586 546054
rect 328822 545818 364586 546054
rect 364822 545818 400586 546054
rect 400822 545818 436586 546054
rect 436822 545818 472586 546054
rect 472822 545818 508586 546054
rect 508822 545818 544586 546054
rect 544822 545818 580586 546054
rect 580822 545818 587342 546054
rect 587578 545818 588680 546054
rect -4756 545734 588680 545818
rect -4756 545498 -3654 545734
rect -3418 545498 4586 545734
rect 4822 545498 40586 545734
rect 40822 545498 76586 545734
rect 76822 545498 112586 545734
rect 112822 545498 148586 545734
rect 148822 545498 184586 545734
rect 184822 545498 220586 545734
rect 220822 545498 256586 545734
rect 256822 545498 292586 545734
rect 292822 545498 328586 545734
rect 328822 545498 364586 545734
rect 364822 545498 400586 545734
rect 400822 545498 436586 545734
rect 436822 545498 472586 545734
rect 472822 545498 508586 545734
rect 508822 545498 544586 545734
rect 544822 545498 580586 545734
rect 580822 545498 587342 545734
rect 587578 545498 588680 545734
rect -4756 545476 588680 545498
rect -3836 545474 -3236 545476
rect 4404 545474 5004 545476
rect 40404 545474 41004 545476
rect 76404 545474 77004 545476
rect 112404 545474 113004 545476
rect 148404 545474 149004 545476
rect 184404 545474 185004 545476
rect 220404 545474 221004 545476
rect 256404 545474 257004 545476
rect 292404 545474 293004 545476
rect 328404 545474 329004 545476
rect 364404 545474 365004 545476
rect 400404 545474 401004 545476
rect 436404 545474 437004 545476
rect 472404 545474 473004 545476
rect 508404 545474 509004 545476
rect 544404 545474 545004 545476
rect 580404 545474 581004 545476
rect 587160 545474 587760 545476
rect -1996 542476 -1396 542478
rect 804 542476 1404 542478
rect 36804 542476 37404 542478
rect 72804 542476 73404 542478
rect 108804 542476 109404 542478
rect 144804 542476 145404 542478
rect 180804 542476 181404 542478
rect 216804 542476 217404 542478
rect 252804 542476 253404 542478
rect 288804 542476 289404 542478
rect 324804 542476 325404 542478
rect 360804 542476 361404 542478
rect 396804 542476 397404 542478
rect 432804 542476 433404 542478
rect 468804 542476 469404 542478
rect 504804 542476 505404 542478
rect 540804 542476 541404 542478
rect 576804 542476 577404 542478
rect 585320 542476 585920 542478
rect -2916 542454 586840 542476
rect -2916 542218 -1814 542454
rect -1578 542218 986 542454
rect 1222 542218 36986 542454
rect 37222 542218 72986 542454
rect 73222 542218 108986 542454
rect 109222 542218 144986 542454
rect 145222 542218 180986 542454
rect 181222 542218 216986 542454
rect 217222 542218 252986 542454
rect 253222 542218 288986 542454
rect 289222 542218 324986 542454
rect 325222 542218 360986 542454
rect 361222 542218 396986 542454
rect 397222 542218 432986 542454
rect 433222 542218 468986 542454
rect 469222 542218 504986 542454
rect 505222 542218 540986 542454
rect 541222 542218 576986 542454
rect 577222 542218 585502 542454
rect 585738 542218 586840 542454
rect -2916 542134 586840 542218
rect -2916 541898 -1814 542134
rect -1578 541898 986 542134
rect 1222 541898 36986 542134
rect 37222 541898 72986 542134
rect 73222 541898 108986 542134
rect 109222 541898 144986 542134
rect 145222 541898 180986 542134
rect 181222 541898 216986 542134
rect 217222 541898 252986 542134
rect 253222 541898 288986 542134
rect 289222 541898 324986 542134
rect 325222 541898 360986 542134
rect 361222 541898 396986 542134
rect 397222 541898 432986 542134
rect 433222 541898 468986 542134
rect 469222 541898 504986 542134
rect 505222 541898 540986 542134
rect 541222 541898 576986 542134
rect 577222 541898 585502 542134
rect 585738 541898 586840 542134
rect -2916 541876 586840 541898
rect -1996 541874 -1396 541876
rect 804 541874 1404 541876
rect 36804 541874 37404 541876
rect 72804 541874 73404 541876
rect 108804 541874 109404 541876
rect 144804 541874 145404 541876
rect 180804 541874 181404 541876
rect 216804 541874 217404 541876
rect 252804 541874 253404 541876
rect 288804 541874 289404 541876
rect 324804 541874 325404 541876
rect 360804 541874 361404 541876
rect 396804 541874 397404 541876
rect 432804 541874 433404 541876
rect 468804 541874 469404 541876
rect 504804 541874 505404 541876
rect 540804 541874 541404 541876
rect 576804 541874 577404 541876
rect 585320 541874 585920 541876
rect -8436 535276 -7836 535278
rect 29604 535276 30204 535278
rect 65604 535276 66204 535278
rect 101604 535276 102204 535278
rect 137604 535276 138204 535278
rect 173604 535276 174204 535278
rect 209604 535276 210204 535278
rect 245604 535276 246204 535278
rect 281604 535276 282204 535278
rect 317604 535276 318204 535278
rect 353604 535276 354204 535278
rect 389604 535276 390204 535278
rect 425604 535276 426204 535278
rect 461604 535276 462204 535278
rect 497604 535276 498204 535278
rect 533604 535276 534204 535278
rect 569604 535276 570204 535278
rect 591760 535276 592360 535278
rect -8436 535254 592360 535276
rect -8436 535018 -8254 535254
rect -8018 535018 29786 535254
rect 30022 535018 65786 535254
rect 66022 535018 101786 535254
rect 102022 535018 137786 535254
rect 138022 535018 173786 535254
rect 174022 535018 209786 535254
rect 210022 535018 245786 535254
rect 246022 535018 281786 535254
rect 282022 535018 317786 535254
rect 318022 535018 353786 535254
rect 354022 535018 389786 535254
rect 390022 535018 425786 535254
rect 426022 535018 461786 535254
rect 462022 535018 497786 535254
rect 498022 535018 533786 535254
rect 534022 535018 569786 535254
rect 570022 535018 591942 535254
rect 592178 535018 592360 535254
rect -8436 534934 592360 535018
rect -8436 534698 -8254 534934
rect -8018 534698 29786 534934
rect 30022 534698 65786 534934
rect 66022 534698 101786 534934
rect 102022 534698 137786 534934
rect 138022 534698 173786 534934
rect 174022 534698 209786 534934
rect 210022 534698 245786 534934
rect 246022 534698 281786 534934
rect 282022 534698 317786 534934
rect 318022 534698 353786 534934
rect 354022 534698 389786 534934
rect 390022 534698 425786 534934
rect 426022 534698 461786 534934
rect 462022 534698 497786 534934
rect 498022 534698 533786 534934
rect 534022 534698 569786 534934
rect 570022 534698 591942 534934
rect 592178 534698 592360 534934
rect -8436 534676 592360 534698
rect -8436 534674 -7836 534676
rect 29604 534674 30204 534676
rect 65604 534674 66204 534676
rect 101604 534674 102204 534676
rect 137604 534674 138204 534676
rect 173604 534674 174204 534676
rect 209604 534674 210204 534676
rect 245604 534674 246204 534676
rect 281604 534674 282204 534676
rect 317604 534674 318204 534676
rect 353604 534674 354204 534676
rect 389604 534674 390204 534676
rect 425604 534674 426204 534676
rect 461604 534674 462204 534676
rect 497604 534674 498204 534676
rect 533604 534674 534204 534676
rect 569604 534674 570204 534676
rect 591760 534674 592360 534676
rect -6596 531676 -5996 531678
rect 26004 531676 26604 531678
rect 62004 531676 62604 531678
rect 98004 531676 98604 531678
rect 134004 531676 134604 531678
rect 170004 531676 170604 531678
rect 206004 531676 206604 531678
rect 242004 531676 242604 531678
rect 278004 531676 278604 531678
rect 314004 531676 314604 531678
rect 350004 531676 350604 531678
rect 386004 531676 386604 531678
rect 422004 531676 422604 531678
rect 458004 531676 458604 531678
rect 494004 531676 494604 531678
rect 530004 531676 530604 531678
rect 566004 531676 566604 531678
rect 589920 531676 590520 531678
rect -6596 531654 590520 531676
rect -6596 531418 -6414 531654
rect -6178 531418 26186 531654
rect 26422 531418 62186 531654
rect 62422 531418 98186 531654
rect 98422 531418 134186 531654
rect 134422 531418 170186 531654
rect 170422 531418 206186 531654
rect 206422 531418 242186 531654
rect 242422 531418 278186 531654
rect 278422 531418 314186 531654
rect 314422 531418 350186 531654
rect 350422 531418 386186 531654
rect 386422 531418 422186 531654
rect 422422 531418 458186 531654
rect 458422 531418 494186 531654
rect 494422 531418 530186 531654
rect 530422 531418 566186 531654
rect 566422 531418 590102 531654
rect 590338 531418 590520 531654
rect -6596 531334 590520 531418
rect -6596 531098 -6414 531334
rect -6178 531098 26186 531334
rect 26422 531098 62186 531334
rect 62422 531098 98186 531334
rect 98422 531098 134186 531334
rect 134422 531098 170186 531334
rect 170422 531098 206186 531334
rect 206422 531098 242186 531334
rect 242422 531098 278186 531334
rect 278422 531098 314186 531334
rect 314422 531098 350186 531334
rect 350422 531098 386186 531334
rect 386422 531098 422186 531334
rect 422422 531098 458186 531334
rect 458422 531098 494186 531334
rect 494422 531098 530186 531334
rect 530422 531098 566186 531334
rect 566422 531098 590102 531334
rect 590338 531098 590520 531334
rect -6596 531076 590520 531098
rect -6596 531074 -5996 531076
rect 26004 531074 26604 531076
rect 62004 531074 62604 531076
rect 98004 531074 98604 531076
rect 134004 531074 134604 531076
rect 170004 531074 170604 531076
rect 206004 531074 206604 531076
rect 242004 531074 242604 531076
rect 278004 531074 278604 531076
rect 314004 531074 314604 531076
rect 350004 531074 350604 531076
rect 386004 531074 386604 531076
rect 422004 531074 422604 531076
rect 458004 531074 458604 531076
rect 494004 531074 494604 531076
rect 530004 531074 530604 531076
rect 566004 531074 566604 531076
rect 589920 531074 590520 531076
rect -4756 528076 -4156 528078
rect 22404 528076 23004 528078
rect 58404 528076 59004 528078
rect 94404 528076 95004 528078
rect 130404 528076 131004 528078
rect 166404 528076 167004 528078
rect 202404 528076 203004 528078
rect 238404 528076 239004 528078
rect 274404 528076 275004 528078
rect 310404 528076 311004 528078
rect 346404 528076 347004 528078
rect 382404 528076 383004 528078
rect 418404 528076 419004 528078
rect 454404 528076 455004 528078
rect 490404 528076 491004 528078
rect 526404 528076 527004 528078
rect 562404 528076 563004 528078
rect 588080 528076 588680 528078
rect -4756 528054 588680 528076
rect -4756 527818 -4574 528054
rect -4338 527818 22586 528054
rect 22822 527818 58586 528054
rect 58822 527818 94586 528054
rect 94822 527818 130586 528054
rect 130822 527818 166586 528054
rect 166822 527818 202586 528054
rect 202822 527818 238586 528054
rect 238822 527818 274586 528054
rect 274822 527818 310586 528054
rect 310822 527818 346586 528054
rect 346822 527818 382586 528054
rect 382822 527818 418586 528054
rect 418822 527818 454586 528054
rect 454822 527818 490586 528054
rect 490822 527818 526586 528054
rect 526822 527818 562586 528054
rect 562822 527818 588262 528054
rect 588498 527818 588680 528054
rect -4756 527734 588680 527818
rect -4756 527498 -4574 527734
rect -4338 527498 22586 527734
rect 22822 527498 58586 527734
rect 58822 527498 94586 527734
rect 94822 527498 130586 527734
rect 130822 527498 166586 527734
rect 166822 527498 202586 527734
rect 202822 527498 238586 527734
rect 238822 527498 274586 527734
rect 274822 527498 310586 527734
rect 310822 527498 346586 527734
rect 346822 527498 382586 527734
rect 382822 527498 418586 527734
rect 418822 527498 454586 527734
rect 454822 527498 490586 527734
rect 490822 527498 526586 527734
rect 526822 527498 562586 527734
rect 562822 527498 588262 527734
rect 588498 527498 588680 527734
rect -4756 527476 588680 527498
rect -4756 527474 -4156 527476
rect 22404 527474 23004 527476
rect 58404 527474 59004 527476
rect 94404 527474 95004 527476
rect 130404 527474 131004 527476
rect 166404 527474 167004 527476
rect 202404 527474 203004 527476
rect 238404 527474 239004 527476
rect 274404 527474 275004 527476
rect 310404 527474 311004 527476
rect 346404 527474 347004 527476
rect 382404 527474 383004 527476
rect 418404 527474 419004 527476
rect 454404 527474 455004 527476
rect 490404 527474 491004 527476
rect 526404 527474 527004 527476
rect 562404 527474 563004 527476
rect 588080 527474 588680 527476
rect -2916 524476 -2316 524478
rect 18804 524476 19404 524478
rect 54804 524476 55404 524478
rect 90804 524476 91404 524478
rect 126804 524476 127404 524478
rect 162804 524476 163404 524478
rect 198804 524476 199404 524478
rect 234804 524476 235404 524478
rect 270804 524476 271404 524478
rect 306804 524476 307404 524478
rect 342804 524476 343404 524478
rect 378804 524476 379404 524478
rect 414804 524476 415404 524478
rect 450804 524476 451404 524478
rect 486804 524476 487404 524478
rect 522804 524476 523404 524478
rect 558804 524476 559404 524478
rect 586240 524476 586840 524478
rect -2916 524454 586840 524476
rect -2916 524218 -2734 524454
rect -2498 524218 18986 524454
rect 19222 524218 54986 524454
rect 55222 524218 90986 524454
rect 91222 524218 126986 524454
rect 127222 524218 162986 524454
rect 163222 524218 198986 524454
rect 199222 524218 234986 524454
rect 235222 524218 270986 524454
rect 271222 524218 306986 524454
rect 307222 524218 342986 524454
rect 343222 524218 378986 524454
rect 379222 524218 414986 524454
rect 415222 524218 450986 524454
rect 451222 524218 486986 524454
rect 487222 524218 522986 524454
rect 523222 524218 558986 524454
rect 559222 524218 586422 524454
rect 586658 524218 586840 524454
rect -2916 524134 586840 524218
rect -2916 523898 -2734 524134
rect -2498 523898 18986 524134
rect 19222 523898 54986 524134
rect 55222 523898 90986 524134
rect 91222 523898 126986 524134
rect 127222 523898 162986 524134
rect 163222 523898 198986 524134
rect 199222 523898 234986 524134
rect 235222 523898 270986 524134
rect 271222 523898 306986 524134
rect 307222 523898 342986 524134
rect 343222 523898 378986 524134
rect 379222 523898 414986 524134
rect 415222 523898 450986 524134
rect 451222 523898 486986 524134
rect 487222 523898 522986 524134
rect 523222 523898 558986 524134
rect 559222 523898 586422 524134
rect 586658 523898 586840 524134
rect -2916 523876 586840 523898
rect -2916 523874 -2316 523876
rect 18804 523874 19404 523876
rect 54804 523874 55404 523876
rect 90804 523874 91404 523876
rect 126804 523874 127404 523876
rect 162804 523874 163404 523876
rect 198804 523874 199404 523876
rect 234804 523874 235404 523876
rect 270804 523874 271404 523876
rect 306804 523874 307404 523876
rect 342804 523874 343404 523876
rect 378804 523874 379404 523876
rect 414804 523874 415404 523876
rect 450804 523874 451404 523876
rect 486804 523874 487404 523876
rect 522804 523874 523404 523876
rect 558804 523874 559404 523876
rect 586240 523874 586840 523876
rect -7516 517276 -6916 517278
rect 11604 517276 12204 517278
rect 47604 517276 48204 517278
rect 83604 517276 84204 517278
rect 119604 517276 120204 517278
rect 155604 517276 156204 517278
rect 191604 517276 192204 517278
rect 227604 517276 228204 517278
rect 263604 517276 264204 517278
rect 299604 517276 300204 517278
rect 335604 517276 336204 517278
rect 371604 517276 372204 517278
rect 407604 517276 408204 517278
rect 443604 517276 444204 517278
rect 479604 517276 480204 517278
rect 515604 517276 516204 517278
rect 551604 517276 552204 517278
rect 590840 517276 591440 517278
rect -8436 517254 592360 517276
rect -8436 517018 -7334 517254
rect -7098 517018 11786 517254
rect 12022 517018 47786 517254
rect 48022 517018 83786 517254
rect 84022 517018 119786 517254
rect 120022 517018 155786 517254
rect 156022 517018 191786 517254
rect 192022 517018 227786 517254
rect 228022 517018 263786 517254
rect 264022 517018 299786 517254
rect 300022 517018 335786 517254
rect 336022 517018 371786 517254
rect 372022 517018 407786 517254
rect 408022 517018 443786 517254
rect 444022 517018 479786 517254
rect 480022 517018 515786 517254
rect 516022 517018 551786 517254
rect 552022 517018 591022 517254
rect 591258 517018 592360 517254
rect -8436 516934 592360 517018
rect -8436 516698 -7334 516934
rect -7098 516698 11786 516934
rect 12022 516698 47786 516934
rect 48022 516698 83786 516934
rect 84022 516698 119786 516934
rect 120022 516698 155786 516934
rect 156022 516698 191786 516934
rect 192022 516698 227786 516934
rect 228022 516698 263786 516934
rect 264022 516698 299786 516934
rect 300022 516698 335786 516934
rect 336022 516698 371786 516934
rect 372022 516698 407786 516934
rect 408022 516698 443786 516934
rect 444022 516698 479786 516934
rect 480022 516698 515786 516934
rect 516022 516698 551786 516934
rect 552022 516698 591022 516934
rect 591258 516698 592360 516934
rect -8436 516676 592360 516698
rect -7516 516674 -6916 516676
rect 11604 516674 12204 516676
rect 47604 516674 48204 516676
rect 83604 516674 84204 516676
rect 119604 516674 120204 516676
rect 155604 516674 156204 516676
rect 191604 516674 192204 516676
rect 227604 516674 228204 516676
rect 263604 516674 264204 516676
rect 299604 516674 300204 516676
rect 335604 516674 336204 516676
rect 371604 516674 372204 516676
rect 407604 516674 408204 516676
rect 443604 516674 444204 516676
rect 479604 516674 480204 516676
rect 515604 516674 516204 516676
rect 551604 516674 552204 516676
rect 590840 516674 591440 516676
rect -5676 513676 -5076 513678
rect 8004 513676 8604 513678
rect 44004 513676 44604 513678
rect 80004 513676 80604 513678
rect 116004 513676 116604 513678
rect 152004 513676 152604 513678
rect 188004 513676 188604 513678
rect 224004 513676 224604 513678
rect 260004 513676 260604 513678
rect 296004 513676 296604 513678
rect 332004 513676 332604 513678
rect 368004 513676 368604 513678
rect 404004 513676 404604 513678
rect 440004 513676 440604 513678
rect 476004 513676 476604 513678
rect 512004 513676 512604 513678
rect 548004 513676 548604 513678
rect 589000 513676 589600 513678
rect -6596 513654 590520 513676
rect -6596 513418 -5494 513654
rect -5258 513418 8186 513654
rect 8422 513418 44186 513654
rect 44422 513418 80186 513654
rect 80422 513418 116186 513654
rect 116422 513418 152186 513654
rect 152422 513418 188186 513654
rect 188422 513418 224186 513654
rect 224422 513418 260186 513654
rect 260422 513418 296186 513654
rect 296422 513418 332186 513654
rect 332422 513418 368186 513654
rect 368422 513418 404186 513654
rect 404422 513418 440186 513654
rect 440422 513418 476186 513654
rect 476422 513418 512186 513654
rect 512422 513418 548186 513654
rect 548422 513418 589182 513654
rect 589418 513418 590520 513654
rect -6596 513334 590520 513418
rect -6596 513098 -5494 513334
rect -5258 513098 8186 513334
rect 8422 513098 44186 513334
rect 44422 513098 80186 513334
rect 80422 513098 116186 513334
rect 116422 513098 152186 513334
rect 152422 513098 188186 513334
rect 188422 513098 224186 513334
rect 224422 513098 260186 513334
rect 260422 513098 296186 513334
rect 296422 513098 332186 513334
rect 332422 513098 368186 513334
rect 368422 513098 404186 513334
rect 404422 513098 440186 513334
rect 440422 513098 476186 513334
rect 476422 513098 512186 513334
rect 512422 513098 548186 513334
rect 548422 513098 589182 513334
rect 589418 513098 590520 513334
rect -6596 513076 590520 513098
rect -5676 513074 -5076 513076
rect 8004 513074 8604 513076
rect 44004 513074 44604 513076
rect 80004 513074 80604 513076
rect 116004 513074 116604 513076
rect 152004 513074 152604 513076
rect 188004 513074 188604 513076
rect 224004 513074 224604 513076
rect 260004 513074 260604 513076
rect 296004 513074 296604 513076
rect 332004 513074 332604 513076
rect 368004 513074 368604 513076
rect 404004 513074 404604 513076
rect 440004 513074 440604 513076
rect 476004 513074 476604 513076
rect 512004 513074 512604 513076
rect 548004 513074 548604 513076
rect 589000 513074 589600 513076
rect -3836 510076 -3236 510078
rect 4404 510076 5004 510078
rect 40404 510076 41004 510078
rect 76404 510076 77004 510078
rect 112404 510076 113004 510078
rect 148404 510076 149004 510078
rect 184404 510076 185004 510078
rect 220404 510076 221004 510078
rect 256404 510076 257004 510078
rect 292404 510076 293004 510078
rect 328404 510076 329004 510078
rect 364404 510076 365004 510078
rect 400404 510076 401004 510078
rect 436404 510076 437004 510078
rect 472404 510076 473004 510078
rect 508404 510076 509004 510078
rect 544404 510076 545004 510078
rect 580404 510076 581004 510078
rect 587160 510076 587760 510078
rect -4756 510054 588680 510076
rect -4756 509818 -3654 510054
rect -3418 509818 4586 510054
rect 4822 509818 40586 510054
rect 40822 509818 76586 510054
rect 76822 509818 112586 510054
rect 112822 509818 148586 510054
rect 148822 509818 184586 510054
rect 184822 509818 220586 510054
rect 220822 509818 256586 510054
rect 256822 509818 292586 510054
rect 292822 509818 328586 510054
rect 328822 509818 364586 510054
rect 364822 509818 400586 510054
rect 400822 509818 436586 510054
rect 436822 509818 472586 510054
rect 472822 509818 508586 510054
rect 508822 509818 544586 510054
rect 544822 509818 580586 510054
rect 580822 509818 587342 510054
rect 587578 509818 588680 510054
rect -4756 509734 588680 509818
rect -4756 509498 -3654 509734
rect -3418 509498 4586 509734
rect 4822 509498 40586 509734
rect 40822 509498 76586 509734
rect 76822 509498 112586 509734
rect 112822 509498 148586 509734
rect 148822 509498 184586 509734
rect 184822 509498 220586 509734
rect 220822 509498 256586 509734
rect 256822 509498 292586 509734
rect 292822 509498 328586 509734
rect 328822 509498 364586 509734
rect 364822 509498 400586 509734
rect 400822 509498 436586 509734
rect 436822 509498 472586 509734
rect 472822 509498 508586 509734
rect 508822 509498 544586 509734
rect 544822 509498 580586 509734
rect 580822 509498 587342 509734
rect 587578 509498 588680 509734
rect -4756 509476 588680 509498
rect -3836 509474 -3236 509476
rect 4404 509474 5004 509476
rect 40404 509474 41004 509476
rect 76404 509474 77004 509476
rect 112404 509474 113004 509476
rect 148404 509474 149004 509476
rect 184404 509474 185004 509476
rect 220404 509474 221004 509476
rect 256404 509474 257004 509476
rect 292404 509474 293004 509476
rect 328404 509474 329004 509476
rect 364404 509474 365004 509476
rect 400404 509474 401004 509476
rect 436404 509474 437004 509476
rect 472404 509474 473004 509476
rect 508404 509474 509004 509476
rect 544404 509474 545004 509476
rect 580404 509474 581004 509476
rect 587160 509474 587760 509476
rect -1996 506476 -1396 506478
rect 804 506476 1404 506478
rect 36804 506476 37404 506478
rect 72804 506476 73404 506478
rect 108804 506476 109404 506478
rect 144804 506476 145404 506478
rect 180804 506476 181404 506478
rect 216804 506476 217404 506478
rect 252804 506476 253404 506478
rect 288804 506476 289404 506478
rect 324804 506476 325404 506478
rect 360804 506476 361404 506478
rect 396804 506476 397404 506478
rect 432804 506476 433404 506478
rect 468804 506476 469404 506478
rect 504804 506476 505404 506478
rect 540804 506476 541404 506478
rect 576804 506476 577404 506478
rect 585320 506476 585920 506478
rect -2916 506454 586840 506476
rect -2916 506218 -1814 506454
rect -1578 506218 986 506454
rect 1222 506218 36986 506454
rect 37222 506218 72986 506454
rect 73222 506218 108986 506454
rect 109222 506218 144986 506454
rect 145222 506218 180986 506454
rect 181222 506218 216986 506454
rect 217222 506218 252986 506454
rect 253222 506218 288986 506454
rect 289222 506218 324986 506454
rect 325222 506218 360986 506454
rect 361222 506218 396986 506454
rect 397222 506218 432986 506454
rect 433222 506218 468986 506454
rect 469222 506218 504986 506454
rect 505222 506218 540986 506454
rect 541222 506218 576986 506454
rect 577222 506218 585502 506454
rect 585738 506218 586840 506454
rect -2916 506134 586840 506218
rect -2916 505898 -1814 506134
rect -1578 505898 986 506134
rect 1222 505898 36986 506134
rect 37222 505898 72986 506134
rect 73222 505898 108986 506134
rect 109222 505898 144986 506134
rect 145222 505898 180986 506134
rect 181222 505898 216986 506134
rect 217222 505898 252986 506134
rect 253222 505898 288986 506134
rect 289222 505898 324986 506134
rect 325222 505898 360986 506134
rect 361222 505898 396986 506134
rect 397222 505898 432986 506134
rect 433222 505898 468986 506134
rect 469222 505898 504986 506134
rect 505222 505898 540986 506134
rect 541222 505898 576986 506134
rect 577222 505898 585502 506134
rect 585738 505898 586840 506134
rect -2916 505876 586840 505898
rect -1996 505874 -1396 505876
rect 804 505874 1404 505876
rect 36804 505874 37404 505876
rect 72804 505874 73404 505876
rect 108804 505874 109404 505876
rect 144804 505874 145404 505876
rect 180804 505874 181404 505876
rect 216804 505874 217404 505876
rect 252804 505874 253404 505876
rect 288804 505874 289404 505876
rect 324804 505874 325404 505876
rect 360804 505874 361404 505876
rect 396804 505874 397404 505876
rect 432804 505874 433404 505876
rect 468804 505874 469404 505876
rect 504804 505874 505404 505876
rect 540804 505874 541404 505876
rect 576804 505874 577404 505876
rect 585320 505874 585920 505876
rect -8436 499276 -7836 499278
rect 29604 499276 30204 499278
rect 65604 499276 66204 499278
rect 101604 499276 102204 499278
rect 137604 499276 138204 499278
rect 173604 499276 174204 499278
rect 209604 499276 210204 499278
rect 245604 499276 246204 499278
rect 281604 499276 282204 499278
rect 317604 499276 318204 499278
rect 353604 499276 354204 499278
rect 389604 499276 390204 499278
rect 425604 499276 426204 499278
rect 461604 499276 462204 499278
rect 497604 499276 498204 499278
rect 533604 499276 534204 499278
rect 569604 499276 570204 499278
rect 591760 499276 592360 499278
rect -8436 499254 592360 499276
rect -8436 499018 -8254 499254
rect -8018 499018 29786 499254
rect 30022 499018 65786 499254
rect 66022 499018 101786 499254
rect 102022 499018 137786 499254
rect 138022 499018 173786 499254
rect 174022 499018 209786 499254
rect 210022 499018 245786 499254
rect 246022 499018 281786 499254
rect 282022 499018 317786 499254
rect 318022 499018 353786 499254
rect 354022 499018 389786 499254
rect 390022 499018 425786 499254
rect 426022 499018 461786 499254
rect 462022 499018 497786 499254
rect 498022 499018 533786 499254
rect 534022 499018 569786 499254
rect 570022 499018 591942 499254
rect 592178 499018 592360 499254
rect -8436 498934 592360 499018
rect -8436 498698 -8254 498934
rect -8018 498698 29786 498934
rect 30022 498698 65786 498934
rect 66022 498698 101786 498934
rect 102022 498698 137786 498934
rect 138022 498698 173786 498934
rect 174022 498698 209786 498934
rect 210022 498698 245786 498934
rect 246022 498698 281786 498934
rect 282022 498698 317786 498934
rect 318022 498698 353786 498934
rect 354022 498698 389786 498934
rect 390022 498698 425786 498934
rect 426022 498698 461786 498934
rect 462022 498698 497786 498934
rect 498022 498698 533786 498934
rect 534022 498698 569786 498934
rect 570022 498698 591942 498934
rect 592178 498698 592360 498934
rect -8436 498676 592360 498698
rect -8436 498674 -7836 498676
rect 29604 498674 30204 498676
rect 65604 498674 66204 498676
rect 101604 498674 102204 498676
rect 137604 498674 138204 498676
rect 173604 498674 174204 498676
rect 209604 498674 210204 498676
rect 245604 498674 246204 498676
rect 281604 498674 282204 498676
rect 317604 498674 318204 498676
rect 353604 498674 354204 498676
rect 389604 498674 390204 498676
rect 425604 498674 426204 498676
rect 461604 498674 462204 498676
rect 497604 498674 498204 498676
rect 533604 498674 534204 498676
rect 569604 498674 570204 498676
rect 591760 498674 592360 498676
rect -6596 495676 -5996 495678
rect 26004 495676 26604 495678
rect 62004 495676 62604 495678
rect 98004 495676 98604 495678
rect 134004 495676 134604 495678
rect 170004 495676 170604 495678
rect 206004 495676 206604 495678
rect 242004 495676 242604 495678
rect 278004 495676 278604 495678
rect 314004 495676 314604 495678
rect 350004 495676 350604 495678
rect 386004 495676 386604 495678
rect 422004 495676 422604 495678
rect 458004 495676 458604 495678
rect 494004 495676 494604 495678
rect 530004 495676 530604 495678
rect 566004 495676 566604 495678
rect 589920 495676 590520 495678
rect -6596 495654 590520 495676
rect -6596 495418 -6414 495654
rect -6178 495418 26186 495654
rect 26422 495418 62186 495654
rect 62422 495418 98186 495654
rect 98422 495418 134186 495654
rect 134422 495418 170186 495654
rect 170422 495418 206186 495654
rect 206422 495418 242186 495654
rect 242422 495418 278186 495654
rect 278422 495418 314186 495654
rect 314422 495418 350186 495654
rect 350422 495418 386186 495654
rect 386422 495418 422186 495654
rect 422422 495418 458186 495654
rect 458422 495418 494186 495654
rect 494422 495418 530186 495654
rect 530422 495418 566186 495654
rect 566422 495418 590102 495654
rect 590338 495418 590520 495654
rect -6596 495334 590520 495418
rect -6596 495098 -6414 495334
rect -6178 495098 26186 495334
rect 26422 495098 62186 495334
rect 62422 495098 98186 495334
rect 98422 495098 134186 495334
rect 134422 495098 170186 495334
rect 170422 495098 206186 495334
rect 206422 495098 242186 495334
rect 242422 495098 278186 495334
rect 278422 495098 314186 495334
rect 314422 495098 350186 495334
rect 350422 495098 386186 495334
rect 386422 495098 422186 495334
rect 422422 495098 458186 495334
rect 458422 495098 494186 495334
rect 494422 495098 530186 495334
rect 530422 495098 566186 495334
rect 566422 495098 590102 495334
rect 590338 495098 590520 495334
rect -6596 495076 590520 495098
rect -6596 495074 -5996 495076
rect 26004 495074 26604 495076
rect 62004 495074 62604 495076
rect 98004 495074 98604 495076
rect 134004 495074 134604 495076
rect 170004 495074 170604 495076
rect 206004 495074 206604 495076
rect 242004 495074 242604 495076
rect 278004 495074 278604 495076
rect 314004 495074 314604 495076
rect 350004 495074 350604 495076
rect 386004 495074 386604 495076
rect 422004 495074 422604 495076
rect 458004 495074 458604 495076
rect 494004 495074 494604 495076
rect 530004 495074 530604 495076
rect 566004 495074 566604 495076
rect 589920 495074 590520 495076
rect -4756 492076 -4156 492078
rect 22404 492076 23004 492078
rect 58404 492076 59004 492078
rect 94404 492076 95004 492078
rect 130404 492076 131004 492078
rect 166404 492076 167004 492078
rect 202404 492076 203004 492078
rect 238404 492076 239004 492078
rect 274404 492076 275004 492078
rect 310404 492076 311004 492078
rect 346404 492076 347004 492078
rect 382404 492076 383004 492078
rect 418404 492076 419004 492078
rect 454404 492076 455004 492078
rect 490404 492076 491004 492078
rect 526404 492076 527004 492078
rect 562404 492076 563004 492078
rect 588080 492076 588680 492078
rect -4756 492054 588680 492076
rect -4756 491818 -4574 492054
rect -4338 491818 22586 492054
rect 22822 491818 58586 492054
rect 58822 491818 94586 492054
rect 94822 491818 130586 492054
rect 130822 491818 166586 492054
rect 166822 491818 202586 492054
rect 202822 491818 238586 492054
rect 238822 491818 274586 492054
rect 274822 491818 310586 492054
rect 310822 491818 346586 492054
rect 346822 491818 382586 492054
rect 382822 491818 418586 492054
rect 418822 491818 454586 492054
rect 454822 491818 490586 492054
rect 490822 491818 526586 492054
rect 526822 491818 562586 492054
rect 562822 491818 588262 492054
rect 588498 491818 588680 492054
rect -4756 491734 588680 491818
rect -4756 491498 -4574 491734
rect -4338 491498 22586 491734
rect 22822 491498 58586 491734
rect 58822 491498 94586 491734
rect 94822 491498 130586 491734
rect 130822 491498 166586 491734
rect 166822 491498 202586 491734
rect 202822 491498 238586 491734
rect 238822 491498 274586 491734
rect 274822 491498 310586 491734
rect 310822 491498 346586 491734
rect 346822 491498 382586 491734
rect 382822 491498 418586 491734
rect 418822 491498 454586 491734
rect 454822 491498 490586 491734
rect 490822 491498 526586 491734
rect 526822 491498 562586 491734
rect 562822 491498 588262 491734
rect 588498 491498 588680 491734
rect -4756 491476 588680 491498
rect -4756 491474 -4156 491476
rect 22404 491474 23004 491476
rect 58404 491474 59004 491476
rect 94404 491474 95004 491476
rect 130404 491474 131004 491476
rect 166404 491474 167004 491476
rect 202404 491474 203004 491476
rect 238404 491474 239004 491476
rect 274404 491474 275004 491476
rect 310404 491474 311004 491476
rect 346404 491474 347004 491476
rect 382404 491474 383004 491476
rect 418404 491474 419004 491476
rect 454404 491474 455004 491476
rect 490404 491474 491004 491476
rect 526404 491474 527004 491476
rect 562404 491474 563004 491476
rect 588080 491474 588680 491476
rect -2916 488476 -2316 488478
rect 18804 488476 19404 488478
rect 54804 488476 55404 488478
rect 90804 488476 91404 488478
rect 126804 488476 127404 488478
rect 162804 488476 163404 488478
rect 198804 488476 199404 488478
rect 234804 488476 235404 488478
rect 270804 488476 271404 488478
rect 306804 488476 307404 488478
rect 342804 488476 343404 488478
rect 378804 488476 379404 488478
rect 414804 488476 415404 488478
rect 450804 488476 451404 488478
rect 486804 488476 487404 488478
rect 522804 488476 523404 488478
rect 558804 488476 559404 488478
rect 586240 488476 586840 488478
rect -2916 488454 586840 488476
rect -2916 488218 -2734 488454
rect -2498 488218 18986 488454
rect 19222 488218 54986 488454
rect 55222 488218 90986 488454
rect 91222 488218 126986 488454
rect 127222 488218 162986 488454
rect 163222 488218 198986 488454
rect 199222 488218 234986 488454
rect 235222 488218 270986 488454
rect 271222 488218 306986 488454
rect 307222 488218 342986 488454
rect 343222 488218 378986 488454
rect 379222 488218 414986 488454
rect 415222 488218 450986 488454
rect 451222 488218 486986 488454
rect 487222 488218 522986 488454
rect 523222 488218 558986 488454
rect 559222 488218 586422 488454
rect 586658 488218 586840 488454
rect -2916 488134 586840 488218
rect -2916 487898 -2734 488134
rect -2498 487898 18986 488134
rect 19222 487898 54986 488134
rect 55222 487898 90986 488134
rect 91222 487898 126986 488134
rect 127222 487898 162986 488134
rect 163222 487898 198986 488134
rect 199222 487898 234986 488134
rect 235222 487898 270986 488134
rect 271222 487898 306986 488134
rect 307222 487898 342986 488134
rect 343222 487898 378986 488134
rect 379222 487898 414986 488134
rect 415222 487898 450986 488134
rect 451222 487898 486986 488134
rect 487222 487898 522986 488134
rect 523222 487898 558986 488134
rect 559222 487898 586422 488134
rect 586658 487898 586840 488134
rect -2916 487876 586840 487898
rect -2916 487874 -2316 487876
rect 18804 487874 19404 487876
rect 54804 487874 55404 487876
rect 90804 487874 91404 487876
rect 126804 487874 127404 487876
rect 162804 487874 163404 487876
rect 198804 487874 199404 487876
rect 234804 487874 235404 487876
rect 270804 487874 271404 487876
rect 306804 487874 307404 487876
rect 342804 487874 343404 487876
rect 378804 487874 379404 487876
rect 414804 487874 415404 487876
rect 450804 487874 451404 487876
rect 486804 487874 487404 487876
rect 522804 487874 523404 487876
rect 558804 487874 559404 487876
rect 586240 487874 586840 487876
rect -7516 481276 -6916 481278
rect 11604 481276 12204 481278
rect 47604 481276 48204 481278
rect 83604 481276 84204 481278
rect 119604 481276 120204 481278
rect 155604 481276 156204 481278
rect 191604 481276 192204 481278
rect 227604 481276 228204 481278
rect 263604 481276 264204 481278
rect 299604 481276 300204 481278
rect 335604 481276 336204 481278
rect 371604 481276 372204 481278
rect 407604 481276 408204 481278
rect 443604 481276 444204 481278
rect 479604 481276 480204 481278
rect 515604 481276 516204 481278
rect 551604 481276 552204 481278
rect 590840 481276 591440 481278
rect -8436 481254 592360 481276
rect -8436 481018 -7334 481254
rect -7098 481018 11786 481254
rect 12022 481018 47786 481254
rect 48022 481018 83786 481254
rect 84022 481018 119786 481254
rect 120022 481018 155786 481254
rect 156022 481018 191786 481254
rect 192022 481018 227786 481254
rect 228022 481018 263786 481254
rect 264022 481018 299786 481254
rect 300022 481018 335786 481254
rect 336022 481018 371786 481254
rect 372022 481018 407786 481254
rect 408022 481018 443786 481254
rect 444022 481018 479786 481254
rect 480022 481018 515786 481254
rect 516022 481018 551786 481254
rect 552022 481018 591022 481254
rect 591258 481018 592360 481254
rect -8436 480934 592360 481018
rect -8436 480698 -7334 480934
rect -7098 480698 11786 480934
rect 12022 480698 47786 480934
rect 48022 480698 83786 480934
rect 84022 480698 119786 480934
rect 120022 480698 155786 480934
rect 156022 480698 191786 480934
rect 192022 480698 227786 480934
rect 228022 480698 263786 480934
rect 264022 480698 299786 480934
rect 300022 480698 335786 480934
rect 336022 480698 371786 480934
rect 372022 480698 407786 480934
rect 408022 480698 443786 480934
rect 444022 480698 479786 480934
rect 480022 480698 515786 480934
rect 516022 480698 551786 480934
rect 552022 480698 591022 480934
rect 591258 480698 592360 480934
rect -8436 480676 592360 480698
rect -7516 480674 -6916 480676
rect 11604 480674 12204 480676
rect 47604 480674 48204 480676
rect 83604 480674 84204 480676
rect 119604 480674 120204 480676
rect 155604 480674 156204 480676
rect 191604 480674 192204 480676
rect 227604 480674 228204 480676
rect 263604 480674 264204 480676
rect 299604 480674 300204 480676
rect 335604 480674 336204 480676
rect 371604 480674 372204 480676
rect 407604 480674 408204 480676
rect 443604 480674 444204 480676
rect 479604 480674 480204 480676
rect 515604 480674 516204 480676
rect 551604 480674 552204 480676
rect 590840 480674 591440 480676
rect -5676 477676 -5076 477678
rect 8004 477676 8604 477678
rect 44004 477676 44604 477678
rect 80004 477676 80604 477678
rect 116004 477676 116604 477678
rect 152004 477676 152604 477678
rect 188004 477676 188604 477678
rect 224004 477676 224604 477678
rect 260004 477676 260604 477678
rect 296004 477676 296604 477678
rect 332004 477676 332604 477678
rect 368004 477676 368604 477678
rect 404004 477676 404604 477678
rect 440004 477676 440604 477678
rect 476004 477676 476604 477678
rect 512004 477676 512604 477678
rect 548004 477676 548604 477678
rect 589000 477676 589600 477678
rect -6596 477654 590520 477676
rect -6596 477418 -5494 477654
rect -5258 477418 8186 477654
rect 8422 477418 44186 477654
rect 44422 477418 80186 477654
rect 80422 477418 116186 477654
rect 116422 477418 152186 477654
rect 152422 477418 188186 477654
rect 188422 477418 224186 477654
rect 224422 477418 260186 477654
rect 260422 477418 296186 477654
rect 296422 477418 332186 477654
rect 332422 477418 368186 477654
rect 368422 477418 404186 477654
rect 404422 477418 440186 477654
rect 440422 477418 476186 477654
rect 476422 477418 512186 477654
rect 512422 477418 548186 477654
rect 548422 477418 589182 477654
rect 589418 477418 590520 477654
rect -6596 477334 590520 477418
rect -6596 477098 -5494 477334
rect -5258 477098 8186 477334
rect 8422 477098 44186 477334
rect 44422 477098 80186 477334
rect 80422 477098 116186 477334
rect 116422 477098 152186 477334
rect 152422 477098 188186 477334
rect 188422 477098 224186 477334
rect 224422 477098 260186 477334
rect 260422 477098 296186 477334
rect 296422 477098 332186 477334
rect 332422 477098 368186 477334
rect 368422 477098 404186 477334
rect 404422 477098 440186 477334
rect 440422 477098 476186 477334
rect 476422 477098 512186 477334
rect 512422 477098 548186 477334
rect 548422 477098 589182 477334
rect 589418 477098 590520 477334
rect -6596 477076 590520 477098
rect -5676 477074 -5076 477076
rect 8004 477074 8604 477076
rect 44004 477074 44604 477076
rect 80004 477074 80604 477076
rect 116004 477074 116604 477076
rect 152004 477074 152604 477076
rect 188004 477074 188604 477076
rect 224004 477074 224604 477076
rect 260004 477074 260604 477076
rect 296004 477074 296604 477076
rect 332004 477074 332604 477076
rect 368004 477074 368604 477076
rect 404004 477074 404604 477076
rect 440004 477074 440604 477076
rect 476004 477074 476604 477076
rect 512004 477074 512604 477076
rect 548004 477074 548604 477076
rect 589000 477074 589600 477076
rect -3836 474076 -3236 474078
rect 4404 474076 5004 474078
rect 40404 474076 41004 474078
rect 76404 474076 77004 474078
rect 112404 474076 113004 474078
rect 148404 474076 149004 474078
rect 184404 474076 185004 474078
rect 220404 474076 221004 474078
rect 256404 474076 257004 474078
rect 292404 474076 293004 474078
rect 328404 474076 329004 474078
rect 364404 474076 365004 474078
rect 400404 474076 401004 474078
rect 436404 474076 437004 474078
rect 472404 474076 473004 474078
rect 508404 474076 509004 474078
rect 544404 474076 545004 474078
rect 580404 474076 581004 474078
rect 587160 474076 587760 474078
rect -4756 474054 588680 474076
rect -4756 473818 -3654 474054
rect -3418 473818 4586 474054
rect 4822 473818 40586 474054
rect 40822 473818 76586 474054
rect 76822 473818 112586 474054
rect 112822 473818 148586 474054
rect 148822 473818 184586 474054
rect 184822 473818 220586 474054
rect 220822 473818 256586 474054
rect 256822 473818 292586 474054
rect 292822 473818 328586 474054
rect 328822 473818 364586 474054
rect 364822 473818 400586 474054
rect 400822 473818 436586 474054
rect 436822 473818 472586 474054
rect 472822 473818 508586 474054
rect 508822 473818 544586 474054
rect 544822 473818 580586 474054
rect 580822 473818 587342 474054
rect 587578 473818 588680 474054
rect -4756 473734 588680 473818
rect -4756 473498 -3654 473734
rect -3418 473498 4586 473734
rect 4822 473498 40586 473734
rect 40822 473498 76586 473734
rect 76822 473498 112586 473734
rect 112822 473498 148586 473734
rect 148822 473498 184586 473734
rect 184822 473498 220586 473734
rect 220822 473498 256586 473734
rect 256822 473498 292586 473734
rect 292822 473498 328586 473734
rect 328822 473498 364586 473734
rect 364822 473498 400586 473734
rect 400822 473498 436586 473734
rect 436822 473498 472586 473734
rect 472822 473498 508586 473734
rect 508822 473498 544586 473734
rect 544822 473498 580586 473734
rect 580822 473498 587342 473734
rect 587578 473498 588680 473734
rect -4756 473476 588680 473498
rect -3836 473474 -3236 473476
rect 4404 473474 5004 473476
rect 40404 473474 41004 473476
rect 76404 473474 77004 473476
rect 112404 473474 113004 473476
rect 148404 473474 149004 473476
rect 184404 473474 185004 473476
rect 220404 473474 221004 473476
rect 256404 473474 257004 473476
rect 292404 473474 293004 473476
rect 328404 473474 329004 473476
rect 364404 473474 365004 473476
rect 400404 473474 401004 473476
rect 436404 473474 437004 473476
rect 472404 473474 473004 473476
rect 508404 473474 509004 473476
rect 544404 473474 545004 473476
rect 580404 473474 581004 473476
rect 587160 473474 587760 473476
rect -1996 470476 -1396 470478
rect 804 470476 1404 470478
rect 36804 470476 37404 470478
rect 72804 470476 73404 470478
rect 108804 470476 109404 470478
rect 144804 470476 145404 470478
rect 180804 470476 181404 470478
rect 216804 470476 217404 470478
rect 252804 470476 253404 470478
rect 288804 470476 289404 470478
rect 324804 470476 325404 470478
rect 360804 470476 361404 470478
rect 396804 470476 397404 470478
rect 432804 470476 433404 470478
rect 468804 470476 469404 470478
rect 504804 470476 505404 470478
rect 540804 470476 541404 470478
rect 576804 470476 577404 470478
rect 585320 470476 585920 470478
rect -2916 470454 586840 470476
rect -2916 470218 -1814 470454
rect -1578 470218 986 470454
rect 1222 470218 36986 470454
rect 37222 470218 72986 470454
rect 73222 470218 108986 470454
rect 109222 470218 144986 470454
rect 145222 470218 180986 470454
rect 181222 470218 216986 470454
rect 217222 470218 252986 470454
rect 253222 470218 288986 470454
rect 289222 470218 324986 470454
rect 325222 470218 360986 470454
rect 361222 470218 396986 470454
rect 397222 470218 432986 470454
rect 433222 470218 468986 470454
rect 469222 470218 504986 470454
rect 505222 470218 540986 470454
rect 541222 470218 576986 470454
rect 577222 470218 585502 470454
rect 585738 470218 586840 470454
rect -2916 470134 586840 470218
rect -2916 469898 -1814 470134
rect -1578 469898 986 470134
rect 1222 469898 36986 470134
rect 37222 469898 72986 470134
rect 73222 469898 108986 470134
rect 109222 469898 144986 470134
rect 145222 469898 180986 470134
rect 181222 469898 216986 470134
rect 217222 469898 252986 470134
rect 253222 469898 288986 470134
rect 289222 469898 324986 470134
rect 325222 469898 360986 470134
rect 361222 469898 396986 470134
rect 397222 469898 432986 470134
rect 433222 469898 468986 470134
rect 469222 469898 504986 470134
rect 505222 469898 540986 470134
rect 541222 469898 576986 470134
rect 577222 469898 585502 470134
rect 585738 469898 586840 470134
rect -2916 469876 586840 469898
rect -1996 469874 -1396 469876
rect 804 469874 1404 469876
rect 36804 469874 37404 469876
rect 72804 469874 73404 469876
rect 108804 469874 109404 469876
rect 144804 469874 145404 469876
rect 180804 469874 181404 469876
rect 216804 469874 217404 469876
rect 252804 469874 253404 469876
rect 288804 469874 289404 469876
rect 324804 469874 325404 469876
rect 360804 469874 361404 469876
rect 396804 469874 397404 469876
rect 432804 469874 433404 469876
rect 468804 469874 469404 469876
rect 504804 469874 505404 469876
rect 540804 469874 541404 469876
rect 576804 469874 577404 469876
rect 585320 469874 585920 469876
rect -8436 463276 -7836 463278
rect 29604 463276 30204 463278
rect 65604 463276 66204 463278
rect 101604 463276 102204 463278
rect 137604 463276 138204 463278
rect 173604 463276 174204 463278
rect 209604 463276 210204 463278
rect 245604 463276 246204 463278
rect 281604 463276 282204 463278
rect 317604 463276 318204 463278
rect 353604 463276 354204 463278
rect 389604 463276 390204 463278
rect 425604 463276 426204 463278
rect 461604 463276 462204 463278
rect 497604 463276 498204 463278
rect 533604 463276 534204 463278
rect 569604 463276 570204 463278
rect 591760 463276 592360 463278
rect -8436 463254 592360 463276
rect -8436 463018 -8254 463254
rect -8018 463018 29786 463254
rect 30022 463018 65786 463254
rect 66022 463018 101786 463254
rect 102022 463018 137786 463254
rect 138022 463018 173786 463254
rect 174022 463018 209786 463254
rect 210022 463018 245786 463254
rect 246022 463018 281786 463254
rect 282022 463018 317786 463254
rect 318022 463018 353786 463254
rect 354022 463018 389786 463254
rect 390022 463018 425786 463254
rect 426022 463018 461786 463254
rect 462022 463018 497786 463254
rect 498022 463018 533786 463254
rect 534022 463018 569786 463254
rect 570022 463018 591942 463254
rect 592178 463018 592360 463254
rect -8436 462934 592360 463018
rect -8436 462698 -8254 462934
rect -8018 462698 29786 462934
rect 30022 462698 65786 462934
rect 66022 462698 101786 462934
rect 102022 462698 137786 462934
rect 138022 462698 173786 462934
rect 174022 462698 209786 462934
rect 210022 462698 245786 462934
rect 246022 462698 281786 462934
rect 282022 462698 317786 462934
rect 318022 462698 353786 462934
rect 354022 462698 389786 462934
rect 390022 462698 425786 462934
rect 426022 462698 461786 462934
rect 462022 462698 497786 462934
rect 498022 462698 533786 462934
rect 534022 462698 569786 462934
rect 570022 462698 591942 462934
rect 592178 462698 592360 462934
rect -8436 462676 592360 462698
rect -8436 462674 -7836 462676
rect 29604 462674 30204 462676
rect 65604 462674 66204 462676
rect 101604 462674 102204 462676
rect 137604 462674 138204 462676
rect 173604 462674 174204 462676
rect 209604 462674 210204 462676
rect 245604 462674 246204 462676
rect 281604 462674 282204 462676
rect 317604 462674 318204 462676
rect 353604 462674 354204 462676
rect 389604 462674 390204 462676
rect 425604 462674 426204 462676
rect 461604 462674 462204 462676
rect 497604 462674 498204 462676
rect 533604 462674 534204 462676
rect 569604 462674 570204 462676
rect 591760 462674 592360 462676
rect -6596 459676 -5996 459678
rect 26004 459676 26604 459678
rect 62004 459676 62604 459678
rect 98004 459676 98604 459678
rect 134004 459676 134604 459678
rect 170004 459676 170604 459678
rect 206004 459676 206604 459678
rect 242004 459676 242604 459678
rect 278004 459676 278604 459678
rect 314004 459676 314604 459678
rect 350004 459676 350604 459678
rect 386004 459676 386604 459678
rect 422004 459676 422604 459678
rect 458004 459676 458604 459678
rect 494004 459676 494604 459678
rect 530004 459676 530604 459678
rect 566004 459676 566604 459678
rect 589920 459676 590520 459678
rect -6596 459654 590520 459676
rect -6596 459418 -6414 459654
rect -6178 459418 26186 459654
rect 26422 459418 62186 459654
rect 62422 459418 98186 459654
rect 98422 459418 134186 459654
rect 134422 459418 170186 459654
rect 170422 459418 206186 459654
rect 206422 459418 242186 459654
rect 242422 459418 278186 459654
rect 278422 459418 314186 459654
rect 314422 459418 350186 459654
rect 350422 459418 386186 459654
rect 386422 459418 422186 459654
rect 422422 459418 458186 459654
rect 458422 459418 494186 459654
rect 494422 459418 530186 459654
rect 530422 459418 566186 459654
rect 566422 459418 590102 459654
rect 590338 459418 590520 459654
rect -6596 459334 590520 459418
rect -6596 459098 -6414 459334
rect -6178 459098 26186 459334
rect 26422 459098 62186 459334
rect 62422 459098 98186 459334
rect 98422 459098 134186 459334
rect 134422 459098 170186 459334
rect 170422 459098 206186 459334
rect 206422 459098 242186 459334
rect 242422 459098 278186 459334
rect 278422 459098 314186 459334
rect 314422 459098 350186 459334
rect 350422 459098 386186 459334
rect 386422 459098 422186 459334
rect 422422 459098 458186 459334
rect 458422 459098 494186 459334
rect 494422 459098 530186 459334
rect 530422 459098 566186 459334
rect 566422 459098 590102 459334
rect 590338 459098 590520 459334
rect -6596 459076 590520 459098
rect -6596 459074 -5996 459076
rect 26004 459074 26604 459076
rect 62004 459074 62604 459076
rect 98004 459074 98604 459076
rect 134004 459074 134604 459076
rect 170004 459074 170604 459076
rect 206004 459074 206604 459076
rect 242004 459074 242604 459076
rect 278004 459074 278604 459076
rect 314004 459074 314604 459076
rect 350004 459074 350604 459076
rect 386004 459074 386604 459076
rect 422004 459074 422604 459076
rect 458004 459074 458604 459076
rect 494004 459074 494604 459076
rect 530004 459074 530604 459076
rect 566004 459074 566604 459076
rect 589920 459074 590520 459076
rect -4756 456076 -4156 456078
rect 22404 456076 23004 456078
rect 58404 456076 59004 456078
rect 94404 456076 95004 456078
rect 130404 456076 131004 456078
rect 166404 456076 167004 456078
rect 202404 456076 203004 456078
rect 238404 456076 239004 456078
rect 274404 456076 275004 456078
rect 310404 456076 311004 456078
rect 346404 456076 347004 456078
rect 382404 456076 383004 456078
rect 418404 456076 419004 456078
rect 454404 456076 455004 456078
rect 490404 456076 491004 456078
rect 526404 456076 527004 456078
rect 562404 456076 563004 456078
rect 588080 456076 588680 456078
rect -4756 456054 588680 456076
rect -4756 455818 -4574 456054
rect -4338 455818 22586 456054
rect 22822 455818 58586 456054
rect 58822 455818 94586 456054
rect 94822 455818 130586 456054
rect 130822 455818 166586 456054
rect 166822 455818 202586 456054
rect 202822 455818 238586 456054
rect 238822 455818 274586 456054
rect 274822 455818 310586 456054
rect 310822 455818 346586 456054
rect 346822 455818 382586 456054
rect 382822 455818 418586 456054
rect 418822 455818 454586 456054
rect 454822 455818 490586 456054
rect 490822 455818 526586 456054
rect 526822 455818 562586 456054
rect 562822 455818 588262 456054
rect 588498 455818 588680 456054
rect -4756 455734 588680 455818
rect -4756 455498 -4574 455734
rect -4338 455498 22586 455734
rect 22822 455498 58586 455734
rect 58822 455498 94586 455734
rect 94822 455498 130586 455734
rect 130822 455498 166586 455734
rect 166822 455498 202586 455734
rect 202822 455498 238586 455734
rect 238822 455498 274586 455734
rect 274822 455498 310586 455734
rect 310822 455498 346586 455734
rect 346822 455498 382586 455734
rect 382822 455498 418586 455734
rect 418822 455498 454586 455734
rect 454822 455498 490586 455734
rect 490822 455498 526586 455734
rect 526822 455498 562586 455734
rect 562822 455498 588262 455734
rect 588498 455498 588680 455734
rect -4756 455476 588680 455498
rect -4756 455474 -4156 455476
rect 22404 455474 23004 455476
rect 58404 455474 59004 455476
rect 94404 455474 95004 455476
rect 130404 455474 131004 455476
rect 166404 455474 167004 455476
rect 202404 455474 203004 455476
rect 238404 455474 239004 455476
rect 274404 455474 275004 455476
rect 310404 455474 311004 455476
rect 346404 455474 347004 455476
rect 382404 455474 383004 455476
rect 418404 455474 419004 455476
rect 454404 455474 455004 455476
rect 490404 455474 491004 455476
rect 526404 455474 527004 455476
rect 562404 455474 563004 455476
rect 588080 455474 588680 455476
rect -2916 452476 -2316 452478
rect 18804 452476 19404 452478
rect 54804 452476 55404 452478
rect 90804 452476 91404 452478
rect 126804 452476 127404 452478
rect 162804 452476 163404 452478
rect 198804 452476 199404 452478
rect 234804 452476 235404 452478
rect 270804 452476 271404 452478
rect 306804 452476 307404 452478
rect 342804 452476 343404 452478
rect 378804 452476 379404 452478
rect 414804 452476 415404 452478
rect 450804 452476 451404 452478
rect 486804 452476 487404 452478
rect 522804 452476 523404 452478
rect 558804 452476 559404 452478
rect 586240 452476 586840 452478
rect -2916 452454 586840 452476
rect -2916 452218 -2734 452454
rect -2498 452218 18986 452454
rect 19222 452218 54986 452454
rect 55222 452218 90986 452454
rect 91222 452218 126986 452454
rect 127222 452218 162986 452454
rect 163222 452218 198986 452454
rect 199222 452218 234986 452454
rect 235222 452218 270986 452454
rect 271222 452218 306986 452454
rect 307222 452218 342986 452454
rect 343222 452218 378986 452454
rect 379222 452218 414986 452454
rect 415222 452218 450986 452454
rect 451222 452218 486986 452454
rect 487222 452218 522986 452454
rect 523222 452218 558986 452454
rect 559222 452218 586422 452454
rect 586658 452218 586840 452454
rect -2916 452134 586840 452218
rect -2916 451898 -2734 452134
rect -2498 451898 18986 452134
rect 19222 451898 54986 452134
rect 55222 451898 90986 452134
rect 91222 451898 126986 452134
rect 127222 451898 162986 452134
rect 163222 451898 198986 452134
rect 199222 451898 234986 452134
rect 235222 451898 270986 452134
rect 271222 451898 306986 452134
rect 307222 451898 342986 452134
rect 343222 451898 378986 452134
rect 379222 451898 414986 452134
rect 415222 451898 450986 452134
rect 451222 451898 486986 452134
rect 487222 451898 522986 452134
rect 523222 451898 558986 452134
rect 559222 451898 586422 452134
rect 586658 451898 586840 452134
rect -2916 451876 586840 451898
rect -2916 451874 -2316 451876
rect 18804 451874 19404 451876
rect 54804 451874 55404 451876
rect 90804 451874 91404 451876
rect 126804 451874 127404 451876
rect 162804 451874 163404 451876
rect 198804 451874 199404 451876
rect 234804 451874 235404 451876
rect 270804 451874 271404 451876
rect 306804 451874 307404 451876
rect 342804 451874 343404 451876
rect 378804 451874 379404 451876
rect 414804 451874 415404 451876
rect 450804 451874 451404 451876
rect 486804 451874 487404 451876
rect 522804 451874 523404 451876
rect 558804 451874 559404 451876
rect 586240 451874 586840 451876
rect -7516 445276 -6916 445278
rect 11604 445276 12204 445278
rect 47604 445276 48204 445278
rect 83604 445276 84204 445278
rect 119604 445276 120204 445278
rect 155604 445276 156204 445278
rect 191604 445276 192204 445278
rect 227604 445276 228204 445278
rect 263604 445276 264204 445278
rect 299604 445276 300204 445278
rect 335604 445276 336204 445278
rect 371604 445276 372204 445278
rect 407604 445276 408204 445278
rect 443604 445276 444204 445278
rect 479604 445276 480204 445278
rect 515604 445276 516204 445278
rect 551604 445276 552204 445278
rect 590840 445276 591440 445278
rect -8436 445254 592360 445276
rect -8436 445018 -7334 445254
rect -7098 445018 11786 445254
rect 12022 445018 47786 445254
rect 48022 445018 83786 445254
rect 84022 445018 119786 445254
rect 120022 445018 155786 445254
rect 156022 445018 191786 445254
rect 192022 445018 227786 445254
rect 228022 445018 263786 445254
rect 264022 445018 299786 445254
rect 300022 445018 335786 445254
rect 336022 445018 371786 445254
rect 372022 445018 407786 445254
rect 408022 445018 443786 445254
rect 444022 445018 479786 445254
rect 480022 445018 515786 445254
rect 516022 445018 551786 445254
rect 552022 445018 591022 445254
rect 591258 445018 592360 445254
rect -8436 444934 592360 445018
rect -8436 444698 -7334 444934
rect -7098 444698 11786 444934
rect 12022 444698 47786 444934
rect 48022 444698 83786 444934
rect 84022 444698 119786 444934
rect 120022 444698 155786 444934
rect 156022 444698 191786 444934
rect 192022 444698 227786 444934
rect 228022 444698 263786 444934
rect 264022 444698 299786 444934
rect 300022 444698 335786 444934
rect 336022 444698 371786 444934
rect 372022 444698 407786 444934
rect 408022 444698 443786 444934
rect 444022 444698 479786 444934
rect 480022 444698 515786 444934
rect 516022 444698 551786 444934
rect 552022 444698 591022 444934
rect 591258 444698 592360 444934
rect -8436 444676 592360 444698
rect -7516 444674 -6916 444676
rect 11604 444674 12204 444676
rect 47604 444674 48204 444676
rect 83604 444674 84204 444676
rect 119604 444674 120204 444676
rect 155604 444674 156204 444676
rect 191604 444674 192204 444676
rect 227604 444674 228204 444676
rect 263604 444674 264204 444676
rect 299604 444674 300204 444676
rect 335604 444674 336204 444676
rect 371604 444674 372204 444676
rect 407604 444674 408204 444676
rect 443604 444674 444204 444676
rect 479604 444674 480204 444676
rect 515604 444674 516204 444676
rect 551604 444674 552204 444676
rect 590840 444674 591440 444676
rect -5676 441676 -5076 441678
rect 8004 441676 8604 441678
rect 44004 441676 44604 441678
rect 80004 441676 80604 441678
rect 116004 441676 116604 441678
rect 152004 441676 152604 441678
rect 188004 441676 188604 441678
rect 224004 441676 224604 441678
rect 260004 441676 260604 441678
rect 296004 441676 296604 441678
rect 332004 441676 332604 441678
rect 368004 441676 368604 441678
rect 404004 441676 404604 441678
rect 440004 441676 440604 441678
rect 476004 441676 476604 441678
rect 512004 441676 512604 441678
rect 548004 441676 548604 441678
rect 589000 441676 589600 441678
rect -6596 441654 590520 441676
rect -6596 441418 -5494 441654
rect -5258 441418 8186 441654
rect 8422 441418 44186 441654
rect 44422 441418 80186 441654
rect 80422 441418 116186 441654
rect 116422 441418 152186 441654
rect 152422 441418 188186 441654
rect 188422 441418 224186 441654
rect 224422 441418 260186 441654
rect 260422 441418 296186 441654
rect 296422 441418 332186 441654
rect 332422 441418 368186 441654
rect 368422 441418 404186 441654
rect 404422 441418 440186 441654
rect 440422 441418 476186 441654
rect 476422 441418 512186 441654
rect 512422 441418 548186 441654
rect 548422 441418 589182 441654
rect 589418 441418 590520 441654
rect -6596 441334 590520 441418
rect -6596 441098 -5494 441334
rect -5258 441098 8186 441334
rect 8422 441098 44186 441334
rect 44422 441098 80186 441334
rect 80422 441098 116186 441334
rect 116422 441098 152186 441334
rect 152422 441098 188186 441334
rect 188422 441098 224186 441334
rect 224422 441098 260186 441334
rect 260422 441098 296186 441334
rect 296422 441098 332186 441334
rect 332422 441098 368186 441334
rect 368422 441098 404186 441334
rect 404422 441098 440186 441334
rect 440422 441098 476186 441334
rect 476422 441098 512186 441334
rect 512422 441098 548186 441334
rect 548422 441098 589182 441334
rect 589418 441098 590520 441334
rect -6596 441076 590520 441098
rect -5676 441074 -5076 441076
rect 8004 441074 8604 441076
rect 44004 441074 44604 441076
rect 80004 441074 80604 441076
rect 116004 441074 116604 441076
rect 152004 441074 152604 441076
rect 188004 441074 188604 441076
rect 224004 441074 224604 441076
rect 260004 441074 260604 441076
rect 296004 441074 296604 441076
rect 332004 441074 332604 441076
rect 368004 441074 368604 441076
rect 404004 441074 404604 441076
rect 440004 441074 440604 441076
rect 476004 441074 476604 441076
rect 512004 441074 512604 441076
rect 548004 441074 548604 441076
rect 589000 441074 589600 441076
rect -3836 438076 -3236 438078
rect 4404 438076 5004 438078
rect 40404 438076 41004 438078
rect 76404 438076 77004 438078
rect 112404 438076 113004 438078
rect 148404 438076 149004 438078
rect 184404 438076 185004 438078
rect 220404 438076 221004 438078
rect 256404 438076 257004 438078
rect 292404 438076 293004 438078
rect 328404 438076 329004 438078
rect 364404 438076 365004 438078
rect 400404 438076 401004 438078
rect 436404 438076 437004 438078
rect 472404 438076 473004 438078
rect 508404 438076 509004 438078
rect 544404 438076 545004 438078
rect 580404 438076 581004 438078
rect 587160 438076 587760 438078
rect -4756 438054 588680 438076
rect -4756 437818 -3654 438054
rect -3418 437818 4586 438054
rect 4822 437818 40586 438054
rect 40822 437818 76586 438054
rect 76822 437818 112586 438054
rect 112822 437818 148586 438054
rect 148822 437818 184586 438054
rect 184822 437818 220586 438054
rect 220822 437818 256586 438054
rect 256822 437818 292586 438054
rect 292822 437818 328586 438054
rect 328822 437818 364586 438054
rect 364822 437818 400586 438054
rect 400822 437818 436586 438054
rect 436822 437818 472586 438054
rect 472822 437818 508586 438054
rect 508822 437818 544586 438054
rect 544822 437818 580586 438054
rect 580822 437818 587342 438054
rect 587578 437818 588680 438054
rect -4756 437734 588680 437818
rect -4756 437498 -3654 437734
rect -3418 437498 4586 437734
rect 4822 437498 40586 437734
rect 40822 437498 76586 437734
rect 76822 437498 112586 437734
rect 112822 437498 148586 437734
rect 148822 437498 184586 437734
rect 184822 437498 220586 437734
rect 220822 437498 256586 437734
rect 256822 437498 292586 437734
rect 292822 437498 328586 437734
rect 328822 437498 364586 437734
rect 364822 437498 400586 437734
rect 400822 437498 436586 437734
rect 436822 437498 472586 437734
rect 472822 437498 508586 437734
rect 508822 437498 544586 437734
rect 544822 437498 580586 437734
rect 580822 437498 587342 437734
rect 587578 437498 588680 437734
rect -4756 437476 588680 437498
rect -3836 437474 -3236 437476
rect 4404 437474 5004 437476
rect 40404 437474 41004 437476
rect 76404 437474 77004 437476
rect 112404 437474 113004 437476
rect 148404 437474 149004 437476
rect 184404 437474 185004 437476
rect 220404 437474 221004 437476
rect 256404 437474 257004 437476
rect 292404 437474 293004 437476
rect 328404 437474 329004 437476
rect 364404 437474 365004 437476
rect 400404 437474 401004 437476
rect 436404 437474 437004 437476
rect 472404 437474 473004 437476
rect 508404 437474 509004 437476
rect 544404 437474 545004 437476
rect 580404 437474 581004 437476
rect 587160 437474 587760 437476
rect -1996 434476 -1396 434478
rect 804 434476 1404 434478
rect 36804 434476 37404 434478
rect 72804 434476 73404 434478
rect 108804 434476 109404 434478
rect 144804 434476 145404 434478
rect 180804 434476 181404 434478
rect 216804 434476 217404 434478
rect 252804 434476 253404 434478
rect 288804 434476 289404 434478
rect 324804 434476 325404 434478
rect 360804 434476 361404 434478
rect 396804 434476 397404 434478
rect 432804 434476 433404 434478
rect 468804 434476 469404 434478
rect 504804 434476 505404 434478
rect 540804 434476 541404 434478
rect 576804 434476 577404 434478
rect 585320 434476 585920 434478
rect -2916 434454 586840 434476
rect -2916 434218 -1814 434454
rect -1578 434218 986 434454
rect 1222 434218 36986 434454
rect 37222 434218 72986 434454
rect 73222 434218 108986 434454
rect 109222 434218 144986 434454
rect 145222 434218 180986 434454
rect 181222 434218 216986 434454
rect 217222 434218 252986 434454
rect 253222 434218 288986 434454
rect 289222 434218 324986 434454
rect 325222 434218 360986 434454
rect 361222 434218 396986 434454
rect 397222 434218 432986 434454
rect 433222 434218 468986 434454
rect 469222 434218 504986 434454
rect 505222 434218 540986 434454
rect 541222 434218 576986 434454
rect 577222 434218 585502 434454
rect 585738 434218 586840 434454
rect -2916 434134 586840 434218
rect -2916 433898 -1814 434134
rect -1578 433898 986 434134
rect 1222 433898 36986 434134
rect 37222 433898 72986 434134
rect 73222 433898 108986 434134
rect 109222 433898 144986 434134
rect 145222 433898 180986 434134
rect 181222 433898 216986 434134
rect 217222 433898 252986 434134
rect 253222 433898 288986 434134
rect 289222 433898 324986 434134
rect 325222 433898 360986 434134
rect 361222 433898 396986 434134
rect 397222 433898 432986 434134
rect 433222 433898 468986 434134
rect 469222 433898 504986 434134
rect 505222 433898 540986 434134
rect 541222 433898 576986 434134
rect 577222 433898 585502 434134
rect 585738 433898 586840 434134
rect -2916 433876 586840 433898
rect -1996 433874 -1396 433876
rect 804 433874 1404 433876
rect 36804 433874 37404 433876
rect 72804 433874 73404 433876
rect 108804 433874 109404 433876
rect 144804 433874 145404 433876
rect 180804 433874 181404 433876
rect 216804 433874 217404 433876
rect 252804 433874 253404 433876
rect 288804 433874 289404 433876
rect 324804 433874 325404 433876
rect 360804 433874 361404 433876
rect 396804 433874 397404 433876
rect 432804 433874 433404 433876
rect 468804 433874 469404 433876
rect 504804 433874 505404 433876
rect 540804 433874 541404 433876
rect 576804 433874 577404 433876
rect 585320 433874 585920 433876
rect -8436 427276 -7836 427278
rect 29604 427276 30204 427278
rect 65604 427276 66204 427278
rect 101604 427276 102204 427278
rect 137604 427276 138204 427278
rect 173604 427276 174204 427278
rect 209604 427276 210204 427278
rect 245604 427276 246204 427278
rect 281604 427276 282204 427278
rect 317604 427276 318204 427278
rect 353604 427276 354204 427278
rect 389604 427276 390204 427278
rect 425604 427276 426204 427278
rect 461604 427276 462204 427278
rect 497604 427276 498204 427278
rect 533604 427276 534204 427278
rect 569604 427276 570204 427278
rect 591760 427276 592360 427278
rect -8436 427254 592360 427276
rect -8436 427018 -8254 427254
rect -8018 427018 29786 427254
rect 30022 427018 65786 427254
rect 66022 427018 101786 427254
rect 102022 427018 137786 427254
rect 138022 427018 173786 427254
rect 174022 427018 209786 427254
rect 210022 427018 245786 427254
rect 246022 427018 281786 427254
rect 282022 427018 317786 427254
rect 318022 427018 353786 427254
rect 354022 427018 389786 427254
rect 390022 427018 425786 427254
rect 426022 427018 461786 427254
rect 462022 427018 497786 427254
rect 498022 427018 533786 427254
rect 534022 427018 569786 427254
rect 570022 427018 591942 427254
rect 592178 427018 592360 427254
rect -8436 426934 592360 427018
rect -8436 426698 -8254 426934
rect -8018 426698 29786 426934
rect 30022 426698 65786 426934
rect 66022 426698 101786 426934
rect 102022 426698 137786 426934
rect 138022 426698 173786 426934
rect 174022 426698 209786 426934
rect 210022 426698 245786 426934
rect 246022 426698 281786 426934
rect 282022 426698 317786 426934
rect 318022 426698 353786 426934
rect 354022 426698 389786 426934
rect 390022 426698 425786 426934
rect 426022 426698 461786 426934
rect 462022 426698 497786 426934
rect 498022 426698 533786 426934
rect 534022 426698 569786 426934
rect 570022 426698 591942 426934
rect 592178 426698 592360 426934
rect -8436 426676 592360 426698
rect -8436 426674 -7836 426676
rect 29604 426674 30204 426676
rect 65604 426674 66204 426676
rect 101604 426674 102204 426676
rect 137604 426674 138204 426676
rect 173604 426674 174204 426676
rect 209604 426674 210204 426676
rect 245604 426674 246204 426676
rect 281604 426674 282204 426676
rect 317604 426674 318204 426676
rect 353604 426674 354204 426676
rect 389604 426674 390204 426676
rect 425604 426674 426204 426676
rect 461604 426674 462204 426676
rect 497604 426674 498204 426676
rect 533604 426674 534204 426676
rect 569604 426674 570204 426676
rect 591760 426674 592360 426676
rect -6596 423676 -5996 423678
rect 26004 423676 26604 423678
rect 62004 423676 62604 423678
rect 98004 423676 98604 423678
rect 134004 423676 134604 423678
rect 170004 423676 170604 423678
rect 206004 423676 206604 423678
rect 242004 423676 242604 423678
rect 278004 423676 278604 423678
rect 314004 423676 314604 423678
rect 350004 423676 350604 423678
rect 386004 423676 386604 423678
rect 422004 423676 422604 423678
rect 458004 423676 458604 423678
rect 494004 423676 494604 423678
rect 530004 423676 530604 423678
rect 566004 423676 566604 423678
rect 589920 423676 590520 423678
rect -6596 423654 590520 423676
rect -6596 423418 -6414 423654
rect -6178 423418 26186 423654
rect 26422 423418 62186 423654
rect 62422 423418 98186 423654
rect 98422 423418 134186 423654
rect 134422 423418 170186 423654
rect 170422 423418 206186 423654
rect 206422 423418 242186 423654
rect 242422 423418 278186 423654
rect 278422 423418 314186 423654
rect 314422 423418 350186 423654
rect 350422 423418 386186 423654
rect 386422 423418 422186 423654
rect 422422 423418 458186 423654
rect 458422 423418 494186 423654
rect 494422 423418 530186 423654
rect 530422 423418 566186 423654
rect 566422 423418 590102 423654
rect 590338 423418 590520 423654
rect -6596 423334 590520 423418
rect -6596 423098 -6414 423334
rect -6178 423098 26186 423334
rect 26422 423098 62186 423334
rect 62422 423098 98186 423334
rect 98422 423098 134186 423334
rect 134422 423098 170186 423334
rect 170422 423098 206186 423334
rect 206422 423098 242186 423334
rect 242422 423098 278186 423334
rect 278422 423098 314186 423334
rect 314422 423098 350186 423334
rect 350422 423098 386186 423334
rect 386422 423098 422186 423334
rect 422422 423098 458186 423334
rect 458422 423098 494186 423334
rect 494422 423098 530186 423334
rect 530422 423098 566186 423334
rect 566422 423098 590102 423334
rect 590338 423098 590520 423334
rect -6596 423076 590520 423098
rect -6596 423074 -5996 423076
rect 26004 423074 26604 423076
rect 62004 423074 62604 423076
rect 98004 423074 98604 423076
rect 134004 423074 134604 423076
rect 170004 423074 170604 423076
rect 206004 423074 206604 423076
rect 242004 423074 242604 423076
rect 278004 423074 278604 423076
rect 314004 423074 314604 423076
rect 350004 423074 350604 423076
rect 386004 423074 386604 423076
rect 422004 423074 422604 423076
rect 458004 423074 458604 423076
rect 494004 423074 494604 423076
rect 530004 423074 530604 423076
rect 566004 423074 566604 423076
rect 589920 423074 590520 423076
rect -4756 420076 -4156 420078
rect 22404 420076 23004 420078
rect 58404 420076 59004 420078
rect 94404 420076 95004 420078
rect 130404 420076 131004 420078
rect 166404 420076 167004 420078
rect 202404 420076 203004 420078
rect 238404 420076 239004 420078
rect 274404 420076 275004 420078
rect 310404 420076 311004 420078
rect 346404 420076 347004 420078
rect 382404 420076 383004 420078
rect 418404 420076 419004 420078
rect 454404 420076 455004 420078
rect 490404 420076 491004 420078
rect 526404 420076 527004 420078
rect 562404 420076 563004 420078
rect 588080 420076 588680 420078
rect -4756 420054 588680 420076
rect -4756 419818 -4574 420054
rect -4338 419818 22586 420054
rect 22822 419818 58586 420054
rect 58822 419818 94586 420054
rect 94822 419818 130586 420054
rect 130822 419818 166586 420054
rect 166822 419818 202586 420054
rect 202822 419818 238586 420054
rect 238822 419818 274586 420054
rect 274822 419818 310586 420054
rect 310822 419818 346586 420054
rect 346822 419818 382586 420054
rect 382822 419818 418586 420054
rect 418822 419818 454586 420054
rect 454822 419818 490586 420054
rect 490822 419818 526586 420054
rect 526822 419818 562586 420054
rect 562822 419818 588262 420054
rect 588498 419818 588680 420054
rect -4756 419734 588680 419818
rect -4756 419498 -4574 419734
rect -4338 419498 22586 419734
rect 22822 419498 58586 419734
rect 58822 419498 94586 419734
rect 94822 419498 130586 419734
rect 130822 419498 166586 419734
rect 166822 419498 202586 419734
rect 202822 419498 238586 419734
rect 238822 419498 274586 419734
rect 274822 419498 310586 419734
rect 310822 419498 346586 419734
rect 346822 419498 382586 419734
rect 382822 419498 418586 419734
rect 418822 419498 454586 419734
rect 454822 419498 490586 419734
rect 490822 419498 526586 419734
rect 526822 419498 562586 419734
rect 562822 419498 588262 419734
rect 588498 419498 588680 419734
rect -4756 419476 588680 419498
rect -4756 419474 -4156 419476
rect 22404 419474 23004 419476
rect 58404 419474 59004 419476
rect 94404 419474 95004 419476
rect 130404 419474 131004 419476
rect 166404 419474 167004 419476
rect 202404 419474 203004 419476
rect 238404 419474 239004 419476
rect 274404 419474 275004 419476
rect 310404 419474 311004 419476
rect 346404 419474 347004 419476
rect 382404 419474 383004 419476
rect 418404 419474 419004 419476
rect 454404 419474 455004 419476
rect 490404 419474 491004 419476
rect 526404 419474 527004 419476
rect 562404 419474 563004 419476
rect 588080 419474 588680 419476
rect -2916 416476 -2316 416478
rect 18804 416476 19404 416478
rect 54804 416476 55404 416478
rect 90804 416476 91404 416478
rect 126804 416476 127404 416478
rect 162804 416476 163404 416478
rect 198804 416476 199404 416478
rect 234804 416476 235404 416478
rect 270804 416476 271404 416478
rect 306804 416476 307404 416478
rect 342804 416476 343404 416478
rect 378804 416476 379404 416478
rect 414804 416476 415404 416478
rect 450804 416476 451404 416478
rect 486804 416476 487404 416478
rect 522804 416476 523404 416478
rect 558804 416476 559404 416478
rect 586240 416476 586840 416478
rect -2916 416454 586840 416476
rect -2916 416218 -2734 416454
rect -2498 416218 18986 416454
rect 19222 416218 54986 416454
rect 55222 416218 90986 416454
rect 91222 416218 126986 416454
rect 127222 416218 162986 416454
rect 163222 416218 198986 416454
rect 199222 416218 234986 416454
rect 235222 416218 270986 416454
rect 271222 416218 306986 416454
rect 307222 416218 342986 416454
rect 343222 416218 378986 416454
rect 379222 416218 414986 416454
rect 415222 416218 450986 416454
rect 451222 416218 486986 416454
rect 487222 416218 522986 416454
rect 523222 416218 558986 416454
rect 559222 416218 586422 416454
rect 586658 416218 586840 416454
rect -2916 416134 586840 416218
rect -2916 415898 -2734 416134
rect -2498 415898 18986 416134
rect 19222 415898 54986 416134
rect 55222 415898 90986 416134
rect 91222 415898 126986 416134
rect 127222 415898 162986 416134
rect 163222 415898 198986 416134
rect 199222 415898 234986 416134
rect 235222 415898 270986 416134
rect 271222 415898 306986 416134
rect 307222 415898 342986 416134
rect 343222 415898 378986 416134
rect 379222 415898 414986 416134
rect 415222 415898 450986 416134
rect 451222 415898 486986 416134
rect 487222 415898 522986 416134
rect 523222 415898 558986 416134
rect 559222 415898 586422 416134
rect 586658 415898 586840 416134
rect -2916 415876 586840 415898
rect -2916 415874 -2316 415876
rect 18804 415874 19404 415876
rect 54804 415874 55404 415876
rect 90804 415874 91404 415876
rect 126804 415874 127404 415876
rect 162804 415874 163404 415876
rect 198804 415874 199404 415876
rect 234804 415874 235404 415876
rect 270804 415874 271404 415876
rect 306804 415874 307404 415876
rect 342804 415874 343404 415876
rect 378804 415874 379404 415876
rect 414804 415874 415404 415876
rect 450804 415874 451404 415876
rect 486804 415874 487404 415876
rect 522804 415874 523404 415876
rect 558804 415874 559404 415876
rect 586240 415874 586840 415876
rect -7516 409276 -6916 409278
rect 11604 409276 12204 409278
rect 47604 409276 48204 409278
rect 83604 409276 84204 409278
rect 119604 409276 120204 409278
rect 155604 409276 156204 409278
rect 191604 409276 192204 409278
rect 227604 409276 228204 409278
rect 263604 409276 264204 409278
rect 299604 409276 300204 409278
rect 335604 409276 336204 409278
rect 371604 409276 372204 409278
rect 407604 409276 408204 409278
rect 443604 409276 444204 409278
rect 479604 409276 480204 409278
rect 515604 409276 516204 409278
rect 551604 409276 552204 409278
rect 590840 409276 591440 409278
rect -8436 409254 592360 409276
rect -8436 409018 -7334 409254
rect -7098 409018 11786 409254
rect 12022 409018 47786 409254
rect 48022 409018 83786 409254
rect 84022 409018 119786 409254
rect 120022 409018 155786 409254
rect 156022 409018 191786 409254
rect 192022 409018 227786 409254
rect 228022 409018 263786 409254
rect 264022 409018 299786 409254
rect 300022 409018 335786 409254
rect 336022 409018 371786 409254
rect 372022 409018 407786 409254
rect 408022 409018 443786 409254
rect 444022 409018 479786 409254
rect 480022 409018 515786 409254
rect 516022 409018 551786 409254
rect 552022 409018 591022 409254
rect 591258 409018 592360 409254
rect -8436 408934 592360 409018
rect -8436 408698 -7334 408934
rect -7098 408698 11786 408934
rect 12022 408698 47786 408934
rect 48022 408698 83786 408934
rect 84022 408698 119786 408934
rect 120022 408698 155786 408934
rect 156022 408698 191786 408934
rect 192022 408698 227786 408934
rect 228022 408698 263786 408934
rect 264022 408698 299786 408934
rect 300022 408698 335786 408934
rect 336022 408698 371786 408934
rect 372022 408698 407786 408934
rect 408022 408698 443786 408934
rect 444022 408698 479786 408934
rect 480022 408698 515786 408934
rect 516022 408698 551786 408934
rect 552022 408698 591022 408934
rect 591258 408698 592360 408934
rect -8436 408676 592360 408698
rect -7516 408674 -6916 408676
rect 11604 408674 12204 408676
rect 47604 408674 48204 408676
rect 83604 408674 84204 408676
rect 119604 408674 120204 408676
rect 155604 408674 156204 408676
rect 191604 408674 192204 408676
rect 227604 408674 228204 408676
rect 263604 408674 264204 408676
rect 299604 408674 300204 408676
rect 335604 408674 336204 408676
rect 371604 408674 372204 408676
rect 407604 408674 408204 408676
rect 443604 408674 444204 408676
rect 479604 408674 480204 408676
rect 515604 408674 516204 408676
rect 551604 408674 552204 408676
rect 590840 408674 591440 408676
rect -5676 405676 -5076 405678
rect 8004 405676 8604 405678
rect 44004 405676 44604 405678
rect 80004 405676 80604 405678
rect 116004 405676 116604 405678
rect 152004 405676 152604 405678
rect 188004 405676 188604 405678
rect 224004 405676 224604 405678
rect 260004 405676 260604 405678
rect 296004 405676 296604 405678
rect 332004 405676 332604 405678
rect 368004 405676 368604 405678
rect 404004 405676 404604 405678
rect 440004 405676 440604 405678
rect 476004 405676 476604 405678
rect 512004 405676 512604 405678
rect 548004 405676 548604 405678
rect 589000 405676 589600 405678
rect -6596 405654 590520 405676
rect -6596 405418 -5494 405654
rect -5258 405418 8186 405654
rect 8422 405418 44186 405654
rect 44422 405418 80186 405654
rect 80422 405418 116186 405654
rect 116422 405418 152186 405654
rect 152422 405418 188186 405654
rect 188422 405418 224186 405654
rect 224422 405418 260186 405654
rect 260422 405418 296186 405654
rect 296422 405418 332186 405654
rect 332422 405418 368186 405654
rect 368422 405418 404186 405654
rect 404422 405418 440186 405654
rect 440422 405418 476186 405654
rect 476422 405418 512186 405654
rect 512422 405418 548186 405654
rect 548422 405418 589182 405654
rect 589418 405418 590520 405654
rect -6596 405334 590520 405418
rect -6596 405098 -5494 405334
rect -5258 405098 8186 405334
rect 8422 405098 44186 405334
rect 44422 405098 80186 405334
rect 80422 405098 116186 405334
rect 116422 405098 152186 405334
rect 152422 405098 188186 405334
rect 188422 405098 224186 405334
rect 224422 405098 260186 405334
rect 260422 405098 296186 405334
rect 296422 405098 332186 405334
rect 332422 405098 368186 405334
rect 368422 405098 404186 405334
rect 404422 405098 440186 405334
rect 440422 405098 476186 405334
rect 476422 405098 512186 405334
rect 512422 405098 548186 405334
rect 548422 405098 589182 405334
rect 589418 405098 590520 405334
rect -6596 405076 590520 405098
rect -5676 405074 -5076 405076
rect 8004 405074 8604 405076
rect 44004 405074 44604 405076
rect 80004 405074 80604 405076
rect 116004 405074 116604 405076
rect 152004 405074 152604 405076
rect 188004 405074 188604 405076
rect 224004 405074 224604 405076
rect 260004 405074 260604 405076
rect 296004 405074 296604 405076
rect 332004 405074 332604 405076
rect 368004 405074 368604 405076
rect 404004 405074 404604 405076
rect 440004 405074 440604 405076
rect 476004 405074 476604 405076
rect 512004 405074 512604 405076
rect 548004 405074 548604 405076
rect 589000 405074 589600 405076
rect -3836 402076 -3236 402078
rect 4404 402076 5004 402078
rect 40404 402076 41004 402078
rect 76404 402076 77004 402078
rect 112404 402076 113004 402078
rect 148404 402076 149004 402078
rect 184404 402076 185004 402078
rect 220404 402076 221004 402078
rect 256404 402076 257004 402078
rect 292404 402076 293004 402078
rect 328404 402076 329004 402078
rect 364404 402076 365004 402078
rect 400404 402076 401004 402078
rect 436404 402076 437004 402078
rect 472404 402076 473004 402078
rect 508404 402076 509004 402078
rect 544404 402076 545004 402078
rect 580404 402076 581004 402078
rect 587160 402076 587760 402078
rect -4756 402054 588680 402076
rect -4756 401818 -3654 402054
rect -3418 401818 4586 402054
rect 4822 401818 40586 402054
rect 40822 401818 76586 402054
rect 76822 401818 112586 402054
rect 112822 401818 148586 402054
rect 148822 401818 184586 402054
rect 184822 401818 220586 402054
rect 220822 401818 256586 402054
rect 256822 401818 292586 402054
rect 292822 401818 328586 402054
rect 328822 401818 364586 402054
rect 364822 401818 400586 402054
rect 400822 401818 436586 402054
rect 436822 401818 472586 402054
rect 472822 401818 508586 402054
rect 508822 401818 544586 402054
rect 544822 401818 580586 402054
rect 580822 401818 587342 402054
rect 587578 401818 588680 402054
rect -4756 401734 588680 401818
rect -4756 401498 -3654 401734
rect -3418 401498 4586 401734
rect 4822 401498 40586 401734
rect 40822 401498 76586 401734
rect 76822 401498 112586 401734
rect 112822 401498 148586 401734
rect 148822 401498 184586 401734
rect 184822 401498 220586 401734
rect 220822 401498 256586 401734
rect 256822 401498 292586 401734
rect 292822 401498 328586 401734
rect 328822 401498 364586 401734
rect 364822 401498 400586 401734
rect 400822 401498 436586 401734
rect 436822 401498 472586 401734
rect 472822 401498 508586 401734
rect 508822 401498 544586 401734
rect 544822 401498 580586 401734
rect 580822 401498 587342 401734
rect 587578 401498 588680 401734
rect -4756 401476 588680 401498
rect -3836 401474 -3236 401476
rect 4404 401474 5004 401476
rect 40404 401474 41004 401476
rect 76404 401474 77004 401476
rect 112404 401474 113004 401476
rect 148404 401474 149004 401476
rect 184404 401474 185004 401476
rect 220404 401474 221004 401476
rect 256404 401474 257004 401476
rect 292404 401474 293004 401476
rect 328404 401474 329004 401476
rect 364404 401474 365004 401476
rect 400404 401474 401004 401476
rect 436404 401474 437004 401476
rect 472404 401474 473004 401476
rect 508404 401474 509004 401476
rect 544404 401474 545004 401476
rect 580404 401474 581004 401476
rect 587160 401474 587760 401476
rect -1996 398476 -1396 398478
rect 804 398476 1404 398478
rect 36804 398476 37404 398478
rect 72804 398476 73404 398478
rect 108804 398476 109404 398478
rect 144804 398476 145404 398478
rect 180804 398476 181404 398478
rect 216804 398476 217404 398478
rect 252804 398476 253404 398478
rect 288804 398476 289404 398478
rect 324804 398476 325404 398478
rect 360804 398476 361404 398478
rect 396804 398476 397404 398478
rect 432804 398476 433404 398478
rect 468804 398476 469404 398478
rect 504804 398476 505404 398478
rect 540804 398476 541404 398478
rect 576804 398476 577404 398478
rect 585320 398476 585920 398478
rect -2916 398454 586840 398476
rect -2916 398218 -1814 398454
rect -1578 398218 986 398454
rect 1222 398218 36986 398454
rect 37222 398218 72986 398454
rect 73222 398218 108986 398454
rect 109222 398218 144986 398454
rect 145222 398218 180986 398454
rect 181222 398218 216986 398454
rect 217222 398218 252986 398454
rect 253222 398218 288986 398454
rect 289222 398218 324986 398454
rect 325222 398218 360986 398454
rect 361222 398218 396986 398454
rect 397222 398218 432986 398454
rect 433222 398218 468986 398454
rect 469222 398218 504986 398454
rect 505222 398218 540986 398454
rect 541222 398218 576986 398454
rect 577222 398218 585502 398454
rect 585738 398218 586840 398454
rect -2916 398134 586840 398218
rect -2916 397898 -1814 398134
rect -1578 397898 986 398134
rect 1222 397898 36986 398134
rect 37222 397898 72986 398134
rect 73222 397898 108986 398134
rect 109222 397898 144986 398134
rect 145222 397898 180986 398134
rect 181222 397898 216986 398134
rect 217222 397898 252986 398134
rect 253222 397898 288986 398134
rect 289222 397898 324986 398134
rect 325222 397898 360986 398134
rect 361222 397898 396986 398134
rect 397222 397898 432986 398134
rect 433222 397898 468986 398134
rect 469222 397898 504986 398134
rect 505222 397898 540986 398134
rect 541222 397898 576986 398134
rect 577222 397898 585502 398134
rect 585738 397898 586840 398134
rect -2916 397876 586840 397898
rect -1996 397874 -1396 397876
rect 804 397874 1404 397876
rect 36804 397874 37404 397876
rect 72804 397874 73404 397876
rect 108804 397874 109404 397876
rect 144804 397874 145404 397876
rect 180804 397874 181404 397876
rect 216804 397874 217404 397876
rect 252804 397874 253404 397876
rect 288804 397874 289404 397876
rect 324804 397874 325404 397876
rect 360804 397874 361404 397876
rect 396804 397874 397404 397876
rect 432804 397874 433404 397876
rect 468804 397874 469404 397876
rect 504804 397874 505404 397876
rect 540804 397874 541404 397876
rect 576804 397874 577404 397876
rect 585320 397874 585920 397876
rect -8436 391276 -7836 391278
rect 29604 391276 30204 391278
rect 65604 391276 66204 391278
rect 101604 391276 102204 391278
rect 137604 391276 138204 391278
rect 173604 391276 174204 391278
rect 209604 391276 210204 391278
rect 245604 391276 246204 391278
rect 281604 391276 282204 391278
rect 317604 391276 318204 391278
rect 353604 391276 354204 391278
rect 389604 391276 390204 391278
rect 425604 391276 426204 391278
rect 461604 391276 462204 391278
rect 497604 391276 498204 391278
rect 533604 391276 534204 391278
rect 569604 391276 570204 391278
rect 591760 391276 592360 391278
rect -8436 391254 592360 391276
rect -8436 391018 -8254 391254
rect -8018 391018 29786 391254
rect 30022 391018 65786 391254
rect 66022 391018 101786 391254
rect 102022 391018 137786 391254
rect 138022 391018 173786 391254
rect 174022 391018 209786 391254
rect 210022 391018 245786 391254
rect 246022 391018 281786 391254
rect 282022 391018 317786 391254
rect 318022 391018 353786 391254
rect 354022 391018 389786 391254
rect 390022 391018 425786 391254
rect 426022 391018 461786 391254
rect 462022 391018 497786 391254
rect 498022 391018 533786 391254
rect 534022 391018 569786 391254
rect 570022 391018 591942 391254
rect 592178 391018 592360 391254
rect -8436 390934 592360 391018
rect -8436 390698 -8254 390934
rect -8018 390698 29786 390934
rect 30022 390698 65786 390934
rect 66022 390698 101786 390934
rect 102022 390698 137786 390934
rect 138022 390698 173786 390934
rect 174022 390698 209786 390934
rect 210022 390698 245786 390934
rect 246022 390698 281786 390934
rect 282022 390698 317786 390934
rect 318022 390698 353786 390934
rect 354022 390698 389786 390934
rect 390022 390698 425786 390934
rect 426022 390698 461786 390934
rect 462022 390698 497786 390934
rect 498022 390698 533786 390934
rect 534022 390698 569786 390934
rect 570022 390698 591942 390934
rect 592178 390698 592360 390934
rect -8436 390676 592360 390698
rect -8436 390674 -7836 390676
rect 29604 390674 30204 390676
rect 65604 390674 66204 390676
rect 101604 390674 102204 390676
rect 137604 390674 138204 390676
rect 173604 390674 174204 390676
rect 209604 390674 210204 390676
rect 245604 390674 246204 390676
rect 281604 390674 282204 390676
rect 317604 390674 318204 390676
rect 353604 390674 354204 390676
rect 389604 390674 390204 390676
rect 425604 390674 426204 390676
rect 461604 390674 462204 390676
rect 497604 390674 498204 390676
rect 533604 390674 534204 390676
rect 569604 390674 570204 390676
rect 591760 390674 592360 390676
rect -6596 387676 -5996 387678
rect 26004 387676 26604 387678
rect 62004 387676 62604 387678
rect 98004 387676 98604 387678
rect 134004 387676 134604 387678
rect 170004 387676 170604 387678
rect 206004 387676 206604 387678
rect 242004 387676 242604 387678
rect 278004 387676 278604 387678
rect 314004 387676 314604 387678
rect 350004 387676 350604 387678
rect 386004 387676 386604 387678
rect 422004 387676 422604 387678
rect 458004 387676 458604 387678
rect 494004 387676 494604 387678
rect 530004 387676 530604 387678
rect 566004 387676 566604 387678
rect 589920 387676 590520 387678
rect -6596 387654 590520 387676
rect -6596 387418 -6414 387654
rect -6178 387418 26186 387654
rect 26422 387418 62186 387654
rect 62422 387418 98186 387654
rect 98422 387418 134186 387654
rect 134422 387418 170186 387654
rect 170422 387418 206186 387654
rect 206422 387418 242186 387654
rect 242422 387418 278186 387654
rect 278422 387418 314186 387654
rect 314422 387418 350186 387654
rect 350422 387418 386186 387654
rect 386422 387418 422186 387654
rect 422422 387418 458186 387654
rect 458422 387418 494186 387654
rect 494422 387418 530186 387654
rect 530422 387418 566186 387654
rect 566422 387418 590102 387654
rect 590338 387418 590520 387654
rect -6596 387334 590520 387418
rect -6596 387098 -6414 387334
rect -6178 387098 26186 387334
rect 26422 387098 62186 387334
rect 62422 387098 98186 387334
rect 98422 387098 134186 387334
rect 134422 387098 170186 387334
rect 170422 387098 206186 387334
rect 206422 387098 242186 387334
rect 242422 387098 278186 387334
rect 278422 387098 314186 387334
rect 314422 387098 350186 387334
rect 350422 387098 386186 387334
rect 386422 387098 422186 387334
rect 422422 387098 458186 387334
rect 458422 387098 494186 387334
rect 494422 387098 530186 387334
rect 530422 387098 566186 387334
rect 566422 387098 590102 387334
rect 590338 387098 590520 387334
rect -6596 387076 590520 387098
rect -6596 387074 -5996 387076
rect 26004 387074 26604 387076
rect 62004 387074 62604 387076
rect 98004 387074 98604 387076
rect 134004 387074 134604 387076
rect 170004 387074 170604 387076
rect 206004 387074 206604 387076
rect 242004 387074 242604 387076
rect 278004 387074 278604 387076
rect 314004 387074 314604 387076
rect 350004 387074 350604 387076
rect 386004 387074 386604 387076
rect 422004 387074 422604 387076
rect 458004 387074 458604 387076
rect 494004 387074 494604 387076
rect 530004 387074 530604 387076
rect 566004 387074 566604 387076
rect 589920 387074 590520 387076
rect -4756 384076 -4156 384078
rect 22404 384076 23004 384078
rect 58404 384076 59004 384078
rect 94404 384076 95004 384078
rect 130404 384076 131004 384078
rect 166404 384076 167004 384078
rect 202404 384076 203004 384078
rect 238404 384076 239004 384078
rect 274404 384076 275004 384078
rect 310404 384076 311004 384078
rect 346404 384076 347004 384078
rect 382404 384076 383004 384078
rect 418404 384076 419004 384078
rect 454404 384076 455004 384078
rect 490404 384076 491004 384078
rect 526404 384076 527004 384078
rect 562404 384076 563004 384078
rect 588080 384076 588680 384078
rect -4756 384054 588680 384076
rect -4756 383818 -4574 384054
rect -4338 383818 22586 384054
rect 22822 383818 58586 384054
rect 58822 383818 94586 384054
rect 94822 383818 130586 384054
rect 130822 383818 166586 384054
rect 166822 383818 202586 384054
rect 202822 383818 238586 384054
rect 238822 383818 274586 384054
rect 274822 383818 310586 384054
rect 310822 383818 346586 384054
rect 346822 383818 382586 384054
rect 382822 383818 418586 384054
rect 418822 383818 454586 384054
rect 454822 383818 490586 384054
rect 490822 383818 526586 384054
rect 526822 383818 562586 384054
rect 562822 383818 588262 384054
rect 588498 383818 588680 384054
rect -4756 383734 588680 383818
rect -4756 383498 -4574 383734
rect -4338 383498 22586 383734
rect 22822 383498 58586 383734
rect 58822 383498 94586 383734
rect 94822 383498 130586 383734
rect 130822 383498 166586 383734
rect 166822 383498 202586 383734
rect 202822 383498 238586 383734
rect 238822 383498 274586 383734
rect 274822 383498 310586 383734
rect 310822 383498 346586 383734
rect 346822 383498 382586 383734
rect 382822 383498 418586 383734
rect 418822 383498 454586 383734
rect 454822 383498 490586 383734
rect 490822 383498 526586 383734
rect 526822 383498 562586 383734
rect 562822 383498 588262 383734
rect 588498 383498 588680 383734
rect -4756 383476 588680 383498
rect -4756 383474 -4156 383476
rect 22404 383474 23004 383476
rect 58404 383474 59004 383476
rect 94404 383474 95004 383476
rect 130404 383474 131004 383476
rect 166404 383474 167004 383476
rect 202404 383474 203004 383476
rect 238404 383474 239004 383476
rect 274404 383474 275004 383476
rect 310404 383474 311004 383476
rect 346404 383474 347004 383476
rect 382404 383474 383004 383476
rect 418404 383474 419004 383476
rect 454404 383474 455004 383476
rect 490404 383474 491004 383476
rect 526404 383474 527004 383476
rect 562404 383474 563004 383476
rect 588080 383474 588680 383476
rect -2916 380476 -2316 380478
rect 18804 380476 19404 380478
rect 54804 380476 55404 380478
rect 90804 380476 91404 380478
rect 126804 380476 127404 380478
rect 162804 380476 163404 380478
rect 198804 380476 199404 380478
rect 234804 380476 235404 380478
rect 270804 380476 271404 380478
rect 306804 380476 307404 380478
rect 342804 380476 343404 380478
rect 378804 380476 379404 380478
rect 414804 380476 415404 380478
rect 450804 380476 451404 380478
rect 486804 380476 487404 380478
rect 522804 380476 523404 380478
rect 558804 380476 559404 380478
rect 586240 380476 586840 380478
rect -2916 380454 586840 380476
rect -2916 380218 -2734 380454
rect -2498 380218 18986 380454
rect 19222 380218 54986 380454
rect 55222 380218 90986 380454
rect 91222 380218 126986 380454
rect 127222 380218 162986 380454
rect 163222 380218 198986 380454
rect 199222 380218 234986 380454
rect 235222 380218 270986 380454
rect 271222 380218 306986 380454
rect 307222 380218 342986 380454
rect 343222 380218 378986 380454
rect 379222 380218 414986 380454
rect 415222 380218 450986 380454
rect 451222 380218 486986 380454
rect 487222 380218 522986 380454
rect 523222 380218 558986 380454
rect 559222 380218 586422 380454
rect 586658 380218 586840 380454
rect -2916 380134 586840 380218
rect -2916 379898 -2734 380134
rect -2498 379898 18986 380134
rect 19222 379898 54986 380134
rect 55222 379898 90986 380134
rect 91222 379898 126986 380134
rect 127222 379898 162986 380134
rect 163222 379898 198986 380134
rect 199222 379898 234986 380134
rect 235222 379898 270986 380134
rect 271222 379898 306986 380134
rect 307222 379898 342986 380134
rect 343222 379898 378986 380134
rect 379222 379898 414986 380134
rect 415222 379898 450986 380134
rect 451222 379898 486986 380134
rect 487222 379898 522986 380134
rect 523222 379898 558986 380134
rect 559222 379898 586422 380134
rect 586658 379898 586840 380134
rect -2916 379876 586840 379898
rect -2916 379874 -2316 379876
rect 18804 379874 19404 379876
rect 54804 379874 55404 379876
rect 90804 379874 91404 379876
rect 126804 379874 127404 379876
rect 162804 379874 163404 379876
rect 198804 379874 199404 379876
rect 234804 379874 235404 379876
rect 270804 379874 271404 379876
rect 306804 379874 307404 379876
rect 342804 379874 343404 379876
rect 378804 379874 379404 379876
rect 414804 379874 415404 379876
rect 450804 379874 451404 379876
rect 486804 379874 487404 379876
rect 522804 379874 523404 379876
rect 558804 379874 559404 379876
rect 586240 379874 586840 379876
rect -7516 373276 -6916 373278
rect 11604 373276 12204 373278
rect 47604 373276 48204 373278
rect 83604 373276 84204 373278
rect 119604 373276 120204 373278
rect 155604 373276 156204 373278
rect 191604 373276 192204 373278
rect 227604 373276 228204 373278
rect 263604 373276 264204 373278
rect 299604 373276 300204 373278
rect 335604 373276 336204 373278
rect 371604 373276 372204 373278
rect 407604 373276 408204 373278
rect 443604 373276 444204 373278
rect 479604 373276 480204 373278
rect 515604 373276 516204 373278
rect 551604 373276 552204 373278
rect 590840 373276 591440 373278
rect -8436 373254 592360 373276
rect -8436 373018 -7334 373254
rect -7098 373018 11786 373254
rect 12022 373018 47786 373254
rect 48022 373018 83786 373254
rect 84022 373018 119786 373254
rect 120022 373018 155786 373254
rect 156022 373018 191786 373254
rect 192022 373018 227786 373254
rect 228022 373018 263786 373254
rect 264022 373018 299786 373254
rect 300022 373018 335786 373254
rect 336022 373018 371786 373254
rect 372022 373018 407786 373254
rect 408022 373018 443786 373254
rect 444022 373018 479786 373254
rect 480022 373018 515786 373254
rect 516022 373018 551786 373254
rect 552022 373018 591022 373254
rect 591258 373018 592360 373254
rect -8436 372934 592360 373018
rect -8436 372698 -7334 372934
rect -7098 372698 11786 372934
rect 12022 372698 47786 372934
rect 48022 372698 83786 372934
rect 84022 372698 119786 372934
rect 120022 372698 155786 372934
rect 156022 372698 191786 372934
rect 192022 372698 227786 372934
rect 228022 372698 263786 372934
rect 264022 372698 299786 372934
rect 300022 372698 335786 372934
rect 336022 372698 371786 372934
rect 372022 372698 407786 372934
rect 408022 372698 443786 372934
rect 444022 372698 479786 372934
rect 480022 372698 515786 372934
rect 516022 372698 551786 372934
rect 552022 372698 591022 372934
rect 591258 372698 592360 372934
rect -8436 372676 592360 372698
rect -7516 372674 -6916 372676
rect 11604 372674 12204 372676
rect 47604 372674 48204 372676
rect 83604 372674 84204 372676
rect 119604 372674 120204 372676
rect 155604 372674 156204 372676
rect 191604 372674 192204 372676
rect 227604 372674 228204 372676
rect 263604 372674 264204 372676
rect 299604 372674 300204 372676
rect 335604 372674 336204 372676
rect 371604 372674 372204 372676
rect 407604 372674 408204 372676
rect 443604 372674 444204 372676
rect 479604 372674 480204 372676
rect 515604 372674 516204 372676
rect 551604 372674 552204 372676
rect 590840 372674 591440 372676
rect -5676 369676 -5076 369678
rect 8004 369676 8604 369678
rect 44004 369676 44604 369678
rect 80004 369676 80604 369678
rect 116004 369676 116604 369678
rect 152004 369676 152604 369678
rect 188004 369676 188604 369678
rect 224004 369676 224604 369678
rect 260004 369676 260604 369678
rect 296004 369676 296604 369678
rect 332004 369676 332604 369678
rect 368004 369676 368604 369678
rect 404004 369676 404604 369678
rect 440004 369676 440604 369678
rect 476004 369676 476604 369678
rect 512004 369676 512604 369678
rect 548004 369676 548604 369678
rect 589000 369676 589600 369678
rect -6596 369654 590520 369676
rect -6596 369418 -5494 369654
rect -5258 369418 8186 369654
rect 8422 369418 44186 369654
rect 44422 369418 80186 369654
rect 80422 369418 116186 369654
rect 116422 369418 152186 369654
rect 152422 369418 188186 369654
rect 188422 369418 224186 369654
rect 224422 369418 260186 369654
rect 260422 369418 296186 369654
rect 296422 369418 332186 369654
rect 332422 369418 368186 369654
rect 368422 369418 404186 369654
rect 404422 369418 440186 369654
rect 440422 369418 476186 369654
rect 476422 369418 512186 369654
rect 512422 369418 548186 369654
rect 548422 369418 589182 369654
rect 589418 369418 590520 369654
rect -6596 369334 590520 369418
rect -6596 369098 -5494 369334
rect -5258 369098 8186 369334
rect 8422 369098 44186 369334
rect 44422 369098 80186 369334
rect 80422 369098 116186 369334
rect 116422 369098 152186 369334
rect 152422 369098 188186 369334
rect 188422 369098 224186 369334
rect 224422 369098 260186 369334
rect 260422 369098 296186 369334
rect 296422 369098 332186 369334
rect 332422 369098 368186 369334
rect 368422 369098 404186 369334
rect 404422 369098 440186 369334
rect 440422 369098 476186 369334
rect 476422 369098 512186 369334
rect 512422 369098 548186 369334
rect 548422 369098 589182 369334
rect 589418 369098 590520 369334
rect -6596 369076 590520 369098
rect -5676 369074 -5076 369076
rect 8004 369074 8604 369076
rect 44004 369074 44604 369076
rect 80004 369074 80604 369076
rect 116004 369074 116604 369076
rect 152004 369074 152604 369076
rect 188004 369074 188604 369076
rect 224004 369074 224604 369076
rect 260004 369074 260604 369076
rect 296004 369074 296604 369076
rect 332004 369074 332604 369076
rect 368004 369074 368604 369076
rect 404004 369074 404604 369076
rect 440004 369074 440604 369076
rect 476004 369074 476604 369076
rect 512004 369074 512604 369076
rect 548004 369074 548604 369076
rect 589000 369074 589600 369076
rect -3836 366076 -3236 366078
rect 4404 366076 5004 366078
rect 40404 366076 41004 366078
rect 76404 366076 77004 366078
rect 112404 366076 113004 366078
rect 148404 366076 149004 366078
rect 184404 366076 185004 366078
rect 220404 366076 221004 366078
rect 256404 366076 257004 366078
rect 292404 366076 293004 366078
rect 328404 366076 329004 366078
rect 364404 366076 365004 366078
rect 400404 366076 401004 366078
rect 436404 366076 437004 366078
rect 472404 366076 473004 366078
rect 508404 366076 509004 366078
rect 544404 366076 545004 366078
rect 580404 366076 581004 366078
rect 587160 366076 587760 366078
rect -4756 366054 588680 366076
rect -4756 365818 -3654 366054
rect -3418 365818 4586 366054
rect 4822 365818 40586 366054
rect 40822 365818 76586 366054
rect 76822 365818 112586 366054
rect 112822 365818 148586 366054
rect 148822 365818 184586 366054
rect 184822 365818 220586 366054
rect 220822 365818 256586 366054
rect 256822 365818 292586 366054
rect 292822 365818 328586 366054
rect 328822 365818 364586 366054
rect 364822 365818 400586 366054
rect 400822 365818 436586 366054
rect 436822 365818 472586 366054
rect 472822 365818 508586 366054
rect 508822 365818 544586 366054
rect 544822 365818 580586 366054
rect 580822 365818 587342 366054
rect 587578 365818 588680 366054
rect -4756 365734 588680 365818
rect -4756 365498 -3654 365734
rect -3418 365498 4586 365734
rect 4822 365498 40586 365734
rect 40822 365498 76586 365734
rect 76822 365498 112586 365734
rect 112822 365498 148586 365734
rect 148822 365498 184586 365734
rect 184822 365498 220586 365734
rect 220822 365498 256586 365734
rect 256822 365498 292586 365734
rect 292822 365498 328586 365734
rect 328822 365498 364586 365734
rect 364822 365498 400586 365734
rect 400822 365498 436586 365734
rect 436822 365498 472586 365734
rect 472822 365498 508586 365734
rect 508822 365498 544586 365734
rect 544822 365498 580586 365734
rect 580822 365498 587342 365734
rect 587578 365498 588680 365734
rect -4756 365476 588680 365498
rect -3836 365474 -3236 365476
rect 4404 365474 5004 365476
rect 40404 365474 41004 365476
rect 76404 365474 77004 365476
rect 112404 365474 113004 365476
rect 148404 365474 149004 365476
rect 184404 365474 185004 365476
rect 220404 365474 221004 365476
rect 256404 365474 257004 365476
rect 292404 365474 293004 365476
rect 328404 365474 329004 365476
rect 364404 365474 365004 365476
rect 400404 365474 401004 365476
rect 436404 365474 437004 365476
rect 472404 365474 473004 365476
rect 508404 365474 509004 365476
rect 544404 365474 545004 365476
rect 580404 365474 581004 365476
rect 587160 365474 587760 365476
rect -1996 362476 -1396 362478
rect 804 362476 1404 362478
rect 36804 362476 37404 362478
rect 72804 362476 73404 362478
rect 108804 362476 109404 362478
rect 144804 362476 145404 362478
rect 180804 362476 181404 362478
rect 216804 362476 217404 362478
rect 252804 362476 253404 362478
rect 288804 362476 289404 362478
rect 324804 362476 325404 362478
rect 360804 362476 361404 362478
rect 396804 362476 397404 362478
rect 432804 362476 433404 362478
rect 468804 362476 469404 362478
rect 504804 362476 505404 362478
rect 540804 362476 541404 362478
rect 576804 362476 577404 362478
rect 585320 362476 585920 362478
rect -2916 362454 586840 362476
rect -2916 362218 -1814 362454
rect -1578 362218 986 362454
rect 1222 362218 36986 362454
rect 37222 362218 72986 362454
rect 73222 362218 108986 362454
rect 109222 362218 144986 362454
rect 145222 362218 180986 362454
rect 181222 362218 216986 362454
rect 217222 362218 252986 362454
rect 253222 362218 288986 362454
rect 289222 362218 324986 362454
rect 325222 362218 360986 362454
rect 361222 362218 396986 362454
rect 397222 362218 432986 362454
rect 433222 362218 468986 362454
rect 469222 362218 504986 362454
rect 505222 362218 540986 362454
rect 541222 362218 576986 362454
rect 577222 362218 585502 362454
rect 585738 362218 586840 362454
rect -2916 362134 586840 362218
rect -2916 361898 -1814 362134
rect -1578 361898 986 362134
rect 1222 361898 36986 362134
rect 37222 361898 72986 362134
rect 73222 361898 108986 362134
rect 109222 361898 144986 362134
rect 145222 361898 180986 362134
rect 181222 361898 216986 362134
rect 217222 361898 252986 362134
rect 253222 361898 288986 362134
rect 289222 361898 324986 362134
rect 325222 361898 360986 362134
rect 361222 361898 396986 362134
rect 397222 361898 432986 362134
rect 433222 361898 468986 362134
rect 469222 361898 504986 362134
rect 505222 361898 540986 362134
rect 541222 361898 576986 362134
rect 577222 361898 585502 362134
rect 585738 361898 586840 362134
rect -2916 361876 586840 361898
rect -1996 361874 -1396 361876
rect 804 361874 1404 361876
rect 36804 361874 37404 361876
rect 72804 361874 73404 361876
rect 108804 361874 109404 361876
rect 144804 361874 145404 361876
rect 180804 361874 181404 361876
rect 216804 361874 217404 361876
rect 252804 361874 253404 361876
rect 288804 361874 289404 361876
rect 324804 361874 325404 361876
rect 360804 361874 361404 361876
rect 396804 361874 397404 361876
rect 432804 361874 433404 361876
rect 468804 361874 469404 361876
rect 504804 361874 505404 361876
rect 540804 361874 541404 361876
rect 576804 361874 577404 361876
rect 585320 361874 585920 361876
rect -8436 355276 -7836 355278
rect 29604 355276 30204 355278
rect 65604 355276 66204 355278
rect 101604 355276 102204 355278
rect 137604 355276 138204 355278
rect 173604 355276 174204 355278
rect 209604 355276 210204 355278
rect 245604 355276 246204 355278
rect 281604 355276 282204 355278
rect 317604 355276 318204 355278
rect 353604 355276 354204 355278
rect 389604 355276 390204 355278
rect 425604 355276 426204 355278
rect 461604 355276 462204 355278
rect 497604 355276 498204 355278
rect 533604 355276 534204 355278
rect 569604 355276 570204 355278
rect 591760 355276 592360 355278
rect -8436 355254 592360 355276
rect -8436 355018 -8254 355254
rect -8018 355018 29786 355254
rect 30022 355018 65786 355254
rect 66022 355018 101786 355254
rect 102022 355018 137786 355254
rect 138022 355018 173786 355254
rect 174022 355018 209786 355254
rect 210022 355018 245786 355254
rect 246022 355018 281786 355254
rect 282022 355018 317786 355254
rect 318022 355018 353786 355254
rect 354022 355018 389786 355254
rect 390022 355018 425786 355254
rect 426022 355018 461786 355254
rect 462022 355018 497786 355254
rect 498022 355018 533786 355254
rect 534022 355018 569786 355254
rect 570022 355018 591942 355254
rect 592178 355018 592360 355254
rect -8436 354934 592360 355018
rect -8436 354698 -8254 354934
rect -8018 354698 29786 354934
rect 30022 354698 65786 354934
rect 66022 354698 101786 354934
rect 102022 354698 137786 354934
rect 138022 354698 173786 354934
rect 174022 354698 209786 354934
rect 210022 354698 245786 354934
rect 246022 354698 281786 354934
rect 282022 354698 317786 354934
rect 318022 354698 353786 354934
rect 354022 354698 389786 354934
rect 390022 354698 425786 354934
rect 426022 354698 461786 354934
rect 462022 354698 497786 354934
rect 498022 354698 533786 354934
rect 534022 354698 569786 354934
rect 570022 354698 591942 354934
rect 592178 354698 592360 354934
rect -8436 354676 592360 354698
rect -8436 354674 -7836 354676
rect 29604 354674 30204 354676
rect 65604 354674 66204 354676
rect 101604 354674 102204 354676
rect 137604 354674 138204 354676
rect 173604 354674 174204 354676
rect 209604 354674 210204 354676
rect 245604 354674 246204 354676
rect 281604 354674 282204 354676
rect 317604 354674 318204 354676
rect 353604 354674 354204 354676
rect 389604 354674 390204 354676
rect 425604 354674 426204 354676
rect 461604 354674 462204 354676
rect 497604 354674 498204 354676
rect 533604 354674 534204 354676
rect 569604 354674 570204 354676
rect 591760 354674 592360 354676
rect -6596 351676 -5996 351678
rect 26004 351676 26604 351678
rect 62004 351676 62604 351678
rect 98004 351676 98604 351678
rect 134004 351676 134604 351678
rect 170004 351676 170604 351678
rect 206004 351676 206604 351678
rect 242004 351676 242604 351678
rect 278004 351676 278604 351678
rect 314004 351676 314604 351678
rect 350004 351676 350604 351678
rect 386004 351676 386604 351678
rect 422004 351676 422604 351678
rect 458004 351676 458604 351678
rect 494004 351676 494604 351678
rect 530004 351676 530604 351678
rect 566004 351676 566604 351678
rect 589920 351676 590520 351678
rect -6596 351654 590520 351676
rect -6596 351418 -6414 351654
rect -6178 351418 26186 351654
rect 26422 351418 62186 351654
rect 62422 351418 98186 351654
rect 98422 351418 134186 351654
rect 134422 351418 170186 351654
rect 170422 351418 206186 351654
rect 206422 351418 242186 351654
rect 242422 351418 278186 351654
rect 278422 351418 314186 351654
rect 314422 351418 350186 351654
rect 350422 351418 386186 351654
rect 386422 351418 422186 351654
rect 422422 351418 458186 351654
rect 458422 351418 494186 351654
rect 494422 351418 530186 351654
rect 530422 351418 566186 351654
rect 566422 351418 590102 351654
rect 590338 351418 590520 351654
rect -6596 351334 590520 351418
rect -6596 351098 -6414 351334
rect -6178 351098 26186 351334
rect 26422 351098 62186 351334
rect 62422 351098 98186 351334
rect 98422 351098 134186 351334
rect 134422 351098 170186 351334
rect 170422 351098 206186 351334
rect 206422 351098 242186 351334
rect 242422 351098 278186 351334
rect 278422 351098 314186 351334
rect 314422 351098 350186 351334
rect 350422 351098 386186 351334
rect 386422 351098 422186 351334
rect 422422 351098 458186 351334
rect 458422 351098 494186 351334
rect 494422 351098 530186 351334
rect 530422 351098 566186 351334
rect 566422 351098 590102 351334
rect 590338 351098 590520 351334
rect -6596 351076 590520 351098
rect -6596 351074 -5996 351076
rect 26004 351074 26604 351076
rect 62004 351074 62604 351076
rect 98004 351074 98604 351076
rect 134004 351074 134604 351076
rect 170004 351074 170604 351076
rect 206004 351074 206604 351076
rect 242004 351074 242604 351076
rect 278004 351074 278604 351076
rect 314004 351074 314604 351076
rect 350004 351074 350604 351076
rect 386004 351074 386604 351076
rect 422004 351074 422604 351076
rect 458004 351074 458604 351076
rect 494004 351074 494604 351076
rect 530004 351074 530604 351076
rect 566004 351074 566604 351076
rect 589920 351074 590520 351076
rect -4756 348076 -4156 348078
rect 22404 348076 23004 348078
rect 58404 348076 59004 348078
rect 94404 348076 95004 348078
rect 130404 348076 131004 348078
rect 166404 348076 167004 348078
rect 202404 348076 203004 348078
rect 238404 348076 239004 348078
rect 274404 348076 275004 348078
rect 310404 348076 311004 348078
rect 346404 348076 347004 348078
rect 382404 348076 383004 348078
rect 418404 348076 419004 348078
rect 454404 348076 455004 348078
rect 490404 348076 491004 348078
rect 526404 348076 527004 348078
rect 562404 348076 563004 348078
rect 588080 348076 588680 348078
rect -4756 348054 588680 348076
rect -4756 347818 -4574 348054
rect -4338 347818 22586 348054
rect 22822 347818 58586 348054
rect 58822 347818 94586 348054
rect 94822 347818 130586 348054
rect 130822 347818 166586 348054
rect 166822 347818 202586 348054
rect 202822 347818 238586 348054
rect 238822 347818 274586 348054
rect 274822 347818 310586 348054
rect 310822 347818 346586 348054
rect 346822 347818 382586 348054
rect 382822 347818 418586 348054
rect 418822 347818 454586 348054
rect 454822 347818 490586 348054
rect 490822 347818 526586 348054
rect 526822 347818 562586 348054
rect 562822 347818 588262 348054
rect 588498 347818 588680 348054
rect -4756 347734 588680 347818
rect -4756 347498 -4574 347734
rect -4338 347498 22586 347734
rect 22822 347498 58586 347734
rect 58822 347498 94586 347734
rect 94822 347498 130586 347734
rect 130822 347498 166586 347734
rect 166822 347498 202586 347734
rect 202822 347498 238586 347734
rect 238822 347498 274586 347734
rect 274822 347498 310586 347734
rect 310822 347498 346586 347734
rect 346822 347498 382586 347734
rect 382822 347498 418586 347734
rect 418822 347498 454586 347734
rect 454822 347498 490586 347734
rect 490822 347498 526586 347734
rect 526822 347498 562586 347734
rect 562822 347498 588262 347734
rect 588498 347498 588680 347734
rect -4756 347476 588680 347498
rect -4756 347474 -4156 347476
rect 22404 347474 23004 347476
rect 58404 347474 59004 347476
rect 94404 347474 95004 347476
rect 130404 347474 131004 347476
rect 166404 347474 167004 347476
rect 202404 347474 203004 347476
rect 238404 347474 239004 347476
rect 274404 347474 275004 347476
rect 310404 347474 311004 347476
rect 346404 347474 347004 347476
rect 382404 347474 383004 347476
rect 418404 347474 419004 347476
rect 454404 347474 455004 347476
rect 490404 347474 491004 347476
rect 526404 347474 527004 347476
rect 562404 347474 563004 347476
rect 588080 347474 588680 347476
rect -2916 344476 -2316 344478
rect 18804 344476 19404 344478
rect 54804 344476 55404 344478
rect 90804 344476 91404 344478
rect 126804 344476 127404 344478
rect 162804 344476 163404 344478
rect 198804 344476 199404 344478
rect 234804 344476 235404 344478
rect 270804 344476 271404 344478
rect 306804 344476 307404 344478
rect 342804 344476 343404 344478
rect 378804 344476 379404 344478
rect 414804 344476 415404 344478
rect 450804 344476 451404 344478
rect 486804 344476 487404 344478
rect 522804 344476 523404 344478
rect 558804 344476 559404 344478
rect 586240 344476 586840 344478
rect -2916 344454 586840 344476
rect -2916 344218 -2734 344454
rect -2498 344218 18986 344454
rect 19222 344218 54986 344454
rect 55222 344218 90986 344454
rect 91222 344218 126986 344454
rect 127222 344218 162986 344454
rect 163222 344218 198986 344454
rect 199222 344218 234986 344454
rect 235222 344218 270986 344454
rect 271222 344218 306986 344454
rect 307222 344218 342986 344454
rect 343222 344218 378986 344454
rect 379222 344218 414986 344454
rect 415222 344218 450986 344454
rect 451222 344218 486986 344454
rect 487222 344218 522986 344454
rect 523222 344218 558986 344454
rect 559222 344218 586422 344454
rect 586658 344218 586840 344454
rect -2916 344134 586840 344218
rect -2916 343898 -2734 344134
rect -2498 343898 18986 344134
rect 19222 343898 54986 344134
rect 55222 343898 90986 344134
rect 91222 343898 126986 344134
rect 127222 343898 162986 344134
rect 163222 343898 198986 344134
rect 199222 343898 234986 344134
rect 235222 343898 270986 344134
rect 271222 343898 306986 344134
rect 307222 343898 342986 344134
rect 343222 343898 378986 344134
rect 379222 343898 414986 344134
rect 415222 343898 450986 344134
rect 451222 343898 486986 344134
rect 487222 343898 522986 344134
rect 523222 343898 558986 344134
rect 559222 343898 586422 344134
rect 586658 343898 586840 344134
rect -2916 343876 586840 343898
rect -2916 343874 -2316 343876
rect 18804 343874 19404 343876
rect 54804 343874 55404 343876
rect 90804 343874 91404 343876
rect 126804 343874 127404 343876
rect 162804 343874 163404 343876
rect 198804 343874 199404 343876
rect 234804 343874 235404 343876
rect 270804 343874 271404 343876
rect 306804 343874 307404 343876
rect 342804 343874 343404 343876
rect 378804 343874 379404 343876
rect 414804 343874 415404 343876
rect 450804 343874 451404 343876
rect 486804 343874 487404 343876
rect 522804 343874 523404 343876
rect 558804 343874 559404 343876
rect 586240 343874 586840 343876
rect -7516 337276 -6916 337278
rect 11604 337276 12204 337278
rect 47604 337276 48204 337278
rect 83604 337276 84204 337278
rect 119604 337276 120204 337278
rect 155604 337276 156204 337278
rect 191604 337276 192204 337278
rect 227604 337276 228204 337278
rect 263604 337276 264204 337278
rect 299604 337276 300204 337278
rect 335604 337276 336204 337278
rect 371604 337276 372204 337278
rect 407604 337276 408204 337278
rect 443604 337276 444204 337278
rect 479604 337276 480204 337278
rect 515604 337276 516204 337278
rect 551604 337276 552204 337278
rect 590840 337276 591440 337278
rect -8436 337254 592360 337276
rect -8436 337018 -7334 337254
rect -7098 337018 11786 337254
rect 12022 337018 47786 337254
rect 48022 337018 83786 337254
rect 84022 337018 119786 337254
rect 120022 337018 155786 337254
rect 156022 337018 191786 337254
rect 192022 337018 227786 337254
rect 228022 337018 263786 337254
rect 264022 337018 299786 337254
rect 300022 337018 335786 337254
rect 336022 337018 371786 337254
rect 372022 337018 407786 337254
rect 408022 337018 443786 337254
rect 444022 337018 479786 337254
rect 480022 337018 515786 337254
rect 516022 337018 551786 337254
rect 552022 337018 591022 337254
rect 591258 337018 592360 337254
rect -8436 336934 592360 337018
rect -8436 336698 -7334 336934
rect -7098 336698 11786 336934
rect 12022 336698 47786 336934
rect 48022 336698 83786 336934
rect 84022 336698 119786 336934
rect 120022 336698 155786 336934
rect 156022 336698 191786 336934
rect 192022 336698 227786 336934
rect 228022 336698 263786 336934
rect 264022 336698 299786 336934
rect 300022 336698 335786 336934
rect 336022 336698 371786 336934
rect 372022 336698 407786 336934
rect 408022 336698 443786 336934
rect 444022 336698 479786 336934
rect 480022 336698 515786 336934
rect 516022 336698 551786 336934
rect 552022 336698 591022 336934
rect 591258 336698 592360 336934
rect -8436 336676 592360 336698
rect -7516 336674 -6916 336676
rect 11604 336674 12204 336676
rect 47604 336674 48204 336676
rect 83604 336674 84204 336676
rect 119604 336674 120204 336676
rect 155604 336674 156204 336676
rect 191604 336674 192204 336676
rect 227604 336674 228204 336676
rect 263604 336674 264204 336676
rect 299604 336674 300204 336676
rect 335604 336674 336204 336676
rect 371604 336674 372204 336676
rect 407604 336674 408204 336676
rect 443604 336674 444204 336676
rect 479604 336674 480204 336676
rect 515604 336674 516204 336676
rect 551604 336674 552204 336676
rect 590840 336674 591440 336676
rect -5676 333676 -5076 333678
rect 8004 333676 8604 333678
rect 44004 333676 44604 333678
rect 80004 333676 80604 333678
rect 116004 333676 116604 333678
rect 152004 333676 152604 333678
rect 188004 333676 188604 333678
rect 224004 333676 224604 333678
rect 260004 333676 260604 333678
rect 296004 333676 296604 333678
rect 332004 333676 332604 333678
rect 368004 333676 368604 333678
rect 404004 333676 404604 333678
rect 440004 333676 440604 333678
rect 476004 333676 476604 333678
rect 512004 333676 512604 333678
rect 548004 333676 548604 333678
rect 589000 333676 589600 333678
rect -6596 333654 590520 333676
rect -6596 333418 -5494 333654
rect -5258 333418 8186 333654
rect 8422 333418 44186 333654
rect 44422 333418 80186 333654
rect 80422 333418 116186 333654
rect 116422 333418 152186 333654
rect 152422 333418 188186 333654
rect 188422 333418 224186 333654
rect 224422 333418 260186 333654
rect 260422 333418 296186 333654
rect 296422 333418 332186 333654
rect 332422 333418 368186 333654
rect 368422 333418 404186 333654
rect 404422 333418 440186 333654
rect 440422 333418 476186 333654
rect 476422 333418 512186 333654
rect 512422 333418 548186 333654
rect 548422 333418 589182 333654
rect 589418 333418 590520 333654
rect -6596 333334 590520 333418
rect -6596 333098 -5494 333334
rect -5258 333098 8186 333334
rect 8422 333098 44186 333334
rect 44422 333098 80186 333334
rect 80422 333098 116186 333334
rect 116422 333098 152186 333334
rect 152422 333098 188186 333334
rect 188422 333098 224186 333334
rect 224422 333098 260186 333334
rect 260422 333098 296186 333334
rect 296422 333098 332186 333334
rect 332422 333098 368186 333334
rect 368422 333098 404186 333334
rect 404422 333098 440186 333334
rect 440422 333098 476186 333334
rect 476422 333098 512186 333334
rect 512422 333098 548186 333334
rect 548422 333098 589182 333334
rect 589418 333098 590520 333334
rect -6596 333076 590520 333098
rect -5676 333074 -5076 333076
rect 8004 333074 8604 333076
rect 44004 333074 44604 333076
rect 80004 333074 80604 333076
rect 116004 333074 116604 333076
rect 152004 333074 152604 333076
rect 188004 333074 188604 333076
rect 224004 333074 224604 333076
rect 260004 333074 260604 333076
rect 296004 333074 296604 333076
rect 332004 333074 332604 333076
rect 368004 333074 368604 333076
rect 404004 333074 404604 333076
rect 440004 333074 440604 333076
rect 476004 333074 476604 333076
rect 512004 333074 512604 333076
rect 548004 333074 548604 333076
rect 589000 333074 589600 333076
rect -3836 330076 -3236 330078
rect 4404 330076 5004 330078
rect 40404 330076 41004 330078
rect 76404 330076 77004 330078
rect 112404 330076 113004 330078
rect 148404 330076 149004 330078
rect 184404 330076 185004 330078
rect 220404 330076 221004 330078
rect 256404 330076 257004 330078
rect 292404 330076 293004 330078
rect 328404 330076 329004 330078
rect 364404 330076 365004 330078
rect 400404 330076 401004 330078
rect 436404 330076 437004 330078
rect 472404 330076 473004 330078
rect 508404 330076 509004 330078
rect 544404 330076 545004 330078
rect 580404 330076 581004 330078
rect 587160 330076 587760 330078
rect -4756 330054 588680 330076
rect -4756 329818 -3654 330054
rect -3418 329818 4586 330054
rect 4822 329818 40586 330054
rect 40822 329818 76586 330054
rect 76822 329818 112586 330054
rect 112822 329818 148586 330054
rect 148822 329818 184586 330054
rect 184822 329818 220586 330054
rect 220822 329818 256586 330054
rect 256822 329818 292586 330054
rect 292822 329818 328586 330054
rect 328822 329818 364586 330054
rect 364822 329818 400586 330054
rect 400822 329818 436586 330054
rect 436822 329818 472586 330054
rect 472822 329818 508586 330054
rect 508822 329818 544586 330054
rect 544822 329818 580586 330054
rect 580822 329818 587342 330054
rect 587578 329818 588680 330054
rect -4756 329734 588680 329818
rect -4756 329498 -3654 329734
rect -3418 329498 4586 329734
rect 4822 329498 40586 329734
rect 40822 329498 76586 329734
rect 76822 329498 112586 329734
rect 112822 329498 148586 329734
rect 148822 329498 184586 329734
rect 184822 329498 220586 329734
rect 220822 329498 256586 329734
rect 256822 329498 292586 329734
rect 292822 329498 328586 329734
rect 328822 329498 364586 329734
rect 364822 329498 400586 329734
rect 400822 329498 436586 329734
rect 436822 329498 472586 329734
rect 472822 329498 508586 329734
rect 508822 329498 544586 329734
rect 544822 329498 580586 329734
rect 580822 329498 587342 329734
rect 587578 329498 588680 329734
rect -4756 329476 588680 329498
rect -3836 329474 -3236 329476
rect 4404 329474 5004 329476
rect 40404 329474 41004 329476
rect 76404 329474 77004 329476
rect 112404 329474 113004 329476
rect 148404 329474 149004 329476
rect 184404 329474 185004 329476
rect 220404 329474 221004 329476
rect 256404 329474 257004 329476
rect 292404 329474 293004 329476
rect 328404 329474 329004 329476
rect 364404 329474 365004 329476
rect 400404 329474 401004 329476
rect 436404 329474 437004 329476
rect 472404 329474 473004 329476
rect 508404 329474 509004 329476
rect 544404 329474 545004 329476
rect 580404 329474 581004 329476
rect 587160 329474 587760 329476
rect -1996 326476 -1396 326478
rect 804 326476 1404 326478
rect 36804 326476 37404 326478
rect 72804 326476 73404 326478
rect 108804 326476 109404 326478
rect 144804 326476 145404 326478
rect 180804 326476 181404 326478
rect 216804 326476 217404 326478
rect 252804 326476 253404 326478
rect 288804 326476 289404 326478
rect 324804 326476 325404 326478
rect 360804 326476 361404 326478
rect 396804 326476 397404 326478
rect 432804 326476 433404 326478
rect 468804 326476 469404 326478
rect 504804 326476 505404 326478
rect 540804 326476 541404 326478
rect 576804 326476 577404 326478
rect 585320 326476 585920 326478
rect -2916 326454 586840 326476
rect -2916 326218 -1814 326454
rect -1578 326218 986 326454
rect 1222 326218 36986 326454
rect 37222 326218 72986 326454
rect 73222 326218 108986 326454
rect 109222 326218 144986 326454
rect 145222 326218 180986 326454
rect 181222 326218 216986 326454
rect 217222 326218 252986 326454
rect 253222 326218 288986 326454
rect 289222 326218 324986 326454
rect 325222 326218 360986 326454
rect 361222 326218 396986 326454
rect 397222 326218 432986 326454
rect 433222 326218 468986 326454
rect 469222 326218 504986 326454
rect 505222 326218 540986 326454
rect 541222 326218 576986 326454
rect 577222 326218 585502 326454
rect 585738 326218 586840 326454
rect -2916 326134 586840 326218
rect -2916 325898 -1814 326134
rect -1578 325898 986 326134
rect 1222 325898 36986 326134
rect 37222 325898 72986 326134
rect 73222 325898 108986 326134
rect 109222 325898 144986 326134
rect 145222 325898 180986 326134
rect 181222 325898 216986 326134
rect 217222 325898 252986 326134
rect 253222 325898 288986 326134
rect 289222 325898 324986 326134
rect 325222 325898 360986 326134
rect 361222 325898 396986 326134
rect 397222 325898 432986 326134
rect 433222 325898 468986 326134
rect 469222 325898 504986 326134
rect 505222 325898 540986 326134
rect 541222 325898 576986 326134
rect 577222 325898 585502 326134
rect 585738 325898 586840 326134
rect -2916 325876 586840 325898
rect -1996 325874 -1396 325876
rect 804 325874 1404 325876
rect 36804 325874 37404 325876
rect 72804 325874 73404 325876
rect 108804 325874 109404 325876
rect 144804 325874 145404 325876
rect 180804 325874 181404 325876
rect 216804 325874 217404 325876
rect 252804 325874 253404 325876
rect 288804 325874 289404 325876
rect 324804 325874 325404 325876
rect 360804 325874 361404 325876
rect 396804 325874 397404 325876
rect 432804 325874 433404 325876
rect 468804 325874 469404 325876
rect 504804 325874 505404 325876
rect 540804 325874 541404 325876
rect 576804 325874 577404 325876
rect 585320 325874 585920 325876
rect -8436 319276 -7836 319278
rect 29604 319276 30204 319278
rect 65604 319276 66204 319278
rect 101604 319276 102204 319278
rect 137604 319276 138204 319278
rect 173604 319276 174204 319278
rect 209604 319276 210204 319278
rect 245604 319276 246204 319278
rect 281604 319276 282204 319278
rect 317604 319276 318204 319278
rect 353604 319276 354204 319278
rect 389604 319276 390204 319278
rect 425604 319276 426204 319278
rect 461604 319276 462204 319278
rect 497604 319276 498204 319278
rect 533604 319276 534204 319278
rect 569604 319276 570204 319278
rect 591760 319276 592360 319278
rect -8436 319254 592360 319276
rect -8436 319018 -8254 319254
rect -8018 319018 29786 319254
rect 30022 319018 65786 319254
rect 66022 319018 101786 319254
rect 102022 319018 137786 319254
rect 138022 319018 173786 319254
rect 174022 319018 209786 319254
rect 210022 319018 245786 319254
rect 246022 319018 281786 319254
rect 282022 319018 317786 319254
rect 318022 319018 353786 319254
rect 354022 319018 389786 319254
rect 390022 319018 425786 319254
rect 426022 319018 461786 319254
rect 462022 319018 497786 319254
rect 498022 319018 533786 319254
rect 534022 319018 569786 319254
rect 570022 319018 591942 319254
rect 592178 319018 592360 319254
rect -8436 318934 592360 319018
rect -8436 318698 -8254 318934
rect -8018 318698 29786 318934
rect 30022 318698 65786 318934
rect 66022 318698 101786 318934
rect 102022 318698 137786 318934
rect 138022 318698 173786 318934
rect 174022 318698 209786 318934
rect 210022 318698 245786 318934
rect 246022 318698 281786 318934
rect 282022 318698 317786 318934
rect 318022 318698 353786 318934
rect 354022 318698 389786 318934
rect 390022 318698 425786 318934
rect 426022 318698 461786 318934
rect 462022 318698 497786 318934
rect 498022 318698 533786 318934
rect 534022 318698 569786 318934
rect 570022 318698 591942 318934
rect 592178 318698 592360 318934
rect -8436 318676 592360 318698
rect -8436 318674 -7836 318676
rect 29604 318674 30204 318676
rect 65604 318674 66204 318676
rect 101604 318674 102204 318676
rect 137604 318674 138204 318676
rect 173604 318674 174204 318676
rect 209604 318674 210204 318676
rect 245604 318674 246204 318676
rect 281604 318674 282204 318676
rect 317604 318674 318204 318676
rect 353604 318674 354204 318676
rect 389604 318674 390204 318676
rect 425604 318674 426204 318676
rect 461604 318674 462204 318676
rect 497604 318674 498204 318676
rect 533604 318674 534204 318676
rect 569604 318674 570204 318676
rect 591760 318674 592360 318676
rect -6596 315676 -5996 315678
rect 26004 315676 26604 315678
rect 62004 315676 62604 315678
rect 98004 315676 98604 315678
rect 134004 315676 134604 315678
rect 170004 315676 170604 315678
rect 206004 315676 206604 315678
rect 242004 315676 242604 315678
rect 278004 315676 278604 315678
rect 314004 315676 314604 315678
rect 350004 315676 350604 315678
rect 386004 315676 386604 315678
rect 422004 315676 422604 315678
rect 458004 315676 458604 315678
rect 494004 315676 494604 315678
rect 530004 315676 530604 315678
rect 566004 315676 566604 315678
rect 589920 315676 590520 315678
rect -6596 315654 590520 315676
rect -6596 315418 -6414 315654
rect -6178 315418 26186 315654
rect 26422 315418 62186 315654
rect 62422 315418 98186 315654
rect 98422 315418 134186 315654
rect 134422 315418 170186 315654
rect 170422 315418 206186 315654
rect 206422 315418 242186 315654
rect 242422 315418 278186 315654
rect 278422 315418 314186 315654
rect 314422 315418 350186 315654
rect 350422 315418 386186 315654
rect 386422 315418 422186 315654
rect 422422 315418 458186 315654
rect 458422 315418 494186 315654
rect 494422 315418 530186 315654
rect 530422 315418 566186 315654
rect 566422 315418 590102 315654
rect 590338 315418 590520 315654
rect -6596 315334 590520 315418
rect -6596 315098 -6414 315334
rect -6178 315098 26186 315334
rect 26422 315098 62186 315334
rect 62422 315098 98186 315334
rect 98422 315098 134186 315334
rect 134422 315098 170186 315334
rect 170422 315098 206186 315334
rect 206422 315098 242186 315334
rect 242422 315098 278186 315334
rect 278422 315098 314186 315334
rect 314422 315098 350186 315334
rect 350422 315098 386186 315334
rect 386422 315098 422186 315334
rect 422422 315098 458186 315334
rect 458422 315098 494186 315334
rect 494422 315098 530186 315334
rect 530422 315098 566186 315334
rect 566422 315098 590102 315334
rect 590338 315098 590520 315334
rect -6596 315076 590520 315098
rect -6596 315074 -5996 315076
rect 26004 315074 26604 315076
rect 62004 315074 62604 315076
rect 98004 315074 98604 315076
rect 134004 315074 134604 315076
rect 170004 315074 170604 315076
rect 206004 315074 206604 315076
rect 242004 315074 242604 315076
rect 278004 315074 278604 315076
rect 314004 315074 314604 315076
rect 350004 315074 350604 315076
rect 386004 315074 386604 315076
rect 422004 315074 422604 315076
rect 458004 315074 458604 315076
rect 494004 315074 494604 315076
rect 530004 315074 530604 315076
rect 566004 315074 566604 315076
rect 589920 315074 590520 315076
rect -4756 312076 -4156 312078
rect 22404 312076 23004 312078
rect 58404 312076 59004 312078
rect 94404 312076 95004 312078
rect 130404 312076 131004 312078
rect 166404 312076 167004 312078
rect 202404 312076 203004 312078
rect 238404 312076 239004 312078
rect 274404 312076 275004 312078
rect 310404 312076 311004 312078
rect 346404 312076 347004 312078
rect 382404 312076 383004 312078
rect 418404 312076 419004 312078
rect 454404 312076 455004 312078
rect 490404 312076 491004 312078
rect 526404 312076 527004 312078
rect 562404 312076 563004 312078
rect 588080 312076 588680 312078
rect -4756 312054 588680 312076
rect -4756 311818 -4574 312054
rect -4338 311818 22586 312054
rect 22822 311818 58586 312054
rect 58822 311818 94586 312054
rect 94822 311818 130586 312054
rect 130822 311818 166586 312054
rect 166822 311818 202586 312054
rect 202822 311818 238586 312054
rect 238822 311818 274586 312054
rect 274822 311818 310586 312054
rect 310822 311818 346586 312054
rect 346822 311818 382586 312054
rect 382822 311818 418586 312054
rect 418822 311818 454586 312054
rect 454822 311818 490586 312054
rect 490822 311818 526586 312054
rect 526822 311818 562586 312054
rect 562822 311818 588262 312054
rect 588498 311818 588680 312054
rect -4756 311734 588680 311818
rect -4756 311498 -4574 311734
rect -4338 311498 22586 311734
rect 22822 311498 58586 311734
rect 58822 311498 94586 311734
rect 94822 311498 130586 311734
rect 130822 311498 166586 311734
rect 166822 311498 202586 311734
rect 202822 311498 238586 311734
rect 238822 311498 274586 311734
rect 274822 311498 310586 311734
rect 310822 311498 346586 311734
rect 346822 311498 382586 311734
rect 382822 311498 418586 311734
rect 418822 311498 454586 311734
rect 454822 311498 490586 311734
rect 490822 311498 526586 311734
rect 526822 311498 562586 311734
rect 562822 311498 588262 311734
rect 588498 311498 588680 311734
rect -4756 311476 588680 311498
rect -4756 311474 -4156 311476
rect 22404 311474 23004 311476
rect 58404 311474 59004 311476
rect 94404 311474 95004 311476
rect 130404 311474 131004 311476
rect 166404 311474 167004 311476
rect 202404 311474 203004 311476
rect 238404 311474 239004 311476
rect 274404 311474 275004 311476
rect 310404 311474 311004 311476
rect 346404 311474 347004 311476
rect 382404 311474 383004 311476
rect 418404 311474 419004 311476
rect 454404 311474 455004 311476
rect 490404 311474 491004 311476
rect 526404 311474 527004 311476
rect 562404 311474 563004 311476
rect 588080 311474 588680 311476
rect -2916 308476 -2316 308478
rect 18804 308476 19404 308478
rect 54804 308476 55404 308478
rect 90804 308476 91404 308478
rect 126804 308476 127404 308478
rect 162804 308476 163404 308478
rect 198804 308476 199404 308478
rect 234804 308476 235404 308478
rect 270804 308476 271404 308478
rect 306804 308476 307404 308478
rect 342804 308476 343404 308478
rect 378804 308476 379404 308478
rect 414804 308476 415404 308478
rect 450804 308476 451404 308478
rect 486804 308476 487404 308478
rect 522804 308476 523404 308478
rect 558804 308476 559404 308478
rect 586240 308476 586840 308478
rect -2916 308454 586840 308476
rect -2916 308218 -2734 308454
rect -2498 308218 18986 308454
rect 19222 308218 54986 308454
rect 55222 308218 90986 308454
rect 91222 308218 126986 308454
rect 127222 308218 162986 308454
rect 163222 308218 198986 308454
rect 199222 308218 234986 308454
rect 235222 308218 270986 308454
rect 271222 308218 306986 308454
rect 307222 308218 342986 308454
rect 343222 308218 378986 308454
rect 379222 308218 414986 308454
rect 415222 308218 450986 308454
rect 451222 308218 486986 308454
rect 487222 308218 522986 308454
rect 523222 308218 558986 308454
rect 559222 308218 586422 308454
rect 586658 308218 586840 308454
rect -2916 308134 586840 308218
rect -2916 307898 -2734 308134
rect -2498 307898 18986 308134
rect 19222 307898 54986 308134
rect 55222 307898 90986 308134
rect 91222 307898 126986 308134
rect 127222 307898 162986 308134
rect 163222 307898 198986 308134
rect 199222 307898 234986 308134
rect 235222 307898 270986 308134
rect 271222 307898 306986 308134
rect 307222 307898 342986 308134
rect 343222 307898 378986 308134
rect 379222 307898 414986 308134
rect 415222 307898 450986 308134
rect 451222 307898 486986 308134
rect 487222 307898 522986 308134
rect 523222 307898 558986 308134
rect 559222 307898 586422 308134
rect 586658 307898 586840 308134
rect -2916 307876 586840 307898
rect -2916 307874 -2316 307876
rect 18804 307874 19404 307876
rect 54804 307874 55404 307876
rect 90804 307874 91404 307876
rect 126804 307874 127404 307876
rect 162804 307874 163404 307876
rect 198804 307874 199404 307876
rect 234804 307874 235404 307876
rect 270804 307874 271404 307876
rect 306804 307874 307404 307876
rect 342804 307874 343404 307876
rect 378804 307874 379404 307876
rect 414804 307874 415404 307876
rect 450804 307874 451404 307876
rect 486804 307874 487404 307876
rect 522804 307874 523404 307876
rect 558804 307874 559404 307876
rect 586240 307874 586840 307876
rect -7516 301276 -6916 301278
rect 11604 301276 12204 301278
rect 47604 301276 48204 301278
rect 83604 301276 84204 301278
rect 119604 301276 120204 301278
rect 155604 301276 156204 301278
rect 191604 301276 192204 301278
rect 227604 301276 228204 301278
rect 263604 301276 264204 301278
rect 299604 301276 300204 301278
rect 335604 301276 336204 301278
rect 371604 301276 372204 301278
rect 407604 301276 408204 301278
rect 443604 301276 444204 301278
rect 479604 301276 480204 301278
rect 515604 301276 516204 301278
rect 551604 301276 552204 301278
rect 590840 301276 591440 301278
rect -8436 301254 592360 301276
rect -8436 301018 -7334 301254
rect -7098 301018 11786 301254
rect 12022 301018 47786 301254
rect 48022 301018 83786 301254
rect 84022 301018 119786 301254
rect 120022 301018 155786 301254
rect 156022 301018 191786 301254
rect 192022 301018 227786 301254
rect 228022 301018 263786 301254
rect 264022 301018 299786 301254
rect 300022 301018 335786 301254
rect 336022 301018 371786 301254
rect 372022 301018 407786 301254
rect 408022 301018 443786 301254
rect 444022 301018 479786 301254
rect 480022 301018 515786 301254
rect 516022 301018 551786 301254
rect 552022 301018 591022 301254
rect 591258 301018 592360 301254
rect -8436 300934 592360 301018
rect -8436 300698 -7334 300934
rect -7098 300698 11786 300934
rect 12022 300698 47786 300934
rect 48022 300698 83786 300934
rect 84022 300698 119786 300934
rect 120022 300698 155786 300934
rect 156022 300698 191786 300934
rect 192022 300698 227786 300934
rect 228022 300698 263786 300934
rect 264022 300698 299786 300934
rect 300022 300698 335786 300934
rect 336022 300698 371786 300934
rect 372022 300698 407786 300934
rect 408022 300698 443786 300934
rect 444022 300698 479786 300934
rect 480022 300698 515786 300934
rect 516022 300698 551786 300934
rect 552022 300698 591022 300934
rect 591258 300698 592360 300934
rect -8436 300676 592360 300698
rect -7516 300674 -6916 300676
rect 11604 300674 12204 300676
rect 47604 300674 48204 300676
rect 83604 300674 84204 300676
rect 119604 300674 120204 300676
rect 155604 300674 156204 300676
rect 191604 300674 192204 300676
rect 227604 300674 228204 300676
rect 263604 300674 264204 300676
rect 299604 300674 300204 300676
rect 335604 300674 336204 300676
rect 371604 300674 372204 300676
rect 407604 300674 408204 300676
rect 443604 300674 444204 300676
rect 479604 300674 480204 300676
rect 515604 300674 516204 300676
rect 551604 300674 552204 300676
rect 590840 300674 591440 300676
rect -5676 297676 -5076 297678
rect 8004 297676 8604 297678
rect 44004 297676 44604 297678
rect 80004 297676 80604 297678
rect 116004 297676 116604 297678
rect 152004 297676 152604 297678
rect 188004 297676 188604 297678
rect 224004 297676 224604 297678
rect 260004 297676 260604 297678
rect 296004 297676 296604 297678
rect 332004 297676 332604 297678
rect 368004 297676 368604 297678
rect 404004 297676 404604 297678
rect 440004 297676 440604 297678
rect 476004 297676 476604 297678
rect 512004 297676 512604 297678
rect 548004 297676 548604 297678
rect 589000 297676 589600 297678
rect -6596 297654 590520 297676
rect -6596 297418 -5494 297654
rect -5258 297418 8186 297654
rect 8422 297418 44186 297654
rect 44422 297418 80186 297654
rect 80422 297418 116186 297654
rect 116422 297418 152186 297654
rect 152422 297418 188186 297654
rect 188422 297418 224186 297654
rect 224422 297418 260186 297654
rect 260422 297418 296186 297654
rect 296422 297418 332186 297654
rect 332422 297418 368186 297654
rect 368422 297418 404186 297654
rect 404422 297418 440186 297654
rect 440422 297418 476186 297654
rect 476422 297418 512186 297654
rect 512422 297418 548186 297654
rect 548422 297418 589182 297654
rect 589418 297418 590520 297654
rect -6596 297334 590520 297418
rect -6596 297098 -5494 297334
rect -5258 297098 8186 297334
rect 8422 297098 44186 297334
rect 44422 297098 80186 297334
rect 80422 297098 116186 297334
rect 116422 297098 152186 297334
rect 152422 297098 188186 297334
rect 188422 297098 224186 297334
rect 224422 297098 260186 297334
rect 260422 297098 296186 297334
rect 296422 297098 332186 297334
rect 332422 297098 368186 297334
rect 368422 297098 404186 297334
rect 404422 297098 440186 297334
rect 440422 297098 476186 297334
rect 476422 297098 512186 297334
rect 512422 297098 548186 297334
rect 548422 297098 589182 297334
rect 589418 297098 590520 297334
rect -6596 297076 590520 297098
rect -5676 297074 -5076 297076
rect 8004 297074 8604 297076
rect 44004 297074 44604 297076
rect 80004 297074 80604 297076
rect 116004 297074 116604 297076
rect 152004 297074 152604 297076
rect 188004 297074 188604 297076
rect 224004 297074 224604 297076
rect 260004 297074 260604 297076
rect 296004 297074 296604 297076
rect 332004 297074 332604 297076
rect 368004 297074 368604 297076
rect 404004 297074 404604 297076
rect 440004 297074 440604 297076
rect 476004 297074 476604 297076
rect 512004 297074 512604 297076
rect 548004 297074 548604 297076
rect 589000 297074 589600 297076
rect -3836 294076 -3236 294078
rect 4404 294076 5004 294078
rect 40404 294076 41004 294078
rect 76404 294076 77004 294078
rect 112404 294076 113004 294078
rect 148404 294076 149004 294078
rect 184404 294076 185004 294078
rect 220404 294076 221004 294078
rect 256404 294076 257004 294078
rect 292404 294076 293004 294078
rect 328404 294076 329004 294078
rect 364404 294076 365004 294078
rect 400404 294076 401004 294078
rect 436404 294076 437004 294078
rect 472404 294076 473004 294078
rect 508404 294076 509004 294078
rect 544404 294076 545004 294078
rect 580404 294076 581004 294078
rect 587160 294076 587760 294078
rect -4756 294054 588680 294076
rect -4756 293818 -3654 294054
rect -3418 293818 4586 294054
rect 4822 293818 40586 294054
rect 40822 293818 76586 294054
rect 76822 293818 112586 294054
rect 112822 293818 148586 294054
rect 148822 293818 184586 294054
rect 184822 293818 220586 294054
rect 220822 293818 256586 294054
rect 256822 293818 292586 294054
rect 292822 293818 328586 294054
rect 328822 293818 364586 294054
rect 364822 293818 400586 294054
rect 400822 293818 436586 294054
rect 436822 293818 472586 294054
rect 472822 293818 508586 294054
rect 508822 293818 544586 294054
rect 544822 293818 580586 294054
rect 580822 293818 587342 294054
rect 587578 293818 588680 294054
rect -4756 293734 588680 293818
rect -4756 293498 -3654 293734
rect -3418 293498 4586 293734
rect 4822 293498 40586 293734
rect 40822 293498 76586 293734
rect 76822 293498 112586 293734
rect 112822 293498 148586 293734
rect 148822 293498 184586 293734
rect 184822 293498 220586 293734
rect 220822 293498 256586 293734
rect 256822 293498 292586 293734
rect 292822 293498 328586 293734
rect 328822 293498 364586 293734
rect 364822 293498 400586 293734
rect 400822 293498 436586 293734
rect 436822 293498 472586 293734
rect 472822 293498 508586 293734
rect 508822 293498 544586 293734
rect 544822 293498 580586 293734
rect 580822 293498 587342 293734
rect 587578 293498 588680 293734
rect -4756 293476 588680 293498
rect -3836 293474 -3236 293476
rect 4404 293474 5004 293476
rect 40404 293474 41004 293476
rect 76404 293474 77004 293476
rect 112404 293474 113004 293476
rect 148404 293474 149004 293476
rect 184404 293474 185004 293476
rect 220404 293474 221004 293476
rect 256404 293474 257004 293476
rect 292404 293474 293004 293476
rect 328404 293474 329004 293476
rect 364404 293474 365004 293476
rect 400404 293474 401004 293476
rect 436404 293474 437004 293476
rect 472404 293474 473004 293476
rect 508404 293474 509004 293476
rect 544404 293474 545004 293476
rect 580404 293474 581004 293476
rect 587160 293474 587760 293476
rect -1996 290476 -1396 290478
rect 804 290476 1404 290478
rect 36804 290476 37404 290478
rect 72804 290476 73404 290478
rect 108804 290476 109404 290478
rect 144804 290476 145404 290478
rect 180804 290476 181404 290478
rect 216804 290476 217404 290478
rect 252804 290476 253404 290478
rect 288804 290476 289404 290478
rect 324804 290476 325404 290478
rect 360804 290476 361404 290478
rect 396804 290476 397404 290478
rect 432804 290476 433404 290478
rect 468804 290476 469404 290478
rect 504804 290476 505404 290478
rect 540804 290476 541404 290478
rect 576804 290476 577404 290478
rect 585320 290476 585920 290478
rect -2916 290454 586840 290476
rect -2916 290218 -1814 290454
rect -1578 290218 986 290454
rect 1222 290218 36986 290454
rect 37222 290218 72986 290454
rect 73222 290218 108986 290454
rect 109222 290218 144986 290454
rect 145222 290218 180986 290454
rect 181222 290218 216986 290454
rect 217222 290218 252986 290454
rect 253222 290218 288986 290454
rect 289222 290218 324986 290454
rect 325222 290218 360986 290454
rect 361222 290218 396986 290454
rect 397222 290218 432986 290454
rect 433222 290218 468986 290454
rect 469222 290218 504986 290454
rect 505222 290218 540986 290454
rect 541222 290218 576986 290454
rect 577222 290218 585502 290454
rect 585738 290218 586840 290454
rect -2916 290134 586840 290218
rect -2916 289898 -1814 290134
rect -1578 289898 986 290134
rect 1222 289898 36986 290134
rect 37222 289898 72986 290134
rect 73222 289898 108986 290134
rect 109222 289898 144986 290134
rect 145222 289898 180986 290134
rect 181222 289898 216986 290134
rect 217222 289898 252986 290134
rect 253222 289898 288986 290134
rect 289222 289898 324986 290134
rect 325222 289898 360986 290134
rect 361222 289898 396986 290134
rect 397222 289898 432986 290134
rect 433222 289898 468986 290134
rect 469222 289898 504986 290134
rect 505222 289898 540986 290134
rect 541222 289898 576986 290134
rect 577222 289898 585502 290134
rect 585738 289898 586840 290134
rect -2916 289876 586840 289898
rect -1996 289874 -1396 289876
rect 804 289874 1404 289876
rect 36804 289874 37404 289876
rect 72804 289874 73404 289876
rect 108804 289874 109404 289876
rect 144804 289874 145404 289876
rect 180804 289874 181404 289876
rect 216804 289874 217404 289876
rect 252804 289874 253404 289876
rect 288804 289874 289404 289876
rect 324804 289874 325404 289876
rect 360804 289874 361404 289876
rect 396804 289874 397404 289876
rect 432804 289874 433404 289876
rect 468804 289874 469404 289876
rect 504804 289874 505404 289876
rect 540804 289874 541404 289876
rect 576804 289874 577404 289876
rect 585320 289874 585920 289876
rect -8436 283276 -7836 283278
rect 29604 283276 30204 283278
rect 65604 283276 66204 283278
rect 101604 283276 102204 283278
rect 137604 283276 138204 283278
rect 173604 283276 174204 283278
rect 209604 283276 210204 283278
rect 245604 283276 246204 283278
rect 281604 283276 282204 283278
rect 317604 283276 318204 283278
rect 353604 283276 354204 283278
rect 389604 283276 390204 283278
rect 425604 283276 426204 283278
rect 461604 283276 462204 283278
rect 497604 283276 498204 283278
rect 533604 283276 534204 283278
rect 569604 283276 570204 283278
rect 591760 283276 592360 283278
rect -8436 283254 592360 283276
rect -8436 283018 -8254 283254
rect -8018 283018 29786 283254
rect 30022 283018 65786 283254
rect 66022 283018 101786 283254
rect 102022 283018 137786 283254
rect 138022 283018 173786 283254
rect 174022 283018 209786 283254
rect 210022 283018 245786 283254
rect 246022 283018 281786 283254
rect 282022 283018 317786 283254
rect 318022 283018 353786 283254
rect 354022 283018 389786 283254
rect 390022 283018 425786 283254
rect 426022 283018 461786 283254
rect 462022 283018 497786 283254
rect 498022 283018 533786 283254
rect 534022 283018 569786 283254
rect 570022 283018 591942 283254
rect 592178 283018 592360 283254
rect -8436 282934 592360 283018
rect -8436 282698 -8254 282934
rect -8018 282698 29786 282934
rect 30022 282698 65786 282934
rect 66022 282698 101786 282934
rect 102022 282698 137786 282934
rect 138022 282698 173786 282934
rect 174022 282698 209786 282934
rect 210022 282698 245786 282934
rect 246022 282698 281786 282934
rect 282022 282698 317786 282934
rect 318022 282698 353786 282934
rect 354022 282698 389786 282934
rect 390022 282698 425786 282934
rect 426022 282698 461786 282934
rect 462022 282698 497786 282934
rect 498022 282698 533786 282934
rect 534022 282698 569786 282934
rect 570022 282698 591942 282934
rect 592178 282698 592360 282934
rect -8436 282676 592360 282698
rect -8436 282674 -7836 282676
rect 29604 282674 30204 282676
rect 65604 282674 66204 282676
rect 101604 282674 102204 282676
rect 137604 282674 138204 282676
rect 173604 282674 174204 282676
rect 209604 282674 210204 282676
rect 245604 282674 246204 282676
rect 281604 282674 282204 282676
rect 317604 282674 318204 282676
rect 353604 282674 354204 282676
rect 389604 282674 390204 282676
rect 425604 282674 426204 282676
rect 461604 282674 462204 282676
rect 497604 282674 498204 282676
rect 533604 282674 534204 282676
rect 569604 282674 570204 282676
rect 591760 282674 592360 282676
rect -6596 279676 -5996 279678
rect 26004 279676 26604 279678
rect 62004 279676 62604 279678
rect 98004 279676 98604 279678
rect 134004 279676 134604 279678
rect 170004 279676 170604 279678
rect 206004 279676 206604 279678
rect 242004 279676 242604 279678
rect 278004 279676 278604 279678
rect 314004 279676 314604 279678
rect 350004 279676 350604 279678
rect 386004 279676 386604 279678
rect 422004 279676 422604 279678
rect 458004 279676 458604 279678
rect 494004 279676 494604 279678
rect 530004 279676 530604 279678
rect 566004 279676 566604 279678
rect 589920 279676 590520 279678
rect -6596 279654 590520 279676
rect -6596 279418 -6414 279654
rect -6178 279418 26186 279654
rect 26422 279418 62186 279654
rect 62422 279418 98186 279654
rect 98422 279418 134186 279654
rect 134422 279418 170186 279654
rect 170422 279418 206186 279654
rect 206422 279418 242186 279654
rect 242422 279418 278186 279654
rect 278422 279418 314186 279654
rect 314422 279418 350186 279654
rect 350422 279418 386186 279654
rect 386422 279418 422186 279654
rect 422422 279418 458186 279654
rect 458422 279418 494186 279654
rect 494422 279418 530186 279654
rect 530422 279418 566186 279654
rect 566422 279418 590102 279654
rect 590338 279418 590520 279654
rect -6596 279334 590520 279418
rect -6596 279098 -6414 279334
rect -6178 279098 26186 279334
rect 26422 279098 62186 279334
rect 62422 279098 98186 279334
rect 98422 279098 134186 279334
rect 134422 279098 170186 279334
rect 170422 279098 206186 279334
rect 206422 279098 242186 279334
rect 242422 279098 278186 279334
rect 278422 279098 314186 279334
rect 314422 279098 350186 279334
rect 350422 279098 386186 279334
rect 386422 279098 422186 279334
rect 422422 279098 458186 279334
rect 458422 279098 494186 279334
rect 494422 279098 530186 279334
rect 530422 279098 566186 279334
rect 566422 279098 590102 279334
rect 590338 279098 590520 279334
rect -6596 279076 590520 279098
rect -6596 279074 -5996 279076
rect 26004 279074 26604 279076
rect 62004 279074 62604 279076
rect 98004 279074 98604 279076
rect 134004 279074 134604 279076
rect 170004 279074 170604 279076
rect 206004 279074 206604 279076
rect 242004 279074 242604 279076
rect 278004 279074 278604 279076
rect 314004 279074 314604 279076
rect 350004 279074 350604 279076
rect 386004 279074 386604 279076
rect 422004 279074 422604 279076
rect 458004 279074 458604 279076
rect 494004 279074 494604 279076
rect 530004 279074 530604 279076
rect 566004 279074 566604 279076
rect 589920 279074 590520 279076
rect -4756 276076 -4156 276078
rect 22404 276076 23004 276078
rect 58404 276076 59004 276078
rect 94404 276076 95004 276078
rect 130404 276076 131004 276078
rect 166404 276076 167004 276078
rect 202404 276076 203004 276078
rect 238404 276076 239004 276078
rect 274404 276076 275004 276078
rect 310404 276076 311004 276078
rect 346404 276076 347004 276078
rect 382404 276076 383004 276078
rect 418404 276076 419004 276078
rect 454404 276076 455004 276078
rect 490404 276076 491004 276078
rect 526404 276076 527004 276078
rect 562404 276076 563004 276078
rect 588080 276076 588680 276078
rect -4756 276054 588680 276076
rect -4756 275818 -4574 276054
rect -4338 275818 22586 276054
rect 22822 275818 58586 276054
rect 58822 275818 94586 276054
rect 94822 275818 130586 276054
rect 130822 275818 166586 276054
rect 166822 275818 202586 276054
rect 202822 275818 238586 276054
rect 238822 275818 274586 276054
rect 274822 275818 310586 276054
rect 310822 275818 346586 276054
rect 346822 275818 382586 276054
rect 382822 275818 418586 276054
rect 418822 275818 454586 276054
rect 454822 275818 490586 276054
rect 490822 275818 526586 276054
rect 526822 275818 562586 276054
rect 562822 275818 588262 276054
rect 588498 275818 588680 276054
rect -4756 275734 588680 275818
rect -4756 275498 -4574 275734
rect -4338 275498 22586 275734
rect 22822 275498 58586 275734
rect 58822 275498 94586 275734
rect 94822 275498 130586 275734
rect 130822 275498 166586 275734
rect 166822 275498 202586 275734
rect 202822 275498 238586 275734
rect 238822 275498 274586 275734
rect 274822 275498 310586 275734
rect 310822 275498 346586 275734
rect 346822 275498 382586 275734
rect 382822 275498 418586 275734
rect 418822 275498 454586 275734
rect 454822 275498 490586 275734
rect 490822 275498 526586 275734
rect 526822 275498 562586 275734
rect 562822 275498 588262 275734
rect 588498 275498 588680 275734
rect -4756 275476 588680 275498
rect -4756 275474 -4156 275476
rect 22404 275474 23004 275476
rect 58404 275474 59004 275476
rect 94404 275474 95004 275476
rect 130404 275474 131004 275476
rect 166404 275474 167004 275476
rect 202404 275474 203004 275476
rect 238404 275474 239004 275476
rect 274404 275474 275004 275476
rect 310404 275474 311004 275476
rect 346404 275474 347004 275476
rect 382404 275474 383004 275476
rect 418404 275474 419004 275476
rect 454404 275474 455004 275476
rect 490404 275474 491004 275476
rect 526404 275474 527004 275476
rect 562404 275474 563004 275476
rect 588080 275474 588680 275476
rect -2916 272476 -2316 272478
rect 18804 272476 19404 272478
rect 54804 272476 55404 272478
rect 90804 272476 91404 272478
rect 126804 272476 127404 272478
rect 162804 272476 163404 272478
rect 198804 272476 199404 272478
rect 234804 272476 235404 272478
rect 270804 272476 271404 272478
rect 306804 272476 307404 272478
rect 342804 272476 343404 272478
rect 378804 272476 379404 272478
rect 414804 272476 415404 272478
rect 450804 272476 451404 272478
rect 486804 272476 487404 272478
rect 522804 272476 523404 272478
rect 558804 272476 559404 272478
rect 586240 272476 586840 272478
rect -2916 272454 586840 272476
rect -2916 272218 -2734 272454
rect -2498 272218 18986 272454
rect 19222 272218 54986 272454
rect 55222 272218 90986 272454
rect 91222 272218 126986 272454
rect 127222 272218 162986 272454
rect 163222 272218 198986 272454
rect 199222 272218 234986 272454
rect 235222 272218 270986 272454
rect 271222 272218 306986 272454
rect 307222 272218 342986 272454
rect 343222 272218 378986 272454
rect 379222 272218 414986 272454
rect 415222 272218 450986 272454
rect 451222 272218 486986 272454
rect 487222 272218 522986 272454
rect 523222 272218 558986 272454
rect 559222 272218 586422 272454
rect 586658 272218 586840 272454
rect -2916 272134 586840 272218
rect -2916 271898 -2734 272134
rect -2498 271898 18986 272134
rect 19222 271898 54986 272134
rect 55222 271898 90986 272134
rect 91222 271898 126986 272134
rect 127222 271898 162986 272134
rect 163222 271898 198986 272134
rect 199222 271898 234986 272134
rect 235222 271898 270986 272134
rect 271222 271898 306986 272134
rect 307222 271898 342986 272134
rect 343222 271898 378986 272134
rect 379222 271898 414986 272134
rect 415222 271898 450986 272134
rect 451222 271898 486986 272134
rect 487222 271898 522986 272134
rect 523222 271898 558986 272134
rect 559222 271898 586422 272134
rect 586658 271898 586840 272134
rect -2916 271876 586840 271898
rect -2916 271874 -2316 271876
rect 18804 271874 19404 271876
rect 54804 271874 55404 271876
rect 90804 271874 91404 271876
rect 126804 271874 127404 271876
rect 162804 271874 163404 271876
rect 198804 271874 199404 271876
rect 234804 271874 235404 271876
rect 270804 271874 271404 271876
rect 306804 271874 307404 271876
rect 342804 271874 343404 271876
rect 378804 271874 379404 271876
rect 414804 271874 415404 271876
rect 450804 271874 451404 271876
rect 486804 271874 487404 271876
rect 522804 271874 523404 271876
rect 558804 271874 559404 271876
rect 586240 271874 586840 271876
rect -7516 265276 -6916 265278
rect 11604 265276 12204 265278
rect 47604 265276 48204 265278
rect 83604 265276 84204 265278
rect 119604 265276 120204 265278
rect 155604 265276 156204 265278
rect 191604 265276 192204 265278
rect 227604 265276 228204 265278
rect 263604 265276 264204 265278
rect 299604 265276 300204 265278
rect 335604 265276 336204 265278
rect 371604 265276 372204 265278
rect 407604 265276 408204 265278
rect 443604 265276 444204 265278
rect 479604 265276 480204 265278
rect 515604 265276 516204 265278
rect 551604 265276 552204 265278
rect 590840 265276 591440 265278
rect -8436 265254 592360 265276
rect -8436 265018 -7334 265254
rect -7098 265018 11786 265254
rect 12022 265018 47786 265254
rect 48022 265018 83786 265254
rect 84022 265018 119786 265254
rect 120022 265018 155786 265254
rect 156022 265018 191786 265254
rect 192022 265018 227786 265254
rect 228022 265018 263786 265254
rect 264022 265018 299786 265254
rect 300022 265018 335786 265254
rect 336022 265018 371786 265254
rect 372022 265018 407786 265254
rect 408022 265018 443786 265254
rect 444022 265018 479786 265254
rect 480022 265018 515786 265254
rect 516022 265018 551786 265254
rect 552022 265018 591022 265254
rect 591258 265018 592360 265254
rect -8436 264934 592360 265018
rect -8436 264698 -7334 264934
rect -7098 264698 11786 264934
rect 12022 264698 47786 264934
rect 48022 264698 83786 264934
rect 84022 264698 119786 264934
rect 120022 264698 155786 264934
rect 156022 264698 191786 264934
rect 192022 264698 227786 264934
rect 228022 264698 263786 264934
rect 264022 264698 299786 264934
rect 300022 264698 335786 264934
rect 336022 264698 371786 264934
rect 372022 264698 407786 264934
rect 408022 264698 443786 264934
rect 444022 264698 479786 264934
rect 480022 264698 515786 264934
rect 516022 264698 551786 264934
rect 552022 264698 591022 264934
rect 591258 264698 592360 264934
rect -8436 264676 592360 264698
rect -7516 264674 -6916 264676
rect 11604 264674 12204 264676
rect 47604 264674 48204 264676
rect 83604 264674 84204 264676
rect 119604 264674 120204 264676
rect 155604 264674 156204 264676
rect 191604 264674 192204 264676
rect 227604 264674 228204 264676
rect 263604 264674 264204 264676
rect 299604 264674 300204 264676
rect 335604 264674 336204 264676
rect 371604 264674 372204 264676
rect 407604 264674 408204 264676
rect 443604 264674 444204 264676
rect 479604 264674 480204 264676
rect 515604 264674 516204 264676
rect 551604 264674 552204 264676
rect 590840 264674 591440 264676
rect -5676 261676 -5076 261678
rect 8004 261676 8604 261678
rect 44004 261676 44604 261678
rect 80004 261676 80604 261678
rect 116004 261676 116604 261678
rect 152004 261676 152604 261678
rect 188004 261676 188604 261678
rect 224004 261676 224604 261678
rect 260004 261676 260604 261678
rect 296004 261676 296604 261678
rect 332004 261676 332604 261678
rect 368004 261676 368604 261678
rect 404004 261676 404604 261678
rect 440004 261676 440604 261678
rect 476004 261676 476604 261678
rect 512004 261676 512604 261678
rect 548004 261676 548604 261678
rect 589000 261676 589600 261678
rect -6596 261654 590520 261676
rect -6596 261418 -5494 261654
rect -5258 261418 8186 261654
rect 8422 261418 44186 261654
rect 44422 261418 80186 261654
rect 80422 261418 116186 261654
rect 116422 261418 152186 261654
rect 152422 261418 188186 261654
rect 188422 261418 224186 261654
rect 224422 261418 260186 261654
rect 260422 261418 296186 261654
rect 296422 261418 332186 261654
rect 332422 261418 368186 261654
rect 368422 261418 404186 261654
rect 404422 261418 440186 261654
rect 440422 261418 476186 261654
rect 476422 261418 512186 261654
rect 512422 261418 548186 261654
rect 548422 261418 589182 261654
rect 589418 261418 590520 261654
rect -6596 261334 590520 261418
rect -6596 261098 -5494 261334
rect -5258 261098 8186 261334
rect 8422 261098 44186 261334
rect 44422 261098 80186 261334
rect 80422 261098 116186 261334
rect 116422 261098 152186 261334
rect 152422 261098 188186 261334
rect 188422 261098 224186 261334
rect 224422 261098 260186 261334
rect 260422 261098 296186 261334
rect 296422 261098 332186 261334
rect 332422 261098 368186 261334
rect 368422 261098 404186 261334
rect 404422 261098 440186 261334
rect 440422 261098 476186 261334
rect 476422 261098 512186 261334
rect 512422 261098 548186 261334
rect 548422 261098 589182 261334
rect 589418 261098 590520 261334
rect -6596 261076 590520 261098
rect -5676 261074 -5076 261076
rect 8004 261074 8604 261076
rect 44004 261074 44604 261076
rect 80004 261074 80604 261076
rect 116004 261074 116604 261076
rect 152004 261074 152604 261076
rect 188004 261074 188604 261076
rect 224004 261074 224604 261076
rect 260004 261074 260604 261076
rect 296004 261074 296604 261076
rect 332004 261074 332604 261076
rect 368004 261074 368604 261076
rect 404004 261074 404604 261076
rect 440004 261074 440604 261076
rect 476004 261074 476604 261076
rect 512004 261074 512604 261076
rect 548004 261074 548604 261076
rect 589000 261074 589600 261076
rect -3836 258076 -3236 258078
rect 4404 258076 5004 258078
rect 40404 258076 41004 258078
rect 76404 258076 77004 258078
rect 112404 258076 113004 258078
rect 148404 258076 149004 258078
rect 184404 258076 185004 258078
rect 220404 258076 221004 258078
rect 256404 258076 257004 258078
rect 292404 258076 293004 258078
rect 328404 258076 329004 258078
rect 364404 258076 365004 258078
rect 400404 258076 401004 258078
rect 436404 258076 437004 258078
rect 472404 258076 473004 258078
rect 508404 258076 509004 258078
rect 544404 258076 545004 258078
rect 580404 258076 581004 258078
rect 587160 258076 587760 258078
rect -4756 258054 588680 258076
rect -4756 257818 -3654 258054
rect -3418 257818 4586 258054
rect 4822 257818 40586 258054
rect 40822 257818 76586 258054
rect 76822 257818 112586 258054
rect 112822 257818 148586 258054
rect 148822 257818 184586 258054
rect 184822 257818 220586 258054
rect 220822 257818 256586 258054
rect 256822 257818 292586 258054
rect 292822 257818 328586 258054
rect 328822 257818 364586 258054
rect 364822 257818 400586 258054
rect 400822 257818 436586 258054
rect 436822 257818 472586 258054
rect 472822 257818 508586 258054
rect 508822 257818 544586 258054
rect 544822 257818 580586 258054
rect 580822 257818 587342 258054
rect 587578 257818 588680 258054
rect -4756 257734 588680 257818
rect -4756 257498 -3654 257734
rect -3418 257498 4586 257734
rect 4822 257498 40586 257734
rect 40822 257498 76586 257734
rect 76822 257498 112586 257734
rect 112822 257498 148586 257734
rect 148822 257498 184586 257734
rect 184822 257498 220586 257734
rect 220822 257498 256586 257734
rect 256822 257498 292586 257734
rect 292822 257498 328586 257734
rect 328822 257498 364586 257734
rect 364822 257498 400586 257734
rect 400822 257498 436586 257734
rect 436822 257498 472586 257734
rect 472822 257498 508586 257734
rect 508822 257498 544586 257734
rect 544822 257498 580586 257734
rect 580822 257498 587342 257734
rect 587578 257498 588680 257734
rect -4756 257476 588680 257498
rect -3836 257474 -3236 257476
rect 4404 257474 5004 257476
rect 40404 257474 41004 257476
rect 76404 257474 77004 257476
rect 112404 257474 113004 257476
rect 148404 257474 149004 257476
rect 184404 257474 185004 257476
rect 220404 257474 221004 257476
rect 256404 257474 257004 257476
rect 292404 257474 293004 257476
rect 328404 257474 329004 257476
rect 364404 257474 365004 257476
rect 400404 257474 401004 257476
rect 436404 257474 437004 257476
rect 472404 257474 473004 257476
rect 508404 257474 509004 257476
rect 544404 257474 545004 257476
rect 580404 257474 581004 257476
rect 587160 257474 587760 257476
rect -1996 254476 -1396 254478
rect 804 254476 1404 254478
rect 36804 254476 37404 254478
rect 72804 254476 73404 254478
rect 108804 254476 109404 254478
rect 144804 254476 145404 254478
rect 180804 254476 181404 254478
rect 216804 254476 217404 254478
rect 252804 254476 253404 254478
rect 288804 254476 289404 254478
rect 324804 254476 325404 254478
rect 360804 254476 361404 254478
rect 396804 254476 397404 254478
rect 432804 254476 433404 254478
rect 468804 254476 469404 254478
rect 504804 254476 505404 254478
rect 540804 254476 541404 254478
rect 576804 254476 577404 254478
rect 585320 254476 585920 254478
rect -2916 254454 586840 254476
rect -2916 254218 -1814 254454
rect -1578 254218 986 254454
rect 1222 254218 36986 254454
rect 37222 254218 72986 254454
rect 73222 254218 108986 254454
rect 109222 254218 144986 254454
rect 145222 254218 180986 254454
rect 181222 254218 216986 254454
rect 217222 254218 252986 254454
rect 253222 254218 288986 254454
rect 289222 254218 324986 254454
rect 325222 254218 360986 254454
rect 361222 254218 396986 254454
rect 397222 254218 432986 254454
rect 433222 254218 468986 254454
rect 469222 254218 504986 254454
rect 505222 254218 540986 254454
rect 541222 254218 576986 254454
rect 577222 254218 585502 254454
rect 585738 254218 586840 254454
rect -2916 254134 586840 254218
rect -2916 253898 -1814 254134
rect -1578 253898 986 254134
rect 1222 253898 36986 254134
rect 37222 253898 72986 254134
rect 73222 253898 108986 254134
rect 109222 253898 144986 254134
rect 145222 253898 180986 254134
rect 181222 253898 216986 254134
rect 217222 253898 252986 254134
rect 253222 253898 288986 254134
rect 289222 253898 324986 254134
rect 325222 253898 360986 254134
rect 361222 253898 396986 254134
rect 397222 253898 432986 254134
rect 433222 253898 468986 254134
rect 469222 253898 504986 254134
rect 505222 253898 540986 254134
rect 541222 253898 576986 254134
rect 577222 253898 585502 254134
rect 585738 253898 586840 254134
rect -2916 253876 586840 253898
rect -1996 253874 -1396 253876
rect 804 253874 1404 253876
rect 36804 253874 37404 253876
rect 72804 253874 73404 253876
rect 108804 253874 109404 253876
rect 144804 253874 145404 253876
rect 180804 253874 181404 253876
rect 216804 253874 217404 253876
rect 252804 253874 253404 253876
rect 288804 253874 289404 253876
rect 324804 253874 325404 253876
rect 360804 253874 361404 253876
rect 396804 253874 397404 253876
rect 432804 253874 433404 253876
rect 468804 253874 469404 253876
rect 504804 253874 505404 253876
rect 540804 253874 541404 253876
rect 576804 253874 577404 253876
rect 585320 253874 585920 253876
rect -8436 247276 -7836 247278
rect 29604 247276 30204 247278
rect 65604 247276 66204 247278
rect 101604 247276 102204 247278
rect 137604 247276 138204 247278
rect 173604 247276 174204 247278
rect 209604 247276 210204 247278
rect 245604 247276 246204 247278
rect 281604 247276 282204 247278
rect 317604 247276 318204 247278
rect 353604 247276 354204 247278
rect 389604 247276 390204 247278
rect 425604 247276 426204 247278
rect 461604 247276 462204 247278
rect 497604 247276 498204 247278
rect 533604 247276 534204 247278
rect 569604 247276 570204 247278
rect 591760 247276 592360 247278
rect -8436 247254 592360 247276
rect -8436 247018 -8254 247254
rect -8018 247018 29786 247254
rect 30022 247018 65786 247254
rect 66022 247018 101786 247254
rect 102022 247018 137786 247254
rect 138022 247018 173786 247254
rect 174022 247018 209786 247254
rect 210022 247018 245786 247254
rect 246022 247018 281786 247254
rect 282022 247018 317786 247254
rect 318022 247018 353786 247254
rect 354022 247018 389786 247254
rect 390022 247018 425786 247254
rect 426022 247018 461786 247254
rect 462022 247018 497786 247254
rect 498022 247018 533786 247254
rect 534022 247018 569786 247254
rect 570022 247018 591942 247254
rect 592178 247018 592360 247254
rect -8436 246934 592360 247018
rect -8436 246698 -8254 246934
rect -8018 246698 29786 246934
rect 30022 246698 65786 246934
rect 66022 246698 101786 246934
rect 102022 246698 137786 246934
rect 138022 246698 173786 246934
rect 174022 246698 209786 246934
rect 210022 246698 245786 246934
rect 246022 246698 281786 246934
rect 282022 246698 317786 246934
rect 318022 246698 353786 246934
rect 354022 246698 389786 246934
rect 390022 246698 425786 246934
rect 426022 246698 461786 246934
rect 462022 246698 497786 246934
rect 498022 246698 533786 246934
rect 534022 246698 569786 246934
rect 570022 246698 591942 246934
rect 592178 246698 592360 246934
rect -8436 246676 592360 246698
rect -8436 246674 -7836 246676
rect 29604 246674 30204 246676
rect 65604 246674 66204 246676
rect 101604 246674 102204 246676
rect 137604 246674 138204 246676
rect 173604 246674 174204 246676
rect 209604 246674 210204 246676
rect 245604 246674 246204 246676
rect 281604 246674 282204 246676
rect 317604 246674 318204 246676
rect 353604 246674 354204 246676
rect 389604 246674 390204 246676
rect 425604 246674 426204 246676
rect 461604 246674 462204 246676
rect 497604 246674 498204 246676
rect 533604 246674 534204 246676
rect 569604 246674 570204 246676
rect 591760 246674 592360 246676
rect -6596 243676 -5996 243678
rect 26004 243676 26604 243678
rect 62004 243676 62604 243678
rect 98004 243676 98604 243678
rect 134004 243676 134604 243678
rect 170004 243676 170604 243678
rect 206004 243676 206604 243678
rect 242004 243676 242604 243678
rect 278004 243676 278604 243678
rect 314004 243676 314604 243678
rect 350004 243676 350604 243678
rect 386004 243676 386604 243678
rect 422004 243676 422604 243678
rect 458004 243676 458604 243678
rect 494004 243676 494604 243678
rect 530004 243676 530604 243678
rect 566004 243676 566604 243678
rect 589920 243676 590520 243678
rect -6596 243654 590520 243676
rect -6596 243418 -6414 243654
rect -6178 243418 26186 243654
rect 26422 243418 62186 243654
rect 62422 243418 98186 243654
rect 98422 243418 134186 243654
rect 134422 243418 170186 243654
rect 170422 243418 206186 243654
rect 206422 243418 242186 243654
rect 242422 243418 278186 243654
rect 278422 243418 314186 243654
rect 314422 243418 350186 243654
rect 350422 243418 386186 243654
rect 386422 243418 422186 243654
rect 422422 243418 458186 243654
rect 458422 243418 494186 243654
rect 494422 243418 530186 243654
rect 530422 243418 566186 243654
rect 566422 243418 590102 243654
rect 590338 243418 590520 243654
rect -6596 243334 590520 243418
rect -6596 243098 -6414 243334
rect -6178 243098 26186 243334
rect 26422 243098 62186 243334
rect 62422 243098 98186 243334
rect 98422 243098 134186 243334
rect 134422 243098 170186 243334
rect 170422 243098 206186 243334
rect 206422 243098 242186 243334
rect 242422 243098 278186 243334
rect 278422 243098 314186 243334
rect 314422 243098 350186 243334
rect 350422 243098 386186 243334
rect 386422 243098 422186 243334
rect 422422 243098 458186 243334
rect 458422 243098 494186 243334
rect 494422 243098 530186 243334
rect 530422 243098 566186 243334
rect 566422 243098 590102 243334
rect 590338 243098 590520 243334
rect -6596 243076 590520 243098
rect -6596 243074 -5996 243076
rect 26004 243074 26604 243076
rect 62004 243074 62604 243076
rect 98004 243074 98604 243076
rect 134004 243074 134604 243076
rect 170004 243074 170604 243076
rect 206004 243074 206604 243076
rect 242004 243074 242604 243076
rect 278004 243074 278604 243076
rect 314004 243074 314604 243076
rect 350004 243074 350604 243076
rect 386004 243074 386604 243076
rect 422004 243074 422604 243076
rect 458004 243074 458604 243076
rect 494004 243074 494604 243076
rect 530004 243074 530604 243076
rect 566004 243074 566604 243076
rect 589920 243074 590520 243076
rect -4756 240076 -4156 240078
rect 22404 240076 23004 240078
rect 58404 240076 59004 240078
rect 94404 240076 95004 240078
rect 130404 240076 131004 240078
rect 166404 240076 167004 240078
rect 202404 240076 203004 240078
rect 238404 240076 239004 240078
rect 274404 240076 275004 240078
rect 310404 240076 311004 240078
rect 346404 240076 347004 240078
rect 382404 240076 383004 240078
rect 418404 240076 419004 240078
rect 454404 240076 455004 240078
rect 490404 240076 491004 240078
rect 526404 240076 527004 240078
rect 562404 240076 563004 240078
rect 588080 240076 588680 240078
rect -4756 240054 588680 240076
rect -4756 239818 -4574 240054
rect -4338 239818 22586 240054
rect 22822 239818 58586 240054
rect 58822 239818 94586 240054
rect 94822 239818 130586 240054
rect 130822 239818 166586 240054
rect 166822 239818 202586 240054
rect 202822 239818 238586 240054
rect 238822 239818 274586 240054
rect 274822 239818 310586 240054
rect 310822 239818 346586 240054
rect 346822 239818 382586 240054
rect 382822 239818 418586 240054
rect 418822 239818 454586 240054
rect 454822 239818 490586 240054
rect 490822 239818 526586 240054
rect 526822 239818 562586 240054
rect 562822 239818 588262 240054
rect 588498 239818 588680 240054
rect -4756 239734 588680 239818
rect -4756 239498 -4574 239734
rect -4338 239498 22586 239734
rect 22822 239498 58586 239734
rect 58822 239498 94586 239734
rect 94822 239498 130586 239734
rect 130822 239498 166586 239734
rect 166822 239498 202586 239734
rect 202822 239498 238586 239734
rect 238822 239498 274586 239734
rect 274822 239498 310586 239734
rect 310822 239498 346586 239734
rect 346822 239498 382586 239734
rect 382822 239498 418586 239734
rect 418822 239498 454586 239734
rect 454822 239498 490586 239734
rect 490822 239498 526586 239734
rect 526822 239498 562586 239734
rect 562822 239498 588262 239734
rect 588498 239498 588680 239734
rect -4756 239476 588680 239498
rect -4756 239474 -4156 239476
rect 22404 239474 23004 239476
rect 58404 239474 59004 239476
rect 94404 239474 95004 239476
rect 130404 239474 131004 239476
rect 166404 239474 167004 239476
rect 202404 239474 203004 239476
rect 238404 239474 239004 239476
rect 274404 239474 275004 239476
rect 310404 239474 311004 239476
rect 346404 239474 347004 239476
rect 382404 239474 383004 239476
rect 418404 239474 419004 239476
rect 454404 239474 455004 239476
rect 490404 239474 491004 239476
rect 526404 239474 527004 239476
rect 562404 239474 563004 239476
rect 588080 239474 588680 239476
rect -2916 236476 -2316 236478
rect 18804 236476 19404 236478
rect 54804 236476 55404 236478
rect 90804 236476 91404 236478
rect 126804 236476 127404 236478
rect 162804 236476 163404 236478
rect 198804 236476 199404 236478
rect 234804 236476 235404 236478
rect 270804 236476 271404 236478
rect 306804 236476 307404 236478
rect 342804 236476 343404 236478
rect 378804 236476 379404 236478
rect 414804 236476 415404 236478
rect 450804 236476 451404 236478
rect 486804 236476 487404 236478
rect 522804 236476 523404 236478
rect 558804 236476 559404 236478
rect 586240 236476 586840 236478
rect -2916 236454 586840 236476
rect -2916 236218 -2734 236454
rect -2498 236218 18986 236454
rect 19222 236218 54986 236454
rect 55222 236218 90986 236454
rect 91222 236218 126986 236454
rect 127222 236218 162986 236454
rect 163222 236218 198986 236454
rect 199222 236218 234986 236454
rect 235222 236218 270986 236454
rect 271222 236218 306986 236454
rect 307222 236218 342986 236454
rect 343222 236218 378986 236454
rect 379222 236218 414986 236454
rect 415222 236218 450986 236454
rect 451222 236218 486986 236454
rect 487222 236218 522986 236454
rect 523222 236218 558986 236454
rect 559222 236218 586422 236454
rect 586658 236218 586840 236454
rect -2916 236134 586840 236218
rect -2916 235898 -2734 236134
rect -2498 235898 18986 236134
rect 19222 235898 54986 236134
rect 55222 235898 90986 236134
rect 91222 235898 126986 236134
rect 127222 235898 162986 236134
rect 163222 235898 198986 236134
rect 199222 235898 234986 236134
rect 235222 235898 270986 236134
rect 271222 235898 306986 236134
rect 307222 235898 342986 236134
rect 343222 235898 378986 236134
rect 379222 235898 414986 236134
rect 415222 235898 450986 236134
rect 451222 235898 486986 236134
rect 487222 235898 522986 236134
rect 523222 235898 558986 236134
rect 559222 235898 586422 236134
rect 586658 235898 586840 236134
rect -2916 235876 586840 235898
rect -2916 235874 -2316 235876
rect 18804 235874 19404 235876
rect 54804 235874 55404 235876
rect 90804 235874 91404 235876
rect 126804 235874 127404 235876
rect 162804 235874 163404 235876
rect 198804 235874 199404 235876
rect 234804 235874 235404 235876
rect 270804 235874 271404 235876
rect 306804 235874 307404 235876
rect 342804 235874 343404 235876
rect 378804 235874 379404 235876
rect 414804 235874 415404 235876
rect 450804 235874 451404 235876
rect 486804 235874 487404 235876
rect 522804 235874 523404 235876
rect 558804 235874 559404 235876
rect 586240 235874 586840 235876
rect -7516 229276 -6916 229278
rect 11604 229276 12204 229278
rect 47604 229276 48204 229278
rect 83604 229276 84204 229278
rect 119604 229276 120204 229278
rect 155604 229276 156204 229278
rect 191604 229276 192204 229278
rect 227604 229276 228204 229278
rect 263604 229276 264204 229278
rect 299604 229276 300204 229278
rect 335604 229276 336204 229278
rect 371604 229276 372204 229278
rect 407604 229276 408204 229278
rect 443604 229276 444204 229278
rect 479604 229276 480204 229278
rect 515604 229276 516204 229278
rect 551604 229276 552204 229278
rect 590840 229276 591440 229278
rect -8436 229254 592360 229276
rect -8436 229018 -7334 229254
rect -7098 229018 11786 229254
rect 12022 229018 47786 229254
rect 48022 229018 83786 229254
rect 84022 229018 119786 229254
rect 120022 229018 155786 229254
rect 156022 229018 191786 229254
rect 192022 229018 227786 229254
rect 228022 229018 263786 229254
rect 264022 229018 299786 229254
rect 300022 229018 335786 229254
rect 336022 229018 371786 229254
rect 372022 229018 407786 229254
rect 408022 229018 443786 229254
rect 444022 229018 479786 229254
rect 480022 229018 515786 229254
rect 516022 229018 551786 229254
rect 552022 229018 591022 229254
rect 591258 229018 592360 229254
rect -8436 228934 592360 229018
rect -8436 228698 -7334 228934
rect -7098 228698 11786 228934
rect 12022 228698 47786 228934
rect 48022 228698 83786 228934
rect 84022 228698 119786 228934
rect 120022 228698 155786 228934
rect 156022 228698 191786 228934
rect 192022 228698 227786 228934
rect 228022 228698 263786 228934
rect 264022 228698 299786 228934
rect 300022 228698 335786 228934
rect 336022 228698 371786 228934
rect 372022 228698 407786 228934
rect 408022 228698 443786 228934
rect 444022 228698 479786 228934
rect 480022 228698 515786 228934
rect 516022 228698 551786 228934
rect 552022 228698 591022 228934
rect 591258 228698 592360 228934
rect -8436 228676 592360 228698
rect -7516 228674 -6916 228676
rect 11604 228674 12204 228676
rect 47604 228674 48204 228676
rect 83604 228674 84204 228676
rect 119604 228674 120204 228676
rect 155604 228674 156204 228676
rect 191604 228674 192204 228676
rect 227604 228674 228204 228676
rect 263604 228674 264204 228676
rect 299604 228674 300204 228676
rect 335604 228674 336204 228676
rect 371604 228674 372204 228676
rect 407604 228674 408204 228676
rect 443604 228674 444204 228676
rect 479604 228674 480204 228676
rect 515604 228674 516204 228676
rect 551604 228674 552204 228676
rect 590840 228674 591440 228676
rect -5676 225676 -5076 225678
rect 8004 225676 8604 225678
rect 44004 225676 44604 225678
rect 80004 225676 80604 225678
rect 116004 225676 116604 225678
rect 152004 225676 152604 225678
rect 188004 225676 188604 225678
rect 224004 225676 224604 225678
rect 260004 225676 260604 225678
rect 296004 225676 296604 225678
rect 332004 225676 332604 225678
rect 368004 225676 368604 225678
rect 404004 225676 404604 225678
rect 440004 225676 440604 225678
rect 476004 225676 476604 225678
rect 512004 225676 512604 225678
rect 548004 225676 548604 225678
rect 589000 225676 589600 225678
rect -6596 225654 590520 225676
rect -6596 225418 -5494 225654
rect -5258 225418 8186 225654
rect 8422 225418 44186 225654
rect 44422 225418 80186 225654
rect 80422 225418 116186 225654
rect 116422 225418 152186 225654
rect 152422 225418 188186 225654
rect 188422 225418 224186 225654
rect 224422 225418 260186 225654
rect 260422 225418 296186 225654
rect 296422 225418 332186 225654
rect 332422 225418 368186 225654
rect 368422 225418 404186 225654
rect 404422 225418 440186 225654
rect 440422 225418 476186 225654
rect 476422 225418 512186 225654
rect 512422 225418 548186 225654
rect 548422 225418 589182 225654
rect 589418 225418 590520 225654
rect -6596 225334 590520 225418
rect -6596 225098 -5494 225334
rect -5258 225098 8186 225334
rect 8422 225098 44186 225334
rect 44422 225098 80186 225334
rect 80422 225098 116186 225334
rect 116422 225098 152186 225334
rect 152422 225098 188186 225334
rect 188422 225098 224186 225334
rect 224422 225098 260186 225334
rect 260422 225098 296186 225334
rect 296422 225098 332186 225334
rect 332422 225098 368186 225334
rect 368422 225098 404186 225334
rect 404422 225098 440186 225334
rect 440422 225098 476186 225334
rect 476422 225098 512186 225334
rect 512422 225098 548186 225334
rect 548422 225098 589182 225334
rect 589418 225098 590520 225334
rect -6596 225076 590520 225098
rect -5676 225074 -5076 225076
rect 8004 225074 8604 225076
rect 44004 225074 44604 225076
rect 80004 225074 80604 225076
rect 116004 225074 116604 225076
rect 152004 225074 152604 225076
rect 188004 225074 188604 225076
rect 224004 225074 224604 225076
rect 260004 225074 260604 225076
rect 296004 225074 296604 225076
rect 332004 225074 332604 225076
rect 368004 225074 368604 225076
rect 404004 225074 404604 225076
rect 440004 225074 440604 225076
rect 476004 225074 476604 225076
rect 512004 225074 512604 225076
rect 548004 225074 548604 225076
rect 589000 225074 589600 225076
rect -3836 222076 -3236 222078
rect 4404 222076 5004 222078
rect 40404 222076 41004 222078
rect 76404 222076 77004 222078
rect 112404 222076 113004 222078
rect 148404 222076 149004 222078
rect 184404 222076 185004 222078
rect 220404 222076 221004 222078
rect 256404 222076 257004 222078
rect 292404 222076 293004 222078
rect 328404 222076 329004 222078
rect 364404 222076 365004 222078
rect 400404 222076 401004 222078
rect 436404 222076 437004 222078
rect 472404 222076 473004 222078
rect 508404 222076 509004 222078
rect 544404 222076 545004 222078
rect 580404 222076 581004 222078
rect 587160 222076 587760 222078
rect -4756 222054 588680 222076
rect -4756 221818 -3654 222054
rect -3418 221818 4586 222054
rect 4822 221818 40586 222054
rect 40822 221818 76586 222054
rect 76822 221818 112586 222054
rect 112822 221818 148586 222054
rect 148822 221818 184586 222054
rect 184822 221818 220586 222054
rect 220822 221818 256586 222054
rect 256822 221818 292586 222054
rect 292822 221818 328586 222054
rect 328822 221818 364586 222054
rect 364822 221818 400586 222054
rect 400822 221818 436586 222054
rect 436822 221818 472586 222054
rect 472822 221818 508586 222054
rect 508822 221818 544586 222054
rect 544822 221818 580586 222054
rect 580822 221818 587342 222054
rect 587578 221818 588680 222054
rect -4756 221734 588680 221818
rect -4756 221498 -3654 221734
rect -3418 221498 4586 221734
rect 4822 221498 40586 221734
rect 40822 221498 76586 221734
rect 76822 221498 112586 221734
rect 112822 221498 148586 221734
rect 148822 221498 184586 221734
rect 184822 221498 220586 221734
rect 220822 221498 256586 221734
rect 256822 221498 292586 221734
rect 292822 221498 328586 221734
rect 328822 221498 364586 221734
rect 364822 221498 400586 221734
rect 400822 221498 436586 221734
rect 436822 221498 472586 221734
rect 472822 221498 508586 221734
rect 508822 221498 544586 221734
rect 544822 221498 580586 221734
rect 580822 221498 587342 221734
rect 587578 221498 588680 221734
rect -4756 221476 588680 221498
rect -3836 221474 -3236 221476
rect 4404 221474 5004 221476
rect 40404 221474 41004 221476
rect 76404 221474 77004 221476
rect 112404 221474 113004 221476
rect 148404 221474 149004 221476
rect 184404 221474 185004 221476
rect 220404 221474 221004 221476
rect 256404 221474 257004 221476
rect 292404 221474 293004 221476
rect 328404 221474 329004 221476
rect 364404 221474 365004 221476
rect 400404 221474 401004 221476
rect 436404 221474 437004 221476
rect 472404 221474 473004 221476
rect 508404 221474 509004 221476
rect 544404 221474 545004 221476
rect 580404 221474 581004 221476
rect 587160 221474 587760 221476
rect -1996 218476 -1396 218478
rect 804 218476 1404 218478
rect 36804 218476 37404 218478
rect 72804 218476 73404 218478
rect 108804 218476 109404 218478
rect 144804 218476 145404 218478
rect 180804 218476 181404 218478
rect 216804 218476 217404 218478
rect 252804 218476 253404 218478
rect 288804 218476 289404 218478
rect 324804 218476 325404 218478
rect 360804 218476 361404 218478
rect 396804 218476 397404 218478
rect 432804 218476 433404 218478
rect 468804 218476 469404 218478
rect 504804 218476 505404 218478
rect 540804 218476 541404 218478
rect 576804 218476 577404 218478
rect 585320 218476 585920 218478
rect -2916 218454 586840 218476
rect -2916 218218 -1814 218454
rect -1578 218218 986 218454
rect 1222 218218 36986 218454
rect 37222 218218 72986 218454
rect 73222 218218 108986 218454
rect 109222 218218 144986 218454
rect 145222 218218 180986 218454
rect 181222 218218 216986 218454
rect 217222 218218 252986 218454
rect 253222 218218 288986 218454
rect 289222 218218 324986 218454
rect 325222 218218 360986 218454
rect 361222 218218 396986 218454
rect 397222 218218 432986 218454
rect 433222 218218 468986 218454
rect 469222 218218 504986 218454
rect 505222 218218 540986 218454
rect 541222 218218 576986 218454
rect 577222 218218 585502 218454
rect 585738 218218 586840 218454
rect -2916 218134 586840 218218
rect -2916 217898 -1814 218134
rect -1578 217898 986 218134
rect 1222 217898 36986 218134
rect 37222 217898 72986 218134
rect 73222 217898 108986 218134
rect 109222 217898 144986 218134
rect 145222 217898 180986 218134
rect 181222 217898 216986 218134
rect 217222 217898 252986 218134
rect 253222 217898 288986 218134
rect 289222 217898 324986 218134
rect 325222 217898 360986 218134
rect 361222 217898 396986 218134
rect 397222 217898 432986 218134
rect 433222 217898 468986 218134
rect 469222 217898 504986 218134
rect 505222 217898 540986 218134
rect 541222 217898 576986 218134
rect 577222 217898 585502 218134
rect 585738 217898 586840 218134
rect -2916 217876 586840 217898
rect -1996 217874 -1396 217876
rect 804 217874 1404 217876
rect 36804 217874 37404 217876
rect 72804 217874 73404 217876
rect 108804 217874 109404 217876
rect 144804 217874 145404 217876
rect 180804 217874 181404 217876
rect 216804 217874 217404 217876
rect 252804 217874 253404 217876
rect 288804 217874 289404 217876
rect 324804 217874 325404 217876
rect 360804 217874 361404 217876
rect 396804 217874 397404 217876
rect 432804 217874 433404 217876
rect 468804 217874 469404 217876
rect 504804 217874 505404 217876
rect 540804 217874 541404 217876
rect 576804 217874 577404 217876
rect 585320 217874 585920 217876
rect -8436 211276 -7836 211278
rect 29604 211276 30204 211278
rect 65604 211276 66204 211278
rect 101604 211276 102204 211278
rect 137604 211276 138204 211278
rect 173604 211276 174204 211278
rect 209604 211276 210204 211278
rect 245604 211276 246204 211278
rect 281604 211276 282204 211278
rect 317604 211276 318204 211278
rect 353604 211276 354204 211278
rect 389604 211276 390204 211278
rect 425604 211276 426204 211278
rect 461604 211276 462204 211278
rect 497604 211276 498204 211278
rect 533604 211276 534204 211278
rect 569604 211276 570204 211278
rect 591760 211276 592360 211278
rect -8436 211254 592360 211276
rect -8436 211018 -8254 211254
rect -8018 211018 29786 211254
rect 30022 211018 65786 211254
rect 66022 211018 101786 211254
rect 102022 211018 137786 211254
rect 138022 211018 173786 211254
rect 174022 211018 209786 211254
rect 210022 211018 245786 211254
rect 246022 211018 281786 211254
rect 282022 211018 317786 211254
rect 318022 211018 353786 211254
rect 354022 211018 389786 211254
rect 390022 211018 425786 211254
rect 426022 211018 461786 211254
rect 462022 211018 497786 211254
rect 498022 211018 533786 211254
rect 534022 211018 569786 211254
rect 570022 211018 591942 211254
rect 592178 211018 592360 211254
rect -8436 210934 592360 211018
rect -8436 210698 -8254 210934
rect -8018 210698 29786 210934
rect 30022 210698 65786 210934
rect 66022 210698 101786 210934
rect 102022 210698 137786 210934
rect 138022 210698 173786 210934
rect 174022 210698 209786 210934
rect 210022 210698 245786 210934
rect 246022 210698 281786 210934
rect 282022 210698 317786 210934
rect 318022 210698 353786 210934
rect 354022 210698 389786 210934
rect 390022 210698 425786 210934
rect 426022 210698 461786 210934
rect 462022 210698 497786 210934
rect 498022 210698 533786 210934
rect 534022 210698 569786 210934
rect 570022 210698 591942 210934
rect 592178 210698 592360 210934
rect -8436 210676 592360 210698
rect -8436 210674 -7836 210676
rect 29604 210674 30204 210676
rect 65604 210674 66204 210676
rect 101604 210674 102204 210676
rect 137604 210674 138204 210676
rect 173604 210674 174204 210676
rect 209604 210674 210204 210676
rect 245604 210674 246204 210676
rect 281604 210674 282204 210676
rect 317604 210674 318204 210676
rect 353604 210674 354204 210676
rect 389604 210674 390204 210676
rect 425604 210674 426204 210676
rect 461604 210674 462204 210676
rect 497604 210674 498204 210676
rect 533604 210674 534204 210676
rect 569604 210674 570204 210676
rect 591760 210674 592360 210676
rect -6596 207676 -5996 207678
rect 26004 207676 26604 207678
rect 62004 207676 62604 207678
rect 98004 207676 98604 207678
rect 134004 207676 134604 207678
rect 170004 207676 170604 207678
rect 206004 207676 206604 207678
rect 242004 207676 242604 207678
rect 278004 207676 278604 207678
rect 314004 207676 314604 207678
rect 350004 207676 350604 207678
rect 386004 207676 386604 207678
rect 422004 207676 422604 207678
rect 458004 207676 458604 207678
rect 494004 207676 494604 207678
rect 530004 207676 530604 207678
rect 566004 207676 566604 207678
rect 589920 207676 590520 207678
rect -6596 207654 590520 207676
rect -6596 207418 -6414 207654
rect -6178 207418 26186 207654
rect 26422 207418 62186 207654
rect 62422 207418 98186 207654
rect 98422 207418 134186 207654
rect 134422 207418 170186 207654
rect 170422 207418 206186 207654
rect 206422 207418 242186 207654
rect 242422 207418 278186 207654
rect 278422 207418 314186 207654
rect 314422 207418 350186 207654
rect 350422 207418 386186 207654
rect 386422 207418 422186 207654
rect 422422 207418 458186 207654
rect 458422 207418 494186 207654
rect 494422 207418 530186 207654
rect 530422 207418 566186 207654
rect 566422 207418 590102 207654
rect 590338 207418 590520 207654
rect -6596 207334 590520 207418
rect -6596 207098 -6414 207334
rect -6178 207098 26186 207334
rect 26422 207098 62186 207334
rect 62422 207098 98186 207334
rect 98422 207098 134186 207334
rect 134422 207098 170186 207334
rect 170422 207098 206186 207334
rect 206422 207098 242186 207334
rect 242422 207098 278186 207334
rect 278422 207098 314186 207334
rect 314422 207098 350186 207334
rect 350422 207098 386186 207334
rect 386422 207098 422186 207334
rect 422422 207098 458186 207334
rect 458422 207098 494186 207334
rect 494422 207098 530186 207334
rect 530422 207098 566186 207334
rect 566422 207098 590102 207334
rect 590338 207098 590520 207334
rect -6596 207076 590520 207098
rect -6596 207074 -5996 207076
rect 26004 207074 26604 207076
rect 62004 207074 62604 207076
rect 98004 207074 98604 207076
rect 134004 207074 134604 207076
rect 170004 207074 170604 207076
rect 206004 207074 206604 207076
rect 242004 207074 242604 207076
rect 278004 207074 278604 207076
rect 314004 207074 314604 207076
rect 350004 207074 350604 207076
rect 386004 207074 386604 207076
rect 422004 207074 422604 207076
rect 458004 207074 458604 207076
rect 494004 207074 494604 207076
rect 530004 207074 530604 207076
rect 566004 207074 566604 207076
rect 589920 207074 590520 207076
rect -4756 204076 -4156 204078
rect 22404 204076 23004 204078
rect 58404 204076 59004 204078
rect 94404 204076 95004 204078
rect 130404 204076 131004 204078
rect 166404 204076 167004 204078
rect 202404 204076 203004 204078
rect 238404 204076 239004 204078
rect 274404 204076 275004 204078
rect 310404 204076 311004 204078
rect 346404 204076 347004 204078
rect 382404 204076 383004 204078
rect 418404 204076 419004 204078
rect 454404 204076 455004 204078
rect 490404 204076 491004 204078
rect 526404 204076 527004 204078
rect 562404 204076 563004 204078
rect 588080 204076 588680 204078
rect -4756 204054 588680 204076
rect -4756 203818 -4574 204054
rect -4338 203818 22586 204054
rect 22822 203818 58586 204054
rect 58822 203818 94586 204054
rect 94822 203818 130586 204054
rect 130822 203818 166586 204054
rect 166822 203818 202586 204054
rect 202822 203818 238586 204054
rect 238822 203818 274586 204054
rect 274822 203818 310586 204054
rect 310822 203818 346586 204054
rect 346822 203818 382586 204054
rect 382822 203818 418586 204054
rect 418822 203818 454586 204054
rect 454822 203818 490586 204054
rect 490822 203818 526586 204054
rect 526822 203818 562586 204054
rect 562822 203818 588262 204054
rect 588498 203818 588680 204054
rect -4756 203734 588680 203818
rect -4756 203498 -4574 203734
rect -4338 203498 22586 203734
rect 22822 203498 58586 203734
rect 58822 203498 94586 203734
rect 94822 203498 130586 203734
rect 130822 203498 166586 203734
rect 166822 203498 202586 203734
rect 202822 203498 238586 203734
rect 238822 203498 274586 203734
rect 274822 203498 310586 203734
rect 310822 203498 346586 203734
rect 346822 203498 382586 203734
rect 382822 203498 418586 203734
rect 418822 203498 454586 203734
rect 454822 203498 490586 203734
rect 490822 203498 526586 203734
rect 526822 203498 562586 203734
rect 562822 203498 588262 203734
rect 588498 203498 588680 203734
rect -4756 203476 588680 203498
rect -4756 203474 -4156 203476
rect 22404 203474 23004 203476
rect 58404 203474 59004 203476
rect 94404 203474 95004 203476
rect 130404 203474 131004 203476
rect 166404 203474 167004 203476
rect 202404 203474 203004 203476
rect 238404 203474 239004 203476
rect 274404 203474 275004 203476
rect 310404 203474 311004 203476
rect 346404 203474 347004 203476
rect 382404 203474 383004 203476
rect 418404 203474 419004 203476
rect 454404 203474 455004 203476
rect 490404 203474 491004 203476
rect 526404 203474 527004 203476
rect 562404 203474 563004 203476
rect 588080 203474 588680 203476
rect -2916 200476 -2316 200478
rect 18804 200476 19404 200478
rect 54804 200476 55404 200478
rect 90804 200476 91404 200478
rect 126804 200476 127404 200478
rect 162804 200476 163404 200478
rect 198804 200476 199404 200478
rect 234804 200476 235404 200478
rect 270804 200476 271404 200478
rect 306804 200476 307404 200478
rect 342804 200476 343404 200478
rect 378804 200476 379404 200478
rect 414804 200476 415404 200478
rect 450804 200476 451404 200478
rect 486804 200476 487404 200478
rect 522804 200476 523404 200478
rect 558804 200476 559404 200478
rect 586240 200476 586840 200478
rect -2916 200454 586840 200476
rect -2916 200218 -2734 200454
rect -2498 200218 18986 200454
rect 19222 200218 54986 200454
rect 55222 200218 90986 200454
rect 91222 200218 126986 200454
rect 127222 200218 162986 200454
rect 163222 200218 198986 200454
rect 199222 200218 234986 200454
rect 235222 200218 270986 200454
rect 271222 200218 306986 200454
rect 307222 200218 342986 200454
rect 343222 200218 378986 200454
rect 379222 200218 414986 200454
rect 415222 200218 450986 200454
rect 451222 200218 486986 200454
rect 487222 200218 522986 200454
rect 523222 200218 558986 200454
rect 559222 200218 586422 200454
rect 586658 200218 586840 200454
rect -2916 200134 586840 200218
rect -2916 199898 -2734 200134
rect -2498 199898 18986 200134
rect 19222 199898 54986 200134
rect 55222 199898 90986 200134
rect 91222 199898 126986 200134
rect 127222 199898 162986 200134
rect 163222 199898 198986 200134
rect 199222 199898 234986 200134
rect 235222 199898 270986 200134
rect 271222 199898 306986 200134
rect 307222 199898 342986 200134
rect 343222 199898 378986 200134
rect 379222 199898 414986 200134
rect 415222 199898 450986 200134
rect 451222 199898 486986 200134
rect 487222 199898 522986 200134
rect 523222 199898 558986 200134
rect 559222 199898 586422 200134
rect 586658 199898 586840 200134
rect -2916 199876 586840 199898
rect -2916 199874 -2316 199876
rect 18804 199874 19404 199876
rect 54804 199874 55404 199876
rect 90804 199874 91404 199876
rect 126804 199874 127404 199876
rect 162804 199874 163404 199876
rect 198804 199874 199404 199876
rect 234804 199874 235404 199876
rect 270804 199874 271404 199876
rect 306804 199874 307404 199876
rect 342804 199874 343404 199876
rect 378804 199874 379404 199876
rect 414804 199874 415404 199876
rect 450804 199874 451404 199876
rect 486804 199874 487404 199876
rect 522804 199874 523404 199876
rect 558804 199874 559404 199876
rect 586240 199874 586840 199876
rect -7516 193276 -6916 193278
rect 11604 193276 12204 193278
rect 47604 193276 48204 193278
rect 83604 193276 84204 193278
rect 119604 193276 120204 193278
rect 155604 193276 156204 193278
rect 191604 193276 192204 193278
rect 227604 193276 228204 193278
rect 263604 193276 264204 193278
rect 299604 193276 300204 193278
rect 335604 193276 336204 193278
rect 371604 193276 372204 193278
rect 407604 193276 408204 193278
rect 443604 193276 444204 193278
rect 479604 193276 480204 193278
rect 515604 193276 516204 193278
rect 551604 193276 552204 193278
rect 590840 193276 591440 193278
rect -8436 193254 592360 193276
rect -8436 193018 -7334 193254
rect -7098 193018 11786 193254
rect 12022 193018 47786 193254
rect 48022 193018 83786 193254
rect 84022 193018 119786 193254
rect 120022 193018 155786 193254
rect 156022 193018 191786 193254
rect 192022 193018 227786 193254
rect 228022 193018 263786 193254
rect 264022 193018 299786 193254
rect 300022 193018 335786 193254
rect 336022 193018 371786 193254
rect 372022 193018 407786 193254
rect 408022 193018 443786 193254
rect 444022 193018 479786 193254
rect 480022 193018 515786 193254
rect 516022 193018 551786 193254
rect 552022 193018 591022 193254
rect 591258 193018 592360 193254
rect -8436 192934 592360 193018
rect -8436 192698 -7334 192934
rect -7098 192698 11786 192934
rect 12022 192698 47786 192934
rect 48022 192698 83786 192934
rect 84022 192698 119786 192934
rect 120022 192698 155786 192934
rect 156022 192698 191786 192934
rect 192022 192698 227786 192934
rect 228022 192698 263786 192934
rect 264022 192698 299786 192934
rect 300022 192698 335786 192934
rect 336022 192698 371786 192934
rect 372022 192698 407786 192934
rect 408022 192698 443786 192934
rect 444022 192698 479786 192934
rect 480022 192698 515786 192934
rect 516022 192698 551786 192934
rect 552022 192698 591022 192934
rect 591258 192698 592360 192934
rect -8436 192676 592360 192698
rect -7516 192674 -6916 192676
rect 11604 192674 12204 192676
rect 47604 192674 48204 192676
rect 83604 192674 84204 192676
rect 119604 192674 120204 192676
rect 155604 192674 156204 192676
rect 191604 192674 192204 192676
rect 227604 192674 228204 192676
rect 263604 192674 264204 192676
rect 299604 192674 300204 192676
rect 335604 192674 336204 192676
rect 371604 192674 372204 192676
rect 407604 192674 408204 192676
rect 443604 192674 444204 192676
rect 479604 192674 480204 192676
rect 515604 192674 516204 192676
rect 551604 192674 552204 192676
rect 590840 192674 591440 192676
rect -5676 189676 -5076 189678
rect 8004 189676 8604 189678
rect 44004 189676 44604 189678
rect 80004 189676 80604 189678
rect 116004 189676 116604 189678
rect 152004 189676 152604 189678
rect 188004 189676 188604 189678
rect 224004 189676 224604 189678
rect 260004 189676 260604 189678
rect 296004 189676 296604 189678
rect 332004 189676 332604 189678
rect 368004 189676 368604 189678
rect 404004 189676 404604 189678
rect 440004 189676 440604 189678
rect 476004 189676 476604 189678
rect 512004 189676 512604 189678
rect 548004 189676 548604 189678
rect 589000 189676 589600 189678
rect -6596 189654 590520 189676
rect -6596 189418 -5494 189654
rect -5258 189418 8186 189654
rect 8422 189418 44186 189654
rect 44422 189418 80186 189654
rect 80422 189418 116186 189654
rect 116422 189418 152186 189654
rect 152422 189418 188186 189654
rect 188422 189418 224186 189654
rect 224422 189418 260186 189654
rect 260422 189418 296186 189654
rect 296422 189418 332186 189654
rect 332422 189418 368186 189654
rect 368422 189418 404186 189654
rect 404422 189418 440186 189654
rect 440422 189418 476186 189654
rect 476422 189418 512186 189654
rect 512422 189418 548186 189654
rect 548422 189418 589182 189654
rect 589418 189418 590520 189654
rect -6596 189334 590520 189418
rect -6596 189098 -5494 189334
rect -5258 189098 8186 189334
rect 8422 189098 44186 189334
rect 44422 189098 80186 189334
rect 80422 189098 116186 189334
rect 116422 189098 152186 189334
rect 152422 189098 188186 189334
rect 188422 189098 224186 189334
rect 224422 189098 260186 189334
rect 260422 189098 296186 189334
rect 296422 189098 332186 189334
rect 332422 189098 368186 189334
rect 368422 189098 404186 189334
rect 404422 189098 440186 189334
rect 440422 189098 476186 189334
rect 476422 189098 512186 189334
rect 512422 189098 548186 189334
rect 548422 189098 589182 189334
rect 589418 189098 590520 189334
rect -6596 189076 590520 189098
rect -5676 189074 -5076 189076
rect 8004 189074 8604 189076
rect 44004 189074 44604 189076
rect 80004 189074 80604 189076
rect 116004 189074 116604 189076
rect 152004 189074 152604 189076
rect 188004 189074 188604 189076
rect 224004 189074 224604 189076
rect 260004 189074 260604 189076
rect 296004 189074 296604 189076
rect 332004 189074 332604 189076
rect 368004 189074 368604 189076
rect 404004 189074 404604 189076
rect 440004 189074 440604 189076
rect 476004 189074 476604 189076
rect 512004 189074 512604 189076
rect 548004 189074 548604 189076
rect 589000 189074 589600 189076
rect -3836 186076 -3236 186078
rect 4404 186076 5004 186078
rect 40404 186076 41004 186078
rect 76404 186076 77004 186078
rect 112404 186076 113004 186078
rect 148404 186076 149004 186078
rect 184404 186076 185004 186078
rect 220404 186076 221004 186078
rect 256404 186076 257004 186078
rect 292404 186076 293004 186078
rect 328404 186076 329004 186078
rect 364404 186076 365004 186078
rect 400404 186076 401004 186078
rect 436404 186076 437004 186078
rect 472404 186076 473004 186078
rect 508404 186076 509004 186078
rect 544404 186076 545004 186078
rect 580404 186076 581004 186078
rect 587160 186076 587760 186078
rect -4756 186054 588680 186076
rect -4756 185818 -3654 186054
rect -3418 185818 4586 186054
rect 4822 185818 40586 186054
rect 40822 185818 76586 186054
rect 76822 185818 112586 186054
rect 112822 185818 148586 186054
rect 148822 185818 184586 186054
rect 184822 185818 220586 186054
rect 220822 185818 256586 186054
rect 256822 185818 292586 186054
rect 292822 185818 328586 186054
rect 328822 185818 364586 186054
rect 364822 185818 400586 186054
rect 400822 185818 436586 186054
rect 436822 185818 472586 186054
rect 472822 185818 508586 186054
rect 508822 185818 544586 186054
rect 544822 185818 580586 186054
rect 580822 185818 587342 186054
rect 587578 185818 588680 186054
rect -4756 185734 588680 185818
rect -4756 185498 -3654 185734
rect -3418 185498 4586 185734
rect 4822 185498 40586 185734
rect 40822 185498 76586 185734
rect 76822 185498 112586 185734
rect 112822 185498 148586 185734
rect 148822 185498 184586 185734
rect 184822 185498 220586 185734
rect 220822 185498 256586 185734
rect 256822 185498 292586 185734
rect 292822 185498 328586 185734
rect 328822 185498 364586 185734
rect 364822 185498 400586 185734
rect 400822 185498 436586 185734
rect 436822 185498 472586 185734
rect 472822 185498 508586 185734
rect 508822 185498 544586 185734
rect 544822 185498 580586 185734
rect 580822 185498 587342 185734
rect 587578 185498 588680 185734
rect -4756 185476 588680 185498
rect -3836 185474 -3236 185476
rect 4404 185474 5004 185476
rect 40404 185474 41004 185476
rect 76404 185474 77004 185476
rect 112404 185474 113004 185476
rect 148404 185474 149004 185476
rect 184404 185474 185004 185476
rect 220404 185474 221004 185476
rect 256404 185474 257004 185476
rect 292404 185474 293004 185476
rect 328404 185474 329004 185476
rect 364404 185474 365004 185476
rect 400404 185474 401004 185476
rect 436404 185474 437004 185476
rect 472404 185474 473004 185476
rect 508404 185474 509004 185476
rect 544404 185474 545004 185476
rect 580404 185474 581004 185476
rect 587160 185474 587760 185476
rect -1996 182476 -1396 182478
rect 804 182476 1404 182478
rect 36804 182476 37404 182478
rect 72804 182476 73404 182478
rect 108804 182476 109404 182478
rect 144804 182476 145404 182478
rect 180804 182476 181404 182478
rect 216804 182476 217404 182478
rect 252804 182476 253404 182478
rect 288804 182476 289404 182478
rect 324804 182476 325404 182478
rect 360804 182476 361404 182478
rect 396804 182476 397404 182478
rect 432804 182476 433404 182478
rect 468804 182476 469404 182478
rect 504804 182476 505404 182478
rect 540804 182476 541404 182478
rect 576804 182476 577404 182478
rect 585320 182476 585920 182478
rect -2916 182454 586840 182476
rect -2916 182218 -1814 182454
rect -1578 182218 986 182454
rect 1222 182218 36986 182454
rect 37222 182218 72986 182454
rect 73222 182218 108986 182454
rect 109222 182218 144986 182454
rect 145222 182218 180986 182454
rect 181222 182218 216986 182454
rect 217222 182218 252986 182454
rect 253222 182218 288986 182454
rect 289222 182218 324986 182454
rect 325222 182218 360986 182454
rect 361222 182218 396986 182454
rect 397222 182218 432986 182454
rect 433222 182218 468986 182454
rect 469222 182218 504986 182454
rect 505222 182218 540986 182454
rect 541222 182218 576986 182454
rect 577222 182218 585502 182454
rect 585738 182218 586840 182454
rect -2916 182134 586840 182218
rect -2916 181898 -1814 182134
rect -1578 181898 986 182134
rect 1222 181898 36986 182134
rect 37222 181898 72986 182134
rect 73222 181898 108986 182134
rect 109222 181898 144986 182134
rect 145222 181898 180986 182134
rect 181222 181898 216986 182134
rect 217222 181898 252986 182134
rect 253222 181898 288986 182134
rect 289222 181898 324986 182134
rect 325222 181898 360986 182134
rect 361222 181898 396986 182134
rect 397222 181898 432986 182134
rect 433222 181898 468986 182134
rect 469222 181898 504986 182134
rect 505222 181898 540986 182134
rect 541222 181898 576986 182134
rect 577222 181898 585502 182134
rect 585738 181898 586840 182134
rect -2916 181876 586840 181898
rect -1996 181874 -1396 181876
rect 804 181874 1404 181876
rect 36804 181874 37404 181876
rect 72804 181874 73404 181876
rect 108804 181874 109404 181876
rect 144804 181874 145404 181876
rect 180804 181874 181404 181876
rect 216804 181874 217404 181876
rect 252804 181874 253404 181876
rect 288804 181874 289404 181876
rect 324804 181874 325404 181876
rect 360804 181874 361404 181876
rect 396804 181874 397404 181876
rect 432804 181874 433404 181876
rect 468804 181874 469404 181876
rect 504804 181874 505404 181876
rect 540804 181874 541404 181876
rect 576804 181874 577404 181876
rect 585320 181874 585920 181876
rect -8436 175276 -7836 175278
rect 29604 175276 30204 175278
rect 65604 175276 66204 175278
rect 101604 175276 102204 175278
rect 137604 175276 138204 175278
rect 173604 175276 174204 175278
rect 209604 175276 210204 175278
rect 245604 175276 246204 175278
rect 281604 175276 282204 175278
rect 317604 175276 318204 175278
rect 353604 175276 354204 175278
rect 389604 175276 390204 175278
rect 425604 175276 426204 175278
rect 461604 175276 462204 175278
rect 497604 175276 498204 175278
rect 533604 175276 534204 175278
rect 569604 175276 570204 175278
rect 591760 175276 592360 175278
rect -8436 175254 592360 175276
rect -8436 175018 -8254 175254
rect -8018 175018 29786 175254
rect 30022 175018 65786 175254
rect 66022 175018 101786 175254
rect 102022 175018 137786 175254
rect 138022 175018 173786 175254
rect 174022 175018 209786 175254
rect 210022 175018 245786 175254
rect 246022 175018 281786 175254
rect 282022 175018 317786 175254
rect 318022 175018 353786 175254
rect 354022 175018 389786 175254
rect 390022 175018 425786 175254
rect 426022 175018 461786 175254
rect 462022 175018 497786 175254
rect 498022 175018 533786 175254
rect 534022 175018 569786 175254
rect 570022 175018 591942 175254
rect 592178 175018 592360 175254
rect -8436 174934 592360 175018
rect -8436 174698 -8254 174934
rect -8018 174698 29786 174934
rect 30022 174698 65786 174934
rect 66022 174698 101786 174934
rect 102022 174698 137786 174934
rect 138022 174698 173786 174934
rect 174022 174698 209786 174934
rect 210022 174698 245786 174934
rect 246022 174698 281786 174934
rect 282022 174698 317786 174934
rect 318022 174698 353786 174934
rect 354022 174698 389786 174934
rect 390022 174698 425786 174934
rect 426022 174698 461786 174934
rect 462022 174698 497786 174934
rect 498022 174698 533786 174934
rect 534022 174698 569786 174934
rect 570022 174698 591942 174934
rect 592178 174698 592360 174934
rect -8436 174676 592360 174698
rect -8436 174674 -7836 174676
rect 29604 174674 30204 174676
rect 65604 174674 66204 174676
rect 101604 174674 102204 174676
rect 137604 174674 138204 174676
rect 173604 174674 174204 174676
rect 209604 174674 210204 174676
rect 245604 174674 246204 174676
rect 281604 174674 282204 174676
rect 317604 174674 318204 174676
rect 353604 174674 354204 174676
rect 389604 174674 390204 174676
rect 425604 174674 426204 174676
rect 461604 174674 462204 174676
rect 497604 174674 498204 174676
rect 533604 174674 534204 174676
rect 569604 174674 570204 174676
rect 591760 174674 592360 174676
rect -6596 171676 -5996 171678
rect 26004 171676 26604 171678
rect 62004 171676 62604 171678
rect 98004 171676 98604 171678
rect 134004 171676 134604 171678
rect 170004 171676 170604 171678
rect 206004 171676 206604 171678
rect 242004 171676 242604 171678
rect 278004 171676 278604 171678
rect 314004 171676 314604 171678
rect 350004 171676 350604 171678
rect 386004 171676 386604 171678
rect 422004 171676 422604 171678
rect 458004 171676 458604 171678
rect 494004 171676 494604 171678
rect 530004 171676 530604 171678
rect 566004 171676 566604 171678
rect 589920 171676 590520 171678
rect -6596 171654 590520 171676
rect -6596 171418 -6414 171654
rect -6178 171418 26186 171654
rect 26422 171418 62186 171654
rect 62422 171418 98186 171654
rect 98422 171418 134186 171654
rect 134422 171418 170186 171654
rect 170422 171418 206186 171654
rect 206422 171418 242186 171654
rect 242422 171418 278186 171654
rect 278422 171418 314186 171654
rect 314422 171418 350186 171654
rect 350422 171418 386186 171654
rect 386422 171418 422186 171654
rect 422422 171418 458186 171654
rect 458422 171418 494186 171654
rect 494422 171418 530186 171654
rect 530422 171418 566186 171654
rect 566422 171418 590102 171654
rect 590338 171418 590520 171654
rect -6596 171334 590520 171418
rect -6596 171098 -6414 171334
rect -6178 171098 26186 171334
rect 26422 171098 62186 171334
rect 62422 171098 98186 171334
rect 98422 171098 134186 171334
rect 134422 171098 170186 171334
rect 170422 171098 206186 171334
rect 206422 171098 242186 171334
rect 242422 171098 278186 171334
rect 278422 171098 314186 171334
rect 314422 171098 350186 171334
rect 350422 171098 386186 171334
rect 386422 171098 422186 171334
rect 422422 171098 458186 171334
rect 458422 171098 494186 171334
rect 494422 171098 530186 171334
rect 530422 171098 566186 171334
rect 566422 171098 590102 171334
rect 590338 171098 590520 171334
rect -6596 171076 590520 171098
rect -6596 171074 -5996 171076
rect 26004 171074 26604 171076
rect 62004 171074 62604 171076
rect 98004 171074 98604 171076
rect 134004 171074 134604 171076
rect 170004 171074 170604 171076
rect 206004 171074 206604 171076
rect 242004 171074 242604 171076
rect 278004 171074 278604 171076
rect 314004 171074 314604 171076
rect 350004 171074 350604 171076
rect 386004 171074 386604 171076
rect 422004 171074 422604 171076
rect 458004 171074 458604 171076
rect 494004 171074 494604 171076
rect 530004 171074 530604 171076
rect 566004 171074 566604 171076
rect 589920 171074 590520 171076
rect -4756 168076 -4156 168078
rect 22404 168076 23004 168078
rect 58404 168076 59004 168078
rect 94404 168076 95004 168078
rect 130404 168076 131004 168078
rect 166404 168076 167004 168078
rect 202404 168076 203004 168078
rect 238404 168076 239004 168078
rect 274404 168076 275004 168078
rect 310404 168076 311004 168078
rect 346404 168076 347004 168078
rect 382404 168076 383004 168078
rect 418404 168076 419004 168078
rect 454404 168076 455004 168078
rect 490404 168076 491004 168078
rect 526404 168076 527004 168078
rect 562404 168076 563004 168078
rect 588080 168076 588680 168078
rect -4756 168054 588680 168076
rect -4756 167818 -4574 168054
rect -4338 167818 22586 168054
rect 22822 167818 58586 168054
rect 58822 167818 94586 168054
rect 94822 167818 130586 168054
rect 130822 167818 166586 168054
rect 166822 167818 202586 168054
rect 202822 167818 238586 168054
rect 238822 167818 274586 168054
rect 274822 167818 310586 168054
rect 310822 167818 346586 168054
rect 346822 167818 382586 168054
rect 382822 167818 418586 168054
rect 418822 167818 454586 168054
rect 454822 167818 490586 168054
rect 490822 167818 526586 168054
rect 526822 167818 562586 168054
rect 562822 167818 588262 168054
rect 588498 167818 588680 168054
rect -4756 167734 588680 167818
rect -4756 167498 -4574 167734
rect -4338 167498 22586 167734
rect 22822 167498 58586 167734
rect 58822 167498 94586 167734
rect 94822 167498 130586 167734
rect 130822 167498 166586 167734
rect 166822 167498 202586 167734
rect 202822 167498 238586 167734
rect 238822 167498 274586 167734
rect 274822 167498 310586 167734
rect 310822 167498 346586 167734
rect 346822 167498 382586 167734
rect 382822 167498 418586 167734
rect 418822 167498 454586 167734
rect 454822 167498 490586 167734
rect 490822 167498 526586 167734
rect 526822 167498 562586 167734
rect 562822 167498 588262 167734
rect 588498 167498 588680 167734
rect -4756 167476 588680 167498
rect -4756 167474 -4156 167476
rect 22404 167474 23004 167476
rect 58404 167474 59004 167476
rect 94404 167474 95004 167476
rect 130404 167474 131004 167476
rect 166404 167474 167004 167476
rect 202404 167474 203004 167476
rect 238404 167474 239004 167476
rect 274404 167474 275004 167476
rect 310404 167474 311004 167476
rect 346404 167474 347004 167476
rect 382404 167474 383004 167476
rect 418404 167474 419004 167476
rect 454404 167474 455004 167476
rect 490404 167474 491004 167476
rect 526404 167474 527004 167476
rect 562404 167474 563004 167476
rect 588080 167474 588680 167476
rect -2916 164476 -2316 164478
rect 18804 164476 19404 164478
rect 54804 164476 55404 164478
rect 90804 164476 91404 164478
rect 126804 164476 127404 164478
rect 162804 164476 163404 164478
rect 198804 164476 199404 164478
rect 234804 164476 235404 164478
rect 270804 164476 271404 164478
rect 306804 164476 307404 164478
rect 342804 164476 343404 164478
rect 378804 164476 379404 164478
rect 414804 164476 415404 164478
rect 450804 164476 451404 164478
rect 486804 164476 487404 164478
rect 522804 164476 523404 164478
rect 558804 164476 559404 164478
rect 586240 164476 586840 164478
rect -2916 164454 586840 164476
rect -2916 164218 -2734 164454
rect -2498 164218 18986 164454
rect 19222 164218 54986 164454
rect 55222 164218 90986 164454
rect 91222 164218 126986 164454
rect 127222 164218 162986 164454
rect 163222 164218 198986 164454
rect 199222 164218 234986 164454
rect 235222 164218 270986 164454
rect 271222 164218 306986 164454
rect 307222 164218 342986 164454
rect 343222 164218 378986 164454
rect 379222 164218 414986 164454
rect 415222 164218 450986 164454
rect 451222 164218 486986 164454
rect 487222 164218 522986 164454
rect 523222 164218 558986 164454
rect 559222 164218 586422 164454
rect 586658 164218 586840 164454
rect -2916 164134 586840 164218
rect -2916 163898 -2734 164134
rect -2498 163898 18986 164134
rect 19222 163898 54986 164134
rect 55222 163898 90986 164134
rect 91222 163898 126986 164134
rect 127222 163898 162986 164134
rect 163222 163898 198986 164134
rect 199222 163898 234986 164134
rect 235222 163898 270986 164134
rect 271222 163898 306986 164134
rect 307222 163898 342986 164134
rect 343222 163898 378986 164134
rect 379222 163898 414986 164134
rect 415222 163898 450986 164134
rect 451222 163898 486986 164134
rect 487222 163898 522986 164134
rect 523222 163898 558986 164134
rect 559222 163898 586422 164134
rect 586658 163898 586840 164134
rect -2916 163876 586840 163898
rect -2916 163874 -2316 163876
rect 18804 163874 19404 163876
rect 54804 163874 55404 163876
rect 90804 163874 91404 163876
rect 126804 163874 127404 163876
rect 162804 163874 163404 163876
rect 198804 163874 199404 163876
rect 234804 163874 235404 163876
rect 270804 163874 271404 163876
rect 306804 163874 307404 163876
rect 342804 163874 343404 163876
rect 378804 163874 379404 163876
rect 414804 163874 415404 163876
rect 450804 163874 451404 163876
rect 486804 163874 487404 163876
rect 522804 163874 523404 163876
rect 558804 163874 559404 163876
rect 586240 163874 586840 163876
rect -7516 157276 -6916 157278
rect 11604 157276 12204 157278
rect 47604 157276 48204 157278
rect 83604 157276 84204 157278
rect 119604 157276 120204 157278
rect 155604 157276 156204 157278
rect 191604 157276 192204 157278
rect 227604 157276 228204 157278
rect 263604 157276 264204 157278
rect 299604 157276 300204 157278
rect 335604 157276 336204 157278
rect 371604 157276 372204 157278
rect 407604 157276 408204 157278
rect 443604 157276 444204 157278
rect 479604 157276 480204 157278
rect 515604 157276 516204 157278
rect 551604 157276 552204 157278
rect 590840 157276 591440 157278
rect -8436 157254 592360 157276
rect -8436 157018 -7334 157254
rect -7098 157018 11786 157254
rect 12022 157018 47786 157254
rect 48022 157018 83786 157254
rect 84022 157018 119786 157254
rect 120022 157018 155786 157254
rect 156022 157018 191786 157254
rect 192022 157018 227786 157254
rect 228022 157018 263786 157254
rect 264022 157018 299786 157254
rect 300022 157018 335786 157254
rect 336022 157018 371786 157254
rect 372022 157018 407786 157254
rect 408022 157018 443786 157254
rect 444022 157018 479786 157254
rect 480022 157018 515786 157254
rect 516022 157018 551786 157254
rect 552022 157018 591022 157254
rect 591258 157018 592360 157254
rect -8436 156934 592360 157018
rect -8436 156698 -7334 156934
rect -7098 156698 11786 156934
rect 12022 156698 47786 156934
rect 48022 156698 83786 156934
rect 84022 156698 119786 156934
rect 120022 156698 155786 156934
rect 156022 156698 191786 156934
rect 192022 156698 227786 156934
rect 228022 156698 263786 156934
rect 264022 156698 299786 156934
rect 300022 156698 335786 156934
rect 336022 156698 371786 156934
rect 372022 156698 407786 156934
rect 408022 156698 443786 156934
rect 444022 156698 479786 156934
rect 480022 156698 515786 156934
rect 516022 156698 551786 156934
rect 552022 156698 591022 156934
rect 591258 156698 592360 156934
rect -8436 156676 592360 156698
rect -7516 156674 -6916 156676
rect 11604 156674 12204 156676
rect 47604 156674 48204 156676
rect 83604 156674 84204 156676
rect 119604 156674 120204 156676
rect 155604 156674 156204 156676
rect 191604 156674 192204 156676
rect 227604 156674 228204 156676
rect 263604 156674 264204 156676
rect 299604 156674 300204 156676
rect 335604 156674 336204 156676
rect 371604 156674 372204 156676
rect 407604 156674 408204 156676
rect 443604 156674 444204 156676
rect 479604 156674 480204 156676
rect 515604 156674 516204 156676
rect 551604 156674 552204 156676
rect 590840 156674 591440 156676
rect -5676 153676 -5076 153678
rect 8004 153676 8604 153678
rect 44004 153676 44604 153678
rect 80004 153676 80604 153678
rect 116004 153676 116604 153678
rect 152004 153676 152604 153678
rect 188004 153676 188604 153678
rect 224004 153676 224604 153678
rect 260004 153676 260604 153678
rect 296004 153676 296604 153678
rect 332004 153676 332604 153678
rect 368004 153676 368604 153678
rect 404004 153676 404604 153678
rect 440004 153676 440604 153678
rect 476004 153676 476604 153678
rect 512004 153676 512604 153678
rect 548004 153676 548604 153678
rect 589000 153676 589600 153678
rect -6596 153654 590520 153676
rect -6596 153418 -5494 153654
rect -5258 153418 8186 153654
rect 8422 153418 44186 153654
rect 44422 153418 80186 153654
rect 80422 153418 116186 153654
rect 116422 153418 152186 153654
rect 152422 153418 188186 153654
rect 188422 153418 224186 153654
rect 224422 153418 260186 153654
rect 260422 153418 296186 153654
rect 296422 153418 332186 153654
rect 332422 153418 368186 153654
rect 368422 153418 404186 153654
rect 404422 153418 440186 153654
rect 440422 153418 476186 153654
rect 476422 153418 512186 153654
rect 512422 153418 548186 153654
rect 548422 153418 589182 153654
rect 589418 153418 590520 153654
rect -6596 153334 590520 153418
rect -6596 153098 -5494 153334
rect -5258 153098 8186 153334
rect 8422 153098 44186 153334
rect 44422 153098 80186 153334
rect 80422 153098 116186 153334
rect 116422 153098 152186 153334
rect 152422 153098 188186 153334
rect 188422 153098 224186 153334
rect 224422 153098 260186 153334
rect 260422 153098 296186 153334
rect 296422 153098 332186 153334
rect 332422 153098 368186 153334
rect 368422 153098 404186 153334
rect 404422 153098 440186 153334
rect 440422 153098 476186 153334
rect 476422 153098 512186 153334
rect 512422 153098 548186 153334
rect 548422 153098 589182 153334
rect 589418 153098 590520 153334
rect -6596 153076 590520 153098
rect -5676 153074 -5076 153076
rect 8004 153074 8604 153076
rect 44004 153074 44604 153076
rect 80004 153074 80604 153076
rect 116004 153074 116604 153076
rect 152004 153074 152604 153076
rect 188004 153074 188604 153076
rect 224004 153074 224604 153076
rect 260004 153074 260604 153076
rect 296004 153074 296604 153076
rect 332004 153074 332604 153076
rect 368004 153074 368604 153076
rect 404004 153074 404604 153076
rect 440004 153074 440604 153076
rect 476004 153074 476604 153076
rect 512004 153074 512604 153076
rect 548004 153074 548604 153076
rect 589000 153074 589600 153076
rect -3836 150076 -3236 150078
rect 4404 150076 5004 150078
rect 40404 150076 41004 150078
rect 76404 150076 77004 150078
rect 112404 150076 113004 150078
rect 148404 150076 149004 150078
rect 184404 150076 185004 150078
rect 220404 150076 221004 150078
rect 256404 150076 257004 150078
rect 292404 150076 293004 150078
rect 328404 150076 329004 150078
rect 364404 150076 365004 150078
rect 400404 150076 401004 150078
rect 436404 150076 437004 150078
rect 472404 150076 473004 150078
rect 508404 150076 509004 150078
rect 544404 150076 545004 150078
rect 580404 150076 581004 150078
rect 587160 150076 587760 150078
rect -4756 150054 588680 150076
rect -4756 149818 -3654 150054
rect -3418 149818 4586 150054
rect 4822 149818 40586 150054
rect 40822 149818 76586 150054
rect 76822 149818 112586 150054
rect 112822 149818 148586 150054
rect 148822 149818 184586 150054
rect 184822 149818 220586 150054
rect 220822 149818 256586 150054
rect 256822 149818 292586 150054
rect 292822 149818 328586 150054
rect 328822 149818 364586 150054
rect 364822 149818 400586 150054
rect 400822 149818 436586 150054
rect 436822 149818 472586 150054
rect 472822 149818 508586 150054
rect 508822 149818 544586 150054
rect 544822 149818 580586 150054
rect 580822 149818 587342 150054
rect 587578 149818 588680 150054
rect -4756 149734 588680 149818
rect -4756 149498 -3654 149734
rect -3418 149498 4586 149734
rect 4822 149498 40586 149734
rect 40822 149498 76586 149734
rect 76822 149498 112586 149734
rect 112822 149498 148586 149734
rect 148822 149498 184586 149734
rect 184822 149498 220586 149734
rect 220822 149498 256586 149734
rect 256822 149498 292586 149734
rect 292822 149498 328586 149734
rect 328822 149498 364586 149734
rect 364822 149498 400586 149734
rect 400822 149498 436586 149734
rect 436822 149498 472586 149734
rect 472822 149498 508586 149734
rect 508822 149498 544586 149734
rect 544822 149498 580586 149734
rect 580822 149498 587342 149734
rect 587578 149498 588680 149734
rect -4756 149476 588680 149498
rect -3836 149474 -3236 149476
rect 4404 149474 5004 149476
rect 40404 149474 41004 149476
rect 76404 149474 77004 149476
rect 112404 149474 113004 149476
rect 148404 149474 149004 149476
rect 184404 149474 185004 149476
rect 220404 149474 221004 149476
rect 256404 149474 257004 149476
rect 292404 149474 293004 149476
rect 328404 149474 329004 149476
rect 364404 149474 365004 149476
rect 400404 149474 401004 149476
rect 436404 149474 437004 149476
rect 472404 149474 473004 149476
rect 508404 149474 509004 149476
rect 544404 149474 545004 149476
rect 580404 149474 581004 149476
rect 587160 149474 587760 149476
rect -1996 146476 -1396 146478
rect 804 146476 1404 146478
rect 36804 146476 37404 146478
rect 72804 146476 73404 146478
rect 108804 146476 109404 146478
rect 144804 146476 145404 146478
rect 180804 146476 181404 146478
rect 216804 146476 217404 146478
rect 252804 146476 253404 146478
rect 288804 146476 289404 146478
rect 324804 146476 325404 146478
rect 360804 146476 361404 146478
rect 396804 146476 397404 146478
rect 432804 146476 433404 146478
rect 468804 146476 469404 146478
rect 504804 146476 505404 146478
rect 540804 146476 541404 146478
rect 576804 146476 577404 146478
rect 585320 146476 585920 146478
rect -2916 146454 586840 146476
rect -2916 146218 -1814 146454
rect -1578 146218 986 146454
rect 1222 146218 36986 146454
rect 37222 146218 72986 146454
rect 73222 146218 108986 146454
rect 109222 146218 144986 146454
rect 145222 146218 180986 146454
rect 181222 146218 216986 146454
rect 217222 146218 252986 146454
rect 253222 146218 288986 146454
rect 289222 146218 324986 146454
rect 325222 146218 360986 146454
rect 361222 146218 396986 146454
rect 397222 146218 432986 146454
rect 433222 146218 468986 146454
rect 469222 146218 504986 146454
rect 505222 146218 540986 146454
rect 541222 146218 576986 146454
rect 577222 146218 585502 146454
rect 585738 146218 586840 146454
rect -2916 146134 586840 146218
rect -2916 145898 -1814 146134
rect -1578 145898 986 146134
rect 1222 145898 36986 146134
rect 37222 145898 72986 146134
rect 73222 145898 108986 146134
rect 109222 145898 144986 146134
rect 145222 145898 180986 146134
rect 181222 145898 216986 146134
rect 217222 145898 252986 146134
rect 253222 145898 288986 146134
rect 289222 145898 324986 146134
rect 325222 145898 360986 146134
rect 361222 145898 396986 146134
rect 397222 145898 432986 146134
rect 433222 145898 468986 146134
rect 469222 145898 504986 146134
rect 505222 145898 540986 146134
rect 541222 145898 576986 146134
rect 577222 145898 585502 146134
rect 585738 145898 586840 146134
rect -2916 145876 586840 145898
rect -1996 145874 -1396 145876
rect 804 145874 1404 145876
rect 36804 145874 37404 145876
rect 72804 145874 73404 145876
rect 108804 145874 109404 145876
rect 144804 145874 145404 145876
rect 180804 145874 181404 145876
rect 216804 145874 217404 145876
rect 252804 145874 253404 145876
rect 288804 145874 289404 145876
rect 324804 145874 325404 145876
rect 360804 145874 361404 145876
rect 396804 145874 397404 145876
rect 432804 145874 433404 145876
rect 468804 145874 469404 145876
rect 504804 145874 505404 145876
rect 540804 145874 541404 145876
rect 576804 145874 577404 145876
rect 585320 145874 585920 145876
rect -8436 139276 -7836 139278
rect 29604 139276 30204 139278
rect 65604 139276 66204 139278
rect 101604 139276 102204 139278
rect 137604 139276 138204 139278
rect 173604 139276 174204 139278
rect 209604 139276 210204 139278
rect 245604 139276 246204 139278
rect 281604 139276 282204 139278
rect 317604 139276 318204 139278
rect 353604 139276 354204 139278
rect 389604 139276 390204 139278
rect 425604 139276 426204 139278
rect 461604 139276 462204 139278
rect 497604 139276 498204 139278
rect 533604 139276 534204 139278
rect 569604 139276 570204 139278
rect 591760 139276 592360 139278
rect -8436 139254 592360 139276
rect -8436 139018 -8254 139254
rect -8018 139018 29786 139254
rect 30022 139018 65786 139254
rect 66022 139018 101786 139254
rect 102022 139018 137786 139254
rect 138022 139018 173786 139254
rect 174022 139018 209786 139254
rect 210022 139018 245786 139254
rect 246022 139018 281786 139254
rect 282022 139018 317786 139254
rect 318022 139018 353786 139254
rect 354022 139018 389786 139254
rect 390022 139018 425786 139254
rect 426022 139018 461786 139254
rect 462022 139018 497786 139254
rect 498022 139018 533786 139254
rect 534022 139018 569786 139254
rect 570022 139018 591942 139254
rect 592178 139018 592360 139254
rect -8436 138934 592360 139018
rect -8436 138698 -8254 138934
rect -8018 138698 29786 138934
rect 30022 138698 65786 138934
rect 66022 138698 101786 138934
rect 102022 138698 137786 138934
rect 138022 138698 173786 138934
rect 174022 138698 209786 138934
rect 210022 138698 245786 138934
rect 246022 138698 281786 138934
rect 282022 138698 317786 138934
rect 318022 138698 353786 138934
rect 354022 138698 389786 138934
rect 390022 138698 425786 138934
rect 426022 138698 461786 138934
rect 462022 138698 497786 138934
rect 498022 138698 533786 138934
rect 534022 138698 569786 138934
rect 570022 138698 591942 138934
rect 592178 138698 592360 138934
rect -8436 138676 592360 138698
rect -8436 138674 -7836 138676
rect 29604 138674 30204 138676
rect 65604 138674 66204 138676
rect 101604 138674 102204 138676
rect 137604 138674 138204 138676
rect 173604 138674 174204 138676
rect 209604 138674 210204 138676
rect 245604 138674 246204 138676
rect 281604 138674 282204 138676
rect 317604 138674 318204 138676
rect 353604 138674 354204 138676
rect 389604 138674 390204 138676
rect 425604 138674 426204 138676
rect 461604 138674 462204 138676
rect 497604 138674 498204 138676
rect 533604 138674 534204 138676
rect 569604 138674 570204 138676
rect 591760 138674 592360 138676
rect -6596 135676 -5996 135678
rect 26004 135676 26604 135678
rect 62004 135676 62604 135678
rect 98004 135676 98604 135678
rect 134004 135676 134604 135678
rect 170004 135676 170604 135678
rect 206004 135676 206604 135678
rect 242004 135676 242604 135678
rect 278004 135676 278604 135678
rect 314004 135676 314604 135678
rect 350004 135676 350604 135678
rect 386004 135676 386604 135678
rect 422004 135676 422604 135678
rect 458004 135676 458604 135678
rect 494004 135676 494604 135678
rect 530004 135676 530604 135678
rect 566004 135676 566604 135678
rect 589920 135676 590520 135678
rect -6596 135654 590520 135676
rect -6596 135418 -6414 135654
rect -6178 135418 26186 135654
rect 26422 135418 62186 135654
rect 62422 135418 98186 135654
rect 98422 135418 134186 135654
rect 134422 135418 170186 135654
rect 170422 135418 206186 135654
rect 206422 135418 242186 135654
rect 242422 135418 278186 135654
rect 278422 135418 314186 135654
rect 314422 135418 350186 135654
rect 350422 135418 386186 135654
rect 386422 135418 422186 135654
rect 422422 135418 458186 135654
rect 458422 135418 494186 135654
rect 494422 135418 530186 135654
rect 530422 135418 566186 135654
rect 566422 135418 590102 135654
rect 590338 135418 590520 135654
rect -6596 135334 590520 135418
rect -6596 135098 -6414 135334
rect -6178 135098 26186 135334
rect 26422 135098 62186 135334
rect 62422 135098 98186 135334
rect 98422 135098 134186 135334
rect 134422 135098 170186 135334
rect 170422 135098 206186 135334
rect 206422 135098 242186 135334
rect 242422 135098 278186 135334
rect 278422 135098 314186 135334
rect 314422 135098 350186 135334
rect 350422 135098 386186 135334
rect 386422 135098 422186 135334
rect 422422 135098 458186 135334
rect 458422 135098 494186 135334
rect 494422 135098 530186 135334
rect 530422 135098 566186 135334
rect 566422 135098 590102 135334
rect 590338 135098 590520 135334
rect -6596 135076 590520 135098
rect -6596 135074 -5996 135076
rect 26004 135074 26604 135076
rect 62004 135074 62604 135076
rect 98004 135074 98604 135076
rect 134004 135074 134604 135076
rect 170004 135074 170604 135076
rect 206004 135074 206604 135076
rect 242004 135074 242604 135076
rect 278004 135074 278604 135076
rect 314004 135074 314604 135076
rect 350004 135074 350604 135076
rect 386004 135074 386604 135076
rect 422004 135074 422604 135076
rect 458004 135074 458604 135076
rect 494004 135074 494604 135076
rect 530004 135074 530604 135076
rect 566004 135074 566604 135076
rect 589920 135074 590520 135076
rect -4756 132076 -4156 132078
rect 22404 132076 23004 132078
rect 58404 132076 59004 132078
rect 94404 132076 95004 132078
rect 130404 132076 131004 132078
rect 166404 132076 167004 132078
rect 202404 132076 203004 132078
rect 238404 132076 239004 132078
rect 274404 132076 275004 132078
rect 310404 132076 311004 132078
rect 346404 132076 347004 132078
rect 382404 132076 383004 132078
rect 418404 132076 419004 132078
rect 454404 132076 455004 132078
rect 490404 132076 491004 132078
rect 526404 132076 527004 132078
rect 562404 132076 563004 132078
rect 588080 132076 588680 132078
rect -4756 132054 588680 132076
rect -4756 131818 -4574 132054
rect -4338 131818 22586 132054
rect 22822 131818 58586 132054
rect 58822 131818 94586 132054
rect 94822 131818 130586 132054
rect 130822 131818 166586 132054
rect 166822 131818 202586 132054
rect 202822 131818 238586 132054
rect 238822 131818 274586 132054
rect 274822 131818 310586 132054
rect 310822 131818 346586 132054
rect 346822 131818 382586 132054
rect 382822 131818 418586 132054
rect 418822 131818 454586 132054
rect 454822 131818 490586 132054
rect 490822 131818 526586 132054
rect 526822 131818 562586 132054
rect 562822 131818 588262 132054
rect 588498 131818 588680 132054
rect -4756 131734 588680 131818
rect -4756 131498 -4574 131734
rect -4338 131498 22586 131734
rect 22822 131498 58586 131734
rect 58822 131498 94586 131734
rect 94822 131498 130586 131734
rect 130822 131498 166586 131734
rect 166822 131498 202586 131734
rect 202822 131498 238586 131734
rect 238822 131498 274586 131734
rect 274822 131498 310586 131734
rect 310822 131498 346586 131734
rect 346822 131498 382586 131734
rect 382822 131498 418586 131734
rect 418822 131498 454586 131734
rect 454822 131498 490586 131734
rect 490822 131498 526586 131734
rect 526822 131498 562586 131734
rect 562822 131498 588262 131734
rect 588498 131498 588680 131734
rect -4756 131476 588680 131498
rect -4756 131474 -4156 131476
rect 22404 131474 23004 131476
rect 58404 131474 59004 131476
rect 94404 131474 95004 131476
rect 130404 131474 131004 131476
rect 166404 131474 167004 131476
rect 202404 131474 203004 131476
rect 238404 131474 239004 131476
rect 274404 131474 275004 131476
rect 310404 131474 311004 131476
rect 346404 131474 347004 131476
rect 382404 131474 383004 131476
rect 418404 131474 419004 131476
rect 454404 131474 455004 131476
rect 490404 131474 491004 131476
rect 526404 131474 527004 131476
rect 562404 131474 563004 131476
rect 588080 131474 588680 131476
rect -2916 128476 -2316 128478
rect 18804 128476 19404 128478
rect 54804 128476 55404 128478
rect 90804 128476 91404 128478
rect 126804 128476 127404 128478
rect 162804 128476 163404 128478
rect 198804 128476 199404 128478
rect 234804 128476 235404 128478
rect 270804 128476 271404 128478
rect 306804 128476 307404 128478
rect 342804 128476 343404 128478
rect 378804 128476 379404 128478
rect 414804 128476 415404 128478
rect 450804 128476 451404 128478
rect 486804 128476 487404 128478
rect 522804 128476 523404 128478
rect 558804 128476 559404 128478
rect 586240 128476 586840 128478
rect -2916 128454 586840 128476
rect -2916 128218 -2734 128454
rect -2498 128218 18986 128454
rect 19222 128218 54986 128454
rect 55222 128218 90986 128454
rect 91222 128218 126986 128454
rect 127222 128218 162986 128454
rect 163222 128218 198986 128454
rect 199222 128218 234986 128454
rect 235222 128218 270986 128454
rect 271222 128218 306986 128454
rect 307222 128218 342986 128454
rect 343222 128218 378986 128454
rect 379222 128218 414986 128454
rect 415222 128218 450986 128454
rect 451222 128218 486986 128454
rect 487222 128218 522986 128454
rect 523222 128218 558986 128454
rect 559222 128218 586422 128454
rect 586658 128218 586840 128454
rect -2916 128134 586840 128218
rect -2916 127898 -2734 128134
rect -2498 127898 18986 128134
rect 19222 127898 54986 128134
rect 55222 127898 90986 128134
rect 91222 127898 126986 128134
rect 127222 127898 162986 128134
rect 163222 127898 198986 128134
rect 199222 127898 234986 128134
rect 235222 127898 270986 128134
rect 271222 127898 306986 128134
rect 307222 127898 342986 128134
rect 343222 127898 378986 128134
rect 379222 127898 414986 128134
rect 415222 127898 450986 128134
rect 451222 127898 486986 128134
rect 487222 127898 522986 128134
rect 523222 127898 558986 128134
rect 559222 127898 586422 128134
rect 586658 127898 586840 128134
rect -2916 127876 586840 127898
rect -2916 127874 -2316 127876
rect 18804 127874 19404 127876
rect 54804 127874 55404 127876
rect 90804 127874 91404 127876
rect 126804 127874 127404 127876
rect 162804 127874 163404 127876
rect 198804 127874 199404 127876
rect 234804 127874 235404 127876
rect 270804 127874 271404 127876
rect 306804 127874 307404 127876
rect 342804 127874 343404 127876
rect 378804 127874 379404 127876
rect 414804 127874 415404 127876
rect 450804 127874 451404 127876
rect 486804 127874 487404 127876
rect 522804 127874 523404 127876
rect 558804 127874 559404 127876
rect 586240 127874 586840 127876
rect -7516 121276 -6916 121278
rect 11604 121276 12204 121278
rect 47604 121276 48204 121278
rect 83604 121276 84204 121278
rect 119604 121276 120204 121278
rect 155604 121276 156204 121278
rect 191604 121276 192204 121278
rect 227604 121276 228204 121278
rect 263604 121276 264204 121278
rect 299604 121276 300204 121278
rect 335604 121276 336204 121278
rect 371604 121276 372204 121278
rect 407604 121276 408204 121278
rect 443604 121276 444204 121278
rect 479604 121276 480204 121278
rect 515604 121276 516204 121278
rect 551604 121276 552204 121278
rect 590840 121276 591440 121278
rect -8436 121254 592360 121276
rect -8436 121018 -7334 121254
rect -7098 121018 11786 121254
rect 12022 121018 47786 121254
rect 48022 121018 83786 121254
rect 84022 121018 119786 121254
rect 120022 121018 155786 121254
rect 156022 121018 191786 121254
rect 192022 121018 227786 121254
rect 228022 121018 263786 121254
rect 264022 121018 299786 121254
rect 300022 121018 335786 121254
rect 336022 121018 371786 121254
rect 372022 121018 407786 121254
rect 408022 121018 443786 121254
rect 444022 121018 479786 121254
rect 480022 121018 515786 121254
rect 516022 121018 551786 121254
rect 552022 121018 591022 121254
rect 591258 121018 592360 121254
rect -8436 120934 592360 121018
rect -8436 120698 -7334 120934
rect -7098 120698 11786 120934
rect 12022 120698 47786 120934
rect 48022 120698 83786 120934
rect 84022 120698 119786 120934
rect 120022 120698 155786 120934
rect 156022 120698 191786 120934
rect 192022 120698 227786 120934
rect 228022 120698 263786 120934
rect 264022 120698 299786 120934
rect 300022 120698 335786 120934
rect 336022 120698 371786 120934
rect 372022 120698 407786 120934
rect 408022 120698 443786 120934
rect 444022 120698 479786 120934
rect 480022 120698 515786 120934
rect 516022 120698 551786 120934
rect 552022 120698 591022 120934
rect 591258 120698 592360 120934
rect -8436 120676 592360 120698
rect -7516 120674 -6916 120676
rect 11604 120674 12204 120676
rect 47604 120674 48204 120676
rect 83604 120674 84204 120676
rect 119604 120674 120204 120676
rect 155604 120674 156204 120676
rect 191604 120674 192204 120676
rect 227604 120674 228204 120676
rect 263604 120674 264204 120676
rect 299604 120674 300204 120676
rect 335604 120674 336204 120676
rect 371604 120674 372204 120676
rect 407604 120674 408204 120676
rect 443604 120674 444204 120676
rect 479604 120674 480204 120676
rect 515604 120674 516204 120676
rect 551604 120674 552204 120676
rect 590840 120674 591440 120676
rect -5676 117676 -5076 117678
rect 8004 117676 8604 117678
rect 44004 117676 44604 117678
rect 80004 117676 80604 117678
rect 116004 117676 116604 117678
rect 152004 117676 152604 117678
rect 188004 117676 188604 117678
rect 224004 117676 224604 117678
rect 260004 117676 260604 117678
rect 296004 117676 296604 117678
rect 332004 117676 332604 117678
rect 368004 117676 368604 117678
rect 404004 117676 404604 117678
rect 440004 117676 440604 117678
rect 476004 117676 476604 117678
rect 512004 117676 512604 117678
rect 548004 117676 548604 117678
rect 589000 117676 589600 117678
rect -6596 117654 590520 117676
rect -6596 117418 -5494 117654
rect -5258 117418 8186 117654
rect 8422 117418 44186 117654
rect 44422 117418 80186 117654
rect 80422 117418 116186 117654
rect 116422 117418 152186 117654
rect 152422 117418 188186 117654
rect 188422 117418 224186 117654
rect 224422 117418 260186 117654
rect 260422 117418 296186 117654
rect 296422 117418 332186 117654
rect 332422 117418 368186 117654
rect 368422 117418 404186 117654
rect 404422 117418 440186 117654
rect 440422 117418 476186 117654
rect 476422 117418 512186 117654
rect 512422 117418 548186 117654
rect 548422 117418 589182 117654
rect 589418 117418 590520 117654
rect -6596 117334 590520 117418
rect -6596 117098 -5494 117334
rect -5258 117098 8186 117334
rect 8422 117098 44186 117334
rect 44422 117098 80186 117334
rect 80422 117098 116186 117334
rect 116422 117098 152186 117334
rect 152422 117098 188186 117334
rect 188422 117098 224186 117334
rect 224422 117098 260186 117334
rect 260422 117098 296186 117334
rect 296422 117098 332186 117334
rect 332422 117098 368186 117334
rect 368422 117098 404186 117334
rect 404422 117098 440186 117334
rect 440422 117098 476186 117334
rect 476422 117098 512186 117334
rect 512422 117098 548186 117334
rect 548422 117098 589182 117334
rect 589418 117098 590520 117334
rect -6596 117076 590520 117098
rect -5676 117074 -5076 117076
rect 8004 117074 8604 117076
rect 44004 117074 44604 117076
rect 80004 117074 80604 117076
rect 116004 117074 116604 117076
rect 152004 117074 152604 117076
rect 188004 117074 188604 117076
rect 224004 117074 224604 117076
rect 260004 117074 260604 117076
rect 296004 117074 296604 117076
rect 332004 117074 332604 117076
rect 368004 117074 368604 117076
rect 404004 117074 404604 117076
rect 440004 117074 440604 117076
rect 476004 117074 476604 117076
rect 512004 117074 512604 117076
rect 548004 117074 548604 117076
rect 589000 117074 589600 117076
rect -3836 114076 -3236 114078
rect 4404 114076 5004 114078
rect 40404 114076 41004 114078
rect 76404 114076 77004 114078
rect 112404 114076 113004 114078
rect 148404 114076 149004 114078
rect 184404 114076 185004 114078
rect 220404 114076 221004 114078
rect 256404 114076 257004 114078
rect 292404 114076 293004 114078
rect 328404 114076 329004 114078
rect 364404 114076 365004 114078
rect 400404 114076 401004 114078
rect 436404 114076 437004 114078
rect 472404 114076 473004 114078
rect 508404 114076 509004 114078
rect 544404 114076 545004 114078
rect 580404 114076 581004 114078
rect 587160 114076 587760 114078
rect -4756 114054 588680 114076
rect -4756 113818 -3654 114054
rect -3418 113818 4586 114054
rect 4822 113818 40586 114054
rect 40822 113818 76586 114054
rect 76822 113818 112586 114054
rect 112822 113818 148586 114054
rect 148822 113818 184586 114054
rect 184822 113818 220586 114054
rect 220822 113818 256586 114054
rect 256822 113818 292586 114054
rect 292822 113818 328586 114054
rect 328822 113818 364586 114054
rect 364822 113818 400586 114054
rect 400822 113818 436586 114054
rect 436822 113818 472586 114054
rect 472822 113818 508586 114054
rect 508822 113818 544586 114054
rect 544822 113818 580586 114054
rect 580822 113818 587342 114054
rect 587578 113818 588680 114054
rect -4756 113734 588680 113818
rect -4756 113498 -3654 113734
rect -3418 113498 4586 113734
rect 4822 113498 40586 113734
rect 40822 113498 76586 113734
rect 76822 113498 112586 113734
rect 112822 113498 148586 113734
rect 148822 113498 184586 113734
rect 184822 113498 220586 113734
rect 220822 113498 256586 113734
rect 256822 113498 292586 113734
rect 292822 113498 328586 113734
rect 328822 113498 364586 113734
rect 364822 113498 400586 113734
rect 400822 113498 436586 113734
rect 436822 113498 472586 113734
rect 472822 113498 508586 113734
rect 508822 113498 544586 113734
rect 544822 113498 580586 113734
rect 580822 113498 587342 113734
rect 587578 113498 588680 113734
rect -4756 113476 588680 113498
rect -3836 113474 -3236 113476
rect 4404 113474 5004 113476
rect 40404 113474 41004 113476
rect 76404 113474 77004 113476
rect 112404 113474 113004 113476
rect 148404 113474 149004 113476
rect 184404 113474 185004 113476
rect 220404 113474 221004 113476
rect 256404 113474 257004 113476
rect 292404 113474 293004 113476
rect 328404 113474 329004 113476
rect 364404 113474 365004 113476
rect 400404 113474 401004 113476
rect 436404 113474 437004 113476
rect 472404 113474 473004 113476
rect 508404 113474 509004 113476
rect 544404 113474 545004 113476
rect 580404 113474 581004 113476
rect 587160 113474 587760 113476
rect -1996 110476 -1396 110478
rect 804 110476 1404 110478
rect 36804 110476 37404 110478
rect 72804 110476 73404 110478
rect 108804 110476 109404 110478
rect 144804 110476 145404 110478
rect 180804 110476 181404 110478
rect 216804 110476 217404 110478
rect 252804 110476 253404 110478
rect 288804 110476 289404 110478
rect 324804 110476 325404 110478
rect 360804 110476 361404 110478
rect 396804 110476 397404 110478
rect 432804 110476 433404 110478
rect 468804 110476 469404 110478
rect 504804 110476 505404 110478
rect 540804 110476 541404 110478
rect 576804 110476 577404 110478
rect 585320 110476 585920 110478
rect -2916 110454 586840 110476
rect -2916 110218 -1814 110454
rect -1578 110218 986 110454
rect 1222 110218 36986 110454
rect 37222 110218 72986 110454
rect 73222 110218 108986 110454
rect 109222 110218 144986 110454
rect 145222 110218 180986 110454
rect 181222 110218 216986 110454
rect 217222 110218 252986 110454
rect 253222 110218 288986 110454
rect 289222 110218 324986 110454
rect 325222 110218 360986 110454
rect 361222 110218 396986 110454
rect 397222 110218 432986 110454
rect 433222 110218 468986 110454
rect 469222 110218 504986 110454
rect 505222 110218 540986 110454
rect 541222 110218 576986 110454
rect 577222 110218 585502 110454
rect 585738 110218 586840 110454
rect -2916 110134 586840 110218
rect -2916 109898 -1814 110134
rect -1578 109898 986 110134
rect 1222 109898 36986 110134
rect 37222 109898 72986 110134
rect 73222 109898 108986 110134
rect 109222 109898 144986 110134
rect 145222 109898 180986 110134
rect 181222 109898 216986 110134
rect 217222 109898 252986 110134
rect 253222 109898 288986 110134
rect 289222 109898 324986 110134
rect 325222 109898 360986 110134
rect 361222 109898 396986 110134
rect 397222 109898 432986 110134
rect 433222 109898 468986 110134
rect 469222 109898 504986 110134
rect 505222 109898 540986 110134
rect 541222 109898 576986 110134
rect 577222 109898 585502 110134
rect 585738 109898 586840 110134
rect -2916 109876 586840 109898
rect -1996 109874 -1396 109876
rect 804 109874 1404 109876
rect 36804 109874 37404 109876
rect 72804 109874 73404 109876
rect 108804 109874 109404 109876
rect 144804 109874 145404 109876
rect 180804 109874 181404 109876
rect 216804 109874 217404 109876
rect 252804 109874 253404 109876
rect 288804 109874 289404 109876
rect 324804 109874 325404 109876
rect 360804 109874 361404 109876
rect 396804 109874 397404 109876
rect 432804 109874 433404 109876
rect 468804 109874 469404 109876
rect 504804 109874 505404 109876
rect 540804 109874 541404 109876
rect 576804 109874 577404 109876
rect 585320 109874 585920 109876
rect -8436 103276 -7836 103278
rect 29604 103276 30204 103278
rect 65604 103276 66204 103278
rect 101604 103276 102204 103278
rect 137604 103276 138204 103278
rect 173604 103276 174204 103278
rect 209604 103276 210204 103278
rect 245604 103276 246204 103278
rect 281604 103276 282204 103278
rect 317604 103276 318204 103278
rect 353604 103276 354204 103278
rect 389604 103276 390204 103278
rect 425604 103276 426204 103278
rect 461604 103276 462204 103278
rect 497604 103276 498204 103278
rect 533604 103276 534204 103278
rect 569604 103276 570204 103278
rect 591760 103276 592360 103278
rect -8436 103254 592360 103276
rect -8436 103018 -8254 103254
rect -8018 103018 29786 103254
rect 30022 103018 65786 103254
rect 66022 103018 101786 103254
rect 102022 103018 137786 103254
rect 138022 103018 173786 103254
rect 174022 103018 209786 103254
rect 210022 103018 245786 103254
rect 246022 103018 281786 103254
rect 282022 103018 317786 103254
rect 318022 103018 353786 103254
rect 354022 103018 389786 103254
rect 390022 103018 425786 103254
rect 426022 103018 461786 103254
rect 462022 103018 497786 103254
rect 498022 103018 533786 103254
rect 534022 103018 569786 103254
rect 570022 103018 591942 103254
rect 592178 103018 592360 103254
rect -8436 102934 592360 103018
rect -8436 102698 -8254 102934
rect -8018 102698 29786 102934
rect 30022 102698 65786 102934
rect 66022 102698 101786 102934
rect 102022 102698 137786 102934
rect 138022 102698 173786 102934
rect 174022 102698 209786 102934
rect 210022 102698 245786 102934
rect 246022 102698 281786 102934
rect 282022 102698 317786 102934
rect 318022 102698 353786 102934
rect 354022 102698 389786 102934
rect 390022 102698 425786 102934
rect 426022 102698 461786 102934
rect 462022 102698 497786 102934
rect 498022 102698 533786 102934
rect 534022 102698 569786 102934
rect 570022 102698 591942 102934
rect 592178 102698 592360 102934
rect -8436 102676 592360 102698
rect -8436 102674 -7836 102676
rect 29604 102674 30204 102676
rect 65604 102674 66204 102676
rect 101604 102674 102204 102676
rect 137604 102674 138204 102676
rect 173604 102674 174204 102676
rect 209604 102674 210204 102676
rect 245604 102674 246204 102676
rect 281604 102674 282204 102676
rect 317604 102674 318204 102676
rect 353604 102674 354204 102676
rect 389604 102674 390204 102676
rect 425604 102674 426204 102676
rect 461604 102674 462204 102676
rect 497604 102674 498204 102676
rect 533604 102674 534204 102676
rect 569604 102674 570204 102676
rect 591760 102674 592360 102676
rect -6596 99676 -5996 99678
rect 26004 99676 26604 99678
rect 62004 99676 62604 99678
rect 98004 99676 98604 99678
rect 134004 99676 134604 99678
rect 170004 99676 170604 99678
rect 206004 99676 206604 99678
rect 242004 99676 242604 99678
rect 278004 99676 278604 99678
rect 314004 99676 314604 99678
rect 350004 99676 350604 99678
rect 386004 99676 386604 99678
rect 422004 99676 422604 99678
rect 458004 99676 458604 99678
rect 494004 99676 494604 99678
rect 530004 99676 530604 99678
rect 566004 99676 566604 99678
rect 589920 99676 590520 99678
rect -6596 99654 590520 99676
rect -6596 99418 -6414 99654
rect -6178 99418 26186 99654
rect 26422 99418 62186 99654
rect 62422 99418 98186 99654
rect 98422 99418 134186 99654
rect 134422 99418 170186 99654
rect 170422 99418 206186 99654
rect 206422 99418 242186 99654
rect 242422 99418 278186 99654
rect 278422 99418 314186 99654
rect 314422 99418 350186 99654
rect 350422 99418 386186 99654
rect 386422 99418 422186 99654
rect 422422 99418 458186 99654
rect 458422 99418 494186 99654
rect 494422 99418 530186 99654
rect 530422 99418 566186 99654
rect 566422 99418 590102 99654
rect 590338 99418 590520 99654
rect -6596 99334 590520 99418
rect -6596 99098 -6414 99334
rect -6178 99098 26186 99334
rect 26422 99098 62186 99334
rect 62422 99098 98186 99334
rect 98422 99098 134186 99334
rect 134422 99098 170186 99334
rect 170422 99098 206186 99334
rect 206422 99098 242186 99334
rect 242422 99098 278186 99334
rect 278422 99098 314186 99334
rect 314422 99098 350186 99334
rect 350422 99098 386186 99334
rect 386422 99098 422186 99334
rect 422422 99098 458186 99334
rect 458422 99098 494186 99334
rect 494422 99098 530186 99334
rect 530422 99098 566186 99334
rect 566422 99098 590102 99334
rect 590338 99098 590520 99334
rect -6596 99076 590520 99098
rect -6596 99074 -5996 99076
rect 26004 99074 26604 99076
rect 62004 99074 62604 99076
rect 98004 99074 98604 99076
rect 134004 99074 134604 99076
rect 170004 99074 170604 99076
rect 206004 99074 206604 99076
rect 242004 99074 242604 99076
rect 278004 99074 278604 99076
rect 314004 99074 314604 99076
rect 350004 99074 350604 99076
rect 386004 99074 386604 99076
rect 422004 99074 422604 99076
rect 458004 99074 458604 99076
rect 494004 99074 494604 99076
rect 530004 99074 530604 99076
rect 566004 99074 566604 99076
rect 589920 99074 590520 99076
rect -4756 96076 -4156 96078
rect 22404 96076 23004 96078
rect 58404 96076 59004 96078
rect 94404 96076 95004 96078
rect 130404 96076 131004 96078
rect 166404 96076 167004 96078
rect 202404 96076 203004 96078
rect 238404 96076 239004 96078
rect 274404 96076 275004 96078
rect 310404 96076 311004 96078
rect 346404 96076 347004 96078
rect 382404 96076 383004 96078
rect 418404 96076 419004 96078
rect 454404 96076 455004 96078
rect 490404 96076 491004 96078
rect 526404 96076 527004 96078
rect 562404 96076 563004 96078
rect 588080 96076 588680 96078
rect -4756 96054 588680 96076
rect -4756 95818 -4574 96054
rect -4338 95818 22586 96054
rect 22822 95818 58586 96054
rect 58822 95818 94586 96054
rect 94822 95818 130586 96054
rect 130822 95818 166586 96054
rect 166822 95818 202586 96054
rect 202822 95818 238586 96054
rect 238822 95818 274586 96054
rect 274822 95818 310586 96054
rect 310822 95818 346586 96054
rect 346822 95818 382586 96054
rect 382822 95818 418586 96054
rect 418822 95818 454586 96054
rect 454822 95818 490586 96054
rect 490822 95818 526586 96054
rect 526822 95818 562586 96054
rect 562822 95818 588262 96054
rect 588498 95818 588680 96054
rect -4756 95734 588680 95818
rect -4756 95498 -4574 95734
rect -4338 95498 22586 95734
rect 22822 95498 58586 95734
rect 58822 95498 94586 95734
rect 94822 95498 130586 95734
rect 130822 95498 166586 95734
rect 166822 95498 202586 95734
rect 202822 95498 238586 95734
rect 238822 95498 274586 95734
rect 274822 95498 310586 95734
rect 310822 95498 346586 95734
rect 346822 95498 382586 95734
rect 382822 95498 418586 95734
rect 418822 95498 454586 95734
rect 454822 95498 490586 95734
rect 490822 95498 526586 95734
rect 526822 95498 562586 95734
rect 562822 95498 588262 95734
rect 588498 95498 588680 95734
rect -4756 95476 588680 95498
rect -4756 95474 -4156 95476
rect 22404 95474 23004 95476
rect 58404 95474 59004 95476
rect 94404 95474 95004 95476
rect 130404 95474 131004 95476
rect 166404 95474 167004 95476
rect 202404 95474 203004 95476
rect 238404 95474 239004 95476
rect 274404 95474 275004 95476
rect 310404 95474 311004 95476
rect 346404 95474 347004 95476
rect 382404 95474 383004 95476
rect 418404 95474 419004 95476
rect 454404 95474 455004 95476
rect 490404 95474 491004 95476
rect 526404 95474 527004 95476
rect 562404 95474 563004 95476
rect 588080 95474 588680 95476
rect -2916 92476 -2316 92478
rect 18804 92476 19404 92478
rect 54804 92476 55404 92478
rect 90804 92476 91404 92478
rect 126804 92476 127404 92478
rect 162804 92476 163404 92478
rect 198804 92476 199404 92478
rect 234804 92476 235404 92478
rect 270804 92476 271404 92478
rect 306804 92476 307404 92478
rect 342804 92476 343404 92478
rect 378804 92476 379404 92478
rect 414804 92476 415404 92478
rect 450804 92476 451404 92478
rect 486804 92476 487404 92478
rect 522804 92476 523404 92478
rect 558804 92476 559404 92478
rect 586240 92476 586840 92478
rect -2916 92454 586840 92476
rect -2916 92218 -2734 92454
rect -2498 92218 18986 92454
rect 19222 92218 54986 92454
rect 55222 92218 90986 92454
rect 91222 92218 126986 92454
rect 127222 92218 162986 92454
rect 163222 92218 198986 92454
rect 199222 92218 234986 92454
rect 235222 92218 270986 92454
rect 271222 92218 306986 92454
rect 307222 92218 342986 92454
rect 343222 92218 378986 92454
rect 379222 92218 414986 92454
rect 415222 92218 450986 92454
rect 451222 92218 486986 92454
rect 487222 92218 522986 92454
rect 523222 92218 558986 92454
rect 559222 92218 586422 92454
rect 586658 92218 586840 92454
rect -2916 92134 586840 92218
rect -2916 91898 -2734 92134
rect -2498 91898 18986 92134
rect 19222 91898 54986 92134
rect 55222 91898 90986 92134
rect 91222 91898 126986 92134
rect 127222 91898 162986 92134
rect 163222 91898 198986 92134
rect 199222 91898 234986 92134
rect 235222 91898 270986 92134
rect 271222 91898 306986 92134
rect 307222 91898 342986 92134
rect 343222 91898 378986 92134
rect 379222 91898 414986 92134
rect 415222 91898 450986 92134
rect 451222 91898 486986 92134
rect 487222 91898 522986 92134
rect 523222 91898 558986 92134
rect 559222 91898 586422 92134
rect 586658 91898 586840 92134
rect -2916 91876 586840 91898
rect -2916 91874 -2316 91876
rect 18804 91874 19404 91876
rect 54804 91874 55404 91876
rect 90804 91874 91404 91876
rect 126804 91874 127404 91876
rect 162804 91874 163404 91876
rect 198804 91874 199404 91876
rect 234804 91874 235404 91876
rect 270804 91874 271404 91876
rect 306804 91874 307404 91876
rect 342804 91874 343404 91876
rect 378804 91874 379404 91876
rect 414804 91874 415404 91876
rect 450804 91874 451404 91876
rect 486804 91874 487404 91876
rect 522804 91874 523404 91876
rect 558804 91874 559404 91876
rect 586240 91874 586840 91876
rect -7516 85276 -6916 85278
rect 11604 85276 12204 85278
rect 47604 85276 48204 85278
rect 83604 85276 84204 85278
rect 119604 85276 120204 85278
rect 155604 85276 156204 85278
rect 191604 85276 192204 85278
rect 227604 85276 228204 85278
rect 263604 85276 264204 85278
rect 299604 85276 300204 85278
rect 335604 85276 336204 85278
rect 371604 85276 372204 85278
rect 407604 85276 408204 85278
rect 443604 85276 444204 85278
rect 479604 85276 480204 85278
rect 515604 85276 516204 85278
rect 551604 85276 552204 85278
rect 590840 85276 591440 85278
rect -8436 85254 592360 85276
rect -8436 85018 -7334 85254
rect -7098 85018 11786 85254
rect 12022 85018 47786 85254
rect 48022 85018 83786 85254
rect 84022 85018 119786 85254
rect 120022 85018 155786 85254
rect 156022 85018 191786 85254
rect 192022 85018 227786 85254
rect 228022 85018 263786 85254
rect 264022 85018 299786 85254
rect 300022 85018 335786 85254
rect 336022 85018 371786 85254
rect 372022 85018 407786 85254
rect 408022 85018 443786 85254
rect 444022 85018 479786 85254
rect 480022 85018 515786 85254
rect 516022 85018 551786 85254
rect 552022 85018 591022 85254
rect 591258 85018 592360 85254
rect -8436 84934 592360 85018
rect -8436 84698 -7334 84934
rect -7098 84698 11786 84934
rect 12022 84698 47786 84934
rect 48022 84698 83786 84934
rect 84022 84698 119786 84934
rect 120022 84698 155786 84934
rect 156022 84698 191786 84934
rect 192022 84698 227786 84934
rect 228022 84698 263786 84934
rect 264022 84698 299786 84934
rect 300022 84698 335786 84934
rect 336022 84698 371786 84934
rect 372022 84698 407786 84934
rect 408022 84698 443786 84934
rect 444022 84698 479786 84934
rect 480022 84698 515786 84934
rect 516022 84698 551786 84934
rect 552022 84698 591022 84934
rect 591258 84698 592360 84934
rect -8436 84676 592360 84698
rect -7516 84674 -6916 84676
rect 11604 84674 12204 84676
rect 47604 84674 48204 84676
rect 83604 84674 84204 84676
rect 119604 84674 120204 84676
rect 155604 84674 156204 84676
rect 191604 84674 192204 84676
rect 227604 84674 228204 84676
rect 263604 84674 264204 84676
rect 299604 84674 300204 84676
rect 335604 84674 336204 84676
rect 371604 84674 372204 84676
rect 407604 84674 408204 84676
rect 443604 84674 444204 84676
rect 479604 84674 480204 84676
rect 515604 84674 516204 84676
rect 551604 84674 552204 84676
rect 590840 84674 591440 84676
rect -5676 81676 -5076 81678
rect 8004 81676 8604 81678
rect 44004 81676 44604 81678
rect 80004 81676 80604 81678
rect 116004 81676 116604 81678
rect 152004 81676 152604 81678
rect 188004 81676 188604 81678
rect 224004 81676 224604 81678
rect 260004 81676 260604 81678
rect 296004 81676 296604 81678
rect 332004 81676 332604 81678
rect 368004 81676 368604 81678
rect 404004 81676 404604 81678
rect 440004 81676 440604 81678
rect 476004 81676 476604 81678
rect 512004 81676 512604 81678
rect 548004 81676 548604 81678
rect 589000 81676 589600 81678
rect -6596 81654 590520 81676
rect -6596 81418 -5494 81654
rect -5258 81418 8186 81654
rect 8422 81418 44186 81654
rect 44422 81418 80186 81654
rect 80422 81418 116186 81654
rect 116422 81418 152186 81654
rect 152422 81418 188186 81654
rect 188422 81418 224186 81654
rect 224422 81418 260186 81654
rect 260422 81418 296186 81654
rect 296422 81418 332186 81654
rect 332422 81418 368186 81654
rect 368422 81418 404186 81654
rect 404422 81418 440186 81654
rect 440422 81418 476186 81654
rect 476422 81418 512186 81654
rect 512422 81418 548186 81654
rect 548422 81418 589182 81654
rect 589418 81418 590520 81654
rect -6596 81334 590520 81418
rect -6596 81098 -5494 81334
rect -5258 81098 8186 81334
rect 8422 81098 44186 81334
rect 44422 81098 80186 81334
rect 80422 81098 116186 81334
rect 116422 81098 152186 81334
rect 152422 81098 188186 81334
rect 188422 81098 224186 81334
rect 224422 81098 260186 81334
rect 260422 81098 296186 81334
rect 296422 81098 332186 81334
rect 332422 81098 368186 81334
rect 368422 81098 404186 81334
rect 404422 81098 440186 81334
rect 440422 81098 476186 81334
rect 476422 81098 512186 81334
rect 512422 81098 548186 81334
rect 548422 81098 589182 81334
rect 589418 81098 590520 81334
rect -6596 81076 590520 81098
rect -5676 81074 -5076 81076
rect 8004 81074 8604 81076
rect 44004 81074 44604 81076
rect 80004 81074 80604 81076
rect 116004 81074 116604 81076
rect 152004 81074 152604 81076
rect 188004 81074 188604 81076
rect 224004 81074 224604 81076
rect 260004 81074 260604 81076
rect 296004 81074 296604 81076
rect 332004 81074 332604 81076
rect 368004 81074 368604 81076
rect 404004 81074 404604 81076
rect 440004 81074 440604 81076
rect 476004 81074 476604 81076
rect 512004 81074 512604 81076
rect 548004 81074 548604 81076
rect 589000 81074 589600 81076
rect -3836 78076 -3236 78078
rect 4404 78076 5004 78078
rect 40404 78076 41004 78078
rect 76404 78076 77004 78078
rect 112404 78076 113004 78078
rect 148404 78076 149004 78078
rect 184404 78076 185004 78078
rect 220404 78076 221004 78078
rect 256404 78076 257004 78078
rect 292404 78076 293004 78078
rect 328404 78076 329004 78078
rect 364404 78076 365004 78078
rect 400404 78076 401004 78078
rect 436404 78076 437004 78078
rect 472404 78076 473004 78078
rect 508404 78076 509004 78078
rect 544404 78076 545004 78078
rect 580404 78076 581004 78078
rect 587160 78076 587760 78078
rect -4756 78054 588680 78076
rect -4756 77818 -3654 78054
rect -3418 77818 4586 78054
rect 4822 77818 40586 78054
rect 40822 77818 76586 78054
rect 76822 77818 112586 78054
rect 112822 77818 148586 78054
rect 148822 77818 184586 78054
rect 184822 77818 220586 78054
rect 220822 77818 256586 78054
rect 256822 77818 292586 78054
rect 292822 77818 328586 78054
rect 328822 77818 364586 78054
rect 364822 77818 400586 78054
rect 400822 77818 436586 78054
rect 436822 77818 472586 78054
rect 472822 77818 508586 78054
rect 508822 77818 544586 78054
rect 544822 77818 580586 78054
rect 580822 77818 587342 78054
rect 587578 77818 588680 78054
rect -4756 77734 588680 77818
rect -4756 77498 -3654 77734
rect -3418 77498 4586 77734
rect 4822 77498 40586 77734
rect 40822 77498 76586 77734
rect 76822 77498 112586 77734
rect 112822 77498 148586 77734
rect 148822 77498 184586 77734
rect 184822 77498 220586 77734
rect 220822 77498 256586 77734
rect 256822 77498 292586 77734
rect 292822 77498 328586 77734
rect 328822 77498 364586 77734
rect 364822 77498 400586 77734
rect 400822 77498 436586 77734
rect 436822 77498 472586 77734
rect 472822 77498 508586 77734
rect 508822 77498 544586 77734
rect 544822 77498 580586 77734
rect 580822 77498 587342 77734
rect 587578 77498 588680 77734
rect -4756 77476 588680 77498
rect -3836 77474 -3236 77476
rect 4404 77474 5004 77476
rect 40404 77474 41004 77476
rect 76404 77474 77004 77476
rect 112404 77474 113004 77476
rect 148404 77474 149004 77476
rect 184404 77474 185004 77476
rect 220404 77474 221004 77476
rect 256404 77474 257004 77476
rect 292404 77474 293004 77476
rect 328404 77474 329004 77476
rect 364404 77474 365004 77476
rect 400404 77474 401004 77476
rect 436404 77474 437004 77476
rect 472404 77474 473004 77476
rect 508404 77474 509004 77476
rect 544404 77474 545004 77476
rect 580404 77474 581004 77476
rect 587160 77474 587760 77476
rect -1996 74476 -1396 74478
rect 804 74476 1404 74478
rect 36804 74476 37404 74478
rect 72804 74476 73404 74478
rect 108804 74476 109404 74478
rect 144804 74476 145404 74478
rect 180804 74476 181404 74478
rect 216804 74476 217404 74478
rect 252804 74476 253404 74478
rect 288804 74476 289404 74478
rect 324804 74476 325404 74478
rect 360804 74476 361404 74478
rect 396804 74476 397404 74478
rect 432804 74476 433404 74478
rect 468804 74476 469404 74478
rect 504804 74476 505404 74478
rect 540804 74476 541404 74478
rect 576804 74476 577404 74478
rect 585320 74476 585920 74478
rect -2916 74454 586840 74476
rect -2916 74218 -1814 74454
rect -1578 74218 986 74454
rect 1222 74218 36986 74454
rect 37222 74218 72986 74454
rect 73222 74218 108986 74454
rect 109222 74218 144986 74454
rect 145222 74218 180986 74454
rect 181222 74218 216986 74454
rect 217222 74218 252986 74454
rect 253222 74218 288986 74454
rect 289222 74218 324986 74454
rect 325222 74218 360986 74454
rect 361222 74218 396986 74454
rect 397222 74218 432986 74454
rect 433222 74218 468986 74454
rect 469222 74218 504986 74454
rect 505222 74218 540986 74454
rect 541222 74218 576986 74454
rect 577222 74218 585502 74454
rect 585738 74218 586840 74454
rect -2916 74134 586840 74218
rect -2916 73898 -1814 74134
rect -1578 73898 986 74134
rect 1222 73898 36986 74134
rect 37222 73898 72986 74134
rect 73222 73898 108986 74134
rect 109222 73898 144986 74134
rect 145222 73898 180986 74134
rect 181222 73898 216986 74134
rect 217222 73898 252986 74134
rect 253222 73898 288986 74134
rect 289222 73898 324986 74134
rect 325222 73898 360986 74134
rect 361222 73898 396986 74134
rect 397222 73898 432986 74134
rect 433222 73898 468986 74134
rect 469222 73898 504986 74134
rect 505222 73898 540986 74134
rect 541222 73898 576986 74134
rect 577222 73898 585502 74134
rect 585738 73898 586840 74134
rect -2916 73876 586840 73898
rect -1996 73874 -1396 73876
rect 804 73874 1404 73876
rect 36804 73874 37404 73876
rect 72804 73874 73404 73876
rect 108804 73874 109404 73876
rect 144804 73874 145404 73876
rect 180804 73874 181404 73876
rect 216804 73874 217404 73876
rect 252804 73874 253404 73876
rect 288804 73874 289404 73876
rect 324804 73874 325404 73876
rect 360804 73874 361404 73876
rect 396804 73874 397404 73876
rect 432804 73874 433404 73876
rect 468804 73874 469404 73876
rect 504804 73874 505404 73876
rect 540804 73874 541404 73876
rect 576804 73874 577404 73876
rect 585320 73874 585920 73876
rect -8436 67276 -7836 67278
rect 29604 67276 30204 67278
rect 65604 67276 66204 67278
rect 101604 67276 102204 67278
rect 137604 67276 138204 67278
rect 173604 67276 174204 67278
rect 209604 67276 210204 67278
rect 245604 67276 246204 67278
rect 281604 67276 282204 67278
rect 317604 67276 318204 67278
rect 353604 67276 354204 67278
rect 389604 67276 390204 67278
rect 425604 67276 426204 67278
rect 461604 67276 462204 67278
rect 497604 67276 498204 67278
rect 533604 67276 534204 67278
rect 569604 67276 570204 67278
rect 591760 67276 592360 67278
rect -8436 67254 592360 67276
rect -8436 67018 -8254 67254
rect -8018 67018 29786 67254
rect 30022 67018 65786 67254
rect 66022 67018 101786 67254
rect 102022 67018 137786 67254
rect 138022 67018 173786 67254
rect 174022 67018 209786 67254
rect 210022 67018 245786 67254
rect 246022 67018 281786 67254
rect 282022 67018 317786 67254
rect 318022 67018 353786 67254
rect 354022 67018 389786 67254
rect 390022 67018 425786 67254
rect 426022 67018 461786 67254
rect 462022 67018 497786 67254
rect 498022 67018 533786 67254
rect 534022 67018 569786 67254
rect 570022 67018 591942 67254
rect 592178 67018 592360 67254
rect -8436 66934 592360 67018
rect -8436 66698 -8254 66934
rect -8018 66698 29786 66934
rect 30022 66698 65786 66934
rect 66022 66698 101786 66934
rect 102022 66698 137786 66934
rect 138022 66698 173786 66934
rect 174022 66698 209786 66934
rect 210022 66698 245786 66934
rect 246022 66698 281786 66934
rect 282022 66698 317786 66934
rect 318022 66698 353786 66934
rect 354022 66698 389786 66934
rect 390022 66698 425786 66934
rect 426022 66698 461786 66934
rect 462022 66698 497786 66934
rect 498022 66698 533786 66934
rect 534022 66698 569786 66934
rect 570022 66698 591942 66934
rect 592178 66698 592360 66934
rect -8436 66676 592360 66698
rect -8436 66674 -7836 66676
rect 29604 66674 30204 66676
rect 65604 66674 66204 66676
rect 101604 66674 102204 66676
rect 137604 66674 138204 66676
rect 173604 66674 174204 66676
rect 209604 66674 210204 66676
rect 245604 66674 246204 66676
rect 281604 66674 282204 66676
rect 317604 66674 318204 66676
rect 353604 66674 354204 66676
rect 389604 66674 390204 66676
rect 425604 66674 426204 66676
rect 461604 66674 462204 66676
rect 497604 66674 498204 66676
rect 533604 66674 534204 66676
rect 569604 66674 570204 66676
rect 591760 66674 592360 66676
rect -6596 63676 -5996 63678
rect 26004 63676 26604 63678
rect 62004 63676 62604 63678
rect 98004 63676 98604 63678
rect 134004 63676 134604 63678
rect 170004 63676 170604 63678
rect 206004 63676 206604 63678
rect 242004 63676 242604 63678
rect 278004 63676 278604 63678
rect 314004 63676 314604 63678
rect 350004 63676 350604 63678
rect 386004 63676 386604 63678
rect 422004 63676 422604 63678
rect 458004 63676 458604 63678
rect 494004 63676 494604 63678
rect 530004 63676 530604 63678
rect 566004 63676 566604 63678
rect 589920 63676 590520 63678
rect -6596 63654 590520 63676
rect -6596 63418 -6414 63654
rect -6178 63418 26186 63654
rect 26422 63418 62186 63654
rect 62422 63418 98186 63654
rect 98422 63418 134186 63654
rect 134422 63418 170186 63654
rect 170422 63418 206186 63654
rect 206422 63418 242186 63654
rect 242422 63418 278186 63654
rect 278422 63418 314186 63654
rect 314422 63418 350186 63654
rect 350422 63418 386186 63654
rect 386422 63418 422186 63654
rect 422422 63418 458186 63654
rect 458422 63418 494186 63654
rect 494422 63418 530186 63654
rect 530422 63418 566186 63654
rect 566422 63418 590102 63654
rect 590338 63418 590520 63654
rect -6596 63334 590520 63418
rect -6596 63098 -6414 63334
rect -6178 63098 26186 63334
rect 26422 63098 62186 63334
rect 62422 63098 98186 63334
rect 98422 63098 134186 63334
rect 134422 63098 170186 63334
rect 170422 63098 206186 63334
rect 206422 63098 242186 63334
rect 242422 63098 278186 63334
rect 278422 63098 314186 63334
rect 314422 63098 350186 63334
rect 350422 63098 386186 63334
rect 386422 63098 422186 63334
rect 422422 63098 458186 63334
rect 458422 63098 494186 63334
rect 494422 63098 530186 63334
rect 530422 63098 566186 63334
rect 566422 63098 590102 63334
rect 590338 63098 590520 63334
rect -6596 63076 590520 63098
rect -6596 63074 -5996 63076
rect 26004 63074 26604 63076
rect 62004 63074 62604 63076
rect 98004 63074 98604 63076
rect 134004 63074 134604 63076
rect 170004 63074 170604 63076
rect 206004 63074 206604 63076
rect 242004 63074 242604 63076
rect 278004 63074 278604 63076
rect 314004 63074 314604 63076
rect 350004 63074 350604 63076
rect 386004 63074 386604 63076
rect 422004 63074 422604 63076
rect 458004 63074 458604 63076
rect 494004 63074 494604 63076
rect 530004 63074 530604 63076
rect 566004 63074 566604 63076
rect 589920 63074 590520 63076
rect -4756 60076 -4156 60078
rect 22404 60076 23004 60078
rect 58404 60076 59004 60078
rect 94404 60076 95004 60078
rect 130404 60076 131004 60078
rect 166404 60076 167004 60078
rect 202404 60076 203004 60078
rect 238404 60076 239004 60078
rect 274404 60076 275004 60078
rect 310404 60076 311004 60078
rect 346404 60076 347004 60078
rect 382404 60076 383004 60078
rect 418404 60076 419004 60078
rect 454404 60076 455004 60078
rect 490404 60076 491004 60078
rect 526404 60076 527004 60078
rect 562404 60076 563004 60078
rect 588080 60076 588680 60078
rect -4756 60054 588680 60076
rect -4756 59818 -4574 60054
rect -4338 59818 22586 60054
rect 22822 59818 58586 60054
rect 58822 59818 94586 60054
rect 94822 59818 130586 60054
rect 130822 59818 166586 60054
rect 166822 59818 202586 60054
rect 202822 59818 238586 60054
rect 238822 59818 274586 60054
rect 274822 59818 310586 60054
rect 310822 59818 346586 60054
rect 346822 59818 382586 60054
rect 382822 59818 418586 60054
rect 418822 59818 454586 60054
rect 454822 59818 490586 60054
rect 490822 59818 526586 60054
rect 526822 59818 562586 60054
rect 562822 59818 588262 60054
rect 588498 59818 588680 60054
rect -4756 59734 588680 59818
rect -4756 59498 -4574 59734
rect -4338 59498 22586 59734
rect 22822 59498 58586 59734
rect 58822 59498 94586 59734
rect 94822 59498 130586 59734
rect 130822 59498 166586 59734
rect 166822 59498 202586 59734
rect 202822 59498 238586 59734
rect 238822 59498 274586 59734
rect 274822 59498 310586 59734
rect 310822 59498 346586 59734
rect 346822 59498 382586 59734
rect 382822 59498 418586 59734
rect 418822 59498 454586 59734
rect 454822 59498 490586 59734
rect 490822 59498 526586 59734
rect 526822 59498 562586 59734
rect 562822 59498 588262 59734
rect 588498 59498 588680 59734
rect -4756 59476 588680 59498
rect -4756 59474 -4156 59476
rect 22404 59474 23004 59476
rect 58404 59474 59004 59476
rect 94404 59474 95004 59476
rect 130404 59474 131004 59476
rect 166404 59474 167004 59476
rect 202404 59474 203004 59476
rect 238404 59474 239004 59476
rect 274404 59474 275004 59476
rect 310404 59474 311004 59476
rect 346404 59474 347004 59476
rect 382404 59474 383004 59476
rect 418404 59474 419004 59476
rect 454404 59474 455004 59476
rect 490404 59474 491004 59476
rect 526404 59474 527004 59476
rect 562404 59474 563004 59476
rect 588080 59474 588680 59476
rect -2916 56476 -2316 56478
rect 18804 56476 19404 56478
rect 54804 56476 55404 56478
rect 90804 56476 91404 56478
rect 126804 56476 127404 56478
rect 162804 56476 163404 56478
rect 198804 56476 199404 56478
rect 234804 56476 235404 56478
rect 270804 56476 271404 56478
rect 306804 56476 307404 56478
rect 342804 56476 343404 56478
rect 378804 56476 379404 56478
rect 414804 56476 415404 56478
rect 450804 56476 451404 56478
rect 486804 56476 487404 56478
rect 522804 56476 523404 56478
rect 558804 56476 559404 56478
rect 586240 56476 586840 56478
rect -2916 56454 586840 56476
rect -2916 56218 -2734 56454
rect -2498 56218 18986 56454
rect 19222 56218 54986 56454
rect 55222 56218 90986 56454
rect 91222 56218 126986 56454
rect 127222 56218 162986 56454
rect 163222 56218 198986 56454
rect 199222 56218 234986 56454
rect 235222 56218 270986 56454
rect 271222 56218 306986 56454
rect 307222 56218 342986 56454
rect 343222 56218 378986 56454
rect 379222 56218 414986 56454
rect 415222 56218 450986 56454
rect 451222 56218 486986 56454
rect 487222 56218 522986 56454
rect 523222 56218 558986 56454
rect 559222 56218 586422 56454
rect 586658 56218 586840 56454
rect -2916 56134 586840 56218
rect -2916 55898 -2734 56134
rect -2498 55898 18986 56134
rect 19222 55898 54986 56134
rect 55222 55898 90986 56134
rect 91222 55898 126986 56134
rect 127222 55898 162986 56134
rect 163222 55898 198986 56134
rect 199222 55898 234986 56134
rect 235222 55898 270986 56134
rect 271222 55898 306986 56134
rect 307222 55898 342986 56134
rect 343222 55898 378986 56134
rect 379222 55898 414986 56134
rect 415222 55898 450986 56134
rect 451222 55898 486986 56134
rect 487222 55898 522986 56134
rect 523222 55898 558986 56134
rect 559222 55898 586422 56134
rect 586658 55898 586840 56134
rect -2916 55876 586840 55898
rect -2916 55874 -2316 55876
rect 18804 55874 19404 55876
rect 54804 55874 55404 55876
rect 90804 55874 91404 55876
rect 126804 55874 127404 55876
rect 162804 55874 163404 55876
rect 198804 55874 199404 55876
rect 234804 55874 235404 55876
rect 270804 55874 271404 55876
rect 306804 55874 307404 55876
rect 342804 55874 343404 55876
rect 378804 55874 379404 55876
rect 414804 55874 415404 55876
rect 450804 55874 451404 55876
rect 486804 55874 487404 55876
rect 522804 55874 523404 55876
rect 558804 55874 559404 55876
rect 586240 55874 586840 55876
rect -7516 49276 -6916 49278
rect 11604 49276 12204 49278
rect 47604 49276 48204 49278
rect 83604 49276 84204 49278
rect 119604 49276 120204 49278
rect 155604 49276 156204 49278
rect 191604 49276 192204 49278
rect 227604 49276 228204 49278
rect 263604 49276 264204 49278
rect 299604 49276 300204 49278
rect 335604 49276 336204 49278
rect 371604 49276 372204 49278
rect 407604 49276 408204 49278
rect 443604 49276 444204 49278
rect 479604 49276 480204 49278
rect 515604 49276 516204 49278
rect 551604 49276 552204 49278
rect 590840 49276 591440 49278
rect -8436 49254 592360 49276
rect -8436 49018 -7334 49254
rect -7098 49018 11786 49254
rect 12022 49018 47786 49254
rect 48022 49018 83786 49254
rect 84022 49018 119786 49254
rect 120022 49018 155786 49254
rect 156022 49018 191786 49254
rect 192022 49018 227786 49254
rect 228022 49018 263786 49254
rect 264022 49018 299786 49254
rect 300022 49018 335786 49254
rect 336022 49018 371786 49254
rect 372022 49018 407786 49254
rect 408022 49018 443786 49254
rect 444022 49018 479786 49254
rect 480022 49018 515786 49254
rect 516022 49018 551786 49254
rect 552022 49018 591022 49254
rect 591258 49018 592360 49254
rect -8436 48934 592360 49018
rect -8436 48698 -7334 48934
rect -7098 48698 11786 48934
rect 12022 48698 47786 48934
rect 48022 48698 83786 48934
rect 84022 48698 119786 48934
rect 120022 48698 155786 48934
rect 156022 48698 191786 48934
rect 192022 48698 227786 48934
rect 228022 48698 263786 48934
rect 264022 48698 299786 48934
rect 300022 48698 335786 48934
rect 336022 48698 371786 48934
rect 372022 48698 407786 48934
rect 408022 48698 443786 48934
rect 444022 48698 479786 48934
rect 480022 48698 515786 48934
rect 516022 48698 551786 48934
rect 552022 48698 591022 48934
rect 591258 48698 592360 48934
rect -8436 48676 592360 48698
rect -7516 48674 -6916 48676
rect 11604 48674 12204 48676
rect 47604 48674 48204 48676
rect 83604 48674 84204 48676
rect 119604 48674 120204 48676
rect 155604 48674 156204 48676
rect 191604 48674 192204 48676
rect 227604 48674 228204 48676
rect 263604 48674 264204 48676
rect 299604 48674 300204 48676
rect 335604 48674 336204 48676
rect 371604 48674 372204 48676
rect 407604 48674 408204 48676
rect 443604 48674 444204 48676
rect 479604 48674 480204 48676
rect 515604 48674 516204 48676
rect 551604 48674 552204 48676
rect 590840 48674 591440 48676
rect -5676 45676 -5076 45678
rect 8004 45676 8604 45678
rect 44004 45676 44604 45678
rect 80004 45676 80604 45678
rect 116004 45676 116604 45678
rect 152004 45676 152604 45678
rect 188004 45676 188604 45678
rect 224004 45676 224604 45678
rect 260004 45676 260604 45678
rect 296004 45676 296604 45678
rect 332004 45676 332604 45678
rect 368004 45676 368604 45678
rect 404004 45676 404604 45678
rect 440004 45676 440604 45678
rect 476004 45676 476604 45678
rect 512004 45676 512604 45678
rect 548004 45676 548604 45678
rect 589000 45676 589600 45678
rect -6596 45654 590520 45676
rect -6596 45418 -5494 45654
rect -5258 45418 8186 45654
rect 8422 45418 44186 45654
rect 44422 45418 80186 45654
rect 80422 45418 116186 45654
rect 116422 45418 152186 45654
rect 152422 45418 188186 45654
rect 188422 45418 224186 45654
rect 224422 45418 260186 45654
rect 260422 45418 296186 45654
rect 296422 45418 332186 45654
rect 332422 45418 368186 45654
rect 368422 45418 404186 45654
rect 404422 45418 440186 45654
rect 440422 45418 476186 45654
rect 476422 45418 512186 45654
rect 512422 45418 548186 45654
rect 548422 45418 589182 45654
rect 589418 45418 590520 45654
rect -6596 45334 590520 45418
rect -6596 45098 -5494 45334
rect -5258 45098 8186 45334
rect 8422 45098 44186 45334
rect 44422 45098 80186 45334
rect 80422 45098 116186 45334
rect 116422 45098 152186 45334
rect 152422 45098 188186 45334
rect 188422 45098 224186 45334
rect 224422 45098 260186 45334
rect 260422 45098 296186 45334
rect 296422 45098 332186 45334
rect 332422 45098 368186 45334
rect 368422 45098 404186 45334
rect 404422 45098 440186 45334
rect 440422 45098 476186 45334
rect 476422 45098 512186 45334
rect 512422 45098 548186 45334
rect 548422 45098 589182 45334
rect 589418 45098 590520 45334
rect -6596 45076 590520 45098
rect -5676 45074 -5076 45076
rect 8004 45074 8604 45076
rect 44004 45074 44604 45076
rect 80004 45074 80604 45076
rect 116004 45074 116604 45076
rect 152004 45074 152604 45076
rect 188004 45074 188604 45076
rect 224004 45074 224604 45076
rect 260004 45074 260604 45076
rect 296004 45074 296604 45076
rect 332004 45074 332604 45076
rect 368004 45074 368604 45076
rect 404004 45074 404604 45076
rect 440004 45074 440604 45076
rect 476004 45074 476604 45076
rect 512004 45074 512604 45076
rect 548004 45074 548604 45076
rect 589000 45074 589600 45076
rect -3836 42076 -3236 42078
rect 4404 42076 5004 42078
rect 40404 42076 41004 42078
rect 76404 42076 77004 42078
rect 112404 42076 113004 42078
rect 148404 42076 149004 42078
rect 184404 42076 185004 42078
rect 220404 42076 221004 42078
rect 256404 42076 257004 42078
rect 292404 42076 293004 42078
rect 328404 42076 329004 42078
rect 364404 42076 365004 42078
rect 400404 42076 401004 42078
rect 436404 42076 437004 42078
rect 472404 42076 473004 42078
rect 508404 42076 509004 42078
rect 544404 42076 545004 42078
rect 580404 42076 581004 42078
rect 587160 42076 587760 42078
rect -4756 42054 588680 42076
rect -4756 41818 -3654 42054
rect -3418 41818 4586 42054
rect 4822 41818 40586 42054
rect 40822 41818 76586 42054
rect 76822 41818 112586 42054
rect 112822 41818 148586 42054
rect 148822 41818 184586 42054
rect 184822 41818 220586 42054
rect 220822 41818 256586 42054
rect 256822 41818 292586 42054
rect 292822 41818 328586 42054
rect 328822 41818 364586 42054
rect 364822 41818 400586 42054
rect 400822 41818 436586 42054
rect 436822 41818 472586 42054
rect 472822 41818 508586 42054
rect 508822 41818 544586 42054
rect 544822 41818 580586 42054
rect 580822 41818 587342 42054
rect 587578 41818 588680 42054
rect -4756 41734 588680 41818
rect -4756 41498 -3654 41734
rect -3418 41498 4586 41734
rect 4822 41498 40586 41734
rect 40822 41498 76586 41734
rect 76822 41498 112586 41734
rect 112822 41498 148586 41734
rect 148822 41498 184586 41734
rect 184822 41498 220586 41734
rect 220822 41498 256586 41734
rect 256822 41498 292586 41734
rect 292822 41498 328586 41734
rect 328822 41498 364586 41734
rect 364822 41498 400586 41734
rect 400822 41498 436586 41734
rect 436822 41498 472586 41734
rect 472822 41498 508586 41734
rect 508822 41498 544586 41734
rect 544822 41498 580586 41734
rect 580822 41498 587342 41734
rect 587578 41498 588680 41734
rect -4756 41476 588680 41498
rect -3836 41474 -3236 41476
rect 4404 41474 5004 41476
rect 40404 41474 41004 41476
rect 76404 41474 77004 41476
rect 112404 41474 113004 41476
rect 148404 41474 149004 41476
rect 184404 41474 185004 41476
rect 220404 41474 221004 41476
rect 256404 41474 257004 41476
rect 292404 41474 293004 41476
rect 328404 41474 329004 41476
rect 364404 41474 365004 41476
rect 400404 41474 401004 41476
rect 436404 41474 437004 41476
rect 472404 41474 473004 41476
rect 508404 41474 509004 41476
rect 544404 41474 545004 41476
rect 580404 41474 581004 41476
rect 587160 41474 587760 41476
rect -1996 38476 -1396 38478
rect 804 38476 1404 38478
rect 36804 38476 37404 38478
rect 72804 38476 73404 38478
rect 108804 38476 109404 38478
rect 144804 38476 145404 38478
rect 180804 38476 181404 38478
rect 216804 38476 217404 38478
rect 252804 38476 253404 38478
rect 288804 38476 289404 38478
rect 324804 38476 325404 38478
rect 360804 38476 361404 38478
rect 396804 38476 397404 38478
rect 432804 38476 433404 38478
rect 468804 38476 469404 38478
rect 504804 38476 505404 38478
rect 540804 38476 541404 38478
rect 576804 38476 577404 38478
rect 585320 38476 585920 38478
rect -2916 38454 586840 38476
rect -2916 38218 -1814 38454
rect -1578 38218 986 38454
rect 1222 38218 36986 38454
rect 37222 38218 72986 38454
rect 73222 38218 108986 38454
rect 109222 38218 144986 38454
rect 145222 38218 180986 38454
rect 181222 38218 216986 38454
rect 217222 38218 252986 38454
rect 253222 38218 288986 38454
rect 289222 38218 324986 38454
rect 325222 38218 360986 38454
rect 361222 38218 396986 38454
rect 397222 38218 432986 38454
rect 433222 38218 468986 38454
rect 469222 38218 504986 38454
rect 505222 38218 540986 38454
rect 541222 38218 576986 38454
rect 577222 38218 585502 38454
rect 585738 38218 586840 38454
rect -2916 38134 586840 38218
rect -2916 37898 -1814 38134
rect -1578 37898 986 38134
rect 1222 37898 36986 38134
rect 37222 37898 72986 38134
rect 73222 37898 108986 38134
rect 109222 37898 144986 38134
rect 145222 37898 180986 38134
rect 181222 37898 216986 38134
rect 217222 37898 252986 38134
rect 253222 37898 288986 38134
rect 289222 37898 324986 38134
rect 325222 37898 360986 38134
rect 361222 37898 396986 38134
rect 397222 37898 432986 38134
rect 433222 37898 468986 38134
rect 469222 37898 504986 38134
rect 505222 37898 540986 38134
rect 541222 37898 576986 38134
rect 577222 37898 585502 38134
rect 585738 37898 586840 38134
rect -2916 37876 586840 37898
rect -1996 37874 -1396 37876
rect 804 37874 1404 37876
rect 36804 37874 37404 37876
rect 72804 37874 73404 37876
rect 108804 37874 109404 37876
rect 144804 37874 145404 37876
rect 180804 37874 181404 37876
rect 216804 37874 217404 37876
rect 252804 37874 253404 37876
rect 288804 37874 289404 37876
rect 324804 37874 325404 37876
rect 360804 37874 361404 37876
rect 396804 37874 397404 37876
rect 432804 37874 433404 37876
rect 468804 37874 469404 37876
rect 504804 37874 505404 37876
rect 540804 37874 541404 37876
rect 576804 37874 577404 37876
rect 585320 37874 585920 37876
rect -8436 31276 -7836 31278
rect 29604 31276 30204 31278
rect 65604 31276 66204 31278
rect 101604 31276 102204 31278
rect 137604 31276 138204 31278
rect 173604 31276 174204 31278
rect 209604 31276 210204 31278
rect 245604 31276 246204 31278
rect 281604 31276 282204 31278
rect 317604 31276 318204 31278
rect 353604 31276 354204 31278
rect 389604 31276 390204 31278
rect 425604 31276 426204 31278
rect 461604 31276 462204 31278
rect 497604 31276 498204 31278
rect 533604 31276 534204 31278
rect 569604 31276 570204 31278
rect 591760 31276 592360 31278
rect -8436 31254 592360 31276
rect -8436 31018 -8254 31254
rect -8018 31018 29786 31254
rect 30022 31018 65786 31254
rect 66022 31018 101786 31254
rect 102022 31018 137786 31254
rect 138022 31018 173786 31254
rect 174022 31018 209786 31254
rect 210022 31018 245786 31254
rect 246022 31018 281786 31254
rect 282022 31018 317786 31254
rect 318022 31018 353786 31254
rect 354022 31018 389786 31254
rect 390022 31018 425786 31254
rect 426022 31018 461786 31254
rect 462022 31018 497786 31254
rect 498022 31018 533786 31254
rect 534022 31018 569786 31254
rect 570022 31018 591942 31254
rect 592178 31018 592360 31254
rect -8436 30934 592360 31018
rect -8436 30698 -8254 30934
rect -8018 30698 29786 30934
rect 30022 30698 65786 30934
rect 66022 30698 101786 30934
rect 102022 30698 137786 30934
rect 138022 30698 173786 30934
rect 174022 30698 209786 30934
rect 210022 30698 245786 30934
rect 246022 30698 281786 30934
rect 282022 30698 317786 30934
rect 318022 30698 353786 30934
rect 354022 30698 389786 30934
rect 390022 30698 425786 30934
rect 426022 30698 461786 30934
rect 462022 30698 497786 30934
rect 498022 30698 533786 30934
rect 534022 30698 569786 30934
rect 570022 30698 591942 30934
rect 592178 30698 592360 30934
rect -8436 30676 592360 30698
rect -8436 30674 -7836 30676
rect 29604 30674 30204 30676
rect 65604 30674 66204 30676
rect 101604 30674 102204 30676
rect 137604 30674 138204 30676
rect 173604 30674 174204 30676
rect 209604 30674 210204 30676
rect 245604 30674 246204 30676
rect 281604 30674 282204 30676
rect 317604 30674 318204 30676
rect 353604 30674 354204 30676
rect 389604 30674 390204 30676
rect 425604 30674 426204 30676
rect 461604 30674 462204 30676
rect 497604 30674 498204 30676
rect 533604 30674 534204 30676
rect 569604 30674 570204 30676
rect 591760 30674 592360 30676
rect -6596 27676 -5996 27678
rect 26004 27676 26604 27678
rect 62004 27676 62604 27678
rect 98004 27676 98604 27678
rect 134004 27676 134604 27678
rect 170004 27676 170604 27678
rect 206004 27676 206604 27678
rect 242004 27676 242604 27678
rect 278004 27676 278604 27678
rect 314004 27676 314604 27678
rect 350004 27676 350604 27678
rect 386004 27676 386604 27678
rect 422004 27676 422604 27678
rect 458004 27676 458604 27678
rect 494004 27676 494604 27678
rect 530004 27676 530604 27678
rect 566004 27676 566604 27678
rect 589920 27676 590520 27678
rect -6596 27654 590520 27676
rect -6596 27418 -6414 27654
rect -6178 27418 26186 27654
rect 26422 27418 62186 27654
rect 62422 27418 98186 27654
rect 98422 27418 134186 27654
rect 134422 27418 170186 27654
rect 170422 27418 206186 27654
rect 206422 27418 242186 27654
rect 242422 27418 278186 27654
rect 278422 27418 314186 27654
rect 314422 27418 350186 27654
rect 350422 27418 386186 27654
rect 386422 27418 422186 27654
rect 422422 27418 458186 27654
rect 458422 27418 494186 27654
rect 494422 27418 530186 27654
rect 530422 27418 566186 27654
rect 566422 27418 590102 27654
rect 590338 27418 590520 27654
rect -6596 27334 590520 27418
rect -6596 27098 -6414 27334
rect -6178 27098 26186 27334
rect 26422 27098 62186 27334
rect 62422 27098 98186 27334
rect 98422 27098 134186 27334
rect 134422 27098 170186 27334
rect 170422 27098 206186 27334
rect 206422 27098 242186 27334
rect 242422 27098 278186 27334
rect 278422 27098 314186 27334
rect 314422 27098 350186 27334
rect 350422 27098 386186 27334
rect 386422 27098 422186 27334
rect 422422 27098 458186 27334
rect 458422 27098 494186 27334
rect 494422 27098 530186 27334
rect 530422 27098 566186 27334
rect 566422 27098 590102 27334
rect 590338 27098 590520 27334
rect -6596 27076 590520 27098
rect -6596 27074 -5996 27076
rect 26004 27074 26604 27076
rect 62004 27074 62604 27076
rect 98004 27074 98604 27076
rect 134004 27074 134604 27076
rect 170004 27074 170604 27076
rect 206004 27074 206604 27076
rect 242004 27074 242604 27076
rect 278004 27074 278604 27076
rect 314004 27074 314604 27076
rect 350004 27074 350604 27076
rect 386004 27074 386604 27076
rect 422004 27074 422604 27076
rect 458004 27074 458604 27076
rect 494004 27074 494604 27076
rect 530004 27074 530604 27076
rect 566004 27074 566604 27076
rect 589920 27074 590520 27076
rect -4756 24076 -4156 24078
rect 22404 24076 23004 24078
rect 58404 24076 59004 24078
rect 94404 24076 95004 24078
rect 130404 24076 131004 24078
rect 166404 24076 167004 24078
rect 202404 24076 203004 24078
rect 238404 24076 239004 24078
rect 274404 24076 275004 24078
rect 310404 24076 311004 24078
rect 346404 24076 347004 24078
rect 382404 24076 383004 24078
rect 418404 24076 419004 24078
rect 454404 24076 455004 24078
rect 490404 24076 491004 24078
rect 526404 24076 527004 24078
rect 562404 24076 563004 24078
rect 588080 24076 588680 24078
rect -4756 24054 588680 24076
rect -4756 23818 -4574 24054
rect -4338 23818 22586 24054
rect 22822 23818 58586 24054
rect 58822 23818 94586 24054
rect 94822 23818 130586 24054
rect 130822 23818 166586 24054
rect 166822 23818 202586 24054
rect 202822 23818 238586 24054
rect 238822 23818 274586 24054
rect 274822 23818 310586 24054
rect 310822 23818 346586 24054
rect 346822 23818 382586 24054
rect 382822 23818 418586 24054
rect 418822 23818 454586 24054
rect 454822 23818 490586 24054
rect 490822 23818 526586 24054
rect 526822 23818 562586 24054
rect 562822 23818 588262 24054
rect 588498 23818 588680 24054
rect -4756 23734 588680 23818
rect -4756 23498 -4574 23734
rect -4338 23498 22586 23734
rect 22822 23498 58586 23734
rect 58822 23498 94586 23734
rect 94822 23498 130586 23734
rect 130822 23498 166586 23734
rect 166822 23498 202586 23734
rect 202822 23498 238586 23734
rect 238822 23498 274586 23734
rect 274822 23498 310586 23734
rect 310822 23498 346586 23734
rect 346822 23498 382586 23734
rect 382822 23498 418586 23734
rect 418822 23498 454586 23734
rect 454822 23498 490586 23734
rect 490822 23498 526586 23734
rect 526822 23498 562586 23734
rect 562822 23498 588262 23734
rect 588498 23498 588680 23734
rect -4756 23476 588680 23498
rect -4756 23474 -4156 23476
rect 22404 23474 23004 23476
rect 58404 23474 59004 23476
rect 94404 23474 95004 23476
rect 130404 23474 131004 23476
rect 166404 23474 167004 23476
rect 202404 23474 203004 23476
rect 238404 23474 239004 23476
rect 274404 23474 275004 23476
rect 310404 23474 311004 23476
rect 346404 23474 347004 23476
rect 382404 23474 383004 23476
rect 418404 23474 419004 23476
rect 454404 23474 455004 23476
rect 490404 23474 491004 23476
rect 526404 23474 527004 23476
rect 562404 23474 563004 23476
rect 588080 23474 588680 23476
rect -2916 20476 -2316 20478
rect 18804 20476 19404 20478
rect 54804 20476 55404 20478
rect 90804 20476 91404 20478
rect 126804 20476 127404 20478
rect 162804 20476 163404 20478
rect 198804 20476 199404 20478
rect 234804 20476 235404 20478
rect 270804 20476 271404 20478
rect 306804 20476 307404 20478
rect 342804 20476 343404 20478
rect 378804 20476 379404 20478
rect 414804 20476 415404 20478
rect 450804 20476 451404 20478
rect 486804 20476 487404 20478
rect 522804 20476 523404 20478
rect 558804 20476 559404 20478
rect 586240 20476 586840 20478
rect -2916 20454 586840 20476
rect -2916 20218 -2734 20454
rect -2498 20218 18986 20454
rect 19222 20218 54986 20454
rect 55222 20218 90986 20454
rect 91222 20218 126986 20454
rect 127222 20218 162986 20454
rect 163222 20218 198986 20454
rect 199222 20218 234986 20454
rect 235222 20218 270986 20454
rect 271222 20218 306986 20454
rect 307222 20218 342986 20454
rect 343222 20218 378986 20454
rect 379222 20218 414986 20454
rect 415222 20218 450986 20454
rect 451222 20218 486986 20454
rect 487222 20218 522986 20454
rect 523222 20218 558986 20454
rect 559222 20218 586422 20454
rect 586658 20218 586840 20454
rect -2916 20134 586840 20218
rect -2916 19898 -2734 20134
rect -2498 19898 18986 20134
rect 19222 19898 54986 20134
rect 55222 19898 90986 20134
rect 91222 19898 126986 20134
rect 127222 19898 162986 20134
rect 163222 19898 198986 20134
rect 199222 19898 234986 20134
rect 235222 19898 270986 20134
rect 271222 19898 306986 20134
rect 307222 19898 342986 20134
rect 343222 19898 378986 20134
rect 379222 19898 414986 20134
rect 415222 19898 450986 20134
rect 451222 19898 486986 20134
rect 487222 19898 522986 20134
rect 523222 19898 558986 20134
rect 559222 19898 586422 20134
rect 586658 19898 586840 20134
rect -2916 19876 586840 19898
rect -2916 19874 -2316 19876
rect 18804 19874 19404 19876
rect 54804 19874 55404 19876
rect 90804 19874 91404 19876
rect 126804 19874 127404 19876
rect 162804 19874 163404 19876
rect 198804 19874 199404 19876
rect 234804 19874 235404 19876
rect 270804 19874 271404 19876
rect 306804 19874 307404 19876
rect 342804 19874 343404 19876
rect 378804 19874 379404 19876
rect 414804 19874 415404 19876
rect 450804 19874 451404 19876
rect 486804 19874 487404 19876
rect 522804 19874 523404 19876
rect 558804 19874 559404 19876
rect 586240 19874 586840 19876
rect -7516 13276 -6916 13278
rect 11604 13276 12204 13278
rect 47604 13276 48204 13278
rect 83604 13276 84204 13278
rect 119604 13276 120204 13278
rect 155604 13276 156204 13278
rect 191604 13276 192204 13278
rect 227604 13276 228204 13278
rect 263604 13276 264204 13278
rect 299604 13276 300204 13278
rect 335604 13276 336204 13278
rect 371604 13276 372204 13278
rect 407604 13276 408204 13278
rect 443604 13276 444204 13278
rect 479604 13276 480204 13278
rect 515604 13276 516204 13278
rect 551604 13276 552204 13278
rect 590840 13276 591440 13278
rect -8436 13254 592360 13276
rect -8436 13018 -7334 13254
rect -7098 13018 11786 13254
rect 12022 13018 47786 13254
rect 48022 13018 83786 13254
rect 84022 13018 119786 13254
rect 120022 13018 155786 13254
rect 156022 13018 191786 13254
rect 192022 13018 227786 13254
rect 228022 13018 263786 13254
rect 264022 13018 299786 13254
rect 300022 13018 335786 13254
rect 336022 13018 371786 13254
rect 372022 13018 407786 13254
rect 408022 13018 443786 13254
rect 444022 13018 479786 13254
rect 480022 13018 515786 13254
rect 516022 13018 551786 13254
rect 552022 13018 591022 13254
rect 591258 13018 592360 13254
rect -8436 12934 592360 13018
rect -8436 12698 -7334 12934
rect -7098 12698 11786 12934
rect 12022 12698 47786 12934
rect 48022 12698 83786 12934
rect 84022 12698 119786 12934
rect 120022 12698 155786 12934
rect 156022 12698 191786 12934
rect 192022 12698 227786 12934
rect 228022 12698 263786 12934
rect 264022 12698 299786 12934
rect 300022 12698 335786 12934
rect 336022 12698 371786 12934
rect 372022 12698 407786 12934
rect 408022 12698 443786 12934
rect 444022 12698 479786 12934
rect 480022 12698 515786 12934
rect 516022 12698 551786 12934
rect 552022 12698 591022 12934
rect 591258 12698 592360 12934
rect -8436 12676 592360 12698
rect -7516 12674 -6916 12676
rect 11604 12674 12204 12676
rect 47604 12674 48204 12676
rect 83604 12674 84204 12676
rect 119604 12674 120204 12676
rect 155604 12674 156204 12676
rect 191604 12674 192204 12676
rect 227604 12674 228204 12676
rect 263604 12674 264204 12676
rect 299604 12674 300204 12676
rect 335604 12674 336204 12676
rect 371604 12674 372204 12676
rect 407604 12674 408204 12676
rect 443604 12674 444204 12676
rect 479604 12674 480204 12676
rect 515604 12674 516204 12676
rect 551604 12674 552204 12676
rect 590840 12674 591440 12676
rect -5676 9676 -5076 9678
rect 8004 9676 8604 9678
rect 44004 9676 44604 9678
rect 80004 9676 80604 9678
rect 116004 9676 116604 9678
rect 152004 9676 152604 9678
rect 188004 9676 188604 9678
rect 224004 9676 224604 9678
rect 260004 9676 260604 9678
rect 296004 9676 296604 9678
rect 332004 9676 332604 9678
rect 368004 9676 368604 9678
rect 404004 9676 404604 9678
rect 440004 9676 440604 9678
rect 476004 9676 476604 9678
rect 512004 9676 512604 9678
rect 548004 9676 548604 9678
rect 589000 9676 589600 9678
rect -6596 9654 590520 9676
rect -6596 9418 -5494 9654
rect -5258 9418 8186 9654
rect 8422 9418 44186 9654
rect 44422 9418 80186 9654
rect 80422 9418 116186 9654
rect 116422 9418 152186 9654
rect 152422 9418 188186 9654
rect 188422 9418 224186 9654
rect 224422 9418 260186 9654
rect 260422 9418 296186 9654
rect 296422 9418 332186 9654
rect 332422 9418 368186 9654
rect 368422 9418 404186 9654
rect 404422 9418 440186 9654
rect 440422 9418 476186 9654
rect 476422 9418 512186 9654
rect 512422 9418 548186 9654
rect 548422 9418 589182 9654
rect 589418 9418 590520 9654
rect -6596 9334 590520 9418
rect -6596 9098 -5494 9334
rect -5258 9098 8186 9334
rect 8422 9098 44186 9334
rect 44422 9098 80186 9334
rect 80422 9098 116186 9334
rect 116422 9098 152186 9334
rect 152422 9098 188186 9334
rect 188422 9098 224186 9334
rect 224422 9098 260186 9334
rect 260422 9098 296186 9334
rect 296422 9098 332186 9334
rect 332422 9098 368186 9334
rect 368422 9098 404186 9334
rect 404422 9098 440186 9334
rect 440422 9098 476186 9334
rect 476422 9098 512186 9334
rect 512422 9098 548186 9334
rect 548422 9098 589182 9334
rect 589418 9098 590520 9334
rect -6596 9076 590520 9098
rect -5676 9074 -5076 9076
rect 8004 9074 8604 9076
rect 44004 9074 44604 9076
rect 80004 9074 80604 9076
rect 116004 9074 116604 9076
rect 152004 9074 152604 9076
rect 188004 9074 188604 9076
rect 224004 9074 224604 9076
rect 260004 9074 260604 9076
rect 296004 9074 296604 9076
rect 332004 9074 332604 9076
rect 368004 9074 368604 9076
rect 404004 9074 404604 9076
rect 440004 9074 440604 9076
rect 476004 9074 476604 9076
rect 512004 9074 512604 9076
rect 548004 9074 548604 9076
rect 589000 9074 589600 9076
rect -3836 6076 -3236 6078
rect 4404 6076 5004 6078
rect 40404 6076 41004 6078
rect 76404 6076 77004 6078
rect 112404 6076 113004 6078
rect 148404 6076 149004 6078
rect 184404 6076 185004 6078
rect 220404 6076 221004 6078
rect 256404 6076 257004 6078
rect 292404 6076 293004 6078
rect 328404 6076 329004 6078
rect 364404 6076 365004 6078
rect 400404 6076 401004 6078
rect 436404 6076 437004 6078
rect 472404 6076 473004 6078
rect 508404 6076 509004 6078
rect 544404 6076 545004 6078
rect 580404 6076 581004 6078
rect 587160 6076 587760 6078
rect -4756 6054 588680 6076
rect -4756 5818 -3654 6054
rect -3418 5818 4586 6054
rect 4822 5818 40586 6054
rect 40822 5818 76586 6054
rect 76822 5818 112586 6054
rect 112822 5818 148586 6054
rect 148822 5818 184586 6054
rect 184822 5818 220586 6054
rect 220822 5818 256586 6054
rect 256822 5818 292586 6054
rect 292822 5818 328586 6054
rect 328822 5818 364586 6054
rect 364822 5818 400586 6054
rect 400822 5818 436586 6054
rect 436822 5818 472586 6054
rect 472822 5818 508586 6054
rect 508822 5818 544586 6054
rect 544822 5818 580586 6054
rect 580822 5818 587342 6054
rect 587578 5818 588680 6054
rect -4756 5734 588680 5818
rect -4756 5498 -3654 5734
rect -3418 5498 4586 5734
rect 4822 5498 40586 5734
rect 40822 5498 76586 5734
rect 76822 5498 112586 5734
rect 112822 5498 148586 5734
rect 148822 5498 184586 5734
rect 184822 5498 220586 5734
rect 220822 5498 256586 5734
rect 256822 5498 292586 5734
rect 292822 5498 328586 5734
rect 328822 5498 364586 5734
rect 364822 5498 400586 5734
rect 400822 5498 436586 5734
rect 436822 5498 472586 5734
rect 472822 5498 508586 5734
rect 508822 5498 544586 5734
rect 544822 5498 580586 5734
rect 580822 5498 587342 5734
rect 587578 5498 588680 5734
rect -4756 5476 588680 5498
rect -3836 5474 -3236 5476
rect 4404 5474 5004 5476
rect 40404 5474 41004 5476
rect 76404 5474 77004 5476
rect 112404 5474 113004 5476
rect 148404 5474 149004 5476
rect 184404 5474 185004 5476
rect 220404 5474 221004 5476
rect 256404 5474 257004 5476
rect 292404 5474 293004 5476
rect 328404 5474 329004 5476
rect 364404 5474 365004 5476
rect 400404 5474 401004 5476
rect 436404 5474 437004 5476
rect 472404 5474 473004 5476
rect 508404 5474 509004 5476
rect 544404 5474 545004 5476
rect 580404 5474 581004 5476
rect 587160 5474 587760 5476
rect -1996 2476 -1396 2478
rect 804 2476 1404 2478
rect 36804 2476 37404 2478
rect 72804 2476 73404 2478
rect 108804 2476 109404 2478
rect 144804 2476 145404 2478
rect 180804 2476 181404 2478
rect 216804 2476 217404 2478
rect 252804 2476 253404 2478
rect 288804 2476 289404 2478
rect 324804 2476 325404 2478
rect 360804 2476 361404 2478
rect 396804 2476 397404 2478
rect 432804 2476 433404 2478
rect 468804 2476 469404 2478
rect 504804 2476 505404 2478
rect 540804 2476 541404 2478
rect 576804 2476 577404 2478
rect 585320 2476 585920 2478
rect -2916 2454 586840 2476
rect -2916 2218 -1814 2454
rect -1578 2218 986 2454
rect 1222 2218 36986 2454
rect 37222 2218 72986 2454
rect 73222 2218 108986 2454
rect 109222 2218 144986 2454
rect 145222 2218 180986 2454
rect 181222 2218 216986 2454
rect 217222 2218 252986 2454
rect 253222 2218 288986 2454
rect 289222 2218 324986 2454
rect 325222 2218 360986 2454
rect 361222 2218 396986 2454
rect 397222 2218 432986 2454
rect 433222 2218 468986 2454
rect 469222 2218 504986 2454
rect 505222 2218 540986 2454
rect 541222 2218 576986 2454
rect 577222 2218 585502 2454
rect 585738 2218 586840 2454
rect -2916 2134 586840 2218
rect -2916 1898 -1814 2134
rect -1578 1898 986 2134
rect 1222 1898 36986 2134
rect 37222 1898 72986 2134
rect 73222 1898 108986 2134
rect 109222 1898 144986 2134
rect 145222 1898 180986 2134
rect 181222 1898 216986 2134
rect 217222 1898 252986 2134
rect 253222 1898 288986 2134
rect 289222 1898 324986 2134
rect 325222 1898 360986 2134
rect 361222 1898 396986 2134
rect 397222 1898 432986 2134
rect 433222 1898 468986 2134
rect 469222 1898 504986 2134
rect 505222 1898 540986 2134
rect 541222 1898 576986 2134
rect 577222 1898 585502 2134
rect 585738 1898 586840 2134
rect -2916 1876 586840 1898
rect -1996 1874 -1396 1876
rect 804 1874 1404 1876
rect 36804 1874 37404 1876
rect 72804 1874 73404 1876
rect 108804 1874 109404 1876
rect 144804 1874 145404 1876
rect 180804 1874 181404 1876
rect 216804 1874 217404 1876
rect 252804 1874 253404 1876
rect 288804 1874 289404 1876
rect 324804 1874 325404 1876
rect 360804 1874 361404 1876
rect 396804 1874 397404 1876
rect 432804 1874 433404 1876
rect 468804 1874 469404 1876
rect 504804 1874 505404 1876
rect 540804 1874 541404 1876
rect 576804 1874 577404 1876
rect 585320 1874 585920 1876
rect -1996 -324 -1396 -322
rect 804 -324 1404 -322
rect 36804 -324 37404 -322
rect 72804 -324 73404 -322
rect 108804 -324 109404 -322
rect 144804 -324 145404 -322
rect 180804 -324 181404 -322
rect 216804 -324 217404 -322
rect 252804 -324 253404 -322
rect 288804 -324 289404 -322
rect 324804 -324 325404 -322
rect 360804 -324 361404 -322
rect 396804 -324 397404 -322
rect 432804 -324 433404 -322
rect 468804 -324 469404 -322
rect 504804 -324 505404 -322
rect 540804 -324 541404 -322
rect 576804 -324 577404 -322
rect 585320 -324 585920 -322
rect -1996 -346 585920 -324
rect -1996 -582 -1814 -346
rect -1578 -582 986 -346
rect 1222 -582 36986 -346
rect 37222 -582 72986 -346
rect 73222 -582 108986 -346
rect 109222 -582 144986 -346
rect 145222 -582 180986 -346
rect 181222 -582 216986 -346
rect 217222 -582 252986 -346
rect 253222 -582 288986 -346
rect 289222 -582 324986 -346
rect 325222 -582 360986 -346
rect 361222 -582 396986 -346
rect 397222 -582 432986 -346
rect 433222 -582 468986 -346
rect 469222 -582 504986 -346
rect 505222 -582 540986 -346
rect 541222 -582 576986 -346
rect 577222 -582 585502 -346
rect 585738 -582 585920 -346
rect -1996 -666 585920 -582
rect -1996 -902 -1814 -666
rect -1578 -902 986 -666
rect 1222 -902 36986 -666
rect 37222 -902 72986 -666
rect 73222 -902 108986 -666
rect 109222 -902 144986 -666
rect 145222 -902 180986 -666
rect 181222 -902 216986 -666
rect 217222 -902 252986 -666
rect 253222 -902 288986 -666
rect 289222 -902 324986 -666
rect 325222 -902 360986 -666
rect 361222 -902 396986 -666
rect 397222 -902 432986 -666
rect 433222 -902 468986 -666
rect 469222 -902 504986 -666
rect 505222 -902 540986 -666
rect 541222 -902 576986 -666
rect 577222 -902 585502 -666
rect 585738 -902 585920 -666
rect -1996 -924 585920 -902
rect -1996 -926 -1396 -924
rect 804 -926 1404 -924
rect 36804 -926 37404 -924
rect 72804 -926 73404 -924
rect 108804 -926 109404 -924
rect 144804 -926 145404 -924
rect 180804 -926 181404 -924
rect 216804 -926 217404 -924
rect 252804 -926 253404 -924
rect 288804 -926 289404 -924
rect 324804 -926 325404 -924
rect 360804 -926 361404 -924
rect 396804 -926 397404 -924
rect 432804 -926 433404 -924
rect 468804 -926 469404 -924
rect 504804 -926 505404 -924
rect 540804 -926 541404 -924
rect 576804 -926 577404 -924
rect 585320 -926 585920 -924
rect -2916 -1244 -2316 -1242
rect 18804 -1244 19404 -1242
rect 54804 -1244 55404 -1242
rect 90804 -1244 91404 -1242
rect 126804 -1244 127404 -1242
rect 162804 -1244 163404 -1242
rect 198804 -1244 199404 -1242
rect 234804 -1244 235404 -1242
rect 270804 -1244 271404 -1242
rect 306804 -1244 307404 -1242
rect 342804 -1244 343404 -1242
rect 378804 -1244 379404 -1242
rect 414804 -1244 415404 -1242
rect 450804 -1244 451404 -1242
rect 486804 -1244 487404 -1242
rect 522804 -1244 523404 -1242
rect 558804 -1244 559404 -1242
rect 586240 -1244 586840 -1242
rect -2916 -1266 586840 -1244
rect -2916 -1502 -2734 -1266
rect -2498 -1502 18986 -1266
rect 19222 -1502 54986 -1266
rect 55222 -1502 90986 -1266
rect 91222 -1502 126986 -1266
rect 127222 -1502 162986 -1266
rect 163222 -1502 198986 -1266
rect 199222 -1502 234986 -1266
rect 235222 -1502 270986 -1266
rect 271222 -1502 306986 -1266
rect 307222 -1502 342986 -1266
rect 343222 -1502 378986 -1266
rect 379222 -1502 414986 -1266
rect 415222 -1502 450986 -1266
rect 451222 -1502 486986 -1266
rect 487222 -1502 522986 -1266
rect 523222 -1502 558986 -1266
rect 559222 -1502 586422 -1266
rect 586658 -1502 586840 -1266
rect -2916 -1586 586840 -1502
rect -2916 -1822 -2734 -1586
rect -2498 -1822 18986 -1586
rect 19222 -1822 54986 -1586
rect 55222 -1822 90986 -1586
rect 91222 -1822 126986 -1586
rect 127222 -1822 162986 -1586
rect 163222 -1822 198986 -1586
rect 199222 -1822 234986 -1586
rect 235222 -1822 270986 -1586
rect 271222 -1822 306986 -1586
rect 307222 -1822 342986 -1586
rect 343222 -1822 378986 -1586
rect 379222 -1822 414986 -1586
rect 415222 -1822 450986 -1586
rect 451222 -1822 486986 -1586
rect 487222 -1822 522986 -1586
rect 523222 -1822 558986 -1586
rect 559222 -1822 586422 -1586
rect 586658 -1822 586840 -1586
rect -2916 -1844 586840 -1822
rect -2916 -1846 -2316 -1844
rect 18804 -1846 19404 -1844
rect 54804 -1846 55404 -1844
rect 90804 -1846 91404 -1844
rect 126804 -1846 127404 -1844
rect 162804 -1846 163404 -1844
rect 198804 -1846 199404 -1844
rect 234804 -1846 235404 -1844
rect 270804 -1846 271404 -1844
rect 306804 -1846 307404 -1844
rect 342804 -1846 343404 -1844
rect 378804 -1846 379404 -1844
rect 414804 -1846 415404 -1844
rect 450804 -1846 451404 -1844
rect 486804 -1846 487404 -1844
rect 522804 -1846 523404 -1844
rect 558804 -1846 559404 -1844
rect 586240 -1846 586840 -1844
rect -3836 -2164 -3236 -2162
rect 4404 -2164 5004 -2162
rect 40404 -2164 41004 -2162
rect 76404 -2164 77004 -2162
rect 112404 -2164 113004 -2162
rect 148404 -2164 149004 -2162
rect 184404 -2164 185004 -2162
rect 220404 -2164 221004 -2162
rect 256404 -2164 257004 -2162
rect 292404 -2164 293004 -2162
rect 328404 -2164 329004 -2162
rect 364404 -2164 365004 -2162
rect 400404 -2164 401004 -2162
rect 436404 -2164 437004 -2162
rect 472404 -2164 473004 -2162
rect 508404 -2164 509004 -2162
rect 544404 -2164 545004 -2162
rect 580404 -2164 581004 -2162
rect 587160 -2164 587760 -2162
rect -3836 -2186 587760 -2164
rect -3836 -2422 -3654 -2186
rect -3418 -2422 4586 -2186
rect 4822 -2422 40586 -2186
rect 40822 -2422 76586 -2186
rect 76822 -2422 112586 -2186
rect 112822 -2422 148586 -2186
rect 148822 -2422 184586 -2186
rect 184822 -2422 220586 -2186
rect 220822 -2422 256586 -2186
rect 256822 -2422 292586 -2186
rect 292822 -2422 328586 -2186
rect 328822 -2422 364586 -2186
rect 364822 -2422 400586 -2186
rect 400822 -2422 436586 -2186
rect 436822 -2422 472586 -2186
rect 472822 -2422 508586 -2186
rect 508822 -2422 544586 -2186
rect 544822 -2422 580586 -2186
rect 580822 -2422 587342 -2186
rect 587578 -2422 587760 -2186
rect -3836 -2506 587760 -2422
rect -3836 -2742 -3654 -2506
rect -3418 -2742 4586 -2506
rect 4822 -2742 40586 -2506
rect 40822 -2742 76586 -2506
rect 76822 -2742 112586 -2506
rect 112822 -2742 148586 -2506
rect 148822 -2742 184586 -2506
rect 184822 -2742 220586 -2506
rect 220822 -2742 256586 -2506
rect 256822 -2742 292586 -2506
rect 292822 -2742 328586 -2506
rect 328822 -2742 364586 -2506
rect 364822 -2742 400586 -2506
rect 400822 -2742 436586 -2506
rect 436822 -2742 472586 -2506
rect 472822 -2742 508586 -2506
rect 508822 -2742 544586 -2506
rect 544822 -2742 580586 -2506
rect 580822 -2742 587342 -2506
rect 587578 -2742 587760 -2506
rect -3836 -2764 587760 -2742
rect -3836 -2766 -3236 -2764
rect 4404 -2766 5004 -2764
rect 40404 -2766 41004 -2764
rect 76404 -2766 77004 -2764
rect 112404 -2766 113004 -2764
rect 148404 -2766 149004 -2764
rect 184404 -2766 185004 -2764
rect 220404 -2766 221004 -2764
rect 256404 -2766 257004 -2764
rect 292404 -2766 293004 -2764
rect 328404 -2766 329004 -2764
rect 364404 -2766 365004 -2764
rect 400404 -2766 401004 -2764
rect 436404 -2766 437004 -2764
rect 472404 -2766 473004 -2764
rect 508404 -2766 509004 -2764
rect 544404 -2766 545004 -2764
rect 580404 -2766 581004 -2764
rect 587160 -2766 587760 -2764
rect -4756 -3084 -4156 -3082
rect 22404 -3084 23004 -3082
rect 58404 -3084 59004 -3082
rect 94404 -3084 95004 -3082
rect 130404 -3084 131004 -3082
rect 166404 -3084 167004 -3082
rect 202404 -3084 203004 -3082
rect 238404 -3084 239004 -3082
rect 274404 -3084 275004 -3082
rect 310404 -3084 311004 -3082
rect 346404 -3084 347004 -3082
rect 382404 -3084 383004 -3082
rect 418404 -3084 419004 -3082
rect 454404 -3084 455004 -3082
rect 490404 -3084 491004 -3082
rect 526404 -3084 527004 -3082
rect 562404 -3084 563004 -3082
rect 588080 -3084 588680 -3082
rect -4756 -3106 588680 -3084
rect -4756 -3342 -4574 -3106
rect -4338 -3342 22586 -3106
rect 22822 -3342 58586 -3106
rect 58822 -3342 94586 -3106
rect 94822 -3342 130586 -3106
rect 130822 -3342 166586 -3106
rect 166822 -3342 202586 -3106
rect 202822 -3342 238586 -3106
rect 238822 -3342 274586 -3106
rect 274822 -3342 310586 -3106
rect 310822 -3342 346586 -3106
rect 346822 -3342 382586 -3106
rect 382822 -3342 418586 -3106
rect 418822 -3342 454586 -3106
rect 454822 -3342 490586 -3106
rect 490822 -3342 526586 -3106
rect 526822 -3342 562586 -3106
rect 562822 -3342 588262 -3106
rect 588498 -3342 588680 -3106
rect -4756 -3426 588680 -3342
rect -4756 -3662 -4574 -3426
rect -4338 -3662 22586 -3426
rect 22822 -3662 58586 -3426
rect 58822 -3662 94586 -3426
rect 94822 -3662 130586 -3426
rect 130822 -3662 166586 -3426
rect 166822 -3662 202586 -3426
rect 202822 -3662 238586 -3426
rect 238822 -3662 274586 -3426
rect 274822 -3662 310586 -3426
rect 310822 -3662 346586 -3426
rect 346822 -3662 382586 -3426
rect 382822 -3662 418586 -3426
rect 418822 -3662 454586 -3426
rect 454822 -3662 490586 -3426
rect 490822 -3662 526586 -3426
rect 526822 -3662 562586 -3426
rect 562822 -3662 588262 -3426
rect 588498 -3662 588680 -3426
rect -4756 -3684 588680 -3662
rect -4756 -3686 -4156 -3684
rect 22404 -3686 23004 -3684
rect 58404 -3686 59004 -3684
rect 94404 -3686 95004 -3684
rect 130404 -3686 131004 -3684
rect 166404 -3686 167004 -3684
rect 202404 -3686 203004 -3684
rect 238404 -3686 239004 -3684
rect 274404 -3686 275004 -3684
rect 310404 -3686 311004 -3684
rect 346404 -3686 347004 -3684
rect 382404 -3686 383004 -3684
rect 418404 -3686 419004 -3684
rect 454404 -3686 455004 -3684
rect 490404 -3686 491004 -3684
rect 526404 -3686 527004 -3684
rect 562404 -3686 563004 -3684
rect 588080 -3686 588680 -3684
rect -5676 -4004 -5076 -4002
rect 8004 -4004 8604 -4002
rect 44004 -4004 44604 -4002
rect 80004 -4004 80604 -4002
rect 116004 -4004 116604 -4002
rect 152004 -4004 152604 -4002
rect 188004 -4004 188604 -4002
rect 224004 -4004 224604 -4002
rect 260004 -4004 260604 -4002
rect 296004 -4004 296604 -4002
rect 332004 -4004 332604 -4002
rect 368004 -4004 368604 -4002
rect 404004 -4004 404604 -4002
rect 440004 -4004 440604 -4002
rect 476004 -4004 476604 -4002
rect 512004 -4004 512604 -4002
rect 548004 -4004 548604 -4002
rect 589000 -4004 589600 -4002
rect -5676 -4026 589600 -4004
rect -5676 -4262 -5494 -4026
rect -5258 -4262 8186 -4026
rect 8422 -4262 44186 -4026
rect 44422 -4262 80186 -4026
rect 80422 -4262 116186 -4026
rect 116422 -4262 152186 -4026
rect 152422 -4262 188186 -4026
rect 188422 -4262 224186 -4026
rect 224422 -4262 260186 -4026
rect 260422 -4262 296186 -4026
rect 296422 -4262 332186 -4026
rect 332422 -4262 368186 -4026
rect 368422 -4262 404186 -4026
rect 404422 -4262 440186 -4026
rect 440422 -4262 476186 -4026
rect 476422 -4262 512186 -4026
rect 512422 -4262 548186 -4026
rect 548422 -4262 589182 -4026
rect 589418 -4262 589600 -4026
rect -5676 -4346 589600 -4262
rect -5676 -4582 -5494 -4346
rect -5258 -4582 8186 -4346
rect 8422 -4582 44186 -4346
rect 44422 -4582 80186 -4346
rect 80422 -4582 116186 -4346
rect 116422 -4582 152186 -4346
rect 152422 -4582 188186 -4346
rect 188422 -4582 224186 -4346
rect 224422 -4582 260186 -4346
rect 260422 -4582 296186 -4346
rect 296422 -4582 332186 -4346
rect 332422 -4582 368186 -4346
rect 368422 -4582 404186 -4346
rect 404422 -4582 440186 -4346
rect 440422 -4582 476186 -4346
rect 476422 -4582 512186 -4346
rect 512422 -4582 548186 -4346
rect 548422 -4582 589182 -4346
rect 589418 -4582 589600 -4346
rect -5676 -4604 589600 -4582
rect -5676 -4606 -5076 -4604
rect 8004 -4606 8604 -4604
rect 44004 -4606 44604 -4604
rect 80004 -4606 80604 -4604
rect 116004 -4606 116604 -4604
rect 152004 -4606 152604 -4604
rect 188004 -4606 188604 -4604
rect 224004 -4606 224604 -4604
rect 260004 -4606 260604 -4604
rect 296004 -4606 296604 -4604
rect 332004 -4606 332604 -4604
rect 368004 -4606 368604 -4604
rect 404004 -4606 404604 -4604
rect 440004 -4606 440604 -4604
rect 476004 -4606 476604 -4604
rect 512004 -4606 512604 -4604
rect 548004 -4606 548604 -4604
rect 589000 -4606 589600 -4604
rect -6596 -4924 -5996 -4922
rect 26004 -4924 26604 -4922
rect 62004 -4924 62604 -4922
rect 98004 -4924 98604 -4922
rect 134004 -4924 134604 -4922
rect 170004 -4924 170604 -4922
rect 206004 -4924 206604 -4922
rect 242004 -4924 242604 -4922
rect 278004 -4924 278604 -4922
rect 314004 -4924 314604 -4922
rect 350004 -4924 350604 -4922
rect 386004 -4924 386604 -4922
rect 422004 -4924 422604 -4922
rect 458004 -4924 458604 -4922
rect 494004 -4924 494604 -4922
rect 530004 -4924 530604 -4922
rect 566004 -4924 566604 -4922
rect 589920 -4924 590520 -4922
rect -6596 -4946 590520 -4924
rect -6596 -5182 -6414 -4946
rect -6178 -5182 26186 -4946
rect 26422 -5182 62186 -4946
rect 62422 -5182 98186 -4946
rect 98422 -5182 134186 -4946
rect 134422 -5182 170186 -4946
rect 170422 -5182 206186 -4946
rect 206422 -5182 242186 -4946
rect 242422 -5182 278186 -4946
rect 278422 -5182 314186 -4946
rect 314422 -5182 350186 -4946
rect 350422 -5182 386186 -4946
rect 386422 -5182 422186 -4946
rect 422422 -5182 458186 -4946
rect 458422 -5182 494186 -4946
rect 494422 -5182 530186 -4946
rect 530422 -5182 566186 -4946
rect 566422 -5182 590102 -4946
rect 590338 -5182 590520 -4946
rect -6596 -5266 590520 -5182
rect -6596 -5502 -6414 -5266
rect -6178 -5502 26186 -5266
rect 26422 -5502 62186 -5266
rect 62422 -5502 98186 -5266
rect 98422 -5502 134186 -5266
rect 134422 -5502 170186 -5266
rect 170422 -5502 206186 -5266
rect 206422 -5502 242186 -5266
rect 242422 -5502 278186 -5266
rect 278422 -5502 314186 -5266
rect 314422 -5502 350186 -5266
rect 350422 -5502 386186 -5266
rect 386422 -5502 422186 -5266
rect 422422 -5502 458186 -5266
rect 458422 -5502 494186 -5266
rect 494422 -5502 530186 -5266
rect 530422 -5502 566186 -5266
rect 566422 -5502 590102 -5266
rect 590338 -5502 590520 -5266
rect -6596 -5524 590520 -5502
rect -6596 -5526 -5996 -5524
rect 26004 -5526 26604 -5524
rect 62004 -5526 62604 -5524
rect 98004 -5526 98604 -5524
rect 134004 -5526 134604 -5524
rect 170004 -5526 170604 -5524
rect 206004 -5526 206604 -5524
rect 242004 -5526 242604 -5524
rect 278004 -5526 278604 -5524
rect 314004 -5526 314604 -5524
rect 350004 -5526 350604 -5524
rect 386004 -5526 386604 -5524
rect 422004 -5526 422604 -5524
rect 458004 -5526 458604 -5524
rect 494004 -5526 494604 -5524
rect 530004 -5526 530604 -5524
rect 566004 -5526 566604 -5524
rect 589920 -5526 590520 -5524
rect -7516 -5844 -6916 -5842
rect 11604 -5844 12204 -5842
rect 47604 -5844 48204 -5842
rect 83604 -5844 84204 -5842
rect 119604 -5844 120204 -5842
rect 155604 -5844 156204 -5842
rect 191604 -5844 192204 -5842
rect 227604 -5844 228204 -5842
rect 263604 -5844 264204 -5842
rect 299604 -5844 300204 -5842
rect 335604 -5844 336204 -5842
rect 371604 -5844 372204 -5842
rect 407604 -5844 408204 -5842
rect 443604 -5844 444204 -5842
rect 479604 -5844 480204 -5842
rect 515604 -5844 516204 -5842
rect 551604 -5844 552204 -5842
rect 590840 -5844 591440 -5842
rect -7516 -5866 591440 -5844
rect -7516 -6102 -7334 -5866
rect -7098 -6102 11786 -5866
rect 12022 -6102 47786 -5866
rect 48022 -6102 83786 -5866
rect 84022 -6102 119786 -5866
rect 120022 -6102 155786 -5866
rect 156022 -6102 191786 -5866
rect 192022 -6102 227786 -5866
rect 228022 -6102 263786 -5866
rect 264022 -6102 299786 -5866
rect 300022 -6102 335786 -5866
rect 336022 -6102 371786 -5866
rect 372022 -6102 407786 -5866
rect 408022 -6102 443786 -5866
rect 444022 -6102 479786 -5866
rect 480022 -6102 515786 -5866
rect 516022 -6102 551786 -5866
rect 552022 -6102 591022 -5866
rect 591258 -6102 591440 -5866
rect -7516 -6186 591440 -6102
rect -7516 -6422 -7334 -6186
rect -7098 -6422 11786 -6186
rect 12022 -6422 47786 -6186
rect 48022 -6422 83786 -6186
rect 84022 -6422 119786 -6186
rect 120022 -6422 155786 -6186
rect 156022 -6422 191786 -6186
rect 192022 -6422 227786 -6186
rect 228022 -6422 263786 -6186
rect 264022 -6422 299786 -6186
rect 300022 -6422 335786 -6186
rect 336022 -6422 371786 -6186
rect 372022 -6422 407786 -6186
rect 408022 -6422 443786 -6186
rect 444022 -6422 479786 -6186
rect 480022 -6422 515786 -6186
rect 516022 -6422 551786 -6186
rect 552022 -6422 591022 -6186
rect 591258 -6422 591440 -6186
rect -7516 -6444 591440 -6422
rect -7516 -6446 -6916 -6444
rect 11604 -6446 12204 -6444
rect 47604 -6446 48204 -6444
rect 83604 -6446 84204 -6444
rect 119604 -6446 120204 -6444
rect 155604 -6446 156204 -6444
rect 191604 -6446 192204 -6444
rect 227604 -6446 228204 -6444
rect 263604 -6446 264204 -6444
rect 299604 -6446 300204 -6444
rect 335604 -6446 336204 -6444
rect 371604 -6446 372204 -6444
rect 407604 -6446 408204 -6444
rect 443604 -6446 444204 -6444
rect 479604 -6446 480204 -6444
rect 515604 -6446 516204 -6444
rect 551604 -6446 552204 -6444
rect 590840 -6446 591440 -6444
rect -8436 -6764 -7836 -6762
rect 29604 -6764 30204 -6762
rect 65604 -6764 66204 -6762
rect 101604 -6764 102204 -6762
rect 137604 -6764 138204 -6762
rect 173604 -6764 174204 -6762
rect 209604 -6764 210204 -6762
rect 245604 -6764 246204 -6762
rect 281604 -6764 282204 -6762
rect 317604 -6764 318204 -6762
rect 353604 -6764 354204 -6762
rect 389604 -6764 390204 -6762
rect 425604 -6764 426204 -6762
rect 461604 -6764 462204 -6762
rect 497604 -6764 498204 -6762
rect 533604 -6764 534204 -6762
rect 569604 -6764 570204 -6762
rect 591760 -6764 592360 -6762
rect -8436 -6786 592360 -6764
rect -8436 -7022 -8254 -6786
rect -8018 -7022 29786 -6786
rect 30022 -7022 65786 -6786
rect 66022 -7022 101786 -6786
rect 102022 -7022 137786 -6786
rect 138022 -7022 173786 -6786
rect 174022 -7022 209786 -6786
rect 210022 -7022 245786 -6786
rect 246022 -7022 281786 -6786
rect 282022 -7022 317786 -6786
rect 318022 -7022 353786 -6786
rect 354022 -7022 389786 -6786
rect 390022 -7022 425786 -6786
rect 426022 -7022 461786 -6786
rect 462022 -7022 497786 -6786
rect 498022 -7022 533786 -6786
rect 534022 -7022 569786 -6786
rect 570022 -7022 591942 -6786
rect 592178 -7022 592360 -6786
rect -8436 -7106 592360 -7022
rect -8436 -7342 -8254 -7106
rect -8018 -7342 29786 -7106
rect 30022 -7342 65786 -7106
rect 66022 -7342 101786 -7106
rect 102022 -7342 137786 -7106
rect 138022 -7342 173786 -7106
rect 174022 -7342 209786 -7106
rect 210022 -7342 245786 -7106
rect 246022 -7342 281786 -7106
rect 282022 -7342 317786 -7106
rect 318022 -7342 353786 -7106
rect 354022 -7342 389786 -7106
rect 390022 -7342 425786 -7106
rect 426022 -7342 461786 -7106
rect 462022 -7342 497786 -7106
rect 498022 -7342 533786 -7106
rect 534022 -7342 569786 -7106
rect 570022 -7342 591942 -7106
rect 592178 -7342 592360 -7106
rect -8436 -7364 592360 -7342
rect -8436 -7366 -7836 -7364
rect 29604 -7366 30204 -7364
rect 65604 -7366 66204 -7364
rect 101604 -7366 102204 -7364
rect 137604 -7366 138204 -7364
rect 173604 -7366 174204 -7364
rect 209604 -7366 210204 -7364
rect 245604 -7366 246204 -7364
rect 281604 -7366 282204 -7364
rect 317604 -7366 318204 -7364
rect 353604 -7366 354204 -7364
rect 389604 -7366 390204 -7364
rect 425604 -7366 426204 -7364
rect 461604 -7366 462204 -7364
rect 497604 -7366 498204 -7364
rect 533604 -7366 534204 -7364
rect 569604 -7366 570204 -7364
rect 591760 -7366 592360 -7364
use user_proj_example  mprj
timestamp 1607592090
transform 1 0 230000 0 1 340000
box 0 0 59856 60000
<< labels >>
rlabel metal3 s 583520 5796 584960 6036 6 analog_io[0]
port 0 nsew default bidirectional
rlabel metal3 s 583520 474996 584960 475236 6 analog_io[10]
port 1 nsew default bidirectional
rlabel metal3 s 583520 521916 584960 522156 6 analog_io[11]
port 2 nsew default bidirectional
rlabel metal3 s 583520 568836 584960 569076 6 analog_io[12]
port 3 nsew default bidirectional
rlabel metal3 s 583520 615756 584960 615996 6 analog_io[13]
port 4 nsew default bidirectional
rlabel metal3 s 583520 662676 584960 662916 6 analog_io[14]
port 5 nsew default bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[15]
port 6 nsew default bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[16]
port 7 nsew default bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[17]
port 8 nsew default bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[18]
port 9 nsew default bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[19]
port 10 nsew default bidirectional
rlabel metal3 s 583520 52716 584960 52956 6 analog_io[1]
port 11 nsew default bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[20]
port 12 nsew default bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[21]
port 13 nsew default bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[22]
port 14 nsew default bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[23]
port 15 nsew default bidirectional
rlabel metal3 s -960 696540 480 696780 4 analog_io[24]
port 16 nsew default bidirectional
rlabel metal3 s -960 639012 480 639252 4 analog_io[25]
port 17 nsew default bidirectional
rlabel metal3 s -960 581620 480 581860 4 analog_io[26]
port 18 nsew default bidirectional
rlabel metal3 s -960 524092 480 524332 4 analog_io[27]
port 19 nsew default bidirectional
rlabel metal3 s -960 466700 480 466940 4 analog_io[28]
port 20 nsew default bidirectional
rlabel metal3 s -960 409172 480 409412 4 analog_io[29]
port 21 nsew default bidirectional
rlabel metal3 s 583520 99636 584960 99876 6 analog_io[2]
port 22 nsew default bidirectional
rlabel metal3 s -960 351780 480 352020 4 analog_io[30]
port 23 nsew default bidirectional
rlabel metal3 s 583520 146556 584960 146796 6 analog_io[3]
port 24 nsew default bidirectional
rlabel metal3 s 583520 193476 584960 193716 6 analog_io[4]
port 25 nsew default bidirectional
rlabel metal3 s 583520 240396 584960 240636 6 analog_io[5]
port 26 nsew default bidirectional
rlabel metal3 s 583520 287316 584960 287556 6 analog_io[6]
port 27 nsew default bidirectional
rlabel metal3 s 583520 334236 584960 334476 6 analog_io[7]
port 28 nsew default bidirectional
rlabel metal3 s 583520 381156 584960 381396 6 analog_io[8]
port 29 nsew default bidirectional
rlabel metal3 s 583520 428076 584960 428316 6 analog_io[9]
port 30 nsew default bidirectional
rlabel metal3 s 583520 17492 584960 17732 6 io_in[0]
port 31 nsew default input
rlabel metal3 s 583520 486692 584960 486932 6 io_in[10]
port 32 nsew default input
rlabel metal3 s 583520 533748 584960 533988 6 io_in[11]
port 33 nsew default input
rlabel metal3 s 583520 580668 584960 580908 6 io_in[12]
port 34 nsew default input
rlabel metal3 s 583520 627588 584960 627828 6 io_in[13]
port 35 nsew default input
rlabel metal3 s 583520 674508 584960 674748 6 io_in[14]
port 36 nsew default input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 37 nsew default input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 38 nsew default input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 39 nsew default input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 40 nsew default input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 41 nsew default input
rlabel metal3 s 583520 64412 584960 64652 6 io_in[1]
port 42 nsew default input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 43 nsew default input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 44 nsew default input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 45 nsew default input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 46 nsew default input
rlabel metal3 s -960 682124 480 682364 4 io_in[24]
port 47 nsew default input
rlabel metal3 s -960 624732 480 624972 4 io_in[25]
port 48 nsew default input
rlabel metal3 s -960 567204 480 567444 4 io_in[26]
port 49 nsew default input
rlabel metal3 s -960 509812 480 510052 4 io_in[27]
port 50 nsew default input
rlabel metal3 s -960 452284 480 452524 4 io_in[28]
port 51 nsew default input
rlabel metal3 s -960 394892 480 395132 4 io_in[29]
port 52 nsew default input
rlabel metal3 s 583520 111332 584960 111572 6 io_in[2]
port 53 nsew default input
rlabel metal3 s -960 337364 480 337604 4 io_in[30]
port 54 nsew default input
rlabel metal3 s -960 294252 480 294492 4 io_in[31]
port 55 nsew default input
rlabel metal3 s -960 251140 480 251380 4 io_in[32]
port 56 nsew default input
rlabel metal3 s -960 208028 480 208268 4 io_in[33]
port 57 nsew default input
rlabel metal3 s -960 164916 480 165156 4 io_in[34]
port 58 nsew default input
rlabel metal3 s -960 121940 480 122180 4 io_in[35]
port 59 nsew default input
rlabel metal3 s -960 78828 480 79068 4 io_in[36]
port 60 nsew default input
rlabel metal3 s -960 35716 480 35956 4 io_in[37]
port 61 nsew default input
rlabel metal3 s 583520 158252 584960 158492 6 io_in[3]
port 62 nsew default input
rlabel metal3 s 583520 205172 584960 205412 6 io_in[4]
port 63 nsew default input
rlabel metal3 s 583520 252092 584960 252332 6 io_in[5]
port 64 nsew default input
rlabel metal3 s 583520 299012 584960 299252 6 io_in[6]
port 65 nsew default input
rlabel metal3 s 583520 345932 584960 346172 6 io_in[7]
port 66 nsew default input
rlabel metal3 s 583520 392852 584960 393092 6 io_in[8]
port 67 nsew default input
rlabel metal3 s 583520 439772 584960 440012 6 io_in[9]
port 68 nsew default input
rlabel metal3 s 583520 40884 584960 41124 6 io_oeb[0]
port 69 nsew default tristate
rlabel metal3 s 583520 510220 584960 510460 6 io_oeb[10]
port 70 nsew default tristate
rlabel metal3 s 583520 557140 584960 557380 6 io_oeb[11]
port 71 nsew default tristate
rlabel metal3 s 583520 604060 584960 604300 6 io_oeb[12]
port 72 nsew default tristate
rlabel metal3 s 583520 650980 584960 651220 6 io_oeb[13]
port 73 nsew default tristate
rlabel metal3 s 583520 697900 584960 698140 6 io_oeb[14]
port 74 nsew default tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 75 nsew default tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 76 nsew default tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 77 nsew default tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 78 nsew default tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 79 nsew default tristate
rlabel metal3 s 583520 87804 584960 88044 6 io_oeb[1]
port 80 nsew default tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 81 nsew default tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 82 nsew default tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 83 nsew default tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 84 nsew default tristate
rlabel metal3 s -960 653428 480 653668 4 io_oeb[24]
port 85 nsew default tristate
rlabel metal3 s -960 595900 480 596140 4 io_oeb[25]
port 86 nsew default tristate
rlabel metal3 s -960 538508 480 538748 4 io_oeb[26]
port 87 nsew default tristate
rlabel metal3 s -960 480980 480 481220 4 io_oeb[27]
port 88 nsew default tristate
rlabel metal3 s -960 423588 480 423828 4 io_oeb[28]
port 89 nsew default tristate
rlabel metal3 s -960 366060 480 366300 4 io_oeb[29]
port 90 nsew default tristate
rlabel metal3 s 583520 134724 584960 134964 6 io_oeb[2]
port 91 nsew default tristate
rlabel metal3 s -960 308668 480 308908 4 io_oeb[30]
port 92 nsew default tristate
rlabel metal3 s -960 265556 480 265796 4 io_oeb[31]
port 93 nsew default tristate
rlabel metal3 s -960 222444 480 222684 4 io_oeb[32]
port 94 nsew default tristate
rlabel metal3 s -960 179332 480 179572 4 io_oeb[33]
port 95 nsew default tristate
rlabel metal3 s -960 136220 480 136460 4 io_oeb[34]
port 96 nsew default tristate
rlabel metal3 s -960 93108 480 93348 4 io_oeb[35]
port 97 nsew default tristate
rlabel metal3 s -960 49996 480 50236 4 io_oeb[36]
port 98 nsew default tristate
rlabel metal3 s -960 7020 480 7260 4 io_oeb[37]
port 99 nsew default tristate
rlabel metal3 s 583520 181780 584960 182020 6 io_oeb[3]
port 100 nsew default tristate
rlabel metal3 s 583520 228700 584960 228940 6 io_oeb[4]
port 101 nsew default tristate
rlabel metal3 s 583520 275620 584960 275860 6 io_oeb[5]
port 102 nsew default tristate
rlabel metal3 s 583520 322540 584960 322780 6 io_oeb[6]
port 103 nsew default tristate
rlabel metal3 s 583520 369460 584960 369700 6 io_oeb[7]
port 104 nsew default tristate
rlabel metal3 s 583520 416380 584960 416620 6 io_oeb[8]
port 105 nsew default tristate
rlabel metal3 s 583520 463300 584960 463540 6 io_oeb[9]
port 106 nsew default tristate
rlabel metal3 s 583520 29188 584960 29428 6 io_out[0]
port 107 nsew default tristate
rlabel metal3 s 583520 498524 584960 498764 6 io_out[10]
port 108 nsew default tristate
rlabel metal3 s 583520 545444 584960 545684 6 io_out[11]
port 109 nsew default tristate
rlabel metal3 s 583520 592364 584960 592604 6 io_out[12]
port 110 nsew default tristate
rlabel metal3 s 583520 639284 584960 639524 6 io_out[13]
port 111 nsew default tristate
rlabel metal3 s 583520 686204 584960 686444 6 io_out[14]
port 112 nsew default tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 113 nsew default tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 114 nsew default tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 115 nsew default tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 116 nsew default tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 117 nsew default tristate
rlabel metal3 s 583520 76108 584960 76348 6 io_out[1]
port 118 nsew default tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 119 nsew default tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 120 nsew default tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 121 nsew default tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 122 nsew default tristate
rlabel metal3 s -960 667844 480 668084 4 io_out[24]
port 123 nsew default tristate
rlabel metal3 s -960 610316 480 610556 4 io_out[25]
port 124 nsew default tristate
rlabel metal3 s -960 552924 480 553164 4 io_out[26]
port 125 nsew default tristate
rlabel metal3 s -960 495396 480 495636 4 io_out[27]
port 126 nsew default tristate
rlabel metal3 s -960 437868 480 438108 4 io_out[28]
port 127 nsew default tristate
rlabel metal3 s -960 380476 480 380716 4 io_out[29]
port 128 nsew default tristate
rlabel metal3 s 583520 123028 584960 123268 6 io_out[2]
port 129 nsew default tristate
rlabel metal3 s -960 322948 480 323188 4 io_out[30]
port 130 nsew default tristate
rlabel metal3 s -960 279972 480 280212 4 io_out[31]
port 131 nsew default tristate
rlabel metal3 s -960 236860 480 237100 4 io_out[32]
port 132 nsew default tristate
rlabel metal3 s -960 193748 480 193988 4 io_out[33]
port 133 nsew default tristate
rlabel metal3 s -960 150636 480 150876 4 io_out[34]
port 134 nsew default tristate
rlabel metal3 s -960 107524 480 107764 4 io_out[35]
port 135 nsew default tristate
rlabel metal3 s -960 64412 480 64652 4 io_out[36]
port 136 nsew default tristate
rlabel metal3 s -960 21300 480 21540 4 io_out[37]
port 137 nsew default tristate
rlabel metal3 s 583520 169948 584960 170188 6 io_out[3]
port 138 nsew default tristate
rlabel metal3 s 583520 216868 584960 217108 6 io_out[4]
port 139 nsew default tristate
rlabel metal3 s 583520 263788 584960 264028 6 io_out[5]
port 140 nsew default tristate
rlabel metal3 s 583520 310708 584960 310948 6 io_out[6]
port 141 nsew default tristate
rlabel metal3 s 583520 357764 584960 358004 6 io_out[7]
port 142 nsew default tristate
rlabel metal3 s 583520 404684 584960 404924 6 io_out[8]
port 143 nsew default tristate
rlabel metal3 s 583520 451604 584960 451844 6 io_out[9]
port 144 nsew default tristate
rlabel metal2 s 126582 -960 126694 480 8 la_data_in[0]
port 145 nsew default input
rlabel metal2 s 483450 -960 483562 480 8 la_data_in[100]
port 146 nsew default input
rlabel metal2 s 486946 -960 487058 480 8 la_data_in[101]
port 147 nsew default input
rlabel metal2 s 490534 -960 490646 480 8 la_data_in[102]
port 148 nsew default input
rlabel metal2 s 494122 -960 494234 480 8 la_data_in[103]
port 149 nsew default input
rlabel metal2 s 497710 -960 497822 480 8 la_data_in[104]
port 150 nsew default input
rlabel metal2 s 501206 -960 501318 480 8 la_data_in[105]
port 151 nsew default input
rlabel metal2 s 504794 -960 504906 480 8 la_data_in[106]
port 152 nsew default input
rlabel metal2 s 508382 -960 508494 480 8 la_data_in[107]
port 153 nsew default input
rlabel metal2 s 511970 -960 512082 480 8 la_data_in[108]
port 154 nsew default input
rlabel metal2 s 515558 -960 515670 480 8 la_data_in[109]
port 155 nsew default input
rlabel metal2 s 162278 -960 162390 480 8 la_data_in[10]
port 156 nsew default input
rlabel metal2 s 519054 -960 519166 480 8 la_data_in[110]
port 157 nsew default input
rlabel metal2 s 522642 -960 522754 480 8 la_data_in[111]
port 158 nsew default input
rlabel metal2 s 526230 -960 526342 480 8 la_data_in[112]
port 159 nsew default input
rlabel metal2 s 529818 -960 529930 480 8 la_data_in[113]
port 160 nsew default input
rlabel metal2 s 533406 -960 533518 480 8 la_data_in[114]
port 161 nsew default input
rlabel metal2 s 536902 -960 537014 480 8 la_data_in[115]
port 162 nsew default input
rlabel metal2 s 540490 -960 540602 480 8 la_data_in[116]
port 163 nsew default input
rlabel metal2 s 544078 -960 544190 480 8 la_data_in[117]
port 164 nsew default input
rlabel metal2 s 547666 -960 547778 480 8 la_data_in[118]
port 165 nsew default input
rlabel metal2 s 551162 -960 551274 480 8 la_data_in[119]
port 166 nsew default input
rlabel metal2 s 165866 -960 165978 480 8 la_data_in[11]
port 167 nsew default input
rlabel metal2 s 554750 -960 554862 480 8 la_data_in[120]
port 168 nsew default input
rlabel metal2 s 558338 -960 558450 480 8 la_data_in[121]
port 169 nsew default input
rlabel metal2 s 561926 -960 562038 480 8 la_data_in[122]
port 170 nsew default input
rlabel metal2 s 565514 -960 565626 480 8 la_data_in[123]
port 171 nsew default input
rlabel metal2 s 569010 -960 569122 480 8 la_data_in[124]
port 172 nsew default input
rlabel metal2 s 572598 -960 572710 480 8 la_data_in[125]
port 173 nsew default input
rlabel metal2 s 576186 -960 576298 480 8 la_data_in[126]
port 174 nsew default input
rlabel metal2 s 579774 -960 579886 480 8 la_data_in[127]
port 175 nsew default input
rlabel metal2 s 169362 -960 169474 480 8 la_data_in[12]
port 176 nsew default input
rlabel metal2 s 172950 -960 173062 480 8 la_data_in[13]
port 177 nsew default input
rlabel metal2 s 176538 -960 176650 480 8 la_data_in[14]
port 178 nsew default input
rlabel metal2 s 180126 -960 180238 480 8 la_data_in[15]
port 179 nsew default input
rlabel metal2 s 183714 -960 183826 480 8 la_data_in[16]
port 180 nsew default input
rlabel metal2 s 187210 -960 187322 480 8 la_data_in[17]
port 181 nsew default input
rlabel metal2 s 190798 -960 190910 480 8 la_data_in[18]
port 182 nsew default input
rlabel metal2 s 194386 -960 194498 480 8 la_data_in[19]
port 183 nsew default input
rlabel metal2 s 130170 -960 130282 480 8 la_data_in[1]
port 184 nsew default input
rlabel metal2 s 197974 -960 198086 480 8 la_data_in[20]
port 185 nsew default input
rlabel metal2 s 201470 -960 201582 480 8 la_data_in[21]
port 186 nsew default input
rlabel metal2 s 205058 -960 205170 480 8 la_data_in[22]
port 187 nsew default input
rlabel metal2 s 208646 -960 208758 480 8 la_data_in[23]
port 188 nsew default input
rlabel metal2 s 212234 -960 212346 480 8 la_data_in[24]
port 189 nsew default input
rlabel metal2 s 215822 -960 215934 480 8 la_data_in[25]
port 190 nsew default input
rlabel metal2 s 219318 -960 219430 480 8 la_data_in[26]
port 191 nsew default input
rlabel metal2 s 222906 -960 223018 480 8 la_data_in[27]
port 192 nsew default input
rlabel metal2 s 226494 -960 226606 480 8 la_data_in[28]
port 193 nsew default input
rlabel metal2 s 230082 -960 230194 480 8 la_data_in[29]
port 194 nsew default input
rlabel metal2 s 133758 -960 133870 480 8 la_data_in[2]
port 195 nsew default input
rlabel metal2 s 233670 -960 233782 480 8 la_data_in[30]
port 196 nsew default input
rlabel metal2 s 237166 -960 237278 480 8 la_data_in[31]
port 197 nsew default input
rlabel metal2 s 240754 -960 240866 480 8 la_data_in[32]
port 198 nsew default input
rlabel metal2 s 244342 -960 244454 480 8 la_data_in[33]
port 199 nsew default input
rlabel metal2 s 247930 -960 248042 480 8 la_data_in[34]
port 200 nsew default input
rlabel metal2 s 251426 -960 251538 480 8 la_data_in[35]
port 201 nsew default input
rlabel metal2 s 255014 -960 255126 480 8 la_data_in[36]
port 202 nsew default input
rlabel metal2 s 258602 -960 258714 480 8 la_data_in[37]
port 203 nsew default input
rlabel metal2 s 262190 -960 262302 480 8 la_data_in[38]
port 204 nsew default input
rlabel metal2 s 265778 -960 265890 480 8 la_data_in[39]
port 205 nsew default input
rlabel metal2 s 137254 -960 137366 480 8 la_data_in[3]
port 206 nsew default input
rlabel metal2 s 269274 -960 269386 480 8 la_data_in[40]
port 207 nsew default input
rlabel metal2 s 272862 -960 272974 480 8 la_data_in[41]
port 208 nsew default input
rlabel metal2 s 276450 -960 276562 480 8 la_data_in[42]
port 209 nsew default input
rlabel metal2 s 280038 -960 280150 480 8 la_data_in[43]
port 210 nsew default input
rlabel metal2 s 283626 -960 283738 480 8 la_data_in[44]
port 211 nsew default input
rlabel metal2 s 287122 -960 287234 480 8 la_data_in[45]
port 212 nsew default input
rlabel metal2 s 290710 -960 290822 480 8 la_data_in[46]
port 213 nsew default input
rlabel metal2 s 294298 -960 294410 480 8 la_data_in[47]
port 214 nsew default input
rlabel metal2 s 297886 -960 297998 480 8 la_data_in[48]
port 215 nsew default input
rlabel metal2 s 301382 -960 301494 480 8 la_data_in[49]
port 216 nsew default input
rlabel metal2 s 140842 -960 140954 480 8 la_data_in[4]
port 217 nsew default input
rlabel metal2 s 304970 -960 305082 480 8 la_data_in[50]
port 218 nsew default input
rlabel metal2 s 308558 -960 308670 480 8 la_data_in[51]
port 219 nsew default input
rlabel metal2 s 312146 -960 312258 480 8 la_data_in[52]
port 220 nsew default input
rlabel metal2 s 315734 -960 315846 480 8 la_data_in[53]
port 221 nsew default input
rlabel metal2 s 319230 -960 319342 480 8 la_data_in[54]
port 222 nsew default input
rlabel metal2 s 322818 -960 322930 480 8 la_data_in[55]
port 223 nsew default input
rlabel metal2 s 326406 -960 326518 480 8 la_data_in[56]
port 224 nsew default input
rlabel metal2 s 329994 -960 330106 480 8 la_data_in[57]
port 225 nsew default input
rlabel metal2 s 333582 -960 333694 480 8 la_data_in[58]
port 226 nsew default input
rlabel metal2 s 337078 -960 337190 480 8 la_data_in[59]
port 227 nsew default input
rlabel metal2 s 144430 -960 144542 480 8 la_data_in[5]
port 228 nsew default input
rlabel metal2 s 340666 -960 340778 480 8 la_data_in[60]
port 229 nsew default input
rlabel metal2 s 344254 -960 344366 480 8 la_data_in[61]
port 230 nsew default input
rlabel metal2 s 347842 -960 347954 480 8 la_data_in[62]
port 231 nsew default input
rlabel metal2 s 351338 -960 351450 480 8 la_data_in[63]
port 232 nsew default input
rlabel metal2 s 354926 -960 355038 480 8 la_data_in[64]
port 233 nsew default input
rlabel metal2 s 358514 -960 358626 480 8 la_data_in[65]
port 234 nsew default input
rlabel metal2 s 362102 -960 362214 480 8 la_data_in[66]
port 235 nsew default input
rlabel metal2 s 365690 -960 365802 480 8 la_data_in[67]
port 236 nsew default input
rlabel metal2 s 369186 -960 369298 480 8 la_data_in[68]
port 237 nsew default input
rlabel metal2 s 372774 -960 372886 480 8 la_data_in[69]
port 238 nsew default input
rlabel metal2 s 148018 -960 148130 480 8 la_data_in[6]
port 239 nsew default input
rlabel metal2 s 376362 -960 376474 480 8 la_data_in[70]
port 240 nsew default input
rlabel metal2 s 379950 -960 380062 480 8 la_data_in[71]
port 241 nsew default input
rlabel metal2 s 383538 -960 383650 480 8 la_data_in[72]
port 242 nsew default input
rlabel metal2 s 387034 -960 387146 480 8 la_data_in[73]
port 243 nsew default input
rlabel metal2 s 390622 -960 390734 480 8 la_data_in[74]
port 244 nsew default input
rlabel metal2 s 394210 -960 394322 480 8 la_data_in[75]
port 245 nsew default input
rlabel metal2 s 397798 -960 397910 480 8 la_data_in[76]
port 246 nsew default input
rlabel metal2 s 401294 -960 401406 480 8 la_data_in[77]
port 247 nsew default input
rlabel metal2 s 404882 -960 404994 480 8 la_data_in[78]
port 248 nsew default input
rlabel metal2 s 408470 -960 408582 480 8 la_data_in[79]
port 249 nsew default input
rlabel metal2 s 151514 -960 151626 480 8 la_data_in[7]
port 250 nsew default input
rlabel metal2 s 412058 -960 412170 480 8 la_data_in[80]
port 251 nsew default input
rlabel metal2 s 415646 -960 415758 480 8 la_data_in[81]
port 252 nsew default input
rlabel metal2 s 419142 -960 419254 480 8 la_data_in[82]
port 253 nsew default input
rlabel metal2 s 422730 -960 422842 480 8 la_data_in[83]
port 254 nsew default input
rlabel metal2 s 426318 -960 426430 480 8 la_data_in[84]
port 255 nsew default input
rlabel metal2 s 429906 -960 430018 480 8 la_data_in[85]
port 256 nsew default input
rlabel metal2 s 433494 -960 433606 480 8 la_data_in[86]
port 257 nsew default input
rlabel metal2 s 436990 -960 437102 480 8 la_data_in[87]
port 258 nsew default input
rlabel metal2 s 440578 -960 440690 480 8 la_data_in[88]
port 259 nsew default input
rlabel metal2 s 444166 -960 444278 480 8 la_data_in[89]
port 260 nsew default input
rlabel metal2 s 155102 -960 155214 480 8 la_data_in[8]
port 261 nsew default input
rlabel metal2 s 447754 -960 447866 480 8 la_data_in[90]
port 262 nsew default input
rlabel metal2 s 451250 -960 451362 480 8 la_data_in[91]
port 263 nsew default input
rlabel metal2 s 454838 -960 454950 480 8 la_data_in[92]
port 264 nsew default input
rlabel metal2 s 458426 -960 458538 480 8 la_data_in[93]
port 265 nsew default input
rlabel metal2 s 462014 -960 462126 480 8 la_data_in[94]
port 266 nsew default input
rlabel metal2 s 465602 -960 465714 480 8 la_data_in[95]
port 267 nsew default input
rlabel metal2 s 469098 -960 469210 480 8 la_data_in[96]
port 268 nsew default input
rlabel metal2 s 472686 -960 472798 480 8 la_data_in[97]
port 269 nsew default input
rlabel metal2 s 476274 -960 476386 480 8 la_data_in[98]
port 270 nsew default input
rlabel metal2 s 479862 -960 479974 480 8 la_data_in[99]
port 271 nsew default input
rlabel metal2 s 158690 -960 158802 480 8 la_data_in[9]
port 272 nsew default input
rlabel metal2 s 127778 -960 127890 480 8 la_data_out[0]
port 273 nsew default tristate
rlabel metal2 s 484554 -960 484666 480 8 la_data_out[100]
port 274 nsew default tristate
rlabel metal2 s 488142 -960 488254 480 8 la_data_out[101]
port 275 nsew default tristate
rlabel metal2 s 491730 -960 491842 480 8 la_data_out[102]
port 276 nsew default tristate
rlabel metal2 s 495318 -960 495430 480 8 la_data_out[103]
port 277 nsew default tristate
rlabel metal2 s 498906 -960 499018 480 8 la_data_out[104]
port 278 nsew default tristate
rlabel metal2 s 502402 -960 502514 480 8 la_data_out[105]
port 279 nsew default tristate
rlabel metal2 s 505990 -960 506102 480 8 la_data_out[106]
port 280 nsew default tristate
rlabel metal2 s 509578 -960 509690 480 8 la_data_out[107]
port 281 nsew default tristate
rlabel metal2 s 513166 -960 513278 480 8 la_data_out[108]
port 282 nsew default tristate
rlabel metal2 s 516754 -960 516866 480 8 la_data_out[109]
port 283 nsew default tristate
rlabel metal2 s 163474 -960 163586 480 8 la_data_out[10]
port 284 nsew default tristate
rlabel metal2 s 520250 -960 520362 480 8 la_data_out[110]
port 285 nsew default tristate
rlabel metal2 s 523838 -960 523950 480 8 la_data_out[111]
port 286 nsew default tristate
rlabel metal2 s 527426 -960 527538 480 8 la_data_out[112]
port 287 nsew default tristate
rlabel metal2 s 531014 -960 531126 480 8 la_data_out[113]
port 288 nsew default tristate
rlabel metal2 s 534510 -960 534622 480 8 la_data_out[114]
port 289 nsew default tristate
rlabel metal2 s 538098 -960 538210 480 8 la_data_out[115]
port 290 nsew default tristate
rlabel metal2 s 541686 -960 541798 480 8 la_data_out[116]
port 291 nsew default tristate
rlabel metal2 s 545274 -960 545386 480 8 la_data_out[117]
port 292 nsew default tristate
rlabel metal2 s 548862 -960 548974 480 8 la_data_out[118]
port 293 nsew default tristate
rlabel metal2 s 552358 -960 552470 480 8 la_data_out[119]
port 294 nsew default tristate
rlabel metal2 s 167062 -960 167174 480 8 la_data_out[11]
port 295 nsew default tristate
rlabel metal2 s 555946 -960 556058 480 8 la_data_out[120]
port 296 nsew default tristate
rlabel metal2 s 559534 -960 559646 480 8 la_data_out[121]
port 297 nsew default tristate
rlabel metal2 s 563122 -960 563234 480 8 la_data_out[122]
port 298 nsew default tristate
rlabel metal2 s 566710 -960 566822 480 8 la_data_out[123]
port 299 nsew default tristate
rlabel metal2 s 570206 -960 570318 480 8 la_data_out[124]
port 300 nsew default tristate
rlabel metal2 s 573794 -960 573906 480 8 la_data_out[125]
port 301 nsew default tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[126]
port 302 nsew default tristate
rlabel metal2 s 580970 -960 581082 480 8 la_data_out[127]
port 303 nsew default tristate
rlabel metal2 s 170558 -960 170670 480 8 la_data_out[12]
port 304 nsew default tristate
rlabel metal2 s 174146 -960 174258 480 8 la_data_out[13]
port 305 nsew default tristate
rlabel metal2 s 177734 -960 177846 480 8 la_data_out[14]
port 306 nsew default tristate
rlabel metal2 s 181322 -960 181434 480 8 la_data_out[15]
port 307 nsew default tristate
rlabel metal2 s 184818 -960 184930 480 8 la_data_out[16]
port 308 nsew default tristate
rlabel metal2 s 188406 -960 188518 480 8 la_data_out[17]
port 309 nsew default tristate
rlabel metal2 s 191994 -960 192106 480 8 la_data_out[18]
port 310 nsew default tristate
rlabel metal2 s 195582 -960 195694 480 8 la_data_out[19]
port 311 nsew default tristate
rlabel metal2 s 131366 -960 131478 480 8 la_data_out[1]
port 312 nsew default tristate
rlabel metal2 s 199170 -960 199282 480 8 la_data_out[20]
port 313 nsew default tristate
rlabel metal2 s 202666 -960 202778 480 8 la_data_out[21]
port 314 nsew default tristate
rlabel metal2 s 206254 -960 206366 480 8 la_data_out[22]
port 315 nsew default tristate
rlabel metal2 s 209842 -960 209954 480 8 la_data_out[23]
port 316 nsew default tristate
rlabel metal2 s 213430 -960 213542 480 8 la_data_out[24]
port 317 nsew default tristate
rlabel metal2 s 217018 -960 217130 480 8 la_data_out[25]
port 318 nsew default tristate
rlabel metal2 s 220514 -960 220626 480 8 la_data_out[26]
port 319 nsew default tristate
rlabel metal2 s 224102 -960 224214 480 8 la_data_out[27]
port 320 nsew default tristate
rlabel metal2 s 227690 -960 227802 480 8 la_data_out[28]
port 321 nsew default tristate
rlabel metal2 s 231278 -960 231390 480 8 la_data_out[29]
port 322 nsew default tristate
rlabel metal2 s 134862 -960 134974 480 8 la_data_out[2]
port 323 nsew default tristate
rlabel metal2 s 234774 -960 234886 480 8 la_data_out[30]
port 324 nsew default tristate
rlabel metal2 s 238362 -960 238474 480 8 la_data_out[31]
port 325 nsew default tristate
rlabel metal2 s 241950 -960 242062 480 8 la_data_out[32]
port 326 nsew default tristate
rlabel metal2 s 245538 -960 245650 480 8 la_data_out[33]
port 327 nsew default tristate
rlabel metal2 s 249126 -960 249238 480 8 la_data_out[34]
port 328 nsew default tristate
rlabel metal2 s 252622 -960 252734 480 8 la_data_out[35]
port 329 nsew default tristate
rlabel metal2 s 256210 -960 256322 480 8 la_data_out[36]
port 330 nsew default tristate
rlabel metal2 s 259798 -960 259910 480 8 la_data_out[37]
port 331 nsew default tristate
rlabel metal2 s 263386 -960 263498 480 8 la_data_out[38]
port 332 nsew default tristate
rlabel metal2 s 266974 -960 267086 480 8 la_data_out[39]
port 333 nsew default tristate
rlabel metal2 s 138450 -960 138562 480 8 la_data_out[3]
port 334 nsew default tristate
rlabel metal2 s 270470 -960 270582 480 8 la_data_out[40]
port 335 nsew default tristate
rlabel metal2 s 274058 -960 274170 480 8 la_data_out[41]
port 336 nsew default tristate
rlabel metal2 s 277646 -960 277758 480 8 la_data_out[42]
port 337 nsew default tristate
rlabel metal2 s 281234 -960 281346 480 8 la_data_out[43]
port 338 nsew default tristate
rlabel metal2 s 284730 -960 284842 480 8 la_data_out[44]
port 339 nsew default tristate
rlabel metal2 s 288318 -960 288430 480 8 la_data_out[45]
port 340 nsew default tristate
rlabel metal2 s 291906 -960 292018 480 8 la_data_out[46]
port 341 nsew default tristate
rlabel metal2 s 295494 -960 295606 480 8 la_data_out[47]
port 342 nsew default tristate
rlabel metal2 s 299082 -960 299194 480 8 la_data_out[48]
port 343 nsew default tristate
rlabel metal2 s 302578 -960 302690 480 8 la_data_out[49]
port 344 nsew default tristate
rlabel metal2 s 142038 -960 142150 480 8 la_data_out[4]
port 345 nsew default tristate
rlabel metal2 s 306166 -960 306278 480 8 la_data_out[50]
port 346 nsew default tristate
rlabel metal2 s 309754 -960 309866 480 8 la_data_out[51]
port 347 nsew default tristate
rlabel metal2 s 313342 -960 313454 480 8 la_data_out[52]
port 348 nsew default tristate
rlabel metal2 s 316930 -960 317042 480 8 la_data_out[53]
port 349 nsew default tristate
rlabel metal2 s 320426 -960 320538 480 8 la_data_out[54]
port 350 nsew default tristate
rlabel metal2 s 324014 -960 324126 480 8 la_data_out[55]
port 351 nsew default tristate
rlabel metal2 s 327602 -960 327714 480 8 la_data_out[56]
port 352 nsew default tristate
rlabel metal2 s 331190 -960 331302 480 8 la_data_out[57]
port 353 nsew default tristate
rlabel metal2 s 334686 -960 334798 480 8 la_data_out[58]
port 354 nsew default tristate
rlabel metal2 s 338274 -960 338386 480 8 la_data_out[59]
port 355 nsew default tristate
rlabel metal2 s 145626 -960 145738 480 8 la_data_out[5]
port 356 nsew default tristate
rlabel metal2 s 341862 -960 341974 480 8 la_data_out[60]
port 357 nsew default tristate
rlabel metal2 s 345450 -960 345562 480 8 la_data_out[61]
port 358 nsew default tristate
rlabel metal2 s 349038 -960 349150 480 8 la_data_out[62]
port 359 nsew default tristate
rlabel metal2 s 352534 -960 352646 480 8 la_data_out[63]
port 360 nsew default tristate
rlabel metal2 s 356122 -960 356234 480 8 la_data_out[64]
port 361 nsew default tristate
rlabel metal2 s 359710 -960 359822 480 8 la_data_out[65]
port 362 nsew default tristate
rlabel metal2 s 363298 -960 363410 480 8 la_data_out[66]
port 363 nsew default tristate
rlabel metal2 s 366886 -960 366998 480 8 la_data_out[67]
port 364 nsew default tristate
rlabel metal2 s 370382 -960 370494 480 8 la_data_out[68]
port 365 nsew default tristate
rlabel metal2 s 373970 -960 374082 480 8 la_data_out[69]
port 366 nsew default tristate
rlabel metal2 s 149214 -960 149326 480 8 la_data_out[6]
port 367 nsew default tristate
rlabel metal2 s 377558 -960 377670 480 8 la_data_out[70]
port 368 nsew default tristate
rlabel metal2 s 381146 -960 381258 480 8 la_data_out[71]
port 369 nsew default tristate
rlabel metal2 s 384642 -960 384754 480 8 la_data_out[72]
port 370 nsew default tristate
rlabel metal2 s 388230 -960 388342 480 8 la_data_out[73]
port 371 nsew default tristate
rlabel metal2 s 391818 -960 391930 480 8 la_data_out[74]
port 372 nsew default tristate
rlabel metal2 s 395406 -960 395518 480 8 la_data_out[75]
port 373 nsew default tristate
rlabel metal2 s 398994 -960 399106 480 8 la_data_out[76]
port 374 nsew default tristate
rlabel metal2 s 402490 -960 402602 480 8 la_data_out[77]
port 375 nsew default tristate
rlabel metal2 s 406078 -960 406190 480 8 la_data_out[78]
port 376 nsew default tristate
rlabel metal2 s 409666 -960 409778 480 8 la_data_out[79]
port 377 nsew default tristate
rlabel metal2 s 152710 -960 152822 480 8 la_data_out[7]
port 378 nsew default tristate
rlabel metal2 s 413254 -960 413366 480 8 la_data_out[80]
port 379 nsew default tristate
rlabel metal2 s 416842 -960 416954 480 8 la_data_out[81]
port 380 nsew default tristate
rlabel metal2 s 420338 -960 420450 480 8 la_data_out[82]
port 381 nsew default tristate
rlabel metal2 s 423926 -960 424038 480 8 la_data_out[83]
port 382 nsew default tristate
rlabel metal2 s 427514 -960 427626 480 8 la_data_out[84]
port 383 nsew default tristate
rlabel metal2 s 431102 -960 431214 480 8 la_data_out[85]
port 384 nsew default tristate
rlabel metal2 s 434598 -960 434710 480 8 la_data_out[86]
port 385 nsew default tristate
rlabel metal2 s 438186 -960 438298 480 8 la_data_out[87]
port 386 nsew default tristate
rlabel metal2 s 441774 -960 441886 480 8 la_data_out[88]
port 387 nsew default tristate
rlabel metal2 s 445362 -960 445474 480 8 la_data_out[89]
port 388 nsew default tristate
rlabel metal2 s 156298 -960 156410 480 8 la_data_out[8]
port 389 nsew default tristate
rlabel metal2 s 448950 -960 449062 480 8 la_data_out[90]
port 390 nsew default tristate
rlabel metal2 s 452446 -960 452558 480 8 la_data_out[91]
port 391 nsew default tristate
rlabel metal2 s 456034 -960 456146 480 8 la_data_out[92]
port 392 nsew default tristate
rlabel metal2 s 459622 -960 459734 480 8 la_data_out[93]
port 393 nsew default tristate
rlabel metal2 s 463210 -960 463322 480 8 la_data_out[94]
port 394 nsew default tristate
rlabel metal2 s 466798 -960 466910 480 8 la_data_out[95]
port 395 nsew default tristate
rlabel metal2 s 470294 -960 470406 480 8 la_data_out[96]
port 396 nsew default tristate
rlabel metal2 s 473882 -960 473994 480 8 la_data_out[97]
port 397 nsew default tristate
rlabel metal2 s 477470 -960 477582 480 8 la_data_out[98]
port 398 nsew default tristate
rlabel metal2 s 481058 -960 481170 480 8 la_data_out[99]
port 399 nsew default tristate
rlabel metal2 s 159886 -960 159998 480 8 la_data_out[9]
port 400 nsew default tristate
rlabel metal2 s 128974 -960 129086 480 8 la_oen[0]
port 401 nsew default input
rlabel metal2 s 485750 -960 485862 480 8 la_oen[100]
port 402 nsew default input
rlabel metal2 s 489338 -960 489450 480 8 la_oen[101]
port 403 nsew default input
rlabel metal2 s 492926 -960 493038 480 8 la_oen[102]
port 404 nsew default input
rlabel metal2 s 496514 -960 496626 480 8 la_oen[103]
port 405 nsew default input
rlabel metal2 s 500102 -960 500214 480 8 la_oen[104]
port 406 nsew default input
rlabel metal2 s 503598 -960 503710 480 8 la_oen[105]
port 407 nsew default input
rlabel metal2 s 507186 -960 507298 480 8 la_oen[106]
port 408 nsew default input
rlabel metal2 s 510774 -960 510886 480 8 la_oen[107]
port 409 nsew default input
rlabel metal2 s 514362 -960 514474 480 8 la_oen[108]
port 410 nsew default input
rlabel metal2 s 517858 -960 517970 480 8 la_oen[109]
port 411 nsew default input
rlabel metal2 s 164670 -960 164782 480 8 la_oen[10]
port 412 nsew default input
rlabel metal2 s 521446 -960 521558 480 8 la_oen[110]
port 413 nsew default input
rlabel metal2 s 525034 -960 525146 480 8 la_oen[111]
port 414 nsew default input
rlabel metal2 s 528622 -960 528734 480 8 la_oen[112]
port 415 nsew default input
rlabel metal2 s 532210 -960 532322 480 8 la_oen[113]
port 416 nsew default input
rlabel metal2 s 535706 -960 535818 480 8 la_oen[114]
port 417 nsew default input
rlabel metal2 s 539294 -960 539406 480 8 la_oen[115]
port 418 nsew default input
rlabel metal2 s 542882 -960 542994 480 8 la_oen[116]
port 419 nsew default input
rlabel metal2 s 546470 -960 546582 480 8 la_oen[117]
port 420 nsew default input
rlabel metal2 s 550058 -960 550170 480 8 la_oen[118]
port 421 nsew default input
rlabel metal2 s 553554 -960 553666 480 8 la_oen[119]
port 422 nsew default input
rlabel metal2 s 168166 -960 168278 480 8 la_oen[11]
port 423 nsew default input
rlabel metal2 s 557142 -960 557254 480 8 la_oen[120]
port 424 nsew default input
rlabel metal2 s 560730 -960 560842 480 8 la_oen[121]
port 425 nsew default input
rlabel metal2 s 564318 -960 564430 480 8 la_oen[122]
port 426 nsew default input
rlabel metal2 s 567814 -960 567926 480 8 la_oen[123]
port 427 nsew default input
rlabel metal2 s 571402 -960 571514 480 8 la_oen[124]
port 428 nsew default input
rlabel metal2 s 574990 -960 575102 480 8 la_oen[125]
port 429 nsew default input
rlabel metal2 s 578578 -960 578690 480 8 la_oen[126]
port 430 nsew default input
rlabel metal2 s 582166 -960 582278 480 8 la_oen[127]
port 431 nsew default input
rlabel metal2 s 171754 -960 171866 480 8 la_oen[12]
port 432 nsew default input
rlabel metal2 s 175342 -960 175454 480 8 la_oen[13]
port 433 nsew default input
rlabel metal2 s 178930 -960 179042 480 8 la_oen[14]
port 434 nsew default input
rlabel metal2 s 182518 -960 182630 480 8 la_oen[15]
port 435 nsew default input
rlabel metal2 s 186014 -960 186126 480 8 la_oen[16]
port 436 nsew default input
rlabel metal2 s 189602 -960 189714 480 8 la_oen[17]
port 437 nsew default input
rlabel metal2 s 193190 -960 193302 480 8 la_oen[18]
port 438 nsew default input
rlabel metal2 s 196778 -960 196890 480 8 la_oen[19]
port 439 nsew default input
rlabel metal2 s 132562 -960 132674 480 8 la_oen[1]
port 440 nsew default input
rlabel metal2 s 200366 -960 200478 480 8 la_oen[20]
port 441 nsew default input
rlabel metal2 s 203862 -960 203974 480 8 la_oen[21]
port 442 nsew default input
rlabel metal2 s 207450 -960 207562 480 8 la_oen[22]
port 443 nsew default input
rlabel metal2 s 211038 -960 211150 480 8 la_oen[23]
port 444 nsew default input
rlabel metal2 s 214626 -960 214738 480 8 la_oen[24]
port 445 nsew default input
rlabel metal2 s 218122 -960 218234 480 8 la_oen[25]
port 446 nsew default input
rlabel metal2 s 221710 -960 221822 480 8 la_oen[26]
port 447 nsew default input
rlabel metal2 s 225298 -960 225410 480 8 la_oen[27]
port 448 nsew default input
rlabel metal2 s 228886 -960 228998 480 8 la_oen[28]
port 449 nsew default input
rlabel metal2 s 232474 -960 232586 480 8 la_oen[29]
port 450 nsew default input
rlabel metal2 s 136058 -960 136170 480 8 la_oen[2]
port 451 nsew default input
rlabel metal2 s 235970 -960 236082 480 8 la_oen[30]
port 452 nsew default input
rlabel metal2 s 239558 -960 239670 480 8 la_oen[31]
port 453 nsew default input
rlabel metal2 s 243146 -960 243258 480 8 la_oen[32]
port 454 nsew default input
rlabel metal2 s 246734 -960 246846 480 8 la_oen[33]
port 455 nsew default input
rlabel metal2 s 250322 -960 250434 480 8 la_oen[34]
port 456 nsew default input
rlabel metal2 s 253818 -960 253930 480 8 la_oen[35]
port 457 nsew default input
rlabel metal2 s 257406 -960 257518 480 8 la_oen[36]
port 458 nsew default input
rlabel metal2 s 260994 -960 261106 480 8 la_oen[37]
port 459 nsew default input
rlabel metal2 s 264582 -960 264694 480 8 la_oen[38]
port 460 nsew default input
rlabel metal2 s 268078 -960 268190 480 8 la_oen[39]
port 461 nsew default input
rlabel metal2 s 139646 -960 139758 480 8 la_oen[3]
port 462 nsew default input
rlabel metal2 s 271666 -960 271778 480 8 la_oen[40]
port 463 nsew default input
rlabel metal2 s 275254 -960 275366 480 8 la_oen[41]
port 464 nsew default input
rlabel metal2 s 278842 -960 278954 480 8 la_oen[42]
port 465 nsew default input
rlabel metal2 s 282430 -960 282542 480 8 la_oen[43]
port 466 nsew default input
rlabel metal2 s 285926 -960 286038 480 8 la_oen[44]
port 467 nsew default input
rlabel metal2 s 289514 -960 289626 480 8 la_oen[45]
port 468 nsew default input
rlabel metal2 s 293102 -960 293214 480 8 la_oen[46]
port 469 nsew default input
rlabel metal2 s 296690 -960 296802 480 8 la_oen[47]
port 470 nsew default input
rlabel metal2 s 300278 -960 300390 480 8 la_oen[48]
port 471 nsew default input
rlabel metal2 s 303774 -960 303886 480 8 la_oen[49]
port 472 nsew default input
rlabel metal2 s 143234 -960 143346 480 8 la_oen[4]
port 473 nsew default input
rlabel metal2 s 307362 -960 307474 480 8 la_oen[50]
port 474 nsew default input
rlabel metal2 s 310950 -960 311062 480 8 la_oen[51]
port 475 nsew default input
rlabel metal2 s 314538 -960 314650 480 8 la_oen[52]
port 476 nsew default input
rlabel metal2 s 318034 -960 318146 480 8 la_oen[53]
port 477 nsew default input
rlabel metal2 s 321622 -960 321734 480 8 la_oen[54]
port 478 nsew default input
rlabel metal2 s 325210 -960 325322 480 8 la_oen[55]
port 479 nsew default input
rlabel metal2 s 328798 -960 328910 480 8 la_oen[56]
port 480 nsew default input
rlabel metal2 s 332386 -960 332498 480 8 la_oen[57]
port 481 nsew default input
rlabel metal2 s 335882 -960 335994 480 8 la_oen[58]
port 482 nsew default input
rlabel metal2 s 339470 -960 339582 480 8 la_oen[59]
port 483 nsew default input
rlabel metal2 s 146822 -960 146934 480 8 la_oen[5]
port 484 nsew default input
rlabel metal2 s 343058 -960 343170 480 8 la_oen[60]
port 485 nsew default input
rlabel metal2 s 346646 -960 346758 480 8 la_oen[61]
port 486 nsew default input
rlabel metal2 s 350234 -960 350346 480 8 la_oen[62]
port 487 nsew default input
rlabel metal2 s 353730 -960 353842 480 8 la_oen[63]
port 488 nsew default input
rlabel metal2 s 357318 -960 357430 480 8 la_oen[64]
port 489 nsew default input
rlabel metal2 s 360906 -960 361018 480 8 la_oen[65]
port 490 nsew default input
rlabel metal2 s 364494 -960 364606 480 8 la_oen[66]
port 491 nsew default input
rlabel metal2 s 367990 -960 368102 480 8 la_oen[67]
port 492 nsew default input
rlabel metal2 s 371578 -960 371690 480 8 la_oen[68]
port 493 nsew default input
rlabel metal2 s 375166 -960 375278 480 8 la_oen[69]
port 494 nsew default input
rlabel metal2 s 150410 -960 150522 480 8 la_oen[6]
port 495 nsew default input
rlabel metal2 s 378754 -960 378866 480 8 la_oen[70]
port 496 nsew default input
rlabel metal2 s 382342 -960 382454 480 8 la_oen[71]
port 497 nsew default input
rlabel metal2 s 385838 -960 385950 480 8 la_oen[72]
port 498 nsew default input
rlabel metal2 s 389426 -960 389538 480 8 la_oen[73]
port 499 nsew default input
rlabel metal2 s 393014 -960 393126 480 8 la_oen[74]
port 500 nsew default input
rlabel metal2 s 396602 -960 396714 480 8 la_oen[75]
port 501 nsew default input
rlabel metal2 s 400190 -960 400302 480 8 la_oen[76]
port 502 nsew default input
rlabel metal2 s 403686 -960 403798 480 8 la_oen[77]
port 503 nsew default input
rlabel metal2 s 407274 -960 407386 480 8 la_oen[78]
port 504 nsew default input
rlabel metal2 s 410862 -960 410974 480 8 la_oen[79]
port 505 nsew default input
rlabel metal2 s 153906 -960 154018 480 8 la_oen[7]
port 506 nsew default input
rlabel metal2 s 414450 -960 414562 480 8 la_oen[80]
port 507 nsew default input
rlabel metal2 s 417946 -960 418058 480 8 la_oen[81]
port 508 nsew default input
rlabel metal2 s 421534 -960 421646 480 8 la_oen[82]
port 509 nsew default input
rlabel metal2 s 425122 -960 425234 480 8 la_oen[83]
port 510 nsew default input
rlabel metal2 s 428710 -960 428822 480 8 la_oen[84]
port 511 nsew default input
rlabel metal2 s 432298 -960 432410 480 8 la_oen[85]
port 512 nsew default input
rlabel metal2 s 435794 -960 435906 480 8 la_oen[86]
port 513 nsew default input
rlabel metal2 s 439382 -960 439494 480 8 la_oen[87]
port 514 nsew default input
rlabel metal2 s 442970 -960 443082 480 8 la_oen[88]
port 515 nsew default input
rlabel metal2 s 446558 -960 446670 480 8 la_oen[89]
port 516 nsew default input
rlabel metal2 s 157494 -960 157606 480 8 la_oen[8]
port 517 nsew default input
rlabel metal2 s 450146 -960 450258 480 8 la_oen[90]
port 518 nsew default input
rlabel metal2 s 453642 -960 453754 480 8 la_oen[91]
port 519 nsew default input
rlabel metal2 s 457230 -960 457342 480 8 la_oen[92]
port 520 nsew default input
rlabel metal2 s 460818 -960 460930 480 8 la_oen[93]
port 521 nsew default input
rlabel metal2 s 464406 -960 464518 480 8 la_oen[94]
port 522 nsew default input
rlabel metal2 s 467902 -960 468014 480 8 la_oen[95]
port 523 nsew default input
rlabel metal2 s 471490 -960 471602 480 8 la_oen[96]
port 524 nsew default input
rlabel metal2 s 475078 -960 475190 480 8 la_oen[97]
port 525 nsew default input
rlabel metal2 s 478666 -960 478778 480 8 la_oen[98]
port 526 nsew default input
rlabel metal2 s 482254 -960 482366 480 8 la_oen[99]
port 527 nsew default input
rlabel metal2 s 161082 -960 161194 480 8 la_oen[9]
port 528 nsew default input
rlabel metal2 s 583362 -960 583474 480 8 user_clock2
port 529 nsew default input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 530 nsew default input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 531 nsew default input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 532 nsew default tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 533 nsew default input
rlabel metal2 s 48106 -960 48218 480 8 wbs_adr_i[10]
port 534 nsew default input
rlabel metal2 s 51602 -960 51714 480 8 wbs_adr_i[11]
port 535 nsew default input
rlabel metal2 s 55190 -960 55302 480 8 wbs_adr_i[12]
port 536 nsew default input
rlabel metal2 s 58778 -960 58890 480 8 wbs_adr_i[13]
port 537 nsew default input
rlabel metal2 s 62366 -960 62478 480 8 wbs_adr_i[14]
port 538 nsew default input
rlabel metal2 s 65954 -960 66066 480 8 wbs_adr_i[15]
port 539 nsew default input
rlabel metal2 s 69450 -960 69562 480 8 wbs_adr_i[16]
port 540 nsew default input
rlabel metal2 s 73038 -960 73150 480 8 wbs_adr_i[17]
port 541 nsew default input
rlabel metal2 s 76626 -960 76738 480 8 wbs_adr_i[18]
port 542 nsew default input
rlabel metal2 s 80214 -960 80326 480 8 wbs_adr_i[19]
port 543 nsew default input
rlabel metal2 s 12410 -960 12522 480 8 wbs_adr_i[1]
port 544 nsew default input
rlabel metal2 s 83802 -960 83914 480 8 wbs_adr_i[20]
port 545 nsew default input
rlabel metal2 s 87298 -960 87410 480 8 wbs_adr_i[21]
port 546 nsew default input
rlabel metal2 s 90886 -960 90998 480 8 wbs_adr_i[22]
port 547 nsew default input
rlabel metal2 s 94474 -960 94586 480 8 wbs_adr_i[23]
port 548 nsew default input
rlabel metal2 s 98062 -960 98174 480 8 wbs_adr_i[24]
port 549 nsew default input
rlabel metal2 s 101558 -960 101670 480 8 wbs_adr_i[25]
port 550 nsew default input
rlabel metal2 s 105146 -960 105258 480 8 wbs_adr_i[26]
port 551 nsew default input
rlabel metal2 s 108734 -960 108846 480 8 wbs_adr_i[27]
port 552 nsew default input
rlabel metal2 s 112322 -960 112434 480 8 wbs_adr_i[28]
port 553 nsew default input
rlabel metal2 s 115910 -960 116022 480 8 wbs_adr_i[29]
port 554 nsew default input
rlabel metal2 s 17194 -960 17306 480 8 wbs_adr_i[2]
port 555 nsew default input
rlabel metal2 s 119406 -960 119518 480 8 wbs_adr_i[30]
port 556 nsew default input
rlabel metal2 s 122994 -960 123106 480 8 wbs_adr_i[31]
port 557 nsew default input
rlabel metal2 s 21886 -960 21998 480 8 wbs_adr_i[3]
port 558 nsew default input
rlabel metal2 s 26670 -960 26782 480 8 wbs_adr_i[4]
port 559 nsew default input
rlabel metal2 s 30258 -960 30370 480 8 wbs_adr_i[5]
port 560 nsew default input
rlabel metal2 s 33846 -960 33958 480 8 wbs_adr_i[6]
port 561 nsew default input
rlabel metal2 s 37342 -960 37454 480 8 wbs_adr_i[7]
port 562 nsew default input
rlabel metal2 s 40930 -960 41042 480 8 wbs_adr_i[8]
port 563 nsew default input
rlabel metal2 s 44518 -960 44630 480 8 wbs_adr_i[9]
port 564 nsew default input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 565 nsew default input
rlabel metal2 s 8822 -960 8934 480 8 wbs_dat_i[0]
port 566 nsew default input
rlabel metal2 s 49302 -960 49414 480 8 wbs_dat_i[10]
port 567 nsew default input
rlabel metal2 s 52798 -960 52910 480 8 wbs_dat_i[11]
port 568 nsew default input
rlabel metal2 s 56386 -960 56498 480 8 wbs_dat_i[12]
port 569 nsew default input
rlabel metal2 s 59974 -960 60086 480 8 wbs_dat_i[13]
port 570 nsew default input
rlabel metal2 s 63562 -960 63674 480 8 wbs_dat_i[14]
port 571 nsew default input
rlabel metal2 s 67150 -960 67262 480 8 wbs_dat_i[15]
port 572 nsew default input
rlabel metal2 s 70646 -960 70758 480 8 wbs_dat_i[16]
port 573 nsew default input
rlabel metal2 s 74234 -960 74346 480 8 wbs_dat_i[17]
port 574 nsew default input
rlabel metal2 s 77822 -960 77934 480 8 wbs_dat_i[18]
port 575 nsew default input
rlabel metal2 s 81410 -960 81522 480 8 wbs_dat_i[19]
port 576 nsew default input
rlabel metal2 s 13606 -960 13718 480 8 wbs_dat_i[1]
port 577 nsew default input
rlabel metal2 s 84906 -960 85018 480 8 wbs_dat_i[20]
port 578 nsew default input
rlabel metal2 s 88494 -960 88606 480 8 wbs_dat_i[21]
port 579 nsew default input
rlabel metal2 s 92082 -960 92194 480 8 wbs_dat_i[22]
port 580 nsew default input
rlabel metal2 s 95670 -960 95782 480 8 wbs_dat_i[23]
port 581 nsew default input
rlabel metal2 s 99258 -960 99370 480 8 wbs_dat_i[24]
port 582 nsew default input
rlabel metal2 s 102754 -960 102866 480 8 wbs_dat_i[25]
port 583 nsew default input
rlabel metal2 s 106342 -960 106454 480 8 wbs_dat_i[26]
port 584 nsew default input
rlabel metal2 s 109930 -960 110042 480 8 wbs_dat_i[27]
port 585 nsew default input
rlabel metal2 s 113518 -960 113630 480 8 wbs_dat_i[28]
port 586 nsew default input
rlabel metal2 s 117106 -960 117218 480 8 wbs_dat_i[29]
port 587 nsew default input
rlabel metal2 s 18298 -960 18410 480 8 wbs_dat_i[2]
port 588 nsew default input
rlabel metal2 s 120602 -960 120714 480 8 wbs_dat_i[30]
port 589 nsew default input
rlabel metal2 s 124190 -960 124302 480 8 wbs_dat_i[31]
port 590 nsew default input
rlabel metal2 s 23082 -960 23194 480 8 wbs_dat_i[3]
port 591 nsew default input
rlabel metal2 s 27866 -960 27978 480 8 wbs_dat_i[4]
port 592 nsew default input
rlabel metal2 s 31454 -960 31566 480 8 wbs_dat_i[5]
port 593 nsew default input
rlabel metal2 s 34950 -960 35062 480 8 wbs_dat_i[6]
port 594 nsew default input
rlabel metal2 s 38538 -960 38650 480 8 wbs_dat_i[7]
port 595 nsew default input
rlabel metal2 s 42126 -960 42238 480 8 wbs_dat_i[8]
port 596 nsew default input
rlabel metal2 s 45714 -960 45826 480 8 wbs_dat_i[9]
port 597 nsew default input
rlabel metal2 s 10018 -960 10130 480 8 wbs_dat_o[0]
port 598 nsew default tristate
rlabel metal2 s 50498 -960 50610 480 8 wbs_dat_o[10]
port 599 nsew default tristate
rlabel metal2 s 53994 -960 54106 480 8 wbs_dat_o[11]
port 600 nsew default tristate
rlabel metal2 s 57582 -960 57694 480 8 wbs_dat_o[12]
port 601 nsew default tristate
rlabel metal2 s 61170 -960 61282 480 8 wbs_dat_o[13]
port 602 nsew default tristate
rlabel metal2 s 64758 -960 64870 480 8 wbs_dat_o[14]
port 603 nsew default tristate
rlabel metal2 s 68254 -960 68366 480 8 wbs_dat_o[15]
port 604 nsew default tristate
rlabel metal2 s 71842 -960 71954 480 8 wbs_dat_o[16]
port 605 nsew default tristate
rlabel metal2 s 75430 -960 75542 480 8 wbs_dat_o[17]
port 606 nsew default tristate
rlabel metal2 s 79018 -960 79130 480 8 wbs_dat_o[18]
port 607 nsew default tristate
rlabel metal2 s 82606 -960 82718 480 8 wbs_dat_o[19]
port 608 nsew default tristate
rlabel metal2 s 14802 -960 14914 480 8 wbs_dat_o[1]
port 609 nsew default tristate
rlabel metal2 s 86102 -960 86214 480 8 wbs_dat_o[20]
port 610 nsew default tristate
rlabel metal2 s 89690 -960 89802 480 8 wbs_dat_o[21]
port 611 nsew default tristate
rlabel metal2 s 93278 -960 93390 480 8 wbs_dat_o[22]
port 612 nsew default tristate
rlabel metal2 s 96866 -960 96978 480 8 wbs_dat_o[23]
port 613 nsew default tristate
rlabel metal2 s 100454 -960 100566 480 8 wbs_dat_o[24]
port 614 nsew default tristate
rlabel metal2 s 103950 -960 104062 480 8 wbs_dat_o[25]
port 615 nsew default tristate
rlabel metal2 s 107538 -960 107650 480 8 wbs_dat_o[26]
port 616 nsew default tristate
rlabel metal2 s 111126 -960 111238 480 8 wbs_dat_o[27]
port 617 nsew default tristate
rlabel metal2 s 114714 -960 114826 480 8 wbs_dat_o[28]
port 618 nsew default tristate
rlabel metal2 s 118210 -960 118322 480 8 wbs_dat_o[29]
port 619 nsew default tristate
rlabel metal2 s 19494 -960 19606 480 8 wbs_dat_o[2]
port 620 nsew default tristate
rlabel metal2 s 121798 -960 121910 480 8 wbs_dat_o[30]
port 621 nsew default tristate
rlabel metal2 s 125386 -960 125498 480 8 wbs_dat_o[31]
port 622 nsew default tristate
rlabel metal2 s 24278 -960 24390 480 8 wbs_dat_o[3]
port 623 nsew default tristate
rlabel metal2 s 29062 -960 29174 480 8 wbs_dat_o[4]
port 624 nsew default tristate
rlabel metal2 s 32650 -960 32762 480 8 wbs_dat_o[5]
port 625 nsew default tristate
rlabel metal2 s 36146 -960 36258 480 8 wbs_dat_o[6]
port 626 nsew default tristate
rlabel metal2 s 39734 -960 39846 480 8 wbs_dat_o[7]
port 627 nsew default tristate
rlabel metal2 s 43322 -960 43434 480 8 wbs_dat_o[8]
port 628 nsew default tristate
rlabel metal2 s 46910 -960 47022 480 8 wbs_dat_o[9]
port 629 nsew default tristate
rlabel metal2 s 11214 -960 11326 480 8 wbs_sel_i[0]
port 630 nsew default input
rlabel metal2 s 15998 -960 16110 480 8 wbs_sel_i[1]
port 631 nsew default input
rlabel metal2 s 20690 -960 20802 480 8 wbs_sel_i[2]
port 632 nsew default input
rlabel metal2 s 25474 -960 25586 480 8 wbs_sel_i[3]
port 633 nsew default input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 634 nsew default input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 635 nsew default input
rlabel metal5 s -1996 -924 585920 -324 8 vccd1
port 636 nsew default input
rlabel metal5 s -2916 -1844 586840 -1244 8 vssd1
port 637 nsew default input
rlabel metal5 s -3836 -2764 587760 -2164 8 vccd2
port 638 nsew default input
rlabel metal5 s -4756 -3684 588680 -3084 8 vssd2
port 639 nsew default input
rlabel metal5 s -5676 -4604 589600 -4004 8 vdda1
port 640 nsew default input
rlabel metal5 s -6596 -5524 590520 -4924 8 vssa1
port 641 nsew default input
rlabel metal5 s -7516 -6444 591440 -5844 8 vdda2
port 642 nsew default input
rlabel metal5 s -8436 -7364 592360 -6764 8 vssa2
port 643 nsew default input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
