`default_nettype none
/*
 *-------------------------------------------------------------
 *
 * user_proj_ls130tw1  (LibreSilicon Testwafer #1)
 *
 */

module AND2X1(
	inout vdd,
	inout gnd,
	inout B,
	inout A,
	inout Y
);
endmodule

module AND2X2(
	inout vdd,
	inout gnd,
	inout B,
	inout A,
	inout Y
);
endmodule 

module OR2X1
(
	inout vdd,
	inout gnd,
	inout B,
	inout A,
	inout Y
);
endmodule

module OR2X2
(
	inout vdd,
	inout gnd,
	inout B,
	inout A,
	inout Y
);
endmodule

module NOR2X1
(
	inout vdd,
	inout gnd,
	inout B,
	inout A,
	inout Y
);
endmodule

module NOR2X2
(
	inout vdd,
	inout gnd,
	inout B,
	inout A,
	inout Y
);
endmodule

module INV(
	inout vdd,
	inout gnd,
	inout A,
	inout Y
);
endmodule

module INVX1(
	inout vdd,
	inout gnd,
	inout A,
	inout Y
);
endmodule
module INVX2(
	inout vdd,
	inout gnd,
	inout A,
	inout Y
);
endmodule
module INVX3(
	inout vdd,
	inout gnd,
	inout A,
	inout Y
);
endmodule
module INVX4(
	inout vdd,
	inout gnd,
	inout A,
	inout Y
);
endmodule

module BUFX1(
	inout vdd,
	inout gnd,
	inout A,
	inout Y
);
endmodule
module BUFX2(
	inout vdd,
	inout gnd,
	inout A,
	inout Y
);
endmodule

module AOI21X1
(
	inout vdd,
	inout gnd,
	inout C,
	inout B,
	inout A,
	inout Y
);
endmodule



