MACRO AOI22X1
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN AOI22X1 0 0 ;
 SITE CORE ;
 SYMMETRY X Y R90 ;
  PIN VDD
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.00000000 2.52500000 4.60000000 2.91500000 ;
    END
  END VDD

  PIN GND
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.00000000 -0.19500000 4.60000000 0.19500000 ;
    END
  END GND

  PIN Y
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        POLYGON 0.34500000 0.60000000 0.34500000 0.83000000 0.57500000 0.83000000 0.57500000 0.78500000 4.02500000 0.78500000 4.02500000 0.83000000 4.25500000 0.83000000 4.25500000 0.60000000 4.02500000 0.60000000 4.02500000 0.64500000 0.57500000 0.64500000 0.57500000 0.60000000 ;
       LAYER metal2 ;
        RECT 1.26500000 1.90000000 1.49500000 2.13000000 ;
    END
  END Y

  PIN C
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 1.72500000 0.99000000 1.95500000 1.35000000 ;
    END
  END C

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        POLYGON 3.56500000 0.99000000 3.56500000 1.22000000 3.61000000 1.22000000 3.61000000 1.51000000 3.56500000 1.51000000 3.56500000 1.74000000 3.79500000 1.74000000 3.79500000 1.51000000 3.75000000 1.51000000 3.75000000 1.22000000 3.79500000 1.22000000 3.79500000 0.99000000 ;
    END
  END B

  PIN D
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.80500000 0.99000000 1.03500000 1.35000000 ;
    END
  END D

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        POLYGON 2.64500000 0.99000000 2.64500000 1.22000000 2.69000000 1.22000000 2.69000000 1.51000000 2.64500000 1.51000000 2.64500000 1.74000000 2.87500000 1.74000000 2.87500000 1.51000000 2.83000000 1.51000000 2.83000000 1.22000000 2.87500000 1.22000000 2.87500000 0.99000000 ;
    END
  END A


END AOI22X1
