magic
tech sky130A
timestamp 1607784144
<< end >>
