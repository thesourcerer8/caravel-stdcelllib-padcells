MACRO NOR3X1
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN NOR3X1 0 0 ;
 SITE CORE ;
 SYMMETRY X Y R90 ;
  PIN VDD
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.00000000 2.48000000 6.44000000 2.96000000 ;
    END
  END VDD

  PIN GND
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.00000000 -0.24000000 6.44000000 0.24000000 ;
    END
  END GND

  PIN Y
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 1.23500000 0.57000000 1.52500000 0.77500000 ;
        RECT 3.07500000 0.57000000 3.36500000 0.77500000 ;
        RECT 0.39000000 0.77500000 6.05000000 0.91500000 ;
        RECT 0.39000000 0.91500000 0.53000000 1.74000000 ;
        RECT 5.91000000 0.91500000 6.05000000 1.74000000 ;
        RECT 0.31500000 1.74000000 0.60500000 2.03000000 ;
        RECT 5.83500000 1.74000000 6.12500000 2.03000000 ;
    END
  END Y

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 2.61500000 1.09000000 2.90500000 1.16500000 ;
        RECT 2.61500000 1.16500000 3.75000000 1.22000000 ;
        RECT 2.61500000 1.22000000 3.82500000 1.30500000 ;
        RECT 2.61500000 1.30500000 2.90500000 1.38000000 ;
        RECT 3.53500000 1.30500000 3.82500000 1.51000000 ;
    END
  END A

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 1.69500000 1.09000000 1.98500000 1.64000000 ;
       LAYER metal2 ;
        RECT 4.45500000 1.35000000 4.74500000 1.64000000 ;
    END
  END B

  PIN C
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.77500000 1.09000000 1.06500000 1.64000000 ;
       LAYER metal2 ;
        RECT 5.37500000 1.35000000 5.66500000 1.64000000 ;
    END
  END C


END NOR3X1
