magic
tech sky130A
timestamp 1607800073
<< end >>
