MACRO BUFX2
 CLASS CORE ;
 ORIGIN 0.0 0.0 ;
 FOREIGN BUFX2 0.0 0.0 ;
 SYMMETRY X Y R90 ;
 SITE unithd ;
  PIN vdd
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 0.00000000 3.96500000 3.12000000 4.35500000 ;
    END
  END vdd

  PIN gnd
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 0.00000000 -0.19500000 3.12000000 0.19500000 ;
    END
  END gnd

  PIN Y
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        POLYGON 2.48500000 0.73000000 2.48500000 0.96000000 2.53000000 0.96000000 2.53000000 3.20000000 2.48500000 3.20000000 2.48500000 3.43000000 2.71500000 3.43000000 2.71500000 3.20000000 2.67000000 3.20000000 2.67000000 0.96000000 2.71500000 0.96000000 2.71500000 0.73000000 ;
    END
  END Y

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 0.92500000 2.81000000 1.15500000 3.04000000 ;
    END
  END A


END BUFX2
