VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO CLKBUF1
  CLASS CORE ;
  FOREIGN CLKBUF1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.280 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 8.280 2.960 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 8.280 0.240 ;
    END
  END gnd
  PIN Y
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 6.760 2.050 7.050 2.310 ;
        RECT 6.760 2.020 7.890 2.050 ;
        RECT 6.830 1.910 7.890 2.020 ;
        RECT 7.750 0.790 7.890 1.910 ;
        RECT 6.830 0.690 7.890 0.790 ;
        RECT 6.760 0.650 7.890 0.690 ;
        RECT 6.760 0.400 7.050 0.650 ;
    END
  END Y
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.780 1.480 1.070 1.770 ;
        RECT 1.700 1.480 1.990 1.770 ;
        RECT 0.850 1.230 0.990 1.480 ;
        RECT 1.770 1.230 1.910 1.480 ;
        RECT 0.780 1.150 1.070 1.230 ;
        RECT 1.700 1.150 1.990 1.230 ;
        RECT 0.780 1.010 1.990 1.150 ;
        RECT 0.780 0.940 1.070 1.010 ;
        RECT 1.700 0.940 1.990 1.010 ;
    END
  END A
END CLKBUF1
END LIBRARY

