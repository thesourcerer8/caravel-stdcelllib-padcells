VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO INVX8
  CLASS CORE ;
  FOREIGN INVX8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.600 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
        RECT 0.000 2.480 4.600 2.960 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
        RECT 0.000 -0.240 4.600 0.240 ;
    END
  END gnd
  PIN Y
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
        RECT 0.320 1.960 0.610 2.030 ;
        RECT 2.160 1.960 2.450 2.030 ;
        RECT 4.000 1.960 4.290 2.030 ;
        RECT 0.320 1.820 4.290 1.960 ;
        RECT 0.320 1.740 0.610 1.820 ;
        RECT 2.160 1.740 2.450 1.820 ;
        RECT 4.000 1.740 4.290 1.820 ;
        RECT 0.390 0.860 0.530 1.740 ;
        RECT 4.070 0.860 4.210 1.740 ;
        RECT 0.320 0.790 0.610 0.860 ;
        RECT 2.160 0.790 2.450 0.860 ;
        RECT 0.320 0.650 2.450 0.790 ;
        RECT 0.320 0.570 0.610 0.650 ;
        RECT 2.160 0.570 2.450 0.650 ;
        RECT 4.000 0.570 4.290 0.860 ;
    END
  END Y
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
        RECT 0.780 1.310 1.070 1.640 ;
        RECT 1.700 1.310 1.990 1.640 ;
        RECT 2.620 1.310 2.910 1.640 ;
        RECT 3.540 1.310 3.830 1.640 ;
        RECT 0.780 1.170 3.830 1.310 ;
        RECT 0.780 1.090 1.070 1.170 ;
        RECT 1.700 1.090 1.990 1.170 ;
        RECT 2.620 1.090 2.910 1.170 ;
        RECT 3.540 1.090 3.830 1.170 ;
    END
  END A
END INVX8
END LIBRARY

