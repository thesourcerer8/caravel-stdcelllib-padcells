MACRO XNOR2X1
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN XNOR2X1 0 0 ;
 SITE CORE ;
 SYMMETRY X Y R90 ;
  PIN VDD
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.00000000 2.52500000 6.44000000 2.91500000 ;
    END
  END VDD

  PIN GND
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.00000000 -0.19500000 6.44000000 0.19500000 ;
    END
  END GND

  PIN Y
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 3.10500000 0.86000000 3.33500000 1.09000000 ;
    END
  END Y

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        POLYGON 0.80500000 0.99000000 0.80500000 1.22000000 1.03500000 1.22000000 1.03500000 1.17500000 1.72500000 1.17500000 1.72500000 1.35000000 1.95500000 1.35000000 1.95500000 0.99000000 1.72500000 0.99000000 1.72500000 1.03500000 1.03500000 1.03500000 1.03500000 0.99000000 ;
    END
  END B

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        POLYGON 5.40500000 0.99000000 5.40500000 1.22000000 5.45000000 1.22000000 5.45000000 1.51000000 5.40500000 1.51000000 5.40500000 1.74000000 5.63500000 1.74000000 5.63500000 1.51000000 5.59000000 1.51000000 5.59000000 1.22000000 5.63500000 1.22000000 5.63500000 0.99000000 ;
       LAYER metal2 ;
        RECT 3.56500000 0.99000000 3.79500000 1.22000000 ;
       LAYER metal2 ;
        RECT 2.64500000 1.90000000 2.87500000 2.13000000 ;
    END
  END A


END XNOR2X1
