MACRO CLKBUF1
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN CLKBUF1 0 0 ;
 SITE CORE ;
 SYMMETRY X Y R90 ;
  PIN VDD
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.00000000 2.48000000 8.28000000 2.96000000 ;
    END
  END VDD

  PIN GND
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.00000000 -0.24000000 8.28000000 0.24000000 ;
    END
  END GND

  PIN Y
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 6.75500000 0.57000000 7.04500000 0.77500000 ;
        RECT 6.75500000 0.77500000 7.89000000 0.86000000 ;
        RECT 6.83000000 0.86000000 7.89000000 0.91500000 ;
        RECT 6.75500000 1.74000000 7.04500000 1.81500000 ;
        RECT 7.75000000 0.91500000 7.89000000 1.81500000 ;
        RECT 6.75500000 1.81500000 7.89000000 1.95500000 ;
        RECT 6.75500000 1.95500000 7.04500000 2.03000000 ;
    END
  END Y

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.77500000 1.09000000 1.06500000 1.42500000 ;
        RECT 1.69500000 1.09000000 1.98500000 1.42500000 ;
        RECT 0.77500000 1.42500000 1.98500000 1.56500000 ;
        RECT 0.77500000 1.56500000 1.06500000 1.64000000 ;
        RECT 1.69500000 1.56500000 1.98500000 1.64000000 ;
    END
  END A


END CLKBUF1
