MACRO AOI22X1
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN AOI22X1 0 0 ;
 SITE CORE ;
 SYMMETRY X Y R90 ;
  PIN VDD
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.00000000 2.48000000 4.60000000 2.96000000 ;
    END
  END VDD

  PIN GND
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.00000000 -0.24000000 4.60000000 0.24000000 ;
    END
  END GND

  PIN Y
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.31500000 0.39500000 0.60500000 0.65000000 ;
        RECT 1.23500000 0.57500000 1.52500000 0.65000000 ;
        RECT 3.99500000 0.39500000 4.28500000 0.65000000 ;
        RECT 0.31500000 0.65000000 4.28500000 0.68500000 ;
        RECT 0.39000000 0.68500000 4.21000000 0.79000000 ;
        RECT 1.23500000 0.79000000 1.52500000 0.86500000 ;
    END
  END Y

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 3.53500000 0.93500000 3.82500000 1.22500000 ;
        RECT 3.61000000 1.22500000 3.75000000 1.47500000 ;
        RECT 3.53500000 1.47500000 3.82500000 1.76500000 ;
    END
  END B

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 2.61500000 0.93500000 2.90500000 1.22500000 ;
        RECT 2.69000000 1.22500000 2.83000000 1.47500000 ;
        RECT 2.61500000 1.47500000 2.90500000 1.76500000 ;
    END
  END A

  PIN D
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.77500000 0.93500000 1.06500000 1.22500000 ;
        RECT 0.85000000 1.22500000 0.99000000 1.47500000 ;
        RECT 0.77500000 1.47500000 1.06500000 1.76500000 ;
    END
  END D

  PIN C
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 1.69500000 0.93500000 1.98500000 1.22500000 ;
        RECT 1.77000000 1.22500000 1.91000000 1.47500000 ;
        RECT 1.69500000 1.47500000 1.98500000 1.76500000 ;
    END
  END C


END AOI22X1
