MACRO OAI22X1
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN OAI22X1 0 0 ;
 SITE CORE ;
 SYMMETRY X Y R90 ;
  PIN VDD
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.00000000 2.48000000 4.60000000 2.96000000 ;
    END
  END VDD

  PIN GND
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.00000000 -0.24000000 4.60000000 0.24000000 ;
    END
  END GND

  PIN Y
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 1.23500000 1.11500000 1.52500000 1.40500000 ;
        RECT 1.31000000 1.40500000 1.45000000 1.91000000 ;
        RECT 1.31000000 1.91000000 4.21000000 2.01500000 ;
        RECT 1.31000000 2.01500000 4.28500000 2.05000000 ;
        RECT 0.31500000 2.01500000 0.60500000 2.09000000 ;
        RECT 1.31000000 2.05000000 1.45000000 2.09000000 ;
        RECT 0.31500000 2.09000000 1.45000000 2.23000000 ;
        RECT 0.31500000 2.23000000 0.60500000 2.30500000 ;
        RECT 3.99500000 2.05000000 4.28500000 2.30500000 ;
    END
  END Y

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 3.53500000 0.93500000 3.82500000 1.22500000 ;
        RECT 3.61000000 1.22500000 3.75000000 1.47500000 ;
        RECT 3.53500000 1.47500000 3.82500000 1.76500000 ;
    END
  END B

  PIN C
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 1.69500000 1.11500000 1.98500000 1.76500000 ;
    END
  END C

  PIN D
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.77500000 1.47500000 1.06500000 1.76500000 ;
    END
  END D

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 2.61500000 0.93500000 2.90500000 1.22500000 ;
        RECT 2.69000000 1.22500000 2.83000000 1.47500000 ;
        RECT 2.61500000 1.47500000 2.90500000 1.76500000 ;
    END
  END A


END OAI22X1
