MACRO TBUFX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN TBUFX2 0 0 ;
 SITE CORE ;
 SYMMETRY X Y R90 ;
  PIN VDD
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.00000000 2.48000000 5.52000000 2.96000000 ;
    END
  END VDD

  PIN GND
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.00000000 -0.24000000 5.52000000 0.24000000 ;
    END
  END GND

  PIN Y
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 3.07500000 0.39500000 3.36500000 0.68500000 ;
    END
  END Y

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 4.45500000 0.93500000 4.74500000 1.22500000 ;
        RECT 4.53000000 1.22500000 4.67000000 1.47500000 ;
        RECT 4.45500000 1.47500000 4.74500000 1.76500000 ;
       LAYER metal2 ;
        RECT 1.69500000 0.93500000 1.98500000 1.22500000 ;
    END
  END A

  PIN EN
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.77500000 0.93500000 1.06500000 1.22500000 ;
       LAYER metal2 ;
        RECT 2.61500000 0.93500000 2.90500000 1.22500000 ;
       LAYER metal2 ;
        RECT 3.53500000 0.93500000 3.82500000 1.22500000 ;
    END
  END EN


END TBUFX2
