MACRO AND2X1
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN AND2X1 0 0 ;
 SITE CORE ;
 SYMMETRY X Y R90 ;
  PIN VDD
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.00000000 2.52500000 3.68000000 2.91500000 ;
    END
  END VDD

  PIN GND
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.00000000 -0.19500000 3.68000000 0.19500000 ;
    END
  END GND

  PIN Y
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        POLYGON 3.10500000 0.60000000 3.10500000 0.83000000 3.15000000 0.83000000 3.15000000 1.90000000 3.10500000 1.90000000 3.10500000 2.13000000 3.33500000 2.13000000 3.33500000 1.90000000 3.29000000 1.90000000 3.29000000 0.83000000 3.33500000 0.83000000 3.33500000 0.60000000 ;
    END
  END Y

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        POLYGON 0.80500000 0.99000000 0.80500000 1.22000000 0.85000000 1.22000000 0.85000000 1.51000000 0.80500000 1.51000000 0.80500000 1.74000000 1.03500000 1.74000000 1.03500000 1.51000000 0.99000000 1.51000000 0.99000000 1.22000000 1.03500000 1.22000000 1.03500000 0.99000000 ;
    END
  END A

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        POLYGON 1.72500000 0.99000000 1.72500000 1.22000000 1.77000000 1.22000000 1.77000000 1.51000000 1.72500000 1.51000000 1.72500000 1.74000000 1.95500000 1.74000000 1.95500000 1.51000000 1.91000000 1.51000000 1.91000000 1.22000000 1.95500000 1.22000000 1.95500000 0.99000000 ;
    END
  END B


END AND2X1
