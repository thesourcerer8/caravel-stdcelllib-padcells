MACRO HAX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN HAX1 0 0 ;
 SITE CORE ;
 SYMMETRY X Y R90 ;
  PIN VDD
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.00000000 2.48000000 10.12000000 2.96000000 ;
    END
  END VDD

  PIN GND
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.00000000 -0.24000000 10.12000000 0.24000000 ;
    END
  END GND

  PIN YC
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 1.23500000 0.39500000 1.52500000 0.65000000 ;
        RECT 0.39000000 0.65000000 1.52500000 0.68500000 ;
        RECT 0.39000000 0.68500000 1.45000000 0.79000000 ;
        RECT 0.39000000 0.79000000 0.53000000 1.91000000 ;
        RECT 0.39000000 1.91000000 1.45000000 2.01500000 ;
        RECT 0.39000000 2.01500000 1.52500000 2.05000000 ;
        RECT 1.23500000 2.05000000 1.52500000 2.30500000 ;
    END
  END YC

  PIN YS
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 8.59500000 0.39500000 8.88500000 0.68500000 ;
    END
  END YS

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 7.21500000 0.93500000 7.50500000 1.22500000 ;
        RECT 7.29000000 1.22500000 7.43000000 1.47500000 ;
        RECT 7.21500000 1.47500000 7.50500000 1.76500000 ;
       LAYER metal2 ;
        RECT 3.53500000 0.93500000 3.82500000 1.22500000 ;
       LAYER metal2 ;
        RECT 3.53500000 1.47500000 3.82500000 1.76500000 ;
    END
  END A

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 2.69000000 0.65000000 5.82000000 0.79000000 ;
        RECT 5.68000000 0.79000000 5.82000000 0.83000000 ;
        RECT 2.69000000 0.79000000 2.83000000 0.93500000 ;
        RECT 5.68000000 0.83000000 6.51000000 0.93500000 ;
        RECT 5.68000000 0.93500000 6.58500000 0.97000000 ;
        RECT 2.61500000 0.93500000 2.90500000 1.22500000 ;
        RECT 6.29500000 0.97000000 6.58500000 1.22500000 ;
        RECT 2.69000000 1.22500000 2.83000000 1.47500000 ;
        RECT 6.37000000 1.22500000 6.51000000 1.47500000 ;
        RECT 2.61500000 1.47500000 2.90500000 1.76500000 ;
        RECT 6.29500000 1.47500000 6.58500000 1.76500000 ;
    END
  END B


END HAX1
