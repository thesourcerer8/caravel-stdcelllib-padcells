MACRO NOR2X1
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN NOR2X1 0 0 ;
 SITE CORE ;
 SYMMETRY X Y R90 ;
  PIN VDD
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.00000000 2.52500000 2.76000000 2.91500000 ;
    END
  END VDD

  PIN GND
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.00000000 -0.19500000 2.76000000 0.19500000 ;
    END
  END GND

  PIN Y
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        POLYGON 0.34500000 0.60000000 0.34500000 0.83000000 0.57500000 0.83000000 0.57500000 0.78500000 2.18500000 0.78500000 2.18500000 0.83000000 2.23000000 0.83000000 2.23000000 1.90000000 2.18500000 1.90000000 2.18500000 2.13000000 2.41500000 2.13000000 2.41500000 1.90000000 2.37000000 1.90000000 2.37000000 0.83000000 2.41500000 0.83000000 2.41500000 0.60000000 2.18500000 0.60000000 2.18500000 0.64500000 0.57500000 0.64500000 0.57500000 0.60000000 ;
    END
  END Y

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        POLYGON 0.80500000 0.99000000 0.80500000 1.22000000 0.85000000 1.22000000 0.85000000 1.51000000 0.80500000 1.51000000 0.80500000 1.74000000 1.03500000 1.74000000 1.03500000 1.51000000 0.99000000 1.51000000 0.99000000 1.22000000 1.03500000 1.22000000 1.03500000 0.99000000 ;
    END
  END A

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        POLYGON 1.72500000 0.99000000 1.72500000 1.22000000 1.77000000 1.22000000 1.77000000 1.51000000 1.72500000 1.51000000 1.72500000 1.74000000 1.95500000 1.74000000 1.95500000 1.51000000 1.91000000 1.51000000 1.91000000 1.22000000 1.95500000 1.22000000 1.95500000 0.99000000 ;
    END
  END B


END NOR2X1
