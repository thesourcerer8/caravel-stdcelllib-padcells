VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO INVX2
  CLASS CORE ;
  FOREIGN INVX2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1.840 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN vdd
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
        RECT 0.000 2.530 1.840 2.920 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
        RECT 0.000 -0.200 1.840 0.200 ;
    END
  END gnd
  PIN Y
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
        RECT 0.350 1.900 0.580 2.130 ;
        RECT 0.390 0.830 0.530 1.900 ;
        RECT 0.350 0.600 0.580 0.830 ;
    END
  END Y
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
        RECT 0.810 1.510 1.040 1.740 ;
        RECT 0.850 1.220 0.990 1.510 ;
        RECT 0.810 0.990 1.040 1.220 ;
    END
  END A
END INVX2
END LIBRARY

