VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO XNOR2X1
  CLASS CORE ;
  FOREIGN XNOR2X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.440 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 6.440 2.960 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 6.440 0.240 ;
    END
  END gnd
  PIN Y
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 3.080 2.230 3.370 2.310 ;
        RECT 3.080 2.090 4.210 2.230 ;
        RECT 3.080 2.020 3.370 2.090 ;
        RECT 3.080 0.610 3.370 0.690 ;
        RECT 4.070 0.610 4.210 2.090 ;
        RECT 3.080 0.470 4.210 0.610 ;
        RECT 3.080 0.400 3.370 0.470 ;
    END
  END Y
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 3.540 0.970 3.830 1.230 ;
        RECT 2.920 0.940 3.830 0.970 ;
        RECT 0.780 0.790 1.070 0.870 ;
        RECT 2.920 0.830 3.750 0.940 ;
        RECT 2.920 0.790 3.060 0.830 ;
        RECT 0.780 0.650 3.060 0.790 ;
        RECT 0.780 0.580 1.070 0.650 ;
    END
  END A
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 1.700 1.480 1.990 1.770 ;
    END
    PORT
      LAYER met1 ;
        RECT 5.380 1.480 5.670 1.770 ;
        RECT 5.450 1.230 5.590 1.480 ;
        RECT 5.380 0.940 5.670 1.230 ;
    END
  END B
END XNOR2X1
END LIBRARY

