MACRO AOI22X1
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN AOI22X1 0 0 ;
 SITE CORE ;
 SYMMETRY X Y R90 ;
  PIN VDD
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.00000000 2.48000000 4.60000000 2.96000000 ;
    END
  END VDD

  PIN GND
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.00000000 -0.24000000 4.60000000 0.24000000 ;
    END
  END GND

  PIN Y
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.31500000 0.57000000 0.60500000 0.77500000 ;
        RECT 1.23500000 0.70000000 1.52500000 0.77500000 ;
        RECT 3.99500000 0.57000000 4.28500000 0.77500000 ;
        RECT 0.31500000 0.77500000 4.28500000 0.86000000 ;
        RECT 0.39000000 0.86000000 4.21000000 0.91500000 ;
        RECT 1.23500000 0.91500000 1.52500000 0.99000000 ;
    END
  END Y

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 3.53500000 1.09000000 3.82500000 1.64000000 ;
    END
  END B

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 2.61500000 1.09000000 2.90500000 1.64000000 ;
    END
  END A

  PIN D
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.77500000 1.09000000 1.06500000 1.64000000 ;
    END
  END D

  PIN C
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 1.69500000 1.09000000 1.98500000 1.64000000 ;
    END
  END C


END AOI22X1
