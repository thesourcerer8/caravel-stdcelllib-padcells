VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO TBUFX2
  CLASS CORE ;
  FOREIGN TBUFX2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 5.520 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
        RECT 0.000 2.530 5.520 2.920 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
        RECT 0.000 -0.200 5.520 0.200 ;
    END
  END gnd
  PIN Y
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
        RECT 3.110 1.900 3.340 2.130 ;
    END
    PORT
      LAYER met2 ;
        RECT 3.110 0.600 3.340 0.830 ;
    END
  END Y
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
        RECT 1.730 1.700 1.960 1.740 ;
        RECT 4.490 1.700 4.720 1.740 ;
        RECT 1.730 1.560 4.720 1.700 ;
        RECT 1.730 1.510 1.960 1.560 ;
        RECT 4.490 1.510 4.720 1.560 ;
        RECT 4.530 1.220 4.670 1.510 ;
        RECT 4.490 0.990 4.720 1.220 ;
    END
  END A
  PIN EN
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
        RECT 0.810 1.510 1.040 1.740 ;
        RECT 0.850 1.220 0.990 1.510 ;
        RECT 0.810 1.180 1.040 1.220 ;
        RECT 2.650 1.180 2.880 1.220 ;
        RECT 3.570 1.180 3.800 1.220 ;
        RECT 0.810 1.040 3.800 1.180 ;
        RECT 0.810 0.990 1.040 1.040 ;
        RECT 2.650 0.990 2.880 1.040 ;
        RECT 3.570 0.990 3.800 1.040 ;
    END
  END EN
END TBUFX2
END LIBRARY

