magic
tech sky130A
magscale 1 2
timestamp 1608117647
<< locali >>
rect 23839 57919 23873 59109
rect 17123 54655 17157 54757
rect 22183 42007 22217 42313
rect 51715 37655 51749 37825
rect 19147 31807 19181 31909
rect 51531 29019 51565 29189
rect 12155 23579 12189 23749
rect 9119 22559 9153 22729
rect 8567 21471 8601 21641
rect 8785 18173 9061 18207
rect 9027 18071 9061 18173
rect 26323 5627 26357 5797
<< viali >>
rect 23839 59109 23873 59143
rect 23839 57885 23873 57919
rect 32487 56729 32521 56763
rect 52451 56729 52485 56763
rect 25127 56661 25161 56695
rect 48679 56253 48713 56287
rect 5071 55573 5105 55607
rect 25495 54825 25529 54859
rect 17123 54757 17157 54791
rect 47851 54689 47885 54723
rect 17123 54621 17157 54655
rect 17399 54485 17433 54519
rect 21631 54485 21665 54519
rect 42423 54485 42457 54519
rect 5715 54077 5749 54111
rect 58339 53601 58373 53635
rect 17031 53193 17065 53227
rect 38283 52989 38317 53023
rect 47575 52989 47609 53023
rect 19239 52309 19273 52343
rect 58431 51901 58465 51935
rect 8751 51221 8785 51255
rect 47667 50677 47701 50711
rect 16479 50133 16513 50167
rect 18319 49045 18353 49079
rect 33499 49045 33533 49079
rect 44631 48637 44665 48671
rect 49231 48637 49265 48671
rect 16847 47957 16881 47991
rect 9947 47617 9981 47651
rect 45735 47549 45769 47583
rect 14639 47413 14673 47447
rect 57695 47413 57729 47447
rect 26783 46937 26817 46971
rect 5347 46461 5381 46495
rect 52083 46461 52117 46495
rect 40767 45373 40801 45407
rect 16847 45033 16881 45067
rect 2311 44693 2345 44727
rect 24483 44693 24517 44727
rect 47667 44693 47701 44727
rect 55855 44693 55889 44727
rect 56959 44693 56993 44727
rect 40123 43401 40157 43435
rect 5715 43197 5749 43231
rect 40675 43197 40709 43231
rect 32763 42653 32797 42687
rect 22183 42313 22217 42347
rect 22459 42313 22493 42347
rect 40215 42313 40249 42347
rect 18227 42177 18261 42211
rect 8751 42109 8785 42143
rect 29635 42177 29669 42211
rect 37639 42109 37673 42143
rect 22183 41973 22217 42007
rect 13535 41633 13569 41667
rect 42239 41429 42273 41463
rect 46287 41021 46321 41055
rect 57879 41021 57913 41055
rect 11879 40341 11913 40375
rect 43711 40341 43745 40375
rect 47023 40137 47057 40171
rect 48771 40069 48805 40103
rect 26967 40001 27001 40035
rect 10959 39253 10993 39287
rect 1851 39049 1885 39083
rect 21447 38913 21481 38947
rect 12615 38845 12649 38879
rect 1667 38165 1701 38199
rect 47851 38165 47885 38199
rect 51715 37825 51749 37859
rect 52083 37825 52117 37859
rect 49783 37757 49817 37791
rect 50519 37757 50553 37791
rect 51715 37621 51749 37655
rect 43619 37281 43653 37315
rect 12983 37077 13017 37111
rect 26691 37077 26725 37111
rect 29267 37077 29301 37111
rect 31107 37077 31141 37111
rect 47391 37077 47425 37111
rect 31659 36669 31693 36703
rect 45275 36669 45309 36703
rect 45643 35989 45677 36023
rect 25771 35581 25805 35615
rect 30647 35105 30681 35139
rect 52911 34901 52945 34935
rect 20803 34629 20837 34663
rect 50795 34561 50829 34595
rect 36535 33813 36569 33847
rect 43619 33813 43653 33847
rect 58431 33813 58465 33847
rect 6543 33473 6577 33507
rect 46287 33405 46321 33439
rect 12431 32725 12465 32759
rect 53095 32385 53129 32419
rect 10407 32317 10441 32351
rect 50887 32317 50921 32351
rect 19147 31909 19181 31943
rect 5071 31841 5105 31875
rect 37179 31841 37213 31875
rect 19147 31773 19181 31807
rect 19423 31773 19457 31807
rect 21907 31773 21941 31807
rect 32395 31773 32429 31807
rect 51623 31773 51657 31807
rect 21171 31229 21205 31263
rect 19331 30753 19365 30787
rect 7371 30549 7405 30583
rect 19699 30549 19733 30583
rect 13259 30209 13293 30243
rect 32579 30209 32613 30243
rect 48219 30141 48253 30175
rect 56959 30141 56993 30175
rect 16019 30005 16053 30039
rect 26691 29461 26725 29495
rect 45735 29461 45769 29495
rect 51439 29189 51473 29223
rect 51531 29189 51565 29223
rect 57879 29121 57913 29155
rect 51531 28985 51565 29019
rect 3783 28577 3817 28611
rect 26691 28373 26725 28407
rect 15467 27285 15501 27319
rect 53371 26945 53405 26979
rect 51899 26877 51933 26911
rect 4243 26401 4277 26435
rect 38559 26401 38593 26435
rect 40215 26401 40249 26435
rect 57143 26333 57177 26367
rect 50335 26265 50369 26299
rect 11419 25993 11453 26027
rect 7923 25789 7957 25823
rect 42791 25789 42825 25823
rect 1391 24769 1425 24803
rect 9855 24225 9889 24259
rect 19699 24021 19733 24055
rect 49231 24021 49265 24055
rect 43527 23817 43561 23851
rect 12155 23749 12189 23783
rect 57511 23749 57545 23783
rect 49599 23613 49633 23647
rect 12155 23545 12189 23579
rect 6911 22933 6945 22967
rect 21263 22933 21297 22967
rect 9119 22729 9153 22763
rect 9119 22525 9153 22559
rect 41503 22525 41537 22559
rect 34419 22049 34453 22083
rect 22551 21845 22585 21879
rect 8567 21641 8601 21675
rect 8567 21437 8601 21471
rect 24391 20961 24425 20995
rect 52083 20893 52117 20927
rect 31567 20825 31601 20859
rect 4059 20553 4093 20587
rect 18503 20417 18537 20451
rect 28623 20349 28657 20383
rect 45827 20349 45861 20383
rect 39571 20009 39605 20043
rect 49599 19873 49633 19907
rect 58155 19669 58189 19703
rect 9855 19329 9889 19363
rect 29451 19329 29485 19363
rect 13167 19261 13201 19295
rect 17307 18581 17341 18615
rect 32211 18241 32245 18275
rect 8751 18173 8785 18207
rect 52819 18173 52853 18207
rect 9027 18037 9061 18071
rect 53463 17493 53497 17527
rect 3967 17085 4001 17119
rect 16663 15997 16697 16031
rect 4243 15317 4277 15351
rect 8935 14909 8969 14943
rect 27151 14909 27185 14943
rect 56683 14909 56717 14943
rect 32211 14025 32245 14059
rect 46287 13889 46321 13923
rect 12615 13821 12649 13855
rect 6543 13345 6577 13379
rect 9855 12869 9889 12903
rect 15191 12733 15225 12767
rect 40675 12733 40709 12767
rect 46103 12597 46137 12631
rect 37915 12053 37949 12087
rect 47207 12053 47241 12087
rect 31199 11101 31233 11135
rect 42147 10557 42181 10591
rect 27519 9945 27553 9979
rect 31015 9877 31049 9911
rect 32119 9469 32153 9503
rect 43527 9469 43561 9503
rect 47483 9469 47517 9503
rect 52451 9469 52485 9503
rect 56683 9333 56717 9367
rect 19515 9129 19549 9163
rect 53647 8789 53681 8823
rect 39755 8585 39789 8619
rect 57511 8517 57545 8551
rect 11235 7701 11269 7735
rect 41595 7701 41629 7735
rect 58431 7701 58465 7735
rect 17583 7497 17617 7531
rect 49691 7497 49725 7531
rect 9855 7293 9889 7327
rect 22091 7293 22125 7327
rect 44999 7293 45033 7327
rect 51807 6749 51841 6783
rect 8383 6681 8417 6715
rect 52451 6613 52485 6647
rect 43159 6273 43193 6307
rect 34511 6205 34545 6239
rect 35799 6205 35833 6239
rect 42791 6205 42825 6239
rect 21907 5797 21941 5831
rect 26323 5797 26357 5831
rect 10315 5661 10349 5695
rect 28163 5729 28197 5763
rect 5715 5593 5749 5627
rect 26323 5593 26357 5627
rect 35707 5525 35741 5559
rect 46195 5185 46229 5219
rect 33775 5117 33809 5151
rect 55119 5117 55153 5151
rect 23839 4233 23873 4267
rect 2127 3553 2161 3587
rect 42331 3553 42365 3587
rect 12523 3349 12557 3383
rect 55303 3349 55337 3383
rect 14915 2261 14949 2295
<< metal1 >>
rect 15084 59100 15090 59152
rect 15142 59140 15148 59152
rect 15360 59140 15366 59152
rect 15142 59112 15366 59140
rect 15142 59100 15148 59112
rect 15360 59100 15366 59112
rect 15418 59100 15424 59152
rect 23824 59140 23830 59152
rect 23785 59112 23830 59140
rect 23824 59100 23830 59112
rect 23882 59100 23888 59152
rect 23824 57916 23830 57928
rect 23785 57888 23830 57916
rect 23824 57876 23830 57888
rect 23882 57876 23888 57928
rect 1086 57690 58862 57712
rect 1086 57638 4228 57690
rect 4280 57638 4292 57690
rect 4344 57638 4356 57690
rect 4408 57638 4420 57690
rect 4472 57638 34948 57690
rect 35000 57638 35012 57690
rect 35064 57638 35076 57690
rect 35128 57638 35140 57690
rect 35192 57638 58862 57690
rect 1086 57616 58862 57638
rect 1086 57146 58862 57168
rect 1086 57094 19588 57146
rect 19640 57094 19652 57146
rect 19704 57094 19716 57146
rect 19768 57094 19780 57146
rect 19832 57094 50308 57146
rect 50360 57094 50372 57146
rect 50424 57094 50436 57146
rect 50488 57094 50500 57146
rect 50552 57094 58862 57146
rect 1086 57072 58862 57094
rect 4964 56720 4970 56772
rect 5022 56760 5028 56772
rect 32475 56763 32533 56769
rect 32475 56760 32487 56763
rect 5022 56732 32487 56760
rect 5022 56720 5028 56732
rect 32475 56729 32487 56732
rect 32521 56729 32533 56763
rect 32475 56723 32533 56729
rect 32656 56720 32662 56772
rect 32714 56760 32720 56772
rect 52439 56763 52497 56769
rect 52439 56760 52451 56763
rect 32714 56732 52451 56760
rect 32714 56720 32720 56732
rect 52439 56729 52451 56732
rect 52485 56729 52497 56763
rect 52439 56723 52497 56729
rect 15084 56652 15090 56704
rect 15142 56692 15148 56704
rect 15268 56692 15274 56704
rect 15142 56664 15274 56692
rect 15142 56652 15148 56664
rect 15268 56652 15274 56664
rect 15326 56652 15332 56704
rect 17844 56652 17850 56704
rect 17902 56692 17908 56704
rect 25115 56695 25173 56701
rect 25115 56692 25127 56695
rect 17902 56664 25127 56692
rect 17902 56652 17908 56664
rect 25115 56661 25127 56664
rect 25161 56661 25173 56695
rect 25115 56655 25173 56661
rect 29988 56652 29994 56704
rect 30046 56692 30052 56704
rect 32196 56692 32202 56704
rect 30046 56664 32202 56692
rect 30046 56652 30052 56664
rect 32196 56652 32202 56664
rect 32254 56652 32260 56704
rect 1086 56602 58862 56624
rect 1086 56550 4228 56602
rect 4280 56550 4292 56602
rect 4344 56550 4356 56602
rect 4408 56550 4420 56602
rect 4472 56550 34948 56602
rect 35000 56550 35012 56602
rect 35064 56550 35076 56602
rect 35128 56550 35140 56602
rect 35192 56550 58862 56602
rect 1086 56528 58862 56550
rect 640 56448 646 56500
rect 698 56488 704 56500
rect 1100 56488 1106 56500
rect 698 56460 1106 56488
rect 698 56448 704 56460
rect 1100 56448 1106 56460
rect 1158 56448 1164 56500
rect 1744 56448 1750 56500
rect 1802 56488 1808 56500
rect 2664 56488 2670 56500
rect 1802 56460 2670 56488
rect 1802 56448 1808 56460
rect 2664 56448 2670 56460
rect 2722 56448 2728 56500
rect 10300 56448 10306 56500
rect 10358 56488 10364 56500
rect 12784 56488 12790 56500
rect 10358 56460 12790 56488
rect 10358 56448 10364 56460
rect 12784 56448 12790 56460
rect 12842 56448 12848 56500
rect 21708 56488 21714 56500
rect 16758 56460 21714 56488
rect 180 56380 186 56432
rect 238 56420 244 56432
rect 1284 56420 1290 56432
rect 238 56392 1290 56420
rect 238 56380 244 56392
rect 1284 56380 1290 56392
rect 1342 56380 1348 56432
rect 1376 56380 1382 56432
rect 1434 56420 1440 56432
rect 2204 56420 2210 56432
rect 1434 56392 2210 56420
rect 1434 56380 1440 56392
rect 2204 56380 2210 56392
rect 2262 56380 2268 56432
rect 2572 56380 2578 56432
rect 2630 56420 2636 56432
rect 16758 56420 16786 56460
rect 21708 56448 21714 56460
rect 21766 56448 21772 56500
rect 24284 56448 24290 56500
rect 24342 56488 24348 56500
rect 29988 56488 29994 56500
rect 24342 56460 29994 56488
rect 24342 56448 24348 56460
rect 29988 56448 29994 56460
rect 30046 56448 30052 56500
rect 33852 56488 33858 56500
rect 31478 56460 33858 56488
rect 17292 56420 17298 56432
rect 2630 56392 16786 56420
rect 16850 56392 17298 56420
rect 2630 56380 2636 56392
rect 1560 56312 1566 56364
rect 1618 56352 1624 56364
rect 16850 56352 16878 56392
rect 17292 56380 17298 56392
rect 17350 56380 17356 56432
rect 21156 56380 21162 56432
rect 21214 56420 21220 56432
rect 21984 56420 21990 56432
rect 21214 56392 21990 56420
rect 21214 56380 21220 56392
rect 21984 56380 21990 56392
rect 22042 56380 22048 56432
rect 22812 56380 22818 56432
rect 22870 56420 22876 56432
rect 28056 56420 28062 56432
rect 22870 56392 28062 56420
rect 22870 56380 22876 56392
rect 28056 56380 28062 56392
rect 28114 56380 28120 56432
rect 28148 56380 28154 56432
rect 28206 56420 28212 56432
rect 30632 56420 30638 56432
rect 28206 56392 30638 56420
rect 28206 56380 28212 56392
rect 30632 56380 30638 56392
rect 30690 56380 30696 56432
rect 31000 56380 31006 56432
rect 31058 56420 31064 56432
rect 31478 56420 31506 56460
rect 33852 56448 33858 56460
rect 33910 56448 33916 56500
rect 33962 56460 40154 56488
rect 32748 56420 32754 56432
rect 31058 56392 31506 56420
rect 31570 56392 32754 56420
rect 31058 56380 31064 56392
rect 1618 56324 16878 56352
rect 1618 56312 1624 56324
rect 16924 56312 16930 56364
rect 16982 56352 16988 56364
rect 24836 56352 24842 56364
rect 16982 56324 24842 56352
rect 16982 56312 16988 56324
rect 24836 56312 24842 56324
rect 24894 56312 24900 56364
rect 24928 56312 24934 56364
rect 24986 56352 24992 56364
rect 29068 56352 29074 56364
rect 24986 56324 29074 56352
rect 24986 56312 24992 56324
rect 29068 56312 29074 56324
rect 29126 56312 29132 56364
rect 29712 56312 29718 56364
rect 29770 56352 29776 56364
rect 31570 56352 31598 56392
rect 32748 56380 32754 56392
rect 32806 56380 32812 56432
rect 33760 56380 33766 56432
rect 33818 56420 33824 56432
rect 33962 56420 33990 56460
rect 33818 56392 33990 56420
rect 33818 56380 33824 56392
rect 35232 56380 35238 56432
rect 35290 56420 35296 56432
rect 40016 56420 40022 56432
rect 35290 56392 40022 56420
rect 35290 56380 35296 56392
rect 40016 56380 40022 56392
rect 40074 56380 40080 56432
rect 40126 56420 40154 56460
rect 40200 56448 40206 56500
rect 40258 56488 40264 56500
rect 41672 56488 41678 56500
rect 40258 56460 41678 56488
rect 40258 56448 40264 56460
rect 41672 56448 41678 56460
rect 41730 56448 41736 56500
rect 44708 56448 44714 56500
rect 44766 56488 44772 56500
rect 48020 56488 48026 56500
rect 44766 56460 48026 56488
rect 44766 56448 44772 56460
rect 48020 56448 48026 56460
rect 48078 56448 48084 56500
rect 48296 56448 48302 56500
rect 48354 56488 48360 56500
rect 49584 56488 49590 56500
rect 48354 56460 49590 56488
rect 48354 56448 48360 56460
rect 49584 56448 49590 56460
rect 49642 56448 49648 56500
rect 40752 56420 40758 56432
rect 40126 56392 40758 56420
rect 40752 56380 40758 56392
rect 40810 56380 40816 56432
rect 40844 56380 40850 56432
rect 40902 56420 40908 56432
rect 45536 56420 45542 56432
rect 40902 56392 45542 56420
rect 40902 56380 40908 56392
rect 45536 56380 45542 56392
rect 45594 56380 45600 56432
rect 46180 56380 46186 56432
rect 46238 56420 46244 56432
rect 51700 56420 51706 56432
rect 46238 56392 51706 56420
rect 46238 56380 46244 56392
rect 51700 56380 51706 56392
rect 51758 56380 51764 56432
rect 29770 56324 31598 56352
rect 29770 56312 29776 56324
rect 31644 56312 31650 56364
rect 31702 56352 31708 56364
rect 38636 56352 38642 56364
rect 31702 56324 38642 56352
rect 31702 56312 31708 56324
rect 38636 56312 38642 56324
rect 38694 56312 38700 56364
rect 49584 56312 49590 56364
rect 49642 56352 49648 56364
rect 53264 56352 53270 56364
rect 49642 56324 53270 56352
rect 49642 56312 49648 56324
rect 53264 56312 53270 56324
rect 53322 56312 53328 56364
rect 3676 56244 3682 56296
rect 3734 56284 3740 56296
rect 35876 56284 35882 56296
rect 3734 56256 35882 56284
rect 3734 56244 3740 56256
rect 35876 56244 35882 56256
rect 35934 56244 35940 56296
rect 35968 56244 35974 56296
rect 36026 56284 36032 56296
rect 40844 56284 40850 56296
rect 36026 56256 40850 56284
rect 36026 56244 36032 56256
rect 40844 56244 40850 56256
rect 40902 56244 40908 56296
rect 40936 56244 40942 56296
rect 40994 56284 41000 56296
rect 45996 56284 46002 56296
rect 40994 56256 46002 56284
rect 40994 56244 41000 56256
rect 45996 56244 46002 56256
rect 46054 56244 46060 56296
rect 48667 56287 48725 56293
rect 48667 56253 48679 56287
rect 48713 56284 48725 56287
rect 57496 56284 57502 56296
rect 48713 56256 57502 56284
rect 48713 56253 48725 56256
rect 48667 56247 48725 56253
rect 57496 56244 57502 56256
rect 57554 56244 57560 56296
rect 10116 56176 10122 56228
rect 10174 56216 10180 56228
rect 13152 56216 13158 56228
rect 10174 56188 13158 56216
rect 10174 56176 10180 56188
rect 13152 56176 13158 56188
rect 13210 56176 13216 56228
rect 14440 56176 14446 56228
rect 14498 56216 14504 56228
rect 20788 56216 20794 56228
rect 14498 56188 20794 56216
rect 14498 56176 14504 56188
rect 20788 56176 20794 56188
rect 20846 56176 20852 56228
rect 20880 56176 20886 56228
rect 20938 56216 20944 56228
rect 20938 56188 45490 56216
rect 20938 56176 20944 56188
rect 11680 56108 11686 56160
rect 11738 56148 11744 56160
rect 16832 56148 16838 56160
rect 11738 56120 16838 56148
rect 11738 56108 11744 56120
rect 16832 56108 16838 56120
rect 16890 56108 16896 56160
rect 17108 56108 17114 56160
rect 17166 56148 17172 56160
rect 41304 56148 41310 56160
rect 17166 56120 41310 56148
rect 17166 56108 17172 56120
rect 41304 56108 41310 56120
rect 41362 56108 41368 56160
rect 41396 56108 41402 56160
rect 41454 56148 41460 56160
rect 45352 56148 45358 56160
rect 41454 56120 45358 56148
rect 41454 56108 41460 56120
rect 45352 56108 45358 56120
rect 45410 56108 45416 56160
rect 45462 56148 45490 56188
rect 45536 56176 45542 56228
rect 45594 56216 45600 56228
rect 45594 56188 48710 56216
rect 45594 56176 45600 56188
rect 48572 56148 48578 56160
rect 45462 56120 48578 56148
rect 48572 56108 48578 56120
rect 48630 56108 48636 56160
rect 48682 56148 48710 56188
rect 49124 56176 49130 56228
rect 49182 56216 49188 56228
rect 52712 56216 52718 56228
rect 49182 56188 52718 56216
rect 49182 56176 49188 56188
rect 52712 56176 52718 56188
rect 52770 56176 52776 56228
rect 54828 56148 54834 56160
rect 48682 56120 54834 56148
rect 54828 56108 54834 56120
rect 54886 56108 54892 56160
rect 1086 56058 58862 56080
rect 1086 56006 19588 56058
rect 19640 56006 19652 56058
rect 19704 56006 19716 56058
rect 19768 56006 19780 56058
rect 19832 56006 50308 56058
rect 50360 56006 50372 56058
rect 50424 56006 50436 56058
rect 50488 56006 50500 56058
rect 50552 56006 58862 56058
rect 1086 55984 58862 56006
rect 4044 55904 4050 55956
rect 4102 55944 4108 55956
rect 4102 55916 17614 55944
rect 4102 55904 4108 55916
rect 17586 55876 17614 55916
rect 17752 55904 17758 55956
rect 17810 55944 17816 55956
rect 41212 55944 41218 55956
rect 17810 55916 41218 55944
rect 17810 55904 17816 55916
rect 41212 55904 41218 55916
rect 41270 55904 41276 55956
rect 41304 55904 41310 55956
rect 41362 55944 41368 55956
rect 44708 55944 44714 55956
rect 41362 55916 44714 55944
rect 41362 55904 41368 55916
rect 44708 55904 44714 55916
rect 44766 55904 44772 55956
rect 45996 55904 46002 55956
rect 46054 55944 46060 55956
rect 59060 55944 59066 55956
rect 46054 55916 59066 55944
rect 46054 55904 46060 55916
rect 59060 55904 59066 55916
rect 59118 55904 59124 55956
rect 31736 55876 31742 55888
rect 17586 55848 31742 55876
rect 31736 55836 31742 55848
rect 31794 55836 31800 55888
rect 31828 55836 31834 55888
rect 31886 55876 31892 55888
rect 35416 55876 35422 55888
rect 31886 55848 35422 55876
rect 31886 55836 31892 55848
rect 35416 55836 35422 55848
rect 35474 55836 35480 55888
rect 36152 55836 36158 55888
rect 36210 55876 36216 55888
rect 40660 55876 40666 55888
rect 36210 55848 40666 55876
rect 36210 55836 36216 55848
rect 40660 55836 40666 55848
rect 40718 55836 40724 55888
rect 40752 55836 40758 55888
rect 40810 55876 40816 55888
rect 42224 55876 42230 55888
rect 40810 55848 42230 55876
rect 40810 55836 40816 55848
rect 42224 55836 42230 55848
rect 42282 55836 42288 55888
rect 42316 55836 42322 55888
rect 42374 55876 42380 55888
rect 46088 55876 46094 55888
rect 42374 55848 46094 55876
rect 42374 55836 42380 55848
rect 46088 55836 46094 55848
rect 46146 55836 46152 55888
rect 46180 55836 46186 55888
rect 46238 55876 46244 55888
rect 55932 55876 55938 55888
rect 46238 55848 55938 55876
rect 46238 55836 46244 55848
rect 55932 55836 55938 55848
rect 55990 55836 55996 55888
rect 6344 55768 6350 55820
rect 6402 55808 6408 55820
rect 16924 55808 16930 55820
rect 6402 55780 16930 55808
rect 6402 55768 6408 55780
rect 16924 55768 16930 55780
rect 16982 55768 16988 55820
rect 17568 55808 17574 55820
rect 17218 55780 17574 55808
rect 11404 55700 11410 55752
rect 11462 55740 11468 55752
rect 17108 55740 17114 55752
rect 11462 55712 17114 55740
rect 11462 55700 11468 55712
rect 17108 55700 17114 55712
rect 17166 55700 17172 55752
rect 1836 55632 1842 55684
rect 1894 55672 1900 55684
rect 2572 55672 2578 55684
rect 1894 55644 2578 55672
rect 1894 55632 1900 55644
rect 2572 55632 2578 55644
rect 2630 55632 2636 55684
rect 8184 55632 8190 55684
rect 8242 55672 8248 55684
rect 17218 55672 17246 55780
rect 17568 55768 17574 55780
rect 17626 55768 17632 55820
rect 17660 55768 17666 55820
rect 17718 55808 17724 55820
rect 22720 55808 22726 55820
rect 17718 55780 22726 55808
rect 17718 55768 17724 55780
rect 22720 55768 22726 55780
rect 22778 55768 22784 55820
rect 22904 55768 22910 55820
rect 22962 55808 22968 55820
rect 24928 55808 24934 55820
rect 22962 55780 24934 55808
rect 22962 55768 22968 55780
rect 24928 55768 24934 55780
rect 24986 55768 24992 55820
rect 25664 55768 25670 55820
rect 25722 55808 25728 55820
rect 25722 55780 26078 55808
rect 25722 55768 25728 55780
rect 17292 55700 17298 55752
rect 17350 55740 17356 55752
rect 24376 55740 24382 55752
rect 17350 55712 24382 55740
rect 17350 55700 17356 55712
rect 24376 55700 24382 55712
rect 24434 55700 24440 55752
rect 25940 55740 25946 55752
rect 24486 55712 25946 55740
rect 8242 55644 17246 55672
rect 8242 55632 8248 55644
rect 17384 55632 17390 55684
rect 17442 55672 17448 55684
rect 20880 55672 20886 55684
rect 17442 55644 20886 55672
rect 17442 55632 17448 55644
rect 20880 55632 20886 55644
rect 20938 55632 20944 55684
rect 21340 55632 21346 55684
rect 21398 55672 21404 55684
rect 24486 55672 24514 55712
rect 25940 55700 25946 55712
rect 25998 55700 26004 55752
rect 26050 55740 26078 55780
rect 26124 55768 26130 55820
rect 26182 55808 26188 55820
rect 28148 55808 28154 55820
rect 26182 55780 28154 55808
rect 26182 55768 26188 55780
rect 28148 55768 28154 55780
rect 28206 55768 28212 55820
rect 28332 55768 28338 55820
rect 28390 55808 28396 55820
rect 51148 55808 51154 55820
rect 28390 55780 51154 55808
rect 28390 55768 28396 55780
rect 51148 55768 51154 55780
rect 51206 55768 51212 55820
rect 41396 55740 41402 55752
rect 26050 55712 41402 55740
rect 41396 55700 41402 55712
rect 41454 55700 41460 55752
rect 41488 55700 41494 55752
rect 41546 55740 41552 55752
rect 49124 55740 49130 55752
rect 41546 55712 49130 55740
rect 41546 55700 41552 55712
rect 49124 55700 49130 55712
rect 49182 55700 49188 55752
rect 49234 55712 49446 55740
rect 21398 55644 24514 55672
rect 21398 55632 21404 55644
rect 25204 55632 25210 55684
rect 25262 55672 25268 55684
rect 34312 55672 34318 55684
rect 25262 55644 34318 55672
rect 25262 55632 25268 55644
rect 34312 55632 34318 55644
rect 34370 55632 34376 55684
rect 35324 55632 35330 55684
rect 35382 55672 35388 55684
rect 49234 55672 49262 55712
rect 35382 55644 49262 55672
rect 49418 55672 49446 55712
rect 59612 55672 59618 55684
rect 49418 55644 59618 55672
rect 35382 55632 35388 55644
rect 59612 55632 59618 55644
rect 59670 55632 59676 55684
rect 5059 55607 5117 55613
rect 5059 55573 5071 55607
rect 5105 55604 5117 55607
rect 30448 55604 30454 55616
rect 5105 55576 30454 55604
rect 5105 55573 5117 55576
rect 5059 55567 5117 55573
rect 30448 55564 30454 55576
rect 30506 55564 30512 55616
rect 31736 55564 31742 55616
rect 31794 55604 31800 55616
rect 36152 55604 36158 55616
rect 31794 55576 36158 55604
rect 31794 55564 31800 55576
rect 36152 55564 36158 55576
rect 36210 55564 36216 55616
rect 39648 55564 39654 55616
rect 39706 55604 39712 55616
rect 42040 55604 42046 55616
rect 39706 55576 42046 55604
rect 39706 55564 39712 55576
rect 42040 55564 42046 55576
rect 42098 55564 42104 55616
rect 42132 55564 42138 55616
rect 42190 55604 42196 55616
rect 43788 55604 43794 55616
rect 42190 55576 43794 55604
rect 42190 55564 42196 55576
rect 43788 55564 43794 55576
rect 43846 55564 43852 55616
rect 43880 55564 43886 55616
rect 43938 55604 43944 55616
rect 48296 55604 48302 55616
rect 43938 55576 48302 55604
rect 43938 55564 43944 55576
rect 48296 55564 48302 55576
rect 48354 55564 48360 55616
rect 1086 55514 58862 55536
rect 1086 55462 4228 55514
rect 4280 55462 4292 55514
rect 4344 55462 4356 55514
rect 4408 55462 4420 55514
rect 4472 55462 34948 55514
rect 35000 55462 35012 55514
rect 35064 55462 35076 55514
rect 35128 55462 35140 55514
rect 35192 55462 58862 55514
rect 1086 55440 58862 55462
rect 4872 55360 4878 55412
rect 4930 55400 4936 55412
rect 7448 55400 7454 55412
rect 4930 55372 7454 55400
rect 4930 55360 4936 55372
rect 7448 55360 7454 55372
rect 7506 55360 7512 55412
rect 9840 55360 9846 55412
rect 9898 55400 9904 55412
rect 9898 55372 17246 55400
rect 9898 55360 9904 55372
rect 6988 55292 6994 55344
rect 7046 55332 7052 55344
rect 7908 55332 7914 55344
rect 7046 55304 7914 55332
rect 7046 55292 7052 55304
rect 7908 55292 7914 55304
rect 7966 55292 7972 55344
rect 8276 55292 8282 55344
rect 8334 55332 8340 55344
rect 9564 55332 9570 55344
rect 8334 55304 9570 55332
rect 8334 55292 8340 55304
rect 9564 55292 9570 55304
rect 9622 55292 9628 55344
rect 13060 55292 13066 55344
rect 13118 55332 13124 55344
rect 17108 55332 17114 55344
rect 13118 55304 17114 55332
rect 13118 55292 13124 55304
rect 17108 55292 17114 55304
rect 17166 55292 17172 55344
rect 2756 55224 2762 55276
rect 2814 55264 2820 55276
rect 3768 55264 3774 55276
rect 2814 55236 3774 55264
rect 2814 55224 2820 55236
rect 3768 55224 3774 55236
rect 3826 55224 3832 55276
rect 4596 55224 4602 55276
rect 4654 55264 4660 55276
rect 4654 55236 5378 55264
rect 4654 55224 4660 55236
rect 5350 55072 5378 55236
rect 7540 55224 7546 55276
rect 7598 55264 7604 55276
rect 8092 55264 8098 55276
rect 7598 55236 8098 55264
rect 7598 55224 7604 55236
rect 8092 55224 8098 55236
rect 8150 55224 8156 55276
rect 13244 55224 13250 55276
rect 13302 55264 13308 55276
rect 13704 55264 13710 55276
rect 13302 55236 13710 55264
rect 13302 55224 13308 55236
rect 13704 55224 13710 55236
rect 13762 55224 13768 55276
rect 17218 55264 17246 55372
rect 17568 55360 17574 55412
rect 17626 55400 17632 55412
rect 17626 55372 20742 55400
rect 17626 55360 17632 55372
rect 18028 55292 18034 55344
rect 18086 55332 18092 55344
rect 19224 55332 19230 55344
rect 18086 55304 19230 55332
rect 18086 55292 18092 55304
rect 19224 55292 19230 55304
rect 19282 55292 19288 55344
rect 19868 55292 19874 55344
rect 19926 55332 19932 55344
rect 20604 55332 20610 55344
rect 19926 55304 20610 55332
rect 19926 55292 19932 55304
rect 20604 55292 20610 55304
rect 20662 55292 20668 55344
rect 20714 55332 20742 55372
rect 20788 55360 20794 55412
rect 20846 55400 20852 55412
rect 23272 55400 23278 55412
rect 20846 55372 23278 55400
rect 20846 55360 20852 55372
rect 23272 55360 23278 55372
rect 23330 55360 23336 55412
rect 31276 55400 31282 55412
rect 24026 55372 31282 55400
rect 24026 55332 24054 55372
rect 31276 55360 31282 55372
rect 31334 55360 31340 55412
rect 35232 55400 35238 55412
rect 31570 55372 35238 55400
rect 20714 55304 24054 55332
rect 24100 55292 24106 55344
rect 24158 55332 24164 55344
rect 26400 55332 26406 55344
rect 24158 55304 26406 55332
rect 24158 55292 24164 55304
rect 26400 55292 26406 55304
rect 26458 55292 26464 55344
rect 27044 55292 27050 55344
rect 27102 55332 27108 55344
rect 31570 55332 31598 55372
rect 35232 55360 35238 55372
rect 35290 55360 35296 55412
rect 35416 55360 35422 55412
rect 35474 55400 35480 55412
rect 40752 55400 40758 55412
rect 35474 55372 40758 55400
rect 35474 55360 35480 55372
rect 40752 55360 40758 55372
rect 40810 55360 40816 55412
rect 41672 55360 41678 55412
rect 41730 55400 41736 55412
rect 54368 55400 54374 55412
rect 41730 55372 54374 55400
rect 41730 55360 41736 55372
rect 54368 55360 54374 55372
rect 54426 55360 54432 55412
rect 27102 55304 31598 55332
rect 27102 55292 27108 55304
rect 38544 55292 38550 55344
rect 38602 55332 38608 55344
rect 40660 55332 40666 55344
rect 38602 55304 40666 55332
rect 38602 55292 38608 55304
rect 40660 55292 40666 55304
rect 40718 55292 40724 55344
rect 41028 55292 41034 55344
rect 41086 55332 41092 55344
rect 56392 55332 56398 55344
rect 41086 55304 56398 55332
rect 41086 55292 41092 55304
rect 56392 55292 56398 55304
rect 56450 55292 56456 55344
rect 25204 55264 25210 55276
rect 17218 55236 25210 55264
rect 25204 55224 25210 55236
rect 25262 55224 25268 55276
rect 25572 55224 25578 55276
rect 25630 55264 25636 55276
rect 25630 55236 41810 55264
rect 25630 55224 25636 55236
rect 24192 55156 24198 55208
rect 24250 55196 24256 55208
rect 26124 55196 26130 55208
rect 24250 55168 26130 55196
rect 24250 55156 24256 55168
rect 26124 55156 26130 55168
rect 26182 55156 26188 55208
rect 32196 55156 32202 55208
rect 32254 55196 32260 55208
rect 41672 55196 41678 55208
rect 32254 55168 41678 55196
rect 32254 55156 32260 55168
rect 41672 55156 41678 55168
rect 41730 55156 41736 55208
rect 41782 55196 41810 55236
rect 43236 55224 43242 55276
rect 43294 55264 43300 55276
rect 44064 55264 44070 55276
rect 43294 55236 44070 55264
rect 43294 55224 43300 55236
rect 44064 55224 44070 55236
rect 44122 55224 44128 55276
rect 44892 55196 44898 55208
rect 41782 55168 44898 55196
rect 44892 55156 44898 55168
rect 44950 55156 44956 55208
rect 5332 55020 5338 55072
rect 5390 55020 5396 55072
rect 1086 54970 58862 54992
rect 1086 54918 19588 54970
rect 19640 54918 19652 54970
rect 19704 54918 19716 54970
rect 19768 54918 19780 54970
rect 19832 54918 50308 54970
rect 50360 54918 50372 54970
rect 50424 54918 50436 54970
rect 50488 54918 50500 54970
rect 50552 54918 58862 54970
rect 1086 54896 58862 54918
rect 16832 54816 16838 54868
rect 16890 54856 16896 54868
rect 25483 54859 25541 54865
rect 25483 54856 25495 54859
rect 16890 54828 25495 54856
rect 16890 54816 16896 54828
rect 25483 54825 25495 54828
rect 25529 54825 25541 54859
rect 25483 54819 25541 54825
rect 8552 54748 8558 54800
rect 8610 54788 8616 54800
rect 17111 54791 17169 54797
rect 17111 54788 17123 54791
rect 8610 54760 17123 54788
rect 8610 54748 8616 54760
rect 17111 54757 17123 54760
rect 17157 54757 17169 54791
rect 17111 54751 17169 54757
rect 21432 54680 21438 54732
rect 21490 54720 21496 54732
rect 27596 54720 27602 54732
rect 21490 54692 27602 54720
rect 21490 54680 21496 54692
rect 27596 54680 27602 54692
rect 27654 54680 27660 54732
rect 38636 54680 38642 54732
rect 38694 54720 38700 54732
rect 47839 54723 47897 54729
rect 47839 54720 47851 54723
rect 38694 54692 47851 54720
rect 38694 54680 38700 54692
rect 47839 54689 47851 54692
rect 47885 54689 47897 54723
rect 47839 54683 47897 54689
rect 17111 54655 17169 54661
rect 17111 54621 17123 54655
rect 17157 54652 17169 54655
rect 19132 54652 19138 54664
rect 17157 54624 19138 54652
rect 17157 54621 17169 54624
rect 17111 54615 17169 54621
rect 19132 54612 19138 54624
rect 19190 54612 19196 54664
rect 17384 54516 17390 54528
rect 17345 54488 17390 54516
rect 17384 54476 17390 54488
rect 17442 54476 17448 54528
rect 19132 54476 19138 54528
rect 19190 54516 19196 54528
rect 21432 54516 21438 54528
rect 19190 54488 21438 54516
rect 19190 54476 19196 54488
rect 21432 54476 21438 54488
rect 21490 54476 21496 54528
rect 21616 54516 21622 54528
rect 21577 54488 21622 54516
rect 21616 54476 21622 54488
rect 21674 54476 21680 54528
rect 27596 54476 27602 54528
rect 27654 54516 27660 54528
rect 38636 54516 38642 54528
rect 27654 54488 38642 54516
rect 27654 54476 27660 54488
rect 38636 54476 38642 54488
rect 38694 54476 38700 54528
rect 42408 54516 42414 54528
rect 42369 54488 42414 54516
rect 42408 54476 42414 54488
rect 42466 54476 42472 54528
rect 1086 54426 58862 54448
rect 1086 54374 4228 54426
rect 4280 54374 4292 54426
rect 4344 54374 4356 54426
rect 4408 54374 4420 54426
rect 4472 54374 34948 54426
rect 35000 54374 35012 54426
rect 35064 54374 35076 54426
rect 35128 54374 35140 54426
rect 35192 54374 58862 54426
rect 1086 54352 58862 54374
rect 17384 54272 17390 54324
rect 17442 54312 17448 54324
rect 50596 54312 50602 54324
rect 17442 54284 50602 54312
rect 17442 54272 17448 54284
rect 50596 54272 50602 54284
rect 50654 54272 50660 54324
rect 14808 54204 14814 54256
rect 14866 54244 14872 54256
rect 42408 54244 42414 54256
rect 14866 54216 42414 54244
rect 14866 54204 14872 54216
rect 42408 54204 42414 54216
rect 42466 54204 42472 54256
rect 21616 54136 21622 54188
rect 21674 54176 21680 54188
rect 43420 54176 43426 54188
rect 21674 54148 43426 54176
rect 21674 54136 21680 54148
rect 43420 54136 43426 54148
rect 43478 54136 43484 54188
rect 5703 54111 5761 54117
rect 5703 54077 5715 54111
rect 5749 54108 5761 54111
rect 47560 54108 47566 54120
rect 5749 54080 47566 54108
rect 5749 54077 5761 54080
rect 5703 54071 5761 54077
rect 47560 54068 47566 54080
rect 47618 54068 47624 54120
rect 1086 53882 58862 53904
rect 1086 53830 19588 53882
rect 19640 53830 19652 53882
rect 19704 53830 19716 53882
rect 19768 53830 19780 53882
rect 19832 53830 50308 53882
rect 50360 53830 50372 53882
rect 50424 53830 50436 53882
rect 50488 53830 50500 53882
rect 50552 53830 58862 53882
rect 1086 53808 58862 53830
rect 58048 53592 58054 53644
rect 58106 53632 58112 53644
rect 58327 53635 58385 53641
rect 58327 53632 58339 53635
rect 58106 53604 58339 53632
rect 58106 53592 58112 53604
rect 58327 53601 58339 53604
rect 58373 53601 58385 53635
rect 58327 53595 58385 53601
rect 1086 53338 58862 53360
rect 1086 53286 4228 53338
rect 4280 53286 4292 53338
rect 4344 53286 4356 53338
rect 4408 53286 4420 53338
rect 4472 53286 34948 53338
rect 35000 53286 35012 53338
rect 35064 53286 35076 53338
rect 35128 53286 35140 53338
rect 35192 53286 58862 53338
rect 1086 53264 58862 53286
rect 17016 53224 17022 53236
rect 16977 53196 17022 53224
rect 17016 53184 17022 53196
rect 17074 53184 17080 53236
rect 15268 53116 15274 53168
rect 15326 53156 15332 53168
rect 15728 53156 15734 53168
rect 15326 53128 15734 53156
rect 15326 53116 15332 53128
rect 15728 53116 15734 53128
rect 15786 53116 15792 53168
rect 26492 53116 26498 53168
rect 26550 53156 26556 53168
rect 26952 53156 26958 53168
rect 26550 53128 26958 53156
rect 26550 53116 26556 53128
rect 26952 53116 26958 53128
rect 27010 53116 27016 53168
rect 15268 52980 15274 53032
rect 15326 53020 15332 53032
rect 15912 53020 15918 53032
rect 15326 52992 15918 53020
rect 15326 52980 15332 52992
rect 15912 52980 15918 52992
rect 15970 52980 15976 53032
rect 18580 52980 18586 53032
rect 18638 53020 18644 53032
rect 38271 53023 38329 53029
rect 38271 53020 38283 53023
rect 18638 52992 38283 53020
rect 18638 52980 18644 52992
rect 38271 52989 38283 52992
rect 38317 52989 38329 53023
rect 47563 53023 47621 53029
rect 47563 53020 47575 53023
rect 38271 52983 38329 52989
rect 38378 52992 47575 53020
rect 33024 52912 33030 52964
rect 33082 52952 33088 52964
rect 38378 52952 38406 52992
rect 47563 52989 47575 52992
rect 47609 52989 47621 53023
rect 47563 52983 47621 52989
rect 33082 52924 38406 52952
rect 33082 52912 33088 52924
rect 1086 52794 58862 52816
rect 1086 52742 19588 52794
rect 19640 52742 19652 52794
rect 19704 52742 19716 52794
rect 19768 52742 19780 52794
rect 19832 52742 50308 52794
rect 50360 52742 50372 52794
rect 50424 52742 50436 52794
rect 50488 52742 50500 52794
rect 50552 52742 58862 52794
rect 1086 52720 58862 52742
rect 19227 52343 19285 52349
rect 19227 52309 19239 52343
rect 19273 52340 19285 52343
rect 20328 52340 20334 52352
rect 19273 52312 20334 52340
rect 19273 52309 19285 52312
rect 19227 52303 19285 52309
rect 20328 52300 20334 52312
rect 20386 52300 20392 52352
rect 1086 52250 58862 52272
rect 1086 52198 4228 52250
rect 4280 52198 4292 52250
rect 4344 52198 4356 52250
rect 4408 52198 4420 52250
rect 4472 52198 34948 52250
rect 35000 52198 35012 52250
rect 35064 52198 35076 52250
rect 35128 52198 35140 52250
rect 35192 52198 58862 52250
rect 1086 52176 58862 52198
rect 30448 51892 30454 51944
rect 30506 51932 30512 51944
rect 32380 51932 32386 51944
rect 30506 51904 32386 51932
rect 30506 51892 30512 51904
rect 32380 51892 32386 51904
rect 32438 51892 32444 51944
rect 38544 51892 38550 51944
rect 38602 51932 38608 51944
rect 58419 51935 58477 51941
rect 58419 51932 58431 51935
rect 38602 51904 58431 51932
rect 38602 51892 38608 51904
rect 58419 51901 58431 51904
rect 58465 51901 58477 51935
rect 58419 51895 58477 51901
rect 1086 51706 58862 51728
rect 1086 51654 19588 51706
rect 19640 51654 19652 51706
rect 19704 51654 19716 51706
rect 19768 51654 19780 51706
rect 19832 51654 50308 51706
rect 50360 51654 50372 51706
rect 50424 51654 50436 51706
rect 50488 51654 50500 51706
rect 50552 51654 58862 51706
rect 1086 51632 58862 51654
rect 48388 51484 48394 51536
rect 48446 51524 48452 51536
rect 49032 51524 49038 51536
rect 48446 51496 49038 51524
rect 48446 51484 48452 51496
rect 49032 51484 49038 51496
rect 49090 51484 49096 51536
rect 8739 51255 8797 51261
rect 8739 51221 8751 51255
rect 8785 51252 8797 51255
rect 35232 51252 35238 51264
rect 8785 51224 35238 51252
rect 8785 51221 8797 51224
rect 8739 51215 8797 51221
rect 35232 51212 35238 51224
rect 35290 51212 35296 51264
rect 1086 51162 58862 51184
rect 1086 51110 4228 51162
rect 4280 51110 4292 51162
rect 4344 51110 4356 51162
rect 4408 51110 4420 51162
rect 4472 51110 34948 51162
rect 35000 51110 35012 51162
rect 35064 51110 35076 51162
rect 35128 51110 35140 51162
rect 35192 51110 58862 51162
rect 1086 51088 58862 51110
rect 1376 50668 1382 50720
rect 1434 50708 1440 50720
rect 47655 50711 47713 50717
rect 47655 50708 47667 50711
rect 1434 50680 47667 50708
rect 1434 50668 1440 50680
rect 47655 50677 47667 50680
rect 47701 50677 47713 50711
rect 47655 50671 47713 50677
rect 1086 50618 58862 50640
rect 1086 50566 19588 50618
rect 19640 50566 19652 50618
rect 19704 50566 19716 50618
rect 19768 50566 19780 50618
rect 19832 50566 50308 50618
rect 50360 50566 50372 50618
rect 50424 50566 50436 50618
rect 50488 50566 50500 50618
rect 50552 50566 58862 50618
rect 1086 50544 58862 50566
rect 16467 50167 16525 50173
rect 16467 50133 16479 50167
rect 16513 50164 16525 50167
rect 42040 50164 42046 50176
rect 16513 50136 42046 50164
rect 16513 50133 16525 50136
rect 16467 50127 16525 50133
rect 42040 50124 42046 50136
rect 42098 50124 42104 50176
rect 1086 50074 58862 50096
rect 1086 50022 4228 50074
rect 4280 50022 4292 50074
rect 4344 50022 4356 50074
rect 4408 50022 4420 50074
rect 4472 50022 34948 50074
rect 35000 50022 35012 50074
rect 35064 50022 35076 50074
rect 35128 50022 35140 50074
rect 35192 50022 58862 50074
rect 1086 50000 58862 50022
rect 1086 49530 58862 49552
rect 1086 49478 19588 49530
rect 19640 49478 19652 49530
rect 19704 49478 19716 49530
rect 19768 49478 19780 49530
rect 19832 49478 50308 49530
rect 50360 49478 50372 49530
rect 50424 49478 50436 49530
rect 50488 49478 50500 49530
rect 50552 49478 58862 49530
rect 1086 49456 58862 49478
rect 18304 49308 18310 49360
rect 18362 49348 18368 49360
rect 19040 49348 19046 49360
rect 18362 49320 19046 49348
rect 18362 49308 18368 49320
rect 19040 49308 19046 49320
rect 19098 49308 19104 49360
rect 12324 49036 12330 49088
rect 12382 49076 12388 49088
rect 18307 49079 18365 49085
rect 18307 49076 18319 49079
rect 12382 49048 18319 49076
rect 12382 49036 12388 49048
rect 18307 49045 18319 49048
rect 18353 49045 18365 49079
rect 18307 49039 18365 49045
rect 33487 49079 33545 49085
rect 33487 49045 33499 49079
rect 33533 49076 33545 49079
rect 39280 49076 39286 49088
rect 33533 49048 39286 49076
rect 33533 49045 33545 49048
rect 33487 49039 33545 49045
rect 39280 49036 39286 49048
rect 39338 49036 39344 49088
rect 1086 48986 58862 49008
rect 1086 48934 4228 48986
rect 4280 48934 4292 48986
rect 4344 48934 4356 48986
rect 4408 48934 4420 48986
rect 4472 48934 34948 48986
rect 35000 48934 35012 48986
rect 35064 48934 35076 48986
rect 35128 48934 35140 48986
rect 35192 48934 58862 48986
rect 1086 48912 58862 48934
rect 8000 48628 8006 48680
rect 8058 48668 8064 48680
rect 44619 48671 44677 48677
rect 44619 48668 44631 48671
rect 8058 48640 44631 48668
rect 8058 48628 8064 48640
rect 44619 48637 44631 48640
rect 44665 48637 44677 48671
rect 44619 48631 44677 48637
rect 49219 48671 49277 48677
rect 49219 48637 49231 48671
rect 49265 48668 49277 48671
rect 53080 48668 53086 48680
rect 49265 48640 53086 48668
rect 49265 48637 49277 48640
rect 49219 48631 49277 48637
rect 53080 48628 53086 48640
rect 53138 48628 53144 48680
rect 1086 48442 58862 48464
rect 1086 48390 19588 48442
rect 19640 48390 19652 48442
rect 19704 48390 19716 48442
rect 19768 48390 19780 48442
rect 19832 48390 50308 48442
rect 50360 48390 50372 48442
rect 50424 48390 50436 48442
rect 50488 48390 50500 48442
rect 50552 48390 58862 48442
rect 1086 48368 58862 48390
rect 29344 48288 29350 48340
rect 29402 48328 29408 48340
rect 30172 48328 30178 48340
rect 29402 48300 30178 48328
rect 29402 48288 29408 48300
rect 30172 48288 30178 48300
rect 30230 48288 30236 48340
rect 31644 48288 31650 48340
rect 31702 48328 31708 48340
rect 32656 48328 32662 48340
rect 31702 48300 32662 48328
rect 31702 48288 31708 48300
rect 32656 48288 32662 48300
rect 32714 48288 32720 48340
rect 39096 48288 39102 48340
rect 39154 48328 39160 48340
rect 39464 48328 39470 48340
rect 39154 48300 39470 48328
rect 39154 48288 39160 48300
rect 39464 48288 39470 48300
rect 39522 48288 39528 48340
rect 6712 47948 6718 48000
rect 6770 47988 6776 48000
rect 16835 47991 16893 47997
rect 16835 47988 16847 47991
rect 6770 47960 16847 47988
rect 6770 47948 6776 47960
rect 16835 47957 16847 47960
rect 16881 47957 16893 47991
rect 16835 47951 16893 47957
rect 1086 47898 58862 47920
rect 1086 47846 4228 47898
rect 4280 47846 4292 47898
rect 4344 47846 4356 47898
rect 4408 47846 4420 47898
rect 4472 47846 34948 47898
rect 35000 47846 35012 47898
rect 35064 47846 35076 47898
rect 35128 47846 35140 47898
rect 35192 47846 58862 47898
rect 1086 47824 58862 47846
rect 9935 47651 9993 47657
rect 9935 47617 9947 47651
rect 9981 47648 9993 47651
rect 19408 47648 19414 47660
rect 9981 47620 19414 47648
rect 9981 47617 9993 47620
rect 9935 47611 9993 47617
rect 19408 47608 19414 47620
rect 19466 47608 19472 47660
rect 3860 47540 3866 47592
rect 3918 47580 3924 47592
rect 45723 47583 45781 47589
rect 45723 47580 45735 47583
rect 3918 47552 45735 47580
rect 3918 47540 3924 47552
rect 45723 47549 45735 47552
rect 45769 47549 45781 47583
rect 45723 47543 45781 47549
rect 14627 47447 14685 47453
rect 14627 47413 14639 47447
rect 14673 47444 14685 47447
rect 24192 47444 24198 47456
rect 14673 47416 24198 47444
rect 14673 47413 14685 47416
rect 14627 47407 14685 47413
rect 24192 47404 24198 47416
rect 24250 47404 24256 47456
rect 44064 47404 44070 47456
rect 44122 47444 44128 47456
rect 57683 47447 57741 47453
rect 57683 47444 57695 47447
rect 44122 47416 57695 47444
rect 44122 47404 44128 47416
rect 57683 47413 57695 47416
rect 57729 47413 57741 47447
rect 57683 47407 57741 47413
rect 1086 47354 58862 47376
rect 1086 47302 19588 47354
rect 19640 47302 19652 47354
rect 19704 47302 19716 47354
rect 19768 47302 19780 47354
rect 19832 47302 50308 47354
rect 50360 47302 50372 47354
rect 50424 47302 50436 47354
rect 50488 47302 50500 47354
rect 50552 47302 58862 47354
rect 1086 47280 58862 47302
rect 8644 47132 8650 47184
rect 8702 47172 8708 47184
rect 9104 47172 9110 47184
rect 8702 47144 9110 47172
rect 8702 47132 8708 47144
rect 9104 47132 9110 47144
rect 9162 47132 9168 47184
rect 24744 46928 24750 46980
rect 24802 46968 24808 46980
rect 26771 46971 26829 46977
rect 26771 46968 26783 46971
rect 24802 46940 26783 46968
rect 24802 46928 24808 46940
rect 26771 46937 26783 46940
rect 26817 46937 26829 46971
rect 26771 46931 26829 46937
rect 26400 46860 26406 46912
rect 26458 46900 26464 46912
rect 26492 46900 26498 46912
rect 26458 46872 26498 46900
rect 26458 46860 26464 46872
rect 26492 46860 26498 46872
rect 26550 46860 26556 46912
rect 29344 46860 29350 46912
rect 29402 46900 29408 46912
rect 29528 46900 29534 46912
rect 29402 46872 29534 46900
rect 29402 46860 29408 46872
rect 29528 46860 29534 46872
rect 29586 46860 29592 46912
rect 48296 46860 48302 46912
rect 48354 46900 48360 46912
rect 48388 46900 48394 46912
rect 48354 46872 48394 46900
rect 48354 46860 48360 46872
rect 48388 46860 48394 46872
rect 48446 46860 48452 46912
rect 1086 46810 58862 46832
rect 1086 46758 4228 46810
rect 4280 46758 4292 46810
rect 4344 46758 4356 46810
rect 4408 46758 4420 46810
rect 4472 46758 34948 46810
rect 35000 46758 35012 46810
rect 35064 46758 35076 46810
rect 35128 46758 35140 46810
rect 35192 46758 58862 46810
rect 1086 46736 58862 46758
rect 5335 46495 5393 46501
rect 5335 46461 5347 46495
rect 5381 46461 5393 46495
rect 5335 46455 5393 46461
rect 5350 46424 5378 46455
rect 46824 46452 46830 46504
rect 46882 46492 46888 46504
rect 52071 46495 52129 46501
rect 52071 46492 52083 46495
rect 46882 46464 52083 46492
rect 46882 46452 46888 46464
rect 52071 46461 52083 46464
rect 52117 46461 52129 46495
rect 52071 46455 52129 46461
rect 50688 46424 50694 46436
rect 5350 46396 50694 46424
rect 50688 46384 50694 46396
rect 50746 46384 50752 46436
rect 1086 46266 58862 46288
rect 1086 46214 19588 46266
rect 19640 46214 19652 46266
rect 19704 46214 19716 46266
rect 19768 46214 19780 46266
rect 19832 46214 50308 46266
rect 50360 46214 50372 46266
rect 50424 46214 50436 46266
rect 50488 46214 50500 46266
rect 50552 46214 58862 46266
rect 1086 46192 58862 46214
rect 1086 45722 58862 45744
rect 1086 45670 4228 45722
rect 4280 45670 4292 45722
rect 4344 45670 4356 45722
rect 4408 45670 4420 45722
rect 4472 45670 34948 45722
rect 35000 45670 35012 45722
rect 35064 45670 35076 45722
rect 35128 45670 35140 45722
rect 35192 45670 58862 45722
rect 1086 45648 58862 45670
rect 34312 45568 34318 45620
rect 34370 45608 34376 45620
rect 34772 45608 34778 45620
rect 34370 45580 34778 45608
rect 34370 45568 34376 45580
rect 34772 45568 34778 45580
rect 34830 45568 34836 45620
rect 8920 45500 8926 45552
rect 8978 45540 8984 45552
rect 9104 45540 9110 45552
rect 8978 45512 9110 45540
rect 8978 45500 8984 45512
rect 9104 45500 9110 45512
rect 9162 45500 9168 45552
rect 14164 45500 14170 45552
rect 14222 45540 14228 45552
rect 14440 45540 14446 45552
rect 14222 45512 14446 45540
rect 14222 45500 14228 45512
rect 14440 45500 14446 45512
rect 14498 45500 14504 45552
rect 39832 45364 39838 45416
rect 39890 45404 39896 45416
rect 40755 45407 40813 45413
rect 40755 45404 40767 45407
rect 39890 45376 40767 45404
rect 39890 45364 39896 45376
rect 40755 45373 40767 45376
rect 40801 45373 40813 45407
rect 40755 45367 40813 45373
rect 1086 45178 58862 45200
rect 1086 45126 19588 45178
rect 19640 45126 19652 45178
rect 19704 45126 19716 45178
rect 19768 45126 19780 45178
rect 19832 45126 50308 45178
rect 50360 45126 50372 45178
rect 50424 45126 50436 45178
rect 50488 45126 50500 45178
rect 50552 45126 58862 45178
rect 1086 45104 58862 45126
rect 16832 45064 16838 45076
rect 16793 45036 16838 45064
rect 16832 45024 16838 45036
rect 16890 45024 16896 45076
rect 2296 44724 2302 44736
rect 2257 44696 2302 44724
rect 2296 44684 2302 44696
rect 2354 44684 2360 44736
rect 24471 44727 24529 44733
rect 24471 44693 24483 44727
rect 24517 44724 24529 44727
rect 26860 44724 26866 44736
rect 24517 44696 26866 44724
rect 24517 44693 24529 44696
rect 24471 44687 24529 44693
rect 26860 44684 26866 44696
rect 26918 44684 26924 44736
rect 37164 44684 37170 44736
rect 37222 44724 37228 44736
rect 47655 44727 47713 44733
rect 47655 44724 47667 44727
rect 37222 44696 47667 44724
rect 37222 44684 37228 44696
rect 47655 44693 47667 44696
rect 47701 44693 47713 44727
rect 47655 44687 47713 44693
rect 50964 44684 50970 44736
rect 51022 44724 51028 44736
rect 55843 44727 55901 44733
rect 55843 44724 55855 44727
rect 51022 44696 55855 44724
rect 51022 44684 51028 44696
rect 55843 44693 55855 44696
rect 55889 44693 55901 44727
rect 56944 44724 56950 44736
rect 56905 44696 56950 44724
rect 55843 44687 55901 44693
rect 56944 44684 56950 44696
rect 57002 44684 57008 44736
rect 1086 44634 58862 44656
rect 1086 44582 4228 44634
rect 4280 44582 4292 44634
rect 4344 44582 4356 44634
rect 4408 44582 4420 44634
rect 4472 44582 34948 44634
rect 35000 44582 35012 44634
rect 35064 44582 35076 44634
rect 35128 44582 35140 44634
rect 35192 44582 58862 44634
rect 1086 44560 58862 44582
rect 23364 44480 23370 44532
rect 23422 44520 23428 44532
rect 56944 44520 56950 44532
rect 23422 44492 56950 44520
rect 23422 44480 23428 44492
rect 56944 44480 56950 44492
rect 57002 44480 57008 44532
rect 2296 44412 2302 44464
rect 2354 44452 2360 44464
rect 39372 44452 39378 44464
rect 2354 44424 39378 44452
rect 2354 44412 2360 44424
rect 39372 44412 39378 44424
rect 39430 44412 39436 44464
rect 1086 44090 58862 44112
rect 1086 44038 19588 44090
rect 19640 44038 19652 44090
rect 19704 44038 19716 44090
rect 19768 44038 19780 44090
rect 19832 44038 50308 44090
rect 50360 44038 50372 44090
rect 50424 44038 50436 44090
rect 50488 44038 50500 44090
rect 50552 44038 58862 44090
rect 1086 44016 58862 44038
rect 1086 43546 58862 43568
rect 1086 43494 4228 43546
rect 4280 43494 4292 43546
rect 4344 43494 4356 43546
rect 4408 43494 4420 43546
rect 4472 43494 34948 43546
rect 35000 43494 35012 43546
rect 35064 43494 35076 43546
rect 35128 43494 35140 43546
rect 35192 43494 58862 43546
rect 1086 43472 58862 43494
rect 40108 43432 40114 43444
rect 40069 43404 40114 43432
rect 40108 43392 40114 43404
rect 40166 43392 40172 43444
rect 4522 43268 5838 43296
rect 2572 43188 2578 43240
rect 2630 43228 2636 43240
rect 4522 43228 4550 43268
rect 2630 43200 4550 43228
rect 5703 43231 5761 43237
rect 2630 43188 2636 43200
rect 5703 43197 5715 43231
rect 5749 43197 5761 43231
rect 5810 43228 5838 43268
rect 40663 43231 40721 43237
rect 40663 43228 40675 43231
rect 5810 43200 40675 43228
rect 5703 43191 5761 43197
rect 40663 43197 40675 43200
rect 40709 43197 40721 43231
rect 40663 43191 40721 43197
rect 5718 43160 5746 43191
rect 40752 43160 40758 43172
rect 5718 43132 40758 43160
rect 40752 43120 40758 43132
rect 40810 43120 40816 43172
rect 1086 43002 58862 43024
rect 1086 42950 19588 43002
rect 19640 42950 19652 43002
rect 19704 42950 19716 43002
rect 19768 42950 19780 43002
rect 19832 42950 50308 43002
rect 50360 42950 50372 43002
rect 50424 42950 50436 43002
rect 50488 42950 50500 43002
rect 50552 42950 58862 43002
rect 1086 42928 58862 42950
rect 16464 42644 16470 42696
rect 16522 42684 16528 42696
rect 32751 42687 32809 42693
rect 32751 42684 32763 42687
rect 16522 42656 32763 42684
rect 16522 42644 16528 42656
rect 32751 42653 32763 42656
rect 32797 42653 32809 42687
rect 32751 42647 32809 42653
rect 1086 42458 58862 42480
rect 1086 42406 4228 42458
rect 4280 42406 4292 42458
rect 4344 42406 4356 42458
rect 4408 42406 4420 42458
rect 4472 42406 34948 42458
rect 35000 42406 35012 42458
rect 35064 42406 35076 42458
rect 35128 42406 35140 42458
rect 35192 42406 58862 42458
rect 1086 42384 58862 42406
rect 22171 42347 22229 42353
rect 22171 42313 22183 42347
rect 22217 42344 22229 42347
rect 22447 42347 22505 42353
rect 22447 42344 22459 42347
rect 22217 42316 22459 42344
rect 22217 42313 22229 42316
rect 22171 42307 22229 42313
rect 22447 42313 22459 42316
rect 22493 42313 22505 42347
rect 22447 42307 22505 42313
rect 40203 42347 40261 42353
rect 40203 42313 40215 42347
rect 40249 42344 40261 42347
rect 42132 42344 42138 42356
rect 40249 42316 42138 42344
rect 40249 42313 40261 42316
rect 40203 42307 40261 42313
rect 42132 42304 42138 42316
rect 42190 42304 42196 42356
rect 13612 42236 13618 42288
rect 13670 42276 13676 42288
rect 13670 42248 26906 42276
rect 13670 42236 13676 42248
rect 18215 42211 18273 42217
rect 18215 42177 18227 42211
rect 18261 42208 18273 42211
rect 18261 42180 22582 42208
rect 18261 42177 18273 42180
rect 18215 42171 18273 42177
rect 8739 42143 8797 42149
rect 8739 42109 8751 42143
rect 8785 42140 8797 42143
rect 17200 42140 17206 42152
rect 8785 42112 17206 42140
rect 8785 42109 8797 42112
rect 8739 42103 8797 42109
rect 17200 42100 17206 42112
rect 17258 42100 17264 42152
rect 22554 42072 22582 42180
rect 26878 42140 26906 42248
rect 29623 42211 29681 42217
rect 29623 42177 29635 42211
rect 29669 42208 29681 42211
rect 31000 42208 31006 42220
rect 29669 42180 31006 42208
rect 29669 42177 29681 42180
rect 29623 42171 29681 42177
rect 31000 42168 31006 42180
rect 31058 42168 31064 42220
rect 37627 42143 37685 42149
rect 37627 42140 37639 42143
rect 26878 42112 37639 42140
rect 37627 42109 37639 42112
rect 37673 42109 37685 42143
rect 37627 42103 37685 42109
rect 37900 42072 37906 42084
rect 22554 42044 37906 42072
rect 37900 42032 37906 42044
rect 37958 42032 37964 42084
rect 3860 41964 3866 42016
rect 3918 42004 3924 42016
rect 22171 42007 22229 42013
rect 22171 42004 22183 42007
rect 3918 41976 22183 42004
rect 3918 41964 3924 41976
rect 22171 41973 22183 41976
rect 22217 41973 22229 42007
rect 22171 41967 22229 41973
rect 1086 41914 58862 41936
rect 1086 41862 19588 41914
rect 19640 41862 19652 41914
rect 19704 41862 19716 41914
rect 19768 41862 19780 41914
rect 19832 41862 50308 41914
rect 50360 41862 50372 41914
rect 50424 41862 50436 41914
rect 50488 41862 50500 41914
rect 50552 41862 58862 41914
rect 1086 41840 58862 41862
rect 17200 41760 17206 41812
rect 17258 41800 17264 41812
rect 27044 41800 27050 41812
rect 17258 41772 27050 41800
rect 17258 41760 17264 41772
rect 27044 41760 27050 41772
rect 27102 41760 27108 41812
rect 13523 41667 13581 41673
rect 13523 41633 13535 41667
rect 13569 41664 13581 41667
rect 13796 41664 13802 41676
rect 13569 41636 13802 41664
rect 13569 41633 13581 41636
rect 13523 41627 13581 41633
rect 13796 41624 13802 41636
rect 13854 41624 13860 41676
rect 42227 41463 42285 41469
rect 42227 41429 42239 41463
rect 42273 41460 42285 41463
rect 43512 41460 43518 41472
rect 42273 41432 43518 41460
rect 42273 41429 42285 41432
rect 42227 41423 42285 41429
rect 43512 41420 43518 41432
rect 43570 41420 43576 41472
rect 1086 41370 58862 41392
rect 1086 41318 4228 41370
rect 4280 41318 4292 41370
rect 4344 41318 4356 41370
rect 4408 41318 4420 41370
rect 4472 41318 34948 41370
rect 35000 41318 35012 41370
rect 35064 41318 35076 41370
rect 35128 41318 35140 41370
rect 35192 41318 58862 41370
rect 1086 41296 58862 41318
rect 38820 41080 38826 41132
rect 38878 41120 38884 41132
rect 39096 41120 39102 41132
rect 38878 41092 39102 41120
rect 38878 41080 38884 41092
rect 39096 41080 39102 41092
rect 39154 41080 39160 41132
rect 43144 41012 43150 41064
rect 43202 41052 43208 41064
rect 46275 41055 46333 41061
rect 46275 41052 46287 41055
rect 43202 41024 46287 41052
rect 43202 41012 43208 41024
rect 46275 41021 46287 41024
rect 46321 41021 46333 41055
rect 46275 41015 46333 41021
rect 50872 41012 50878 41064
rect 50930 41052 50936 41064
rect 57867 41055 57925 41061
rect 57867 41052 57879 41055
rect 50930 41024 57879 41052
rect 50930 41012 50936 41024
rect 57867 41021 57879 41024
rect 57913 41021 57925 41055
rect 57867 41015 57925 41021
rect 1086 40826 58862 40848
rect 1086 40774 19588 40826
rect 19640 40774 19652 40826
rect 19704 40774 19716 40826
rect 19768 40774 19780 40826
rect 19832 40774 50308 40826
rect 50360 40774 50372 40826
rect 50424 40774 50436 40826
rect 50488 40774 50500 40826
rect 50552 40774 58862 40826
rect 1086 40752 58862 40774
rect 3676 40400 3682 40452
rect 3734 40440 3740 40452
rect 3734 40412 12002 40440
rect 3734 40400 3740 40412
rect 11864 40372 11870 40384
rect 11825 40344 11870 40372
rect 11864 40332 11870 40344
rect 11922 40332 11928 40384
rect 11974 40372 12002 40412
rect 43699 40375 43757 40381
rect 43699 40372 43711 40375
rect 11974 40344 43711 40372
rect 43699 40341 43711 40344
rect 43745 40341 43757 40375
rect 43699 40335 43757 40341
rect 1086 40282 58862 40304
rect 1086 40230 4228 40282
rect 4280 40230 4292 40282
rect 4344 40230 4356 40282
rect 4408 40230 4420 40282
rect 4472 40230 34948 40282
rect 35000 40230 35012 40282
rect 35064 40230 35076 40282
rect 35128 40230 35140 40282
rect 35192 40230 58862 40282
rect 1086 40208 58862 40230
rect 11864 40128 11870 40180
rect 11922 40168 11928 40180
rect 24192 40168 24198 40180
rect 11922 40140 24198 40168
rect 11922 40128 11928 40140
rect 24192 40128 24198 40140
rect 24250 40128 24256 40180
rect 38452 40128 38458 40180
rect 38510 40168 38516 40180
rect 47011 40171 47069 40177
rect 47011 40168 47023 40171
rect 38510 40140 47023 40168
rect 38510 40128 38516 40140
rect 47011 40137 47023 40140
rect 47057 40137 47069 40171
rect 47011 40131 47069 40137
rect 23272 40060 23278 40112
rect 23330 40100 23336 40112
rect 48759 40103 48817 40109
rect 48759 40100 48771 40103
rect 23330 40072 48771 40100
rect 23330 40060 23336 40072
rect 48759 40069 48771 40072
rect 48805 40069 48817 40103
rect 48759 40063 48817 40069
rect 26952 40032 26958 40044
rect 26913 40004 26958 40032
rect 26952 39992 26958 40004
rect 27010 39992 27016 40044
rect 1086 39738 58862 39760
rect 1086 39686 19588 39738
rect 19640 39686 19652 39738
rect 19704 39686 19716 39738
rect 19768 39686 19780 39738
rect 19832 39686 50308 39738
rect 50360 39686 50372 39738
rect 50424 39686 50436 39738
rect 50488 39686 50500 39738
rect 50552 39686 58862 39738
rect 1086 39664 58862 39686
rect 10947 39287 11005 39293
rect 10947 39253 10959 39287
rect 10993 39284 11005 39287
rect 42132 39284 42138 39296
rect 10993 39256 42138 39284
rect 10993 39253 11005 39256
rect 10947 39247 11005 39253
rect 42132 39244 42138 39256
rect 42190 39244 42196 39296
rect 1086 39194 58862 39216
rect 1086 39142 4228 39194
rect 4280 39142 4292 39194
rect 4344 39142 4356 39194
rect 4408 39142 4420 39194
rect 4472 39142 34948 39194
rect 35000 39142 35012 39194
rect 35064 39142 35076 39194
rect 35128 39142 35140 39194
rect 35192 39142 58862 39194
rect 1086 39120 58862 39142
rect 1836 39080 1842 39092
rect 1797 39052 1842 39080
rect 1836 39040 1842 39052
rect 1894 39040 1900 39092
rect 4780 38904 4786 38956
rect 4838 38944 4844 38956
rect 21435 38947 21493 38953
rect 21435 38944 21447 38947
rect 4838 38916 21447 38944
rect 4838 38904 4844 38916
rect 21435 38913 21447 38916
rect 21481 38913 21493 38947
rect 21435 38907 21493 38913
rect 12603 38879 12661 38885
rect 12603 38845 12615 38879
rect 12649 38876 12661 38879
rect 16280 38876 16286 38888
rect 12649 38848 16286 38876
rect 12649 38845 12661 38848
rect 12603 38839 12661 38845
rect 16280 38836 16286 38848
rect 16338 38836 16344 38888
rect 1086 38650 58862 38672
rect 1086 38598 19588 38650
rect 19640 38598 19652 38650
rect 19704 38598 19716 38650
rect 19768 38598 19780 38650
rect 19832 38598 50308 38650
rect 50360 38598 50372 38650
rect 50424 38598 50436 38650
rect 50488 38598 50500 38650
rect 50552 38598 58862 38650
rect 1086 38576 58862 38598
rect 1655 38199 1713 38205
rect 1655 38165 1667 38199
rect 1701 38196 1713 38199
rect 28240 38196 28246 38208
rect 1701 38168 28246 38196
rect 1701 38165 1713 38168
rect 1655 38159 1713 38165
rect 28240 38156 28246 38168
rect 28298 38156 28304 38208
rect 47836 38196 47842 38208
rect 47797 38168 47842 38196
rect 47836 38156 47842 38168
rect 47894 38156 47900 38208
rect 1086 38106 58862 38128
rect 1086 38054 4228 38106
rect 4280 38054 4292 38106
rect 4344 38054 4356 38106
rect 4408 38054 4420 38106
rect 4472 38054 34948 38106
rect 35000 38054 35012 38106
rect 35064 38054 35076 38106
rect 35128 38054 35140 38106
rect 35192 38054 58862 38106
rect 1086 38032 58862 38054
rect 51703 37859 51761 37865
rect 51703 37825 51715 37859
rect 51749 37856 51761 37859
rect 52071 37859 52129 37865
rect 52071 37856 52083 37859
rect 51749 37828 52083 37856
rect 51749 37825 51761 37828
rect 51703 37819 51761 37825
rect 52071 37825 52083 37828
rect 52117 37825 52129 37859
rect 52071 37819 52129 37825
rect 49492 37748 49498 37800
rect 49550 37788 49556 37800
rect 49771 37791 49829 37797
rect 49771 37788 49783 37791
rect 49550 37760 49783 37788
rect 49550 37748 49556 37760
rect 49771 37757 49783 37760
rect 49817 37757 49829 37791
rect 49771 37751 49829 37757
rect 50507 37791 50565 37797
rect 50507 37757 50519 37791
rect 50553 37757 50565 37791
rect 50507 37751 50565 37757
rect 21892 37680 21898 37732
rect 21950 37720 21956 37732
rect 50522 37720 50550 37751
rect 21950 37692 50550 37720
rect 21950 37680 21956 37692
rect 8552 37612 8558 37664
rect 8610 37652 8616 37664
rect 51703 37655 51761 37661
rect 51703 37652 51715 37655
rect 8610 37624 51715 37652
rect 8610 37612 8616 37624
rect 51703 37621 51715 37624
rect 51749 37621 51761 37655
rect 51703 37615 51761 37621
rect 1086 37562 58862 37584
rect 1086 37510 19588 37562
rect 19640 37510 19652 37562
rect 19704 37510 19716 37562
rect 19768 37510 19780 37562
rect 19832 37510 50308 37562
rect 50360 37510 50372 37562
rect 50424 37510 50436 37562
rect 50488 37510 50500 37562
rect 50552 37510 58862 37562
rect 1086 37488 58862 37510
rect 3492 37272 3498 37324
rect 3550 37312 3556 37324
rect 4780 37312 4786 37324
rect 3550 37284 4786 37312
rect 3550 37272 3556 37284
rect 4780 37272 4786 37284
rect 4838 37272 4844 37324
rect 12048 37272 12054 37324
rect 12106 37312 12112 37324
rect 19132 37312 19138 37324
rect 12106 37284 19138 37312
rect 12106 37272 12112 37284
rect 19132 37272 19138 37284
rect 19190 37272 19196 37324
rect 26400 37272 26406 37324
rect 26458 37312 26464 37324
rect 26492 37312 26498 37324
rect 26458 37284 26498 37312
rect 26458 37272 26464 37284
rect 26492 37272 26498 37284
rect 26550 37272 26556 37324
rect 27504 37272 27510 37324
rect 27562 37312 27568 37324
rect 43607 37315 43665 37321
rect 43607 37312 43619 37315
rect 27562 37284 43619 37312
rect 27562 37272 27568 37284
rect 43607 37281 43619 37284
rect 43653 37281 43665 37315
rect 43607 37275 43665 37281
rect 48296 37272 48302 37324
rect 48354 37312 48360 37324
rect 48388 37312 48394 37324
rect 48354 37284 48394 37312
rect 48354 37272 48360 37284
rect 48388 37272 48394 37284
rect 48446 37272 48452 37324
rect 49768 37272 49774 37324
rect 49826 37312 49832 37324
rect 49860 37312 49866 37324
rect 49826 37284 49866 37312
rect 49826 37272 49832 37284
rect 49860 37272 49866 37284
rect 49918 37272 49924 37324
rect 27780 37204 27786 37256
rect 27838 37244 27844 37256
rect 27838 37216 37302 37244
rect 27838 37204 27844 37216
rect 12968 37108 12974 37120
rect 12929 37080 12974 37108
rect 12968 37068 12974 37080
rect 13026 37068 13032 37120
rect 26676 37108 26682 37120
rect 26637 37080 26682 37108
rect 26676 37068 26682 37080
rect 26734 37068 26740 37120
rect 29252 37108 29258 37120
rect 29213 37080 29258 37108
rect 29252 37068 29258 37080
rect 29310 37068 29316 37120
rect 31092 37108 31098 37120
rect 31053 37080 31098 37108
rect 31092 37068 31098 37080
rect 31150 37068 31156 37120
rect 37274 37108 37302 37216
rect 47836 37204 47842 37256
rect 47894 37244 47900 37256
rect 48020 37244 48026 37256
rect 47894 37216 48026 37244
rect 47894 37204 47900 37216
rect 48020 37204 48026 37216
rect 48078 37204 48084 37256
rect 42776 37136 42782 37188
rect 42834 37176 42840 37188
rect 43144 37176 43150 37188
rect 42834 37148 43150 37176
rect 42834 37136 42840 37148
rect 43144 37136 43150 37148
rect 43202 37136 43208 37188
rect 47379 37111 47437 37117
rect 47379 37108 47391 37111
rect 37274 37080 47391 37108
rect 47379 37077 47391 37080
rect 47425 37077 47437 37111
rect 47379 37071 47437 37077
rect 1086 37018 58862 37040
rect 1086 36966 4228 37018
rect 4280 36966 4292 37018
rect 4344 36966 4356 37018
rect 4408 36966 4420 37018
rect 4472 36966 34948 37018
rect 35000 36966 35012 37018
rect 35064 36966 35076 37018
rect 35128 36966 35140 37018
rect 35192 36966 58862 37018
rect 1086 36944 58862 36966
rect 14992 36864 14998 36916
rect 15050 36904 15056 36916
rect 26676 36904 26682 36916
rect 15050 36876 26682 36904
rect 15050 36864 15056 36876
rect 26676 36864 26682 36876
rect 26734 36864 26740 36916
rect 29252 36864 29258 36916
rect 29310 36904 29316 36916
rect 46272 36904 46278 36916
rect 29310 36876 46278 36904
rect 29310 36864 29316 36876
rect 46272 36864 46278 36876
rect 46330 36864 46336 36916
rect 31647 36703 31705 36709
rect 31647 36669 31659 36703
rect 31693 36669 31705 36703
rect 31647 36663 31705 36669
rect 31662 36632 31690 36663
rect 37072 36660 37078 36712
rect 37130 36700 37136 36712
rect 45263 36703 45321 36709
rect 45263 36700 45275 36703
rect 37130 36672 45275 36700
rect 37130 36660 37136 36672
rect 45263 36669 45275 36672
rect 45309 36669 45321 36703
rect 45263 36663 45321 36669
rect 50780 36632 50786 36644
rect 31662 36604 50786 36632
rect 50780 36592 50786 36604
rect 50838 36592 50844 36644
rect 1086 36474 58862 36496
rect 1086 36422 19588 36474
rect 19640 36422 19652 36474
rect 19704 36422 19716 36474
rect 19768 36422 19780 36474
rect 19832 36422 50308 36474
rect 50360 36422 50372 36474
rect 50424 36422 50436 36474
rect 50488 36422 50500 36474
rect 50552 36422 58862 36474
rect 1086 36400 58862 36422
rect 13520 35980 13526 36032
rect 13578 36020 13584 36032
rect 45631 36023 45689 36029
rect 45631 36020 45643 36023
rect 13578 35992 45643 36020
rect 13578 35980 13584 35992
rect 45631 35989 45643 35992
rect 45677 35989 45689 36023
rect 45631 35983 45689 35989
rect 1086 35930 58862 35952
rect 1086 35878 4228 35930
rect 4280 35878 4292 35930
rect 4344 35878 4356 35930
rect 4408 35878 4420 35930
rect 4472 35878 34948 35930
rect 35000 35878 35012 35930
rect 35064 35878 35076 35930
rect 35128 35878 35140 35930
rect 35192 35878 58862 35930
rect 1086 35856 58862 35878
rect 12232 35572 12238 35624
rect 12290 35612 12296 35624
rect 25759 35615 25817 35621
rect 25759 35612 25771 35615
rect 12290 35584 25771 35612
rect 12290 35572 12296 35584
rect 25759 35581 25771 35584
rect 25805 35581 25817 35615
rect 25759 35575 25817 35581
rect 1086 35386 58862 35408
rect 1086 35334 19588 35386
rect 19640 35334 19652 35386
rect 19704 35334 19716 35386
rect 19768 35334 19780 35386
rect 19832 35334 50308 35386
rect 50360 35334 50372 35386
rect 50424 35334 50436 35386
rect 50488 35334 50500 35386
rect 50552 35334 58862 35386
rect 1086 35312 58862 35334
rect 30635 35139 30693 35145
rect 30635 35105 30647 35139
rect 30681 35136 30693 35139
rect 32564 35136 32570 35148
rect 30681 35108 32570 35136
rect 30681 35105 30693 35108
rect 30635 35099 30693 35105
rect 32564 35096 32570 35108
rect 32622 35096 32628 35148
rect 52896 34932 52902 34944
rect 52857 34904 52902 34932
rect 52896 34892 52902 34904
rect 52954 34892 52960 34944
rect 1086 34842 58862 34864
rect 1086 34790 4228 34842
rect 4280 34790 4292 34842
rect 4344 34790 4356 34842
rect 4408 34790 4420 34842
rect 4472 34790 34948 34842
rect 35000 34790 35012 34842
rect 35064 34790 35076 34842
rect 35128 34790 35140 34842
rect 35192 34790 58862 34842
rect 1086 34768 58862 34790
rect 2480 34688 2486 34740
rect 2538 34728 2544 34740
rect 52896 34728 52902 34740
rect 2538 34700 52902 34728
rect 2538 34688 2544 34700
rect 52896 34688 52902 34700
rect 52954 34688 52960 34740
rect 20791 34663 20849 34669
rect 20791 34629 20803 34663
rect 20837 34660 20849 34663
rect 25572 34660 25578 34672
rect 20837 34632 25578 34660
rect 20837 34629 20849 34632
rect 20791 34623 20849 34629
rect 25572 34620 25578 34632
rect 25630 34620 25636 34672
rect 10852 34552 10858 34604
rect 10910 34592 10916 34604
rect 50783 34595 50841 34601
rect 50783 34592 50795 34595
rect 10910 34564 50795 34592
rect 10910 34552 10916 34564
rect 50783 34561 50795 34564
rect 50829 34561 50841 34595
rect 50783 34555 50841 34561
rect 1086 34298 58862 34320
rect 1086 34246 19588 34298
rect 19640 34246 19652 34298
rect 19704 34246 19716 34298
rect 19768 34246 19780 34298
rect 19832 34246 50308 34298
rect 50360 34246 50372 34298
rect 50424 34246 50436 34298
rect 50488 34246 50500 34298
rect 50552 34246 58862 34298
rect 1086 34224 58862 34246
rect 21800 33804 21806 33856
rect 21858 33844 21864 33856
rect 36523 33847 36581 33853
rect 36523 33844 36535 33847
rect 21858 33816 36535 33844
rect 21858 33804 21864 33816
rect 36523 33813 36535 33816
rect 36569 33813 36581 33847
rect 43604 33844 43610 33856
rect 43565 33816 43610 33844
rect 36523 33807 36581 33813
rect 43604 33804 43610 33816
rect 43662 33804 43668 33856
rect 58416 33844 58422 33856
rect 58377 33816 58422 33844
rect 58416 33804 58422 33816
rect 58474 33804 58480 33856
rect 1086 33754 58862 33776
rect 1086 33702 4228 33754
rect 4280 33702 4292 33754
rect 4344 33702 4356 33754
rect 4408 33702 4420 33754
rect 4472 33702 34948 33754
rect 35000 33702 35012 33754
rect 35064 33702 35076 33754
rect 35128 33702 35140 33754
rect 35192 33702 58862 33754
rect 1086 33680 58862 33702
rect 35784 33600 35790 33652
rect 35842 33640 35848 33652
rect 43604 33640 43610 33652
rect 35842 33612 43610 33640
rect 35842 33600 35848 33612
rect 43604 33600 43610 33612
rect 43662 33600 43668 33652
rect 32932 33532 32938 33584
rect 32990 33572 32996 33584
rect 58416 33572 58422 33584
rect 32990 33544 58422 33572
rect 32990 33532 32996 33544
rect 58416 33532 58422 33544
rect 58474 33532 58480 33584
rect 6531 33507 6589 33513
rect 6531 33473 6543 33507
rect 6577 33504 6589 33507
rect 22812 33504 22818 33516
rect 6577 33476 22818 33504
rect 6577 33473 6589 33476
rect 6531 33467 6589 33473
rect 22812 33464 22818 33476
rect 22870 33464 22876 33516
rect 2388 33396 2394 33448
rect 2446 33436 2452 33448
rect 46275 33439 46333 33445
rect 46275 33436 46287 33439
rect 2446 33408 46287 33436
rect 2446 33396 2452 33408
rect 46275 33405 46287 33408
rect 46321 33405 46333 33439
rect 46275 33399 46333 33405
rect 1086 33210 58862 33232
rect 1086 33158 19588 33210
rect 19640 33158 19652 33210
rect 19704 33158 19716 33210
rect 19768 33158 19780 33210
rect 19832 33158 50308 33210
rect 50360 33158 50372 33210
rect 50424 33158 50436 33210
rect 50488 33158 50500 33210
rect 50552 33158 58862 33210
rect 1086 33136 58862 33158
rect 12419 32759 12477 32765
rect 12419 32725 12431 32759
rect 12465 32756 12477 32759
rect 50136 32756 50142 32768
rect 12465 32728 50142 32756
rect 12465 32725 12477 32728
rect 12419 32719 12477 32725
rect 50136 32716 50142 32728
rect 50194 32716 50200 32768
rect 1086 32666 58862 32688
rect 1086 32614 4228 32666
rect 4280 32614 4292 32666
rect 4344 32614 4356 32666
rect 4408 32614 4420 32666
rect 4472 32614 34948 32666
rect 35000 32614 35012 32666
rect 35064 32614 35076 32666
rect 35128 32614 35140 32666
rect 35192 32614 58862 32666
rect 1086 32592 58862 32614
rect 39832 32376 39838 32428
rect 39890 32416 39896 32428
rect 53083 32419 53141 32425
rect 53083 32416 53095 32419
rect 39890 32388 53095 32416
rect 39890 32376 39896 32388
rect 53083 32385 53095 32388
rect 53129 32385 53141 32419
rect 53083 32379 53141 32385
rect 10395 32351 10453 32357
rect 10395 32317 10407 32351
rect 10441 32348 10453 32351
rect 14532 32348 14538 32360
rect 10441 32320 14538 32348
rect 10441 32317 10453 32320
rect 10395 32311 10453 32317
rect 14532 32308 14538 32320
rect 14590 32308 14596 32360
rect 50875 32351 50933 32357
rect 50875 32317 50887 32351
rect 50921 32348 50933 32351
rect 54000 32348 54006 32360
rect 50921 32320 54006 32348
rect 50921 32317 50933 32320
rect 50875 32311 50933 32317
rect 54000 32308 54006 32320
rect 54058 32308 54064 32360
rect 1086 32122 58862 32144
rect 1086 32070 19588 32122
rect 19640 32070 19652 32122
rect 19704 32070 19716 32122
rect 19768 32070 19780 32122
rect 19832 32070 50308 32122
rect 50360 32070 50372 32122
rect 50424 32070 50436 32122
rect 50488 32070 50500 32122
rect 50552 32070 58862 32122
rect 1086 32048 58862 32070
rect 37992 32008 37998 32020
rect 5074 31980 37998 32008
rect 5074 31881 5102 31980
rect 37992 31968 37998 31980
rect 38050 31968 38056 32020
rect 38102 31980 51746 32008
rect 10760 31900 10766 31952
rect 10818 31940 10824 31952
rect 19135 31943 19193 31949
rect 19135 31940 19147 31943
rect 10818 31912 19147 31940
rect 10818 31900 10824 31912
rect 19135 31909 19147 31912
rect 19181 31909 19193 31943
rect 19135 31903 19193 31909
rect 31552 31900 31558 31952
rect 31610 31940 31616 31952
rect 38102 31940 38130 31980
rect 31610 31912 38130 31940
rect 31610 31900 31616 31912
rect 5059 31875 5117 31881
rect 5059 31841 5071 31875
rect 5105 31841 5117 31875
rect 5059 31835 5117 31841
rect 9288 31832 9294 31884
rect 9346 31872 9352 31884
rect 37167 31875 37225 31881
rect 37167 31872 37179 31875
rect 9346 31844 37179 31872
rect 9346 31832 9352 31844
rect 37167 31841 37179 31844
rect 37213 31841 37225 31875
rect 37167 31835 37225 31841
rect 19135 31807 19193 31813
rect 19135 31773 19147 31807
rect 19181 31804 19193 31807
rect 19411 31807 19469 31813
rect 19411 31804 19423 31807
rect 19181 31776 19423 31804
rect 19181 31773 19193 31776
rect 19135 31767 19193 31773
rect 19411 31773 19423 31776
rect 19457 31773 19469 31807
rect 19411 31767 19469 31773
rect 21895 31807 21953 31813
rect 21895 31773 21907 31807
rect 21941 31804 21953 31807
rect 24284 31804 24290 31816
rect 21941 31776 24290 31804
rect 21941 31773 21953 31776
rect 21895 31767 21953 31773
rect 24284 31764 24290 31776
rect 24342 31764 24348 31816
rect 32383 31807 32441 31813
rect 32383 31773 32395 31807
rect 32429 31804 32441 31807
rect 40844 31804 40850 31816
rect 32429 31776 40850 31804
rect 32429 31773 32441 31776
rect 32383 31767 32441 31773
rect 40844 31764 40850 31776
rect 40902 31764 40908 31816
rect 51611 31807 51669 31813
rect 51611 31773 51623 31807
rect 51657 31804 51669 31807
rect 51718 31804 51746 31980
rect 51657 31776 51746 31804
rect 51657 31773 51669 31776
rect 51611 31767 51669 31773
rect 23456 31696 23462 31748
rect 23514 31736 23520 31748
rect 23640 31736 23646 31748
rect 23514 31708 23646 31736
rect 23514 31696 23520 31708
rect 23640 31696 23646 31708
rect 23698 31696 23704 31748
rect 1086 31578 58862 31600
rect 1086 31526 4228 31578
rect 4280 31526 4292 31578
rect 4344 31526 4356 31578
rect 4408 31526 4420 31578
rect 4472 31526 34948 31578
rect 35000 31526 35012 31578
rect 35064 31526 35076 31578
rect 35128 31526 35140 31578
rect 35192 31526 58862 31578
rect 1086 31504 58862 31526
rect 8736 31260 8742 31272
rect 8616 31232 8742 31260
rect 8616 31178 8644 31232
rect 8736 31220 8742 31232
rect 8794 31220 8800 31272
rect 21159 31263 21217 31269
rect 9182 31232 9426 31260
rect 9398 31192 9426 31232
rect 21159 31229 21171 31263
rect 21205 31260 21217 31263
rect 36520 31260 36526 31272
rect 21205 31232 36526 31260
rect 21205 31229 21217 31232
rect 21159 31223 21217 31229
rect 36520 31220 36526 31232
rect 36578 31220 36584 31272
rect 17200 31192 17206 31204
rect 9398 31164 17206 31192
rect 17200 31152 17206 31164
rect 17258 31152 17264 31204
rect 5240 31084 5246 31136
rect 5298 31124 5304 31136
rect 5424 31124 5430 31136
rect 5298 31096 5430 31124
rect 5298 31084 5304 31096
rect 5424 31084 5430 31096
rect 5482 31084 5488 31136
rect 8828 31084 8834 31136
rect 8886 31084 8892 31136
rect 9012 31084 9018 31136
rect 9070 31124 9076 31136
rect 25572 31124 25578 31136
rect 9070 31096 25578 31124
rect 9070 31084 9076 31096
rect 25572 31084 25578 31096
rect 25630 31084 25636 31136
rect 1086 31034 58862 31056
rect 1086 30982 19588 31034
rect 19640 30982 19652 31034
rect 19704 30982 19716 31034
rect 19768 30982 19780 31034
rect 19832 30982 50308 31034
rect 50360 30982 50372 31034
rect 50424 30982 50436 31034
rect 50488 30982 50500 31034
rect 50552 30982 58862 31034
rect 1086 30960 58862 30982
rect 17200 30880 17206 30932
rect 17258 30920 17264 30932
rect 28792 30920 28798 30932
rect 17258 30892 28798 30920
rect 17258 30880 17264 30892
rect 28792 30880 28798 30892
rect 28850 30880 28856 30932
rect 8736 30812 8742 30864
rect 8794 30852 8800 30864
rect 28700 30852 28706 30864
rect 8794 30824 28706 30852
rect 8794 30812 8800 30824
rect 28700 30812 28706 30824
rect 28758 30812 28764 30864
rect 19319 30787 19377 30793
rect 19319 30753 19331 30787
rect 19365 30784 19377 30787
rect 22720 30784 22726 30796
rect 19365 30756 22726 30784
rect 19365 30753 19377 30756
rect 19319 30747 19377 30753
rect 22720 30744 22726 30756
rect 22778 30744 22784 30796
rect 7356 30580 7362 30592
rect 7317 30552 7362 30580
rect 7356 30540 7362 30552
rect 7414 30540 7420 30592
rect 19687 30583 19745 30589
rect 19687 30549 19699 30583
rect 19733 30580 19745 30583
rect 21156 30580 21162 30592
rect 19733 30552 21162 30580
rect 19733 30549 19745 30552
rect 19687 30543 19745 30549
rect 21156 30540 21162 30552
rect 21214 30540 21220 30592
rect 1086 30490 58862 30512
rect 1086 30438 4228 30490
rect 4280 30438 4292 30490
rect 4344 30438 4356 30490
rect 4408 30438 4420 30490
rect 4472 30438 34948 30490
rect 35000 30438 35012 30490
rect 35064 30438 35076 30490
rect 35128 30438 35140 30490
rect 35192 30438 58862 30490
rect 1086 30416 58862 30438
rect 25664 30308 25670 30320
rect 13262 30280 25670 30308
rect 13262 30249 13290 30280
rect 25664 30268 25670 30280
rect 25722 30268 25728 30320
rect 13247 30243 13305 30249
rect 13247 30209 13259 30243
rect 13293 30209 13305 30243
rect 13247 30203 13305 30209
rect 14900 30200 14906 30252
rect 14958 30240 14964 30252
rect 32567 30243 32625 30249
rect 32567 30240 32579 30243
rect 14958 30212 32579 30240
rect 14958 30200 14964 30212
rect 32567 30209 32579 30212
rect 32613 30209 32625 30243
rect 32567 30203 32625 30209
rect 46198 30212 48342 30240
rect 8460 30132 8466 30184
rect 8518 30132 8524 30184
rect 9182 30144 9334 30172
rect 8478 30056 8506 30132
rect 9306 30104 9334 30144
rect 12140 30132 12146 30184
rect 12198 30172 12204 30184
rect 46198 30172 46226 30212
rect 12198 30144 46226 30172
rect 48207 30175 48265 30181
rect 12198 30132 12204 30144
rect 48207 30141 48219 30175
rect 48253 30141 48265 30175
rect 48314 30172 48342 30212
rect 56947 30175 57005 30181
rect 56947 30172 56959 30175
rect 48314 30144 56959 30172
rect 48207 30135 48265 30141
rect 56947 30141 56959 30144
rect 56993 30141 57005 30175
rect 56947 30135 57005 30141
rect 12876 30104 12882 30116
rect 9306 30076 12882 30104
rect 12876 30064 12882 30076
rect 12934 30064 12940 30116
rect 15838 30076 16142 30104
rect 8828 29996 8834 30048
rect 8886 29996 8892 30048
rect 9012 29996 9018 30048
rect 9070 30036 9076 30048
rect 15838 30036 15866 30076
rect 16004 30036 16010 30048
rect 9070 30008 15866 30036
rect 15965 30008 16010 30036
rect 9070 29996 9076 30008
rect 16004 29996 16010 30008
rect 16062 29996 16068 30048
rect 16114 30036 16142 30076
rect 26124 30064 26130 30116
rect 26182 30104 26188 30116
rect 48222 30104 48250 30135
rect 26182 30076 48250 30104
rect 26182 30064 26188 30076
rect 24284 30036 24290 30048
rect 16114 30008 24290 30036
rect 24284 29996 24290 30008
rect 24342 29996 24348 30048
rect 1086 29946 58862 29968
rect 1086 29894 19588 29946
rect 19640 29894 19652 29946
rect 19704 29894 19716 29946
rect 19768 29894 19780 29946
rect 19832 29894 50308 29946
rect 50360 29894 50372 29946
rect 50424 29894 50436 29946
rect 50488 29894 50500 29946
rect 50552 29894 58862 29946
rect 1086 29872 58862 29894
rect 12876 29792 12882 29844
rect 12934 29832 12940 29844
rect 27228 29832 27234 29844
rect 12934 29804 27234 29832
rect 12934 29792 12940 29804
rect 27228 29792 27234 29804
rect 27286 29792 27292 29844
rect 1100 29724 1106 29776
rect 1158 29764 1164 29776
rect 16004 29764 16010 29776
rect 1158 29736 16010 29764
rect 1158 29724 1164 29736
rect 16004 29724 16010 29736
rect 16062 29724 16068 29776
rect 8460 29656 8466 29708
rect 8518 29696 8524 29708
rect 27596 29696 27602 29708
rect 8518 29668 27602 29696
rect 8518 29656 8524 29668
rect 27596 29656 27602 29668
rect 27654 29656 27660 29708
rect 26676 29492 26682 29504
rect 26637 29464 26682 29492
rect 26676 29452 26682 29464
rect 26734 29452 26740 29504
rect 45723 29495 45781 29501
rect 45723 29461 45735 29495
rect 45769 29492 45781 29495
rect 48940 29492 48946 29504
rect 45769 29464 48946 29492
rect 45769 29461 45781 29464
rect 45723 29455 45781 29461
rect 48940 29452 48946 29464
rect 48998 29452 49004 29504
rect 1086 29402 58862 29424
rect 1086 29350 4228 29402
rect 4280 29350 4292 29402
rect 4344 29350 4356 29402
rect 4408 29350 4420 29402
rect 4472 29350 34948 29402
rect 35000 29350 35012 29402
rect 35064 29350 35076 29402
rect 35128 29350 35140 29402
rect 35192 29350 58862 29402
rect 1086 29328 58862 29350
rect 25112 29288 25118 29300
rect 8800 29260 25118 29288
rect 8552 29152 8558 29164
rect 7834 29124 8558 29152
rect 3492 29044 3498 29096
rect 3550 29084 3556 29096
rect 3550 29062 3630 29084
rect 3550 29056 3590 29062
rect 3550 29044 3556 29056
rect 3584 29010 3590 29056
rect 3642 29010 3648 29062
rect 7834 29028 7862 29124
rect 8552 29112 8558 29124
rect 8610 29112 8616 29164
rect 8800 29070 8828 29260
rect 25112 29248 25118 29260
rect 25170 29248 25176 29300
rect 26676 29248 26682 29300
rect 26734 29288 26740 29300
rect 51700 29288 51706 29300
rect 26734 29260 51706 29288
rect 26734 29248 26740 29260
rect 51700 29248 51706 29260
rect 51758 29248 51764 29300
rect 51427 29223 51485 29229
rect 51427 29189 51439 29223
rect 51473 29220 51485 29223
rect 51519 29223 51577 29229
rect 51519 29220 51531 29223
rect 51473 29192 51531 29220
rect 51473 29189 51485 29192
rect 51427 29183 51485 29189
rect 51519 29189 51531 29192
rect 51565 29189 51577 29223
rect 51519 29183 51577 29189
rect 34312 29112 34318 29164
rect 34370 29152 34376 29164
rect 57867 29155 57925 29161
rect 57867 29152 57879 29155
rect 34370 29124 57879 29152
rect 34370 29112 34376 29124
rect 57867 29121 57879 29124
rect 57913 29121 57925 29155
rect 57867 29115 57925 29121
rect 27320 29084 27326 29096
rect 8998 29056 27326 29084
rect 27320 29044 27326 29056
rect 27378 29044 27384 29096
rect 7816 28976 7822 29028
rect 7874 28976 7880 29028
rect 15544 28976 15550 29028
rect 15602 29016 15608 29028
rect 15636 29016 15642 29028
rect 15602 28988 15642 29016
rect 15602 28976 15608 28988
rect 15636 28976 15642 28988
rect 15694 28976 15700 29028
rect 34404 28976 34410 29028
rect 34462 29016 34468 29028
rect 51519 29019 51577 29025
rect 51519 29016 51531 29019
rect 34462 28988 51531 29016
rect 34462 28976 34468 28988
rect 51519 28985 51531 28988
rect 51565 28985 51577 29019
rect 51519 28979 51577 28985
rect 22720 28948 22726 28960
rect 8722 28920 22726 28948
rect 22720 28908 22726 28920
rect 22778 28908 22784 28960
rect 1086 28858 58862 28880
rect 1086 28806 19588 28858
rect 19640 28806 19652 28858
rect 19704 28806 19716 28858
rect 19768 28806 19780 28858
rect 19832 28806 50308 28858
rect 50360 28806 50372 28858
rect 50424 28806 50436 28858
rect 50488 28806 50500 28858
rect 50552 28806 58862 28858
rect 1086 28784 58862 28806
rect 3768 28608 3774 28620
rect 3729 28580 3774 28608
rect 3768 28568 3774 28580
rect 3826 28568 3832 28620
rect 26679 28407 26737 28413
rect 26679 28373 26691 28407
rect 26725 28404 26737 28407
rect 36796 28404 36802 28416
rect 26725 28376 36802 28404
rect 26725 28373 26737 28376
rect 26679 28367 26737 28373
rect 36796 28364 36802 28376
rect 36854 28364 36860 28416
rect 1086 28314 58862 28336
rect 1086 28262 4228 28314
rect 4280 28262 4292 28314
rect 4344 28262 4356 28314
rect 4408 28262 4420 28314
rect 4472 28262 34948 28314
rect 35000 28262 35012 28314
rect 35064 28262 35076 28314
rect 35128 28262 35140 28314
rect 35192 28262 58862 28314
rect 1086 28240 58862 28262
rect 28056 28160 28062 28212
rect 28114 28200 28120 28212
rect 28240 28200 28246 28212
rect 28114 28172 28246 28200
rect 28114 28160 28120 28172
rect 28240 28160 28246 28172
rect 28298 28160 28304 28212
rect 8552 28064 8558 28076
rect 8446 28036 8558 28064
rect 8552 28024 8558 28036
rect 8610 28024 8616 28076
rect 8920 28024 8926 28076
rect 8978 28064 8984 28076
rect 25388 28064 25394 28076
rect 8978 28036 25394 28064
rect 8978 28024 8984 28036
rect 25388 28024 25394 28036
rect 25446 28024 25452 28076
rect 8828 27956 8834 28008
rect 8886 27996 8892 28008
rect 25848 27996 25854 28008
rect 8886 27968 25854 27996
rect 8886 27956 8892 27968
rect 25848 27956 25854 27968
rect 25906 27956 25912 28008
rect 8478 27860 8506 27948
rect 8552 27860 8558 27872
rect 8478 27832 8558 27860
rect 8552 27820 8558 27832
rect 8610 27820 8616 27872
rect 21432 27860 21438 27872
rect 8722 27832 21438 27860
rect 21432 27820 21438 27832
rect 21490 27820 21496 27872
rect 1086 27770 58862 27792
rect 1086 27718 19588 27770
rect 19640 27718 19652 27770
rect 19704 27718 19716 27770
rect 19768 27718 19780 27770
rect 19832 27718 50308 27770
rect 50360 27718 50372 27770
rect 50424 27718 50436 27770
rect 50488 27718 50500 27770
rect 50552 27718 58862 27770
rect 1086 27696 58862 27718
rect 5332 27616 5338 27668
rect 5390 27616 5396 27668
rect 28056 27616 28062 27668
rect 28114 27656 28120 27668
rect 28148 27656 28154 27668
rect 28114 27628 28154 27656
rect 28114 27616 28120 27628
rect 28148 27616 28154 27628
rect 28206 27616 28212 27668
rect 34496 27616 34502 27668
rect 34554 27656 34560 27668
rect 34772 27656 34778 27668
rect 34554 27628 34778 27656
rect 34554 27616 34560 27628
rect 34772 27616 34778 27628
rect 34830 27616 34836 27668
rect 38728 27616 38734 27668
rect 38786 27656 38792 27668
rect 38820 27656 38826 27668
rect 38786 27628 38826 27656
rect 38786 27616 38792 27628
rect 38820 27616 38826 27628
rect 38878 27616 38884 27668
rect 47836 27616 47842 27668
rect 47894 27656 47900 27668
rect 48020 27656 48026 27668
rect 47894 27628 48026 27656
rect 47894 27616 47900 27628
rect 48020 27616 48026 27628
rect 48078 27616 48084 27668
rect 3400 27548 3406 27600
rect 3458 27588 3464 27600
rect 3584 27588 3590 27600
rect 3458 27560 3590 27588
rect 3458 27548 3464 27560
rect 3584 27548 3590 27560
rect 3642 27548 3648 27600
rect 5350 27464 5378 27616
rect 14808 27548 14814 27600
rect 14866 27588 14872 27600
rect 14900 27588 14906 27600
rect 14866 27560 14906 27588
rect 14866 27548 14872 27560
rect 14900 27548 14906 27560
rect 14958 27548 14964 27600
rect 18212 27548 18218 27600
rect 18270 27588 18276 27600
rect 18304 27588 18310 27600
rect 18270 27560 18310 27588
rect 18270 27548 18276 27560
rect 18304 27548 18310 27560
rect 18362 27548 18368 27600
rect 26492 27548 26498 27600
rect 26550 27588 26556 27600
rect 26584 27588 26590 27600
rect 26550 27560 26590 27588
rect 26550 27548 26556 27560
rect 26584 27548 26590 27560
rect 26642 27548 26648 27600
rect 5332 27412 5338 27464
rect 5390 27412 5396 27464
rect 15455 27319 15513 27325
rect 15455 27285 15467 27319
rect 15501 27316 15513 27319
rect 17200 27316 17206 27328
rect 15501 27288 17206 27316
rect 15501 27285 15513 27288
rect 15455 27279 15513 27285
rect 17200 27276 17206 27288
rect 17258 27276 17264 27328
rect 1086 27226 58862 27248
rect 1086 27174 4228 27226
rect 4280 27174 4292 27226
rect 4344 27174 4356 27226
rect 4408 27174 4420 27226
rect 4472 27174 34948 27226
rect 35000 27174 35012 27226
rect 35064 27174 35076 27226
rect 35128 27174 35140 27226
rect 35192 27174 58862 27226
rect 1086 27152 58862 27174
rect 7632 26936 7638 26988
rect 7690 26976 7696 26988
rect 7908 26976 7914 26988
rect 7690 26948 7914 26976
rect 7690 26936 7696 26948
rect 7908 26936 7914 26948
rect 7966 26936 7972 26988
rect 8552 26976 8558 26988
rect 8446 26948 8558 26976
rect 8552 26936 8558 26948
rect 8610 26936 8616 26988
rect 8828 26936 8834 26988
rect 8886 26976 8892 26988
rect 23640 26976 23646 26988
rect 8886 26948 23646 26976
rect 8886 26936 8892 26948
rect 23640 26936 23646 26948
rect 23698 26936 23704 26988
rect 53359 26979 53417 26985
rect 53359 26976 53371 26979
rect 51810 26948 53371 26976
rect 8460 26908 8466 26920
rect 8262 26880 8466 26908
rect 8460 26868 8466 26880
rect 8518 26868 8524 26920
rect 8920 26868 8926 26920
rect 8978 26908 8984 26920
rect 24376 26908 24382 26920
rect 8978 26880 24382 26908
rect 8978 26868 8984 26880
rect 24376 26868 24382 26880
rect 24434 26868 24440 26920
rect 46732 26868 46738 26920
rect 46790 26908 46796 26920
rect 51810 26908 51838 26948
rect 53359 26945 53371 26948
rect 53405 26945 53417 26979
rect 53359 26939 53417 26945
rect 46790 26880 51838 26908
rect 51887 26911 51945 26917
rect 46790 26868 46796 26880
rect 51887 26877 51899 26911
rect 51933 26908 51945 26911
rect 55840 26908 55846 26920
rect 51933 26880 55846 26908
rect 51933 26877 51945 26880
rect 51887 26871 51945 26877
rect 55840 26868 55846 26880
rect 55898 26868 55904 26920
rect 21524 26772 21530 26784
rect 8722 26744 21530 26772
rect 21524 26732 21530 26744
rect 21582 26732 21588 26784
rect 1086 26682 58862 26704
rect 1086 26630 19588 26682
rect 19640 26630 19652 26682
rect 19704 26630 19716 26682
rect 19768 26630 19780 26682
rect 19832 26630 50308 26682
rect 50360 26630 50372 26682
rect 50424 26630 50436 26682
rect 50488 26630 50500 26682
rect 50552 26630 58862 26682
rect 1086 26608 58862 26630
rect 4231 26435 4289 26441
rect 4231 26401 4243 26435
rect 4277 26432 4289 26435
rect 5516 26432 5522 26444
rect 4277 26404 5522 26432
rect 4277 26401 4289 26404
rect 4231 26395 4289 26401
rect 5516 26392 5522 26404
rect 5574 26392 5580 26444
rect 36980 26392 36986 26444
rect 37038 26432 37044 26444
rect 38547 26435 38605 26441
rect 38547 26432 38559 26435
rect 37038 26404 38559 26432
rect 37038 26392 37044 26404
rect 38547 26401 38559 26404
rect 38593 26401 38605 26435
rect 38547 26395 38605 26401
rect 40203 26435 40261 26441
rect 40203 26401 40215 26435
rect 40249 26432 40261 26435
rect 50044 26432 50050 26444
rect 40249 26404 50050 26432
rect 40249 26401 40261 26404
rect 40203 26395 40261 26401
rect 50044 26392 50050 26404
rect 50102 26392 50108 26444
rect 20604 26324 20610 26376
rect 20662 26364 20668 26376
rect 57131 26367 57189 26373
rect 57131 26364 57143 26367
rect 20662 26336 57143 26364
rect 20662 26324 20668 26336
rect 57131 26333 57143 26336
rect 57177 26333 57189 26367
rect 57131 26327 57189 26333
rect 6620 26256 6626 26308
rect 6678 26296 6684 26308
rect 50323 26299 50381 26305
rect 50323 26296 50335 26299
rect 6678 26268 50335 26296
rect 6678 26256 6684 26268
rect 50323 26265 50335 26268
rect 50369 26265 50381 26299
rect 50323 26259 50381 26265
rect 25664 26188 25670 26240
rect 25722 26228 25728 26240
rect 25756 26228 25762 26240
rect 25722 26200 25762 26228
rect 25722 26188 25728 26200
rect 25756 26188 25762 26200
rect 25814 26188 25820 26240
rect 39740 26188 39746 26240
rect 39798 26228 39804 26240
rect 39924 26228 39930 26240
rect 39798 26200 39930 26228
rect 39798 26188 39804 26200
rect 39924 26188 39930 26200
rect 39982 26188 39988 26240
rect 1086 26138 58862 26160
rect 1086 26086 4228 26138
rect 4280 26086 4292 26138
rect 4344 26086 4356 26138
rect 4408 26086 4420 26138
rect 4472 26086 34948 26138
rect 35000 26086 35012 26138
rect 35064 26086 35076 26138
rect 35128 26086 35140 26138
rect 35192 26086 58862 26138
rect 1086 26064 58862 26086
rect 8552 26024 8558 26036
rect 8248 25996 8558 26024
rect 8248 25908 8276 25996
rect 8552 25984 8558 25996
rect 8610 25984 8616 26036
rect 11404 26024 11410 26036
rect 11365 25996 11410 26024
rect 11404 25984 11410 25996
rect 11462 25984 11468 26036
rect 8552 25888 8558 25900
rect 8446 25860 8558 25888
rect 8552 25848 8558 25860
rect 8610 25848 8616 25900
rect 7724 25780 7730 25832
rect 7782 25820 7788 25832
rect 7911 25823 7969 25829
rect 7911 25820 7923 25823
rect 7782 25792 7923 25820
rect 7782 25780 7788 25792
rect 7911 25789 7923 25792
rect 7957 25789 7969 25823
rect 7911 25783 7969 25789
rect 35692 25780 35698 25832
rect 35750 25820 35756 25832
rect 42779 25823 42837 25829
rect 42779 25820 42791 25823
rect 35750 25792 42791 25820
rect 35750 25780 35756 25792
rect 42779 25789 42791 25792
rect 42825 25789 42837 25823
rect 42779 25783 42837 25789
rect 8920 25712 8926 25764
rect 8978 25752 8984 25764
rect 22904 25752 22910 25764
rect 8978 25724 22910 25752
rect 8978 25712 8984 25724
rect 22904 25712 22910 25724
rect 22962 25712 22968 25764
rect 8690 25644 8696 25696
rect 8748 25644 8754 25696
rect 8828 25644 8834 25696
rect 8886 25684 8892 25696
rect 22536 25684 22542 25696
rect 8886 25656 22542 25684
rect 8886 25644 8892 25656
rect 22536 25644 22542 25656
rect 22594 25644 22600 25696
rect 1086 25594 58862 25616
rect 1086 25542 19588 25594
rect 19640 25542 19652 25594
rect 19704 25542 19716 25594
rect 19768 25542 19780 25594
rect 19832 25542 50308 25594
rect 50360 25542 50372 25594
rect 50424 25542 50436 25594
rect 50488 25542 50500 25594
rect 50552 25542 58862 25594
rect 1086 25520 58862 25542
rect 8690 25440 8696 25492
rect 8748 25480 8754 25492
rect 20052 25480 20058 25492
rect 8748 25452 20058 25480
rect 8748 25440 8754 25452
rect 20052 25440 20058 25452
rect 20110 25440 20116 25492
rect 7724 25372 7730 25424
rect 7782 25412 7788 25424
rect 32564 25412 32570 25424
rect 7782 25384 32570 25412
rect 7782 25372 7788 25384
rect 32564 25372 32570 25384
rect 32622 25372 32628 25424
rect 8276 25100 8282 25152
rect 8334 25140 8340 25152
rect 12416 25140 12422 25152
rect 8334 25112 12422 25140
rect 8334 25100 8340 25112
rect 12416 25100 12422 25112
rect 12474 25100 12480 25152
rect 1086 25050 58862 25072
rect 1086 24998 4228 25050
rect 4280 24998 4292 25050
rect 4344 24998 4356 25050
rect 4408 24998 4420 25050
rect 4472 24998 34948 25050
rect 35000 24998 35012 25050
rect 35064 24998 35076 25050
rect 35128 24998 35140 25050
rect 35192 24998 58862 25050
rect 1086 24976 58862 24998
rect 8276 24896 8282 24948
rect 8334 24896 8340 24948
rect 12416 24896 12422 24948
rect 12474 24936 12480 24948
rect 19960 24936 19966 24948
rect 12474 24908 19966 24936
rect 12474 24896 12480 24908
rect 19960 24896 19966 24908
rect 20018 24896 20024 24948
rect 8604 24812 8656 24818
rect 1379 24803 1437 24809
rect 1379 24769 1391 24803
rect 1425 24800 1437 24803
rect 1560 24800 1566 24812
rect 1425 24772 1566 24800
rect 1425 24769 1437 24772
rect 1379 24763 1437 24769
rect 1560 24760 1566 24772
rect 1618 24760 1624 24812
rect 8248 24596 8276 24786
rect 8920 24760 8926 24812
rect 8978 24800 8984 24812
rect 8978 24772 10162 24800
rect 8978 24760 8984 24772
rect 8604 24754 8656 24760
rect 10134 24732 10162 24772
rect 10208 24760 10214 24812
rect 10266 24800 10272 24812
rect 21064 24800 21070 24812
rect 10266 24772 21070 24800
rect 10266 24760 10272 24772
rect 21064 24760 21070 24772
rect 21122 24760 21128 24812
rect 22076 24732 22082 24744
rect 8432 24676 8460 24718
rect 8814 24704 10070 24732
rect 10134 24704 22082 24732
rect 8432 24636 8466 24676
rect 8460 24624 8466 24636
rect 8518 24624 8524 24676
rect 10042 24664 10070 24704
rect 22076 24692 22082 24704
rect 22134 24692 22140 24744
rect 21708 24664 21714 24676
rect 10042 24636 21714 24664
rect 21708 24624 21714 24636
rect 21766 24624 21772 24676
rect 10208 24596 10214 24608
rect 8248 24568 10214 24596
rect 10208 24556 10214 24568
rect 10266 24556 10272 24608
rect 1086 24506 58862 24528
rect 1086 24454 19588 24506
rect 19640 24454 19652 24506
rect 19704 24454 19716 24506
rect 19768 24454 19780 24506
rect 19832 24454 50308 24506
rect 50360 24454 50372 24506
rect 50424 24454 50436 24506
rect 50488 24454 50500 24506
rect 50552 24454 58862 24506
rect 1086 24432 58862 24454
rect 8460 24352 8466 24404
rect 8518 24392 8524 24404
rect 20788 24392 20794 24404
rect 8518 24364 20794 24392
rect 8518 24352 8524 24364
rect 20788 24352 20794 24364
rect 20846 24352 20852 24404
rect 9840 24256 9846 24268
rect 9801 24228 9846 24256
rect 9840 24216 9846 24228
rect 9898 24216 9904 24268
rect 51056 24148 51062 24200
rect 51114 24148 51120 24200
rect 3768 24080 3774 24132
rect 3826 24120 3832 24132
rect 34220 24120 34226 24132
rect 3826 24092 34226 24120
rect 3826 24080 3832 24092
rect 34220 24080 34226 24092
rect 34278 24080 34284 24132
rect 51074 24064 51102 24148
rect 16464 24012 16470 24064
rect 16522 24052 16528 24064
rect 19687 24055 19745 24061
rect 19687 24052 19699 24055
rect 16522 24024 19699 24052
rect 16522 24012 16528 24024
rect 19687 24021 19699 24024
rect 19733 24021 19745 24055
rect 19687 24015 19745 24021
rect 31552 24012 31558 24064
rect 31610 24052 31616 24064
rect 49219 24055 49277 24061
rect 49219 24052 49231 24055
rect 31610 24024 49231 24052
rect 31610 24012 31616 24024
rect 49219 24021 49231 24024
rect 49265 24021 49277 24055
rect 49219 24015 49277 24021
rect 51056 24012 51062 24064
rect 51114 24012 51120 24064
rect 1086 23962 58862 23984
rect 1086 23910 4228 23962
rect 4280 23910 4292 23962
rect 4344 23910 4356 23962
rect 4408 23910 4420 23962
rect 4472 23910 34948 23962
rect 35000 23910 35012 23962
rect 35064 23910 35076 23962
rect 35128 23910 35140 23962
rect 35192 23910 58862 23962
rect 1086 23888 58862 23910
rect 8644 23808 8650 23860
rect 8702 23808 8708 23860
rect 8828 23808 8834 23860
rect 8886 23848 8892 23860
rect 18580 23848 18586 23860
rect 8886 23820 18586 23848
rect 8886 23808 8892 23820
rect 18580 23808 18586 23820
rect 18638 23808 18644 23860
rect 34220 23808 34226 23860
rect 34278 23848 34284 23860
rect 43515 23851 43573 23857
rect 43515 23848 43527 23851
rect 34278 23820 43527 23848
rect 34278 23808 34284 23820
rect 43515 23817 43527 23820
rect 43561 23817 43573 23851
rect 43515 23811 43573 23817
rect 8598 23706 8604 23758
rect 8656 23706 8662 23758
rect 9472 23740 9478 23792
rect 9530 23780 9536 23792
rect 12143 23783 12201 23789
rect 12143 23780 12155 23783
rect 9530 23752 12155 23780
rect 9530 23740 9536 23752
rect 12143 23749 12155 23752
rect 12189 23749 12201 23783
rect 57499 23783 57557 23789
rect 57499 23780 57511 23783
rect 12143 23743 12201 23749
rect 46198 23752 57511 23780
rect 8736 23672 8742 23724
rect 8794 23712 8800 23724
rect 20420 23712 20426 23724
rect 8794 23684 20426 23712
rect 8794 23672 8800 23684
rect 20420 23672 20426 23684
rect 20478 23672 20484 23724
rect 8460 23644 8466 23656
rect 8446 23616 8466 23644
rect 8460 23604 8466 23616
rect 8518 23604 8524 23656
rect 8828 23604 8834 23656
rect 8886 23644 8892 23656
rect 19868 23644 19874 23656
rect 8886 23616 19874 23644
rect 8886 23604 8892 23616
rect 19868 23604 19874 23616
rect 19926 23604 19932 23656
rect 46198 23644 46226 23752
rect 57499 23749 57511 23752
rect 57545 23749 57557 23783
rect 57499 23743 57557 23749
rect 26878 23616 46226 23644
rect 49587 23647 49645 23653
rect 8248 23508 8276 23596
rect 12143 23579 12201 23585
rect 12143 23545 12155 23579
rect 12189 23576 12201 23579
rect 12189 23548 20374 23576
rect 12189 23545 12201 23548
rect 12143 23539 12201 23545
rect 8460 23508 8466 23520
rect 8248 23480 8466 23508
rect 8460 23468 8466 23480
rect 8518 23468 8524 23520
rect 11772 23468 11778 23520
rect 11830 23508 11836 23520
rect 20236 23508 20242 23520
rect 11830 23480 20242 23508
rect 11830 23468 11836 23480
rect 20236 23468 20242 23480
rect 20294 23468 20300 23520
rect 20346 23508 20374 23548
rect 26878 23508 26906 23616
rect 49587 23613 49599 23647
rect 49633 23613 49645 23647
rect 49587 23607 49645 23613
rect 30264 23536 30270 23588
rect 30322 23576 30328 23588
rect 49602 23576 49630 23607
rect 30322 23548 49630 23576
rect 30322 23536 30328 23548
rect 20346 23480 26906 23508
rect 1086 23418 58862 23440
rect 1086 23366 19588 23418
rect 19640 23366 19652 23418
rect 19704 23366 19716 23418
rect 19768 23366 19780 23418
rect 19832 23366 50308 23418
rect 50360 23366 50372 23418
rect 50424 23366 50436 23418
rect 50488 23366 50500 23418
rect 50552 23366 58862 23418
rect 1086 23344 58862 23366
rect 6899 22967 6957 22973
rect 6899 22933 6911 22967
rect 6945 22964 6957 22967
rect 9656 22964 9662 22976
rect 6945 22936 9662 22964
rect 6945 22933 6957 22936
rect 6899 22927 6957 22933
rect 9656 22924 9662 22936
rect 9714 22924 9720 22976
rect 20604 22924 20610 22976
rect 20662 22964 20668 22976
rect 21251 22967 21309 22973
rect 21251 22964 21263 22967
rect 20662 22936 21263 22964
rect 20662 22924 20668 22936
rect 21251 22933 21263 22936
rect 21297 22933 21309 22967
rect 21251 22927 21309 22933
rect 1086 22874 58862 22896
rect 1086 22822 4228 22874
rect 4280 22822 4292 22874
rect 4344 22822 4356 22874
rect 4408 22822 4420 22874
rect 4472 22822 34948 22874
rect 35000 22822 35012 22874
rect 35064 22822 35076 22874
rect 35128 22822 35140 22874
rect 35192 22822 58862 22874
rect 1086 22800 58862 22822
rect 9107 22763 9165 22769
rect 9107 22760 9119 22763
rect 8800 22732 9119 22760
rect 8800 22610 8828 22732
rect 9107 22729 9119 22732
rect 9153 22729 9165 22763
rect 18672 22760 18678 22772
rect 9274 22732 18678 22760
rect 9107 22723 9165 22729
rect 18672 22720 18678 22732
rect 18730 22720 18736 22772
rect 18028 22624 18034 22636
rect 8998 22596 9058 22624
rect 9182 22596 18034 22624
rect 9030 22420 9058 22596
rect 18028 22584 18034 22596
rect 18086 22584 18092 22636
rect 9107 22559 9165 22565
rect 9107 22525 9119 22559
rect 9153 22556 9165 22559
rect 18764 22556 18770 22568
rect 9153 22528 18770 22556
rect 9153 22525 9165 22528
rect 9107 22519 9165 22525
rect 18764 22516 18770 22528
rect 18822 22516 18828 22568
rect 41488 22556 41494 22568
rect 41449 22528 41494 22556
rect 41488 22516 41494 22528
rect 41546 22516 41552 22568
rect 18120 22420 18126 22432
rect 9030 22392 18126 22420
rect 18120 22380 18126 22392
rect 18178 22380 18184 22432
rect 1086 22330 58862 22352
rect 1086 22278 19588 22330
rect 19640 22278 19652 22330
rect 19704 22278 19716 22330
rect 19768 22278 19780 22330
rect 19832 22278 50308 22330
rect 50360 22278 50372 22330
rect 50424 22278 50436 22330
rect 50488 22278 50500 22330
rect 50552 22278 58862 22330
rect 1086 22256 58862 22278
rect 9656 22176 9662 22228
rect 9714 22216 9720 22228
rect 28424 22216 28430 22228
rect 9714 22188 28430 22216
rect 9714 22176 9720 22188
rect 28424 22176 28430 22188
rect 28482 22176 28488 22228
rect 34407 22083 34465 22089
rect 34407 22049 34419 22083
rect 34453 22080 34465 22083
rect 35416 22080 35422 22092
rect 34453 22052 35422 22080
rect 34453 22049 34465 22052
rect 34407 22043 34465 22049
rect 35416 22040 35422 22052
rect 35474 22040 35480 22092
rect 9380 21836 9386 21888
rect 9438 21876 9444 21888
rect 22539 21879 22597 21885
rect 22539 21876 22551 21879
rect 9438 21848 22551 21876
rect 9438 21836 9444 21848
rect 22539 21845 22551 21848
rect 22585 21845 22597 21879
rect 22539 21839 22597 21845
rect 1086 21786 58862 21808
rect 1086 21734 4228 21786
rect 4280 21734 4292 21786
rect 4344 21734 4356 21786
rect 4408 21734 4420 21786
rect 4472 21734 34948 21786
rect 35000 21734 35012 21786
rect 35064 21734 35076 21786
rect 35128 21734 35140 21786
rect 35192 21734 58862 21786
rect 1086 21712 58862 21734
rect 8555 21675 8613 21681
rect 8555 21672 8567 21675
rect 8248 21644 8567 21672
rect 8248 21556 8276 21644
rect 8555 21641 8567 21644
rect 8601 21641 8613 21675
rect 8555 21635 8613 21641
rect 17292 21536 17298 21548
rect 8446 21508 17298 21536
rect 17292 21496 17298 21508
rect 17350 21496 17356 21548
rect 8555 21471 8613 21477
rect 8555 21437 8567 21471
rect 8601 21468 8613 21471
rect 16924 21468 16930 21480
rect 8601 21440 16930 21468
rect 8601 21437 8613 21440
rect 8555 21431 8613 21437
rect 16924 21428 16930 21440
rect 16982 21428 16988 21480
rect 8460 21292 8466 21344
rect 8518 21292 8524 21344
rect 8644 21292 8650 21344
rect 8702 21332 8708 21344
rect 17384 21332 17390 21344
rect 8702 21304 17390 21332
rect 8702 21292 8708 21304
rect 17384 21292 17390 21304
rect 17442 21292 17448 21344
rect 1086 21242 58862 21264
rect 1086 21190 19588 21242
rect 19640 21190 19652 21242
rect 19704 21190 19716 21242
rect 19768 21190 19780 21242
rect 19832 21190 50308 21242
rect 50360 21190 50372 21242
rect 50424 21190 50436 21242
rect 50488 21190 50500 21242
rect 50552 21190 58862 21242
rect 1086 21168 58862 21190
rect 24379 20995 24437 21001
rect 24379 20961 24391 20995
rect 24425 20992 24437 20995
rect 28332 20992 28338 21004
rect 24425 20964 28338 20992
rect 24425 20961 24437 20964
rect 24379 20955 24437 20961
rect 28332 20952 28338 20964
rect 28390 20952 28396 21004
rect 7724 20884 7730 20936
rect 7782 20924 7788 20936
rect 52071 20927 52129 20933
rect 52071 20924 52083 20927
rect 7782 20896 52083 20924
rect 7782 20884 7788 20896
rect 52071 20893 52083 20896
rect 52117 20893 52129 20927
rect 52071 20887 52129 20893
rect 31555 20859 31613 20865
rect 31555 20825 31567 20859
rect 31601 20856 31613 20859
rect 43604 20856 43610 20868
rect 31601 20828 43610 20856
rect 31601 20825 31613 20828
rect 31555 20819 31613 20825
rect 43604 20816 43610 20828
rect 43662 20816 43668 20868
rect 1086 20698 58862 20720
rect 1086 20646 4228 20698
rect 4280 20646 4292 20698
rect 4344 20646 4356 20698
rect 4408 20646 4420 20698
rect 4472 20646 34948 20698
rect 35000 20646 35012 20698
rect 35064 20646 35076 20698
rect 35128 20646 35140 20698
rect 35192 20646 58862 20698
rect 1086 20624 58862 20646
rect 4044 20584 4050 20596
rect 4005 20556 4050 20584
rect 4044 20544 4050 20556
rect 4102 20544 4108 20596
rect 8460 20544 8466 20596
rect 8518 20544 8524 20596
rect 8644 20544 8650 20596
rect 8702 20584 8708 20596
rect 16832 20584 16838 20596
rect 8702 20556 16838 20584
rect 8702 20544 8708 20556
rect 16832 20544 16838 20556
rect 16890 20544 16896 20596
rect 31570 20488 31782 20516
rect 18491 20451 18549 20457
rect 18491 20417 18503 20451
rect 18537 20448 18549 20451
rect 31570 20448 31598 20488
rect 18537 20420 31598 20448
rect 31754 20448 31782 20488
rect 51792 20448 51798 20460
rect 31754 20420 51798 20448
rect 18537 20417 18549 20420
rect 18491 20411 18549 20417
rect 51792 20408 51798 20420
rect 51850 20408 51856 20460
rect 15544 20380 15550 20392
rect 8630 20352 15550 20380
rect 15544 20340 15550 20352
rect 15602 20340 15608 20392
rect 28608 20380 28614 20392
rect 28569 20352 28614 20380
rect 28608 20340 28614 20352
rect 28666 20340 28672 20392
rect 45815 20383 45873 20389
rect 45815 20349 45827 20383
rect 45861 20349 45873 20383
rect 45815 20343 45873 20349
rect 8248 20256 8276 20332
rect 8248 20216 8282 20256
rect 8276 20204 8282 20216
rect 8334 20204 8340 20256
rect 8432 20244 8460 20332
rect 15820 20312 15826 20324
rect 11330 20284 15826 20312
rect 11330 20244 11358 20284
rect 15820 20272 15826 20284
rect 15878 20272 15884 20324
rect 38360 20272 38366 20324
rect 38418 20312 38424 20324
rect 45830 20312 45858 20343
rect 38418 20284 45858 20312
rect 38418 20272 38424 20284
rect 8432 20216 11358 20244
rect 11404 20204 11410 20256
rect 11462 20244 11468 20256
rect 14624 20244 14630 20256
rect 11462 20216 14630 20244
rect 11462 20204 11468 20216
rect 14624 20204 14630 20216
rect 14682 20204 14688 20256
rect 1086 20154 58862 20176
rect 1086 20102 19588 20154
rect 19640 20102 19652 20154
rect 19704 20102 19716 20154
rect 19768 20102 19780 20154
rect 19832 20102 50308 20154
rect 50360 20102 50372 20154
rect 50424 20102 50436 20154
rect 50488 20102 50500 20154
rect 50552 20102 58862 20154
rect 1086 20080 58862 20102
rect 8276 20000 8282 20052
rect 8334 20040 8340 20052
rect 11404 20040 11410 20052
rect 8334 20012 11410 20040
rect 8334 20000 8340 20012
rect 11404 20000 11410 20012
rect 11462 20000 11468 20052
rect 28608 20040 28614 20052
rect 12250 20012 28614 20040
rect 5148 19932 5154 19984
rect 5206 19972 5212 19984
rect 12250 19972 12278 20012
rect 28608 20000 28614 20012
rect 28666 20000 28672 20052
rect 39556 20040 39562 20052
rect 39517 20012 39562 20040
rect 39556 20000 39562 20012
rect 39614 20000 39620 20052
rect 5206 19944 12278 19972
rect 5206 19932 5212 19944
rect 49584 19904 49590 19916
rect 49545 19876 49590 19904
rect 49584 19864 49590 19876
rect 49642 19864 49648 19916
rect 8460 19660 8466 19712
rect 8518 19700 8524 19712
rect 15912 19700 15918 19712
rect 8518 19672 15918 19700
rect 8518 19660 8524 19672
rect 15912 19660 15918 19672
rect 15970 19660 15976 19712
rect 16372 19660 16378 19712
rect 16430 19700 16436 19712
rect 58143 19703 58201 19709
rect 58143 19700 58155 19703
rect 16430 19672 58155 19700
rect 16430 19660 16436 19672
rect 58143 19669 58155 19672
rect 58189 19669 58201 19703
rect 58143 19663 58201 19669
rect 1086 19610 58862 19632
rect 1086 19558 4228 19610
rect 4280 19558 4292 19610
rect 4344 19558 4356 19610
rect 4408 19558 4420 19610
rect 4472 19558 34948 19610
rect 35000 19558 35012 19610
rect 35064 19558 35076 19610
rect 35128 19558 35140 19610
rect 35192 19558 58862 19610
rect 1086 19536 58862 19558
rect 8460 19456 8466 19508
rect 8518 19456 8524 19508
rect 34772 19428 34778 19440
rect 34606 19400 34778 19428
rect 34606 19372 34634 19400
rect 34772 19388 34778 19400
rect 34830 19388 34836 19440
rect 9843 19363 9901 19369
rect 7448 19252 7454 19304
rect 7506 19292 7512 19304
rect 7816 19292 7822 19338
rect 7506 19286 7822 19292
rect 7874 19286 7880 19338
rect 9843 19329 9855 19363
rect 9889 19360 9901 19363
rect 21340 19360 21346 19372
rect 9889 19332 21346 19360
rect 9889 19329 9901 19332
rect 9843 19323 9901 19329
rect 21340 19320 21346 19332
rect 21398 19320 21404 19372
rect 29252 19320 29258 19372
rect 29310 19360 29316 19372
rect 29344 19360 29350 19372
rect 29310 19332 29350 19360
rect 29310 19320 29316 19332
rect 29344 19320 29350 19332
rect 29402 19320 29408 19372
rect 29439 19363 29497 19369
rect 29439 19329 29451 19363
rect 29485 19360 29497 19363
rect 32656 19360 32662 19372
rect 29485 19332 32662 19360
rect 29485 19329 29497 19332
rect 29439 19323 29497 19329
rect 32656 19320 32662 19332
rect 32714 19320 32720 19372
rect 34588 19320 34594 19372
rect 34646 19320 34652 19372
rect 7506 19264 7862 19286
rect 7506 19252 7512 19264
rect 8000 19252 8006 19304
rect 8058 19292 8064 19304
rect 13152 19292 13158 19304
rect 8058 19264 8262 19292
rect 8058 19252 8064 19264
rect 8414 19218 8420 19270
rect 8472 19218 8478 19270
rect 13113 19264 13158 19292
rect 13152 19252 13158 19264
rect 13210 19252 13216 19304
rect 20972 19252 20978 19304
rect 21030 19292 21036 19304
rect 21064 19292 21070 19304
rect 21030 19264 21070 19292
rect 21030 19252 21036 19264
rect 21064 19252 21070 19264
rect 21122 19252 21128 19304
rect 22904 19252 22910 19304
rect 22962 19292 22968 19304
rect 23088 19292 23094 19304
rect 22962 19264 23094 19292
rect 22962 19252 22968 19264
rect 23088 19252 23094 19264
rect 23146 19252 23152 19304
rect 23640 19252 23646 19304
rect 23698 19292 23704 19304
rect 23916 19292 23922 19304
rect 23698 19264 23922 19292
rect 23698 19252 23704 19264
rect 23916 19252 23922 19264
rect 23974 19252 23980 19304
rect 36888 19252 36894 19304
rect 36946 19292 36952 19304
rect 37072 19292 37078 19304
rect 36946 19264 37078 19292
rect 36946 19252 36952 19264
rect 37072 19252 37078 19264
rect 37130 19252 37136 19304
rect 48388 19252 48394 19304
rect 48446 19252 48452 19304
rect 52068 19252 52074 19304
rect 52126 19292 52132 19304
rect 56668 19292 56674 19304
rect 52126 19264 56674 19292
rect 52126 19252 52132 19264
rect 56668 19252 56674 19264
rect 56726 19252 56732 19304
rect 48406 19168 48434 19252
rect 8920 19116 8926 19168
rect 8978 19156 8984 19168
rect 13152 19156 13158 19168
rect 8978 19128 13158 19156
rect 8978 19116 8984 19128
rect 13152 19116 13158 19128
rect 13210 19116 13216 19168
rect 48388 19116 48394 19168
rect 48446 19116 48452 19168
rect 1086 19066 58862 19088
rect 1086 19014 19588 19066
rect 19640 19014 19652 19066
rect 19704 19014 19716 19066
rect 19768 19014 19780 19066
rect 19832 19014 50308 19066
rect 50360 19014 50372 19066
rect 50424 19014 50436 19066
rect 50488 19014 50500 19066
rect 50552 19014 58862 19066
rect 1086 18992 58862 19014
rect 8460 18912 8466 18964
rect 8518 18952 8524 18964
rect 13336 18952 13342 18964
rect 8518 18924 13342 18952
rect 8518 18912 8524 18924
rect 13336 18912 13342 18924
rect 13394 18912 13400 18964
rect 7632 18640 7638 18692
rect 7690 18680 7696 18692
rect 26768 18680 26774 18692
rect 7690 18652 26774 18680
rect 7690 18640 7696 18652
rect 26768 18640 26774 18652
rect 26826 18640 26832 18692
rect 8644 18572 8650 18624
rect 8702 18612 8708 18624
rect 12784 18612 12790 18624
rect 8702 18584 12790 18612
rect 8702 18572 8708 18584
rect 12784 18572 12790 18584
rect 12842 18572 12848 18624
rect 17295 18615 17353 18621
rect 17295 18581 17307 18615
rect 17341 18612 17353 18615
rect 28332 18612 28338 18624
rect 17341 18584 28338 18612
rect 17341 18581 17353 18584
rect 17295 18575 17353 18581
rect 28332 18572 28338 18584
rect 28390 18572 28396 18624
rect 1086 18522 58862 18544
rect 1086 18470 4228 18522
rect 4280 18470 4292 18522
rect 4344 18470 4356 18522
rect 4408 18470 4420 18522
rect 4472 18470 34948 18522
rect 35000 18470 35012 18522
rect 35064 18470 35076 18522
rect 35128 18470 35140 18522
rect 35192 18470 58862 18522
rect 1086 18448 58862 18470
rect 8828 18368 8834 18420
rect 8886 18368 8892 18420
rect 9012 18368 9018 18420
rect 9070 18408 9076 18420
rect 14164 18408 14170 18420
rect 9070 18380 14170 18408
rect 9070 18368 9076 18380
rect 14164 18368 14170 18380
rect 14222 18368 14228 18420
rect 8644 18272 8650 18284
rect 8446 18244 8650 18272
rect 8644 18232 8650 18244
rect 8702 18232 8708 18284
rect 8754 18244 8814 18272
rect 8754 18213 8782 18244
rect 26768 18232 26774 18284
rect 26826 18272 26832 18284
rect 32199 18275 32257 18281
rect 32199 18272 32211 18275
rect 26826 18244 32211 18272
rect 26826 18232 26832 18244
rect 32199 18241 32211 18244
rect 32245 18241 32257 18275
rect 32199 18235 32257 18241
rect 8739 18207 8797 18213
rect 8739 18173 8751 18207
rect 8785 18173 8797 18207
rect 12600 18204 12606 18216
rect 8998 18176 12606 18204
rect 8739 18167 8797 18173
rect 12600 18164 12606 18176
rect 12658 18164 12664 18216
rect 23180 18164 23186 18216
rect 23238 18204 23244 18216
rect 52807 18207 52865 18213
rect 52807 18204 52819 18207
rect 23238 18176 52819 18204
rect 23238 18164 23244 18176
rect 52807 18173 52819 18176
rect 52853 18173 52865 18207
rect 52807 18167 52865 18173
rect 9015 18071 9073 18077
rect 9015 18037 9027 18071
rect 9061 18068 9073 18071
rect 12876 18068 12882 18080
rect 9061 18040 12882 18068
rect 9061 18037 9073 18040
rect 9015 18031 9073 18037
rect 12876 18028 12882 18040
rect 12934 18028 12940 18080
rect 23456 18028 23462 18080
rect 23514 18068 23520 18080
rect 23548 18068 23554 18080
rect 23514 18040 23554 18068
rect 23514 18028 23520 18040
rect 23548 18028 23554 18040
rect 23606 18028 23612 18080
rect 1086 17978 58862 18000
rect 1086 17926 19588 17978
rect 19640 17926 19652 17978
rect 19704 17926 19716 17978
rect 19768 17926 19780 17978
rect 19832 17926 50308 17978
rect 50360 17926 50372 17978
rect 50424 17926 50436 17978
rect 50488 17926 50500 17978
rect 50552 17926 58862 17978
rect 1086 17904 58862 17926
rect 8828 17620 8834 17672
rect 8886 17660 8892 17672
rect 52068 17660 52074 17672
rect 8886 17632 52074 17660
rect 8886 17620 8892 17632
rect 52068 17620 52074 17632
rect 52126 17620 52132 17672
rect 8736 17552 8742 17604
rect 8794 17592 8800 17604
rect 55380 17592 55386 17604
rect 8794 17564 55386 17592
rect 8794 17552 8800 17564
rect 55380 17552 55386 17564
rect 55438 17552 55444 17604
rect 5056 17484 5062 17536
rect 5114 17524 5120 17536
rect 53451 17527 53509 17533
rect 53451 17524 53463 17527
rect 5114 17496 53463 17524
rect 5114 17484 5120 17496
rect 53451 17493 53463 17496
rect 53497 17493 53509 17527
rect 53451 17487 53509 17493
rect 1086 17434 58862 17456
rect 1086 17382 4228 17434
rect 4280 17382 4292 17434
rect 4344 17382 4356 17434
rect 4408 17382 4420 17434
rect 4472 17382 34948 17434
rect 35000 17382 35012 17434
rect 35064 17382 35076 17434
rect 35128 17382 35140 17434
rect 35192 17382 58862 17434
rect 1086 17360 58862 17382
rect 8828 17320 8834 17332
rect 8800 17280 8834 17320
rect 8886 17280 8892 17332
rect 8800 17204 8828 17280
rect 9104 17246 9110 17298
rect 9162 17246 9168 17298
rect 9564 17212 9570 17264
rect 9622 17252 9628 17264
rect 35324 17252 35330 17264
rect 9622 17224 35330 17252
rect 9622 17212 9628 17224
rect 35324 17212 35330 17224
rect 35382 17212 35388 17264
rect 3955 17119 4013 17125
rect 3955 17085 3967 17119
rect 4001 17116 4013 17119
rect 8000 17116 8006 17128
rect 4001 17088 8006 17116
rect 4001 17085 4013 17088
rect 3955 17079 4013 17085
rect 8000 17076 8006 17088
rect 8058 17076 8064 17128
rect 8736 17116 8742 17128
rect 8446 17088 8742 17116
rect 8736 17076 8742 17088
rect 8794 17076 8800 17128
rect 1086 16890 58862 16912
rect 1086 16838 19588 16890
rect 19640 16838 19652 16890
rect 19704 16838 19716 16890
rect 19768 16838 19780 16890
rect 19832 16838 50308 16890
rect 50360 16838 50372 16890
rect 50424 16838 50436 16890
rect 50488 16838 50500 16890
rect 50552 16838 58862 16890
rect 1086 16816 58862 16838
rect 8000 16736 8006 16788
rect 8058 16776 8064 16788
rect 51884 16776 51890 16788
rect 8058 16748 51890 16776
rect 8058 16736 8064 16748
rect 51884 16736 51890 16748
rect 51942 16736 51948 16788
rect 25756 16600 25762 16652
rect 25814 16640 25820 16652
rect 25940 16640 25946 16652
rect 25814 16612 25946 16640
rect 25814 16600 25820 16612
rect 25940 16600 25946 16612
rect 25998 16600 26004 16652
rect 39648 16600 39654 16652
rect 39706 16640 39712 16652
rect 39924 16640 39930 16652
rect 39706 16612 39930 16640
rect 39706 16600 39712 16612
rect 39924 16600 39930 16612
rect 39982 16600 39988 16652
rect 8644 16396 8650 16448
rect 8702 16436 8708 16448
rect 51056 16436 51062 16448
rect 8702 16408 51062 16436
rect 8702 16396 8708 16408
rect 51056 16396 51062 16408
rect 51114 16396 51120 16448
rect 1086 16346 58862 16368
rect 1086 16294 4228 16346
rect 4280 16294 4292 16346
rect 4344 16294 4356 16346
rect 4408 16294 4420 16346
rect 4472 16294 34948 16346
rect 35000 16294 35012 16346
rect 35064 16294 35076 16346
rect 35128 16294 35140 16346
rect 35192 16294 58862 16346
rect 1086 16272 58862 16294
rect 8736 16192 8742 16244
rect 8794 16192 8800 16244
rect 8644 16074 8650 16126
rect 8702 16074 8708 16126
rect 16648 16028 16654 16040
rect 16609 16000 16654 16028
rect 16648 15988 16654 16000
rect 16706 15988 16712 16040
rect 8736 15852 8742 15904
rect 8794 15892 8800 15904
rect 33852 15892 33858 15904
rect 8794 15864 33858 15892
rect 8794 15852 8800 15864
rect 33852 15852 33858 15864
rect 33910 15852 33916 15904
rect 1086 15802 58862 15824
rect 1086 15750 19588 15802
rect 19640 15750 19652 15802
rect 19704 15750 19716 15802
rect 19768 15750 19780 15802
rect 19832 15750 50308 15802
rect 50360 15750 50372 15802
rect 50424 15750 50436 15802
rect 50488 15750 50500 15802
rect 50552 15750 58862 15802
rect 1086 15728 58862 15750
rect 1100 15648 1106 15700
rect 1158 15688 1164 15700
rect 16648 15688 16654 15700
rect 1158 15660 16654 15688
rect 1158 15648 1164 15660
rect 16648 15648 16654 15660
rect 16706 15648 16712 15700
rect 4231 15351 4289 15357
rect 4231 15317 4243 15351
rect 4277 15348 4289 15351
rect 44800 15348 44806 15360
rect 4277 15320 44806 15348
rect 4277 15317 4289 15320
rect 4231 15311 4289 15317
rect 44800 15308 44806 15320
rect 44858 15308 44864 15360
rect 1086 15258 58862 15280
rect 1086 15206 4228 15258
rect 4280 15206 4292 15258
rect 4344 15206 4356 15258
rect 4408 15206 4420 15258
rect 4472 15206 34948 15258
rect 35000 15206 35012 15258
rect 35064 15206 35076 15258
rect 35128 15206 35140 15258
rect 35192 15206 58862 15258
rect 1086 15184 58862 15206
rect 8460 15104 8466 15156
rect 8518 15104 8524 15156
rect 8644 15104 8650 15156
rect 8702 15144 8708 15156
rect 25480 15144 25486 15156
rect 8702 15116 25486 15144
rect 8702 15104 8708 15116
rect 25480 15104 25486 15116
rect 25538 15104 25544 15156
rect 8644 14968 8650 15020
rect 8702 15008 8708 15020
rect 8702 14980 27274 15008
rect 8702 14968 8708 14980
rect 8923 14943 8981 14949
rect 8276 14866 8282 14918
rect 8334 14866 8340 14918
rect 8923 14909 8935 14943
rect 8969 14940 8981 14943
rect 27136 14940 27142 14952
rect 8969 14912 23962 14940
rect 27097 14912 27142 14940
rect 8969 14909 8981 14912
rect 8923 14903 8981 14909
rect 23934 14872 23962 14912
rect 27136 14900 27142 14912
rect 27194 14900 27200 14952
rect 27246 14940 27274 14980
rect 48388 14940 48394 14952
rect 27246 14912 48394 14940
rect 48388 14900 48394 14912
rect 48446 14900 48452 14952
rect 56671 14943 56729 14949
rect 56671 14909 56683 14943
rect 56717 14909 56729 14943
rect 56671 14903 56729 14909
rect 29712 14872 29718 14884
rect 23934 14844 29718 14872
rect 29712 14832 29718 14844
rect 29770 14832 29776 14884
rect 31460 14832 31466 14884
rect 31518 14872 31524 14884
rect 56686 14872 56714 14903
rect 31518 14844 56714 14872
rect 31518 14832 31524 14844
rect 1086 14714 58862 14736
rect 1086 14662 19588 14714
rect 19640 14662 19652 14714
rect 19704 14662 19716 14714
rect 19768 14662 19780 14714
rect 19832 14662 50308 14714
rect 50360 14662 50372 14714
rect 50424 14662 50436 14714
rect 50488 14662 50500 14714
rect 50552 14662 58862 14714
rect 1086 14640 58862 14662
rect 5240 14492 5246 14544
rect 5298 14532 5304 14544
rect 5424 14532 5430 14544
rect 5298 14504 5430 14532
rect 5298 14492 5304 14504
rect 5424 14492 5430 14504
rect 5482 14492 5488 14544
rect 16832 14492 16838 14544
rect 16890 14532 16896 14544
rect 17016 14532 17022 14544
rect 16890 14504 17022 14532
rect 16890 14492 16896 14504
rect 17016 14492 17022 14504
rect 17074 14492 17080 14544
rect 1086 14170 58862 14192
rect 1086 14118 4228 14170
rect 4280 14118 4292 14170
rect 4344 14118 4356 14170
rect 4408 14118 4420 14170
rect 4472 14118 34948 14170
rect 35000 14118 35012 14170
rect 35064 14118 35076 14170
rect 35128 14118 35140 14170
rect 35192 14118 58862 14170
rect 1086 14096 58862 14118
rect 8828 14016 8834 14068
rect 8886 14056 8892 14068
rect 32196 14056 32202 14068
rect 8886 14028 12002 14056
rect 32157 14028 32202 14056
rect 8886 14016 8892 14028
rect 11974 13988 12002 14028
rect 32196 14016 32202 14028
rect 32254 14016 32260 14068
rect 45720 13988 45726 14000
rect 11974 13960 45726 13988
rect 45720 13948 45726 13960
rect 45778 13948 45784 14000
rect 8000 13880 8006 13932
rect 8058 13920 8064 13932
rect 13060 13920 13066 13932
rect 8058 13892 8262 13920
rect 8354 13892 13066 13920
rect 8058 13880 8064 13892
rect 13060 13880 13066 13892
rect 13118 13880 13124 13932
rect 13428 13880 13434 13932
rect 13486 13920 13492 13932
rect 46275 13923 46333 13929
rect 46275 13920 46287 13923
rect 13486 13892 46287 13920
rect 13486 13880 13492 13892
rect 46275 13889 46287 13892
rect 46321 13889 46333 13923
rect 46275 13883 46333 13889
rect 12603 13855 12661 13861
rect 12603 13821 12615 13855
rect 12649 13852 12661 13855
rect 20144 13852 20150 13864
rect 12649 13824 20150 13852
rect 12649 13821 12661 13824
rect 12603 13815 12661 13821
rect 20144 13812 20150 13824
rect 20202 13812 20208 13864
rect 1086 13626 58862 13648
rect 1086 13574 19588 13626
rect 19640 13574 19652 13626
rect 19704 13574 19716 13626
rect 19768 13574 19780 13626
rect 19832 13574 50308 13626
rect 50360 13574 50372 13626
rect 50424 13574 50436 13626
rect 50488 13574 50500 13626
rect 50552 13574 58862 13626
rect 1086 13552 58862 13574
rect 6528 13376 6534 13388
rect 6489 13348 6534 13376
rect 6528 13336 6534 13348
rect 6586 13336 6592 13388
rect 1086 13082 58862 13104
rect 1086 13030 4228 13082
rect 4280 13030 4292 13082
rect 4344 13030 4356 13082
rect 4408 13030 4420 13082
rect 4472 13030 34948 13082
rect 35000 13030 35012 13082
rect 35064 13030 35076 13082
rect 35128 13030 35140 13082
rect 35192 13030 58862 13082
rect 1086 13008 58862 13030
rect 8138 12928 8144 12980
rect 8196 12928 8202 12980
rect 9843 12903 9901 12909
rect 9843 12869 9855 12903
rect 9889 12900 9901 12903
rect 18948 12900 18954 12912
rect 9889 12872 18954 12900
rect 9889 12869 9901 12872
rect 9843 12863 9901 12869
rect 18948 12860 18954 12872
rect 19006 12860 19012 12912
rect 42960 12832 42966 12844
rect 8262 12804 42966 12832
rect 42960 12792 42966 12804
rect 43018 12792 43024 12844
rect 8920 12724 8926 12776
rect 8978 12764 8984 12776
rect 15179 12767 15237 12773
rect 15179 12764 15191 12767
rect 8978 12736 15191 12764
rect 8978 12724 8984 12736
rect 15179 12733 15191 12736
rect 15225 12733 15237 12767
rect 15179 12727 15237 12733
rect 40663 12767 40721 12773
rect 40663 12733 40675 12767
rect 40709 12764 40721 12767
rect 51976 12764 51982 12776
rect 40709 12736 51982 12764
rect 40709 12733 40721 12736
rect 40663 12727 40721 12733
rect 51976 12724 51982 12736
rect 52034 12724 52040 12776
rect 21984 12588 21990 12640
rect 22042 12628 22048 12640
rect 46091 12631 46149 12637
rect 46091 12628 46103 12631
rect 22042 12600 46103 12628
rect 22042 12588 22048 12600
rect 46091 12597 46103 12600
rect 46137 12597 46149 12631
rect 46091 12591 46149 12597
rect 1086 12538 58862 12560
rect 1086 12486 19588 12538
rect 19640 12486 19652 12538
rect 19704 12486 19716 12538
rect 19768 12486 19780 12538
rect 19832 12486 50308 12538
rect 50360 12486 50372 12538
rect 50424 12486 50436 12538
rect 50488 12486 50500 12538
rect 50552 12486 58862 12538
rect 1086 12464 58862 12486
rect 5792 12044 5798 12096
rect 5850 12084 5856 12096
rect 37903 12087 37961 12093
rect 37903 12084 37915 12087
rect 5850 12056 37915 12084
rect 5850 12044 5856 12056
rect 37903 12053 37915 12056
rect 37949 12053 37961 12087
rect 47192 12084 47198 12096
rect 47153 12056 47198 12084
rect 37903 12047 37961 12053
rect 47192 12044 47198 12056
rect 47250 12044 47256 12096
rect 1086 11994 58862 12016
rect 1086 11942 4228 11994
rect 4280 11942 4292 11994
rect 4344 11942 4356 11994
rect 4408 11942 4420 11994
rect 4472 11942 34948 11994
rect 35000 11942 35012 11994
rect 35064 11942 35076 11994
rect 35128 11942 35140 11994
rect 35192 11942 58862 11994
rect 1086 11920 58862 11942
rect 35324 11840 35330 11892
rect 35382 11880 35388 11892
rect 47192 11880 47198 11892
rect 35382 11852 47198 11880
rect 35382 11840 35388 11852
rect 47192 11840 47198 11852
rect 47250 11840 47256 11892
rect 8230 11602 8236 11654
rect 8288 11602 8294 11654
rect 8460 11636 8466 11688
rect 8518 11676 8524 11688
rect 38728 11676 38734 11688
rect 8518 11648 38734 11676
rect 8518 11636 8524 11648
rect 38728 11636 38734 11648
rect 38786 11636 38792 11688
rect 33760 11540 33766 11552
rect 8354 11512 33766 11540
rect 33760 11500 33766 11512
rect 33818 11500 33824 11552
rect 1086 11450 58862 11472
rect 1086 11398 19588 11450
rect 19640 11398 19652 11450
rect 19704 11398 19716 11450
rect 19768 11398 19780 11450
rect 19832 11398 50308 11450
rect 50360 11398 50372 11450
rect 50424 11398 50436 11450
rect 50488 11398 50500 11450
rect 50552 11398 58862 11450
rect 1086 11376 58862 11398
rect 9196 11160 9202 11212
rect 9254 11200 9260 11212
rect 9380 11200 9386 11212
rect 9254 11172 9386 11200
rect 9254 11160 9260 11172
rect 9380 11160 9386 11172
rect 9438 11160 9444 11212
rect 31184 11132 31190 11144
rect 31145 11104 31190 11132
rect 31184 11092 31190 11104
rect 31242 11092 31248 11144
rect 31110 11036 31322 11064
rect 9288 10956 9294 11008
rect 9346 10996 9352 11008
rect 31110 10996 31138 11036
rect 9346 10968 31138 10996
rect 31294 10996 31322 11036
rect 33300 10996 33306 11008
rect 31294 10968 33306 10996
rect 9346 10956 9352 10968
rect 33300 10956 33306 10968
rect 33358 10956 33364 11008
rect 1086 10906 58862 10928
rect 1086 10854 4228 10906
rect 4280 10854 4292 10906
rect 4344 10854 4356 10906
rect 4408 10854 4420 10906
rect 4472 10854 34948 10906
rect 35000 10854 35012 10906
rect 35064 10854 35076 10906
rect 35128 10854 35140 10906
rect 35192 10854 58862 10906
rect 1086 10832 58862 10854
rect 38636 10792 38642 10804
rect 8524 10764 38642 10792
rect 8524 10588 8552 10764
rect 38636 10752 38642 10764
rect 38694 10752 38700 10804
rect 13244 10588 13250 10600
rect 8294 10560 8552 10588
rect 9550 10560 13250 10588
rect 8294 10472 8322 10560
rect 13244 10548 13250 10560
rect 13302 10548 13308 10600
rect 42135 10591 42193 10597
rect 42135 10557 42147 10591
rect 42181 10588 42193 10591
rect 52068 10588 52074 10600
rect 42181 10560 52074 10588
rect 42181 10557 42193 10560
rect 42135 10551 42193 10557
rect 52068 10548 52074 10560
rect 52126 10548 52132 10600
rect 9288 10480 9294 10532
rect 9346 10480 9352 10532
rect 37256 10452 37262 10464
rect 9826 10424 37262 10452
rect 37256 10412 37262 10424
rect 37314 10412 37320 10464
rect 1086 10362 58862 10384
rect 1086 10310 19588 10362
rect 19640 10310 19652 10362
rect 19704 10310 19716 10362
rect 19768 10310 19780 10362
rect 19832 10310 50308 10362
rect 50360 10310 50372 10362
rect 50424 10310 50436 10362
rect 50488 10310 50500 10362
rect 50552 10310 58862 10362
rect 1086 10288 58862 10310
rect 13244 10208 13250 10260
rect 13302 10248 13308 10260
rect 34588 10248 34594 10260
rect 13302 10220 34594 10248
rect 13302 10208 13308 10220
rect 34588 10208 34594 10220
rect 34646 10208 34652 10260
rect 27507 9979 27565 9985
rect 27507 9945 27519 9979
rect 27553 9976 27565 9979
rect 32840 9976 32846 9988
rect 27553 9948 32846 9976
rect 27553 9945 27565 9948
rect 27507 9939 27565 9945
rect 32840 9936 32846 9948
rect 32898 9936 32904 9988
rect 31003 9911 31061 9917
rect 31003 9877 31015 9911
rect 31049 9908 31061 9911
rect 32748 9908 32754 9920
rect 31049 9880 32754 9908
rect 31049 9877 31061 9880
rect 31003 9871 31061 9877
rect 32748 9868 32754 9880
rect 32806 9868 32812 9920
rect 1086 9818 58862 9840
rect 1086 9766 4228 9818
rect 4280 9766 4292 9818
rect 4344 9766 4356 9818
rect 4408 9766 4420 9818
rect 4472 9766 34948 9818
rect 35000 9766 35012 9818
rect 35064 9766 35076 9818
rect 35128 9766 35140 9818
rect 35192 9766 58862 9818
rect 1086 9744 58862 9766
rect 3216 9664 3222 9716
rect 3274 9704 3280 9716
rect 3492 9704 3498 9716
rect 3274 9676 3498 9704
rect 3274 9664 3280 9676
rect 3492 9664 3498 9676
rect 3550 9664 3556 9716
rect 7448 9664 7454 9716
rect 7506 9704 7512 9716
rect 7816 9704 7822 9716
rect 7506 9676 7822 9704
rect 7506 9664 7512 9676
rect 7816 9664 7822 9676
rect 7874 9664 7880 9716
rect 36888 9664 36894 9716
rect 36946 9704 36952 9716
rect 37072 9704 37078 9716
rect 36946 9676 37078 9704
rect 36946 9664 36952 9676
rect 37072 9664 37078 9676
rect 37130 9664 37136 9716
rect 32107 9503 32165 9509
rect 8368 9426 8374 9478
rect 8426 9426 8432 9478
rect 32107 9469 32119 9503
rect 32153 9500 32165 9503
rect 41120 9500 41126 9512
rect 32153 9472 41126 9500
rect 32153 9469 32165 9472
rect 32107 9463 32165 9469
rect 41120 9460 41126 9472
rect 41178 9460 41184 9512
rect 43512 9500 43518 9512
rect 43473 9472 43518 9500
rect 43512 9460 43518 9472
rect 43570 9460 43576 9512
rect 47468 9500 47474 9512
rect 47429 9472 47474 9500
rect 47468 9460 47474 9472
rect 47526 9460 47532 9512
rect 52439 9503 52497 9509
rect 52439 9469 52451 9503
rect 52485 9500 52497 9503
rect 54920 9500 54926 9512
rect 52485 9472 54926 9500
rect 52485 9469 52497 9472
rect 52439 9463 52497 9469
rect 54920 9460 54926 9472
rect 54978 9460 54984 9512
rect 29620 9432 29626 9444
rect 9490 9404 29626 9432
rect 9490 9384 9518 9404
rect 29620 9392 29626 9404
rect 29678 9392 29684 9444
rect 13704 9324 13710 9376
rect 13762 9364 13768 9376
rect 56671 9367 56729 9373
rect 56671 9364 56683 9367
rect 13762 9336 56683 9364
rect 13762 9324 13768 9336
rect 56671 9333 56683 9336
rect 56717 9333 56729 9367
rect 56671 9327 56729 9333
rect 1086 9274 58862 9296
rect 1086 9222 19588 9274
rect 19640 9222 19652 9274
rect 19704 9222 19716 9274
rect 19768 9222 19780 9274
rect 19832 9222 50308 9274
rect 50360 9222 50372 9274
rect 50424 9222 50436 9274
rect 50488 9222 50500 9274
rect 50552 9222 58862 9274
rect 1086 9200 58862 9222
rect 19224 9120 19230 9172
rect 19282 9160 19288 9172
rect 19503 9163 19561 9169
rect 19503 9160 19515 9163
rect 19282 9132 19515 9160
rect 19282 9120 19288 9132
rect 19503 9129 19515 9132
rect 19549 9129 19561 9163
rect 19503 9123 19561 9129
rect 25204 9120 25210 9172
rect 25262 9160 25268 9172
rect 43512 9160 43518 9172
rect 25262 9132 43518 9160
rect 25262 9120 25268 9132
rect 43512 9120 43518 9132
rect 43570 9120 43576 9172
rect 3952 9052 3958 9104
rect 4010 9092 4016 9104
rect 47468 9092 47474 9104
rect 4010 9064 47474 9092
rect 4010 9052 4016 9064
rect 47468 9052 47474 9064
rect 47526 9052 47532 9104
rect 8368 8984 8374 9036
rect 8426 9024 8432 9036
rect 29252 9024 29258 9036
rect 8426 8996 29258 9024
rect 8426 8984 8432 8996
rect 29252 8984 29258 8996
rect 29310 8984 29316 9036
rect 5240 8780 5246 8832
rect 5298 8820 5304 8832
rect 39740 8820 39746 8832
rect 5298 8792 39746 8820
rect 5298 8780 5304 8792
rect 39740 8780 39746 8792
rect 39798 8780 39804 8832
rect 49676 8780 49682 8832
rect 49734 8820 49740 8832
rect 53635 8823 53693 8829
rect 53635 8820 53647 8823
rect 49734 8792 53647 8820
rect 49734 8780 49740 8792
rect 53635 8789 53647 8792
rect 53681 8789 53693 8823
rect 53635 8783 53693 8789
rect 1086 8730 58862 8752
rect 1086 8678 4228 8730
rect 4280 8678 4292 8730
rect 4344 8678 4356 8730
rect 4408 8678 4420 8730
rect 4472 8678 34948 8730
rect 35000 8678 35012 8730
rect 35064 8678 35076 8730
rect 35128 8678 35140 8730
rect 35192 8678 58862 8730
rect 1086 8656 58862 8678
rect 39740 8616 39746 8628
rect 39701 8588 39746 8616
rect 8570 8480 8598 8568
rect 8828 8508 8834 8560
rect 8886 8548 8892 8560
rect 17770 8554 17890 8582
rect 39740 8576 39746 8588
rect 39798 8576 39804 8628
rect 17770 8548 17798 8554
rect 8886 8520 17798 8548
rect 17862 8548 17890 8554
rect 26584 8548 26590 8560
rect 17862 8520 26590 8548
rect 8886 8508 8892 8520
rect 26584 8508 26590 8520
rect 26642 8508 26648 8560
rect 48296 8508 48302 8560
rect 48354 8548 48360 8560
rect 57499 8551 57557 8557
rect 57499 8548 57511 8551
rect 48354 8520 57511 8548
rect 48354 8508 48360 8520
rect 57499 8517 57511 8520
rect 57545 8517 57557 8551
rect 57499 8511 57557 8517
rect 27412 8480 27418 8492
rect 8570 8452 27418 8480
rect 27412 8440 27418 8452
rect 27470 8440 27476 8492
rect 27504 8440 27510 8492
rect 27562 8480 27568 8492
rect 29068 8480 29074 8492
rect 27562 8452 29074 8480
rect 27562 8440 27568 8452
rect 29068 8440 29074 8452
rect 29126 8440 29132 8492
rect 8552 8412 8558 8424
rect 8262 8384 8558 8412
rect 8552 8372 8558 8384
rect 8610 8372 8616 8424
rect 10576 8372 10582 8424
rect 10634 8412 10640 8424
rect 48204 8412 48210 8424
rect 10634 8384 48210 8412
rect 10634 8372 10640 8384
rect 48204 8372 48210 8384
rect 48262 8372 48268 8424
rect 20144 8304 20150 8356
rect 20202 8344 20208 8356
rect 20512 8344 20518 8356
rect 20202 8316 20518 8344
rect 20202 8304 20208 8316
rect 20512 8304 20518 8316
rect 20570 8304 20576 8356
rect 25664 8304 25670 8356
rect 25722 8344 25728 8356
rect 25940 8344 25946 8356
rect 25722 8316 25946 8344
rect 25722 8304 25728 8316
rect 25940 8304 25946 8316
rect 25998 8304 26004 8356
rect 20052 8236 20058 8288
rect 20110 8276 20116 8288
rect 23732 8276 23738 8288
rect 20110 8248 23738 8276
rect 20110 8236 20116 8248
rect 23732 8236 23738 8248
rect 23790 8236 23796 8288
rect 28148 8236 28154 8288
rect 28206 8276 28212 8288
rect 35416 8276 35422 8288
rect 28206 8248 35422 8276
rect 28206 8236 28212 8248
rect 35416 8236 35422 8248
rect 35474 8236 35480 8288
rect 1086 8186 58862 8208
rect 1086 8134 19588 8186
rect 19640 8134 19652 8186
rect 19704 8134 19716 8186
rect 19768 8134 19780 8186
rect 19832 8134 50308 8186
rect 50360 8134 50372 8186
rect 50424 8134 50436 8186
rect 50488 8134 50500 8186
rect 50552 8134 58862 8186
rect 1086 8112 58862 8134
rect 14532 7896 14538 7948
rect 14590 7936 14596 7948
rect 14716 7936 14722 7948
rect 14590 7908 14722 7936
rect 14590 7896 14596 7908
rect 14716 7896 14722 7908
rect 14774 7896 14780 7948
rect 17936 7760 17942 7812
rect 17994 7800 18000 7812
rect 18120 7800 18126 7812
rect 17994 7772 18126 7800
rect 17994 7760 18000 7772
rect 18120 7760 18126 7772
rect 18178 7760 18184 7812
rect 26676 7760 26682 7812
rect 26734 7800 26740 7812
rect 26734 7772 57910 7800
rect 26734 7760 26740 7772
rect 11223 7735 11281 7741
rect 11223 7701 11235 7735
rect 11269 7732 11281 7735
rect 24836 7732 24842 7744
rect 11269 7704 24842 7732
rect 11269 7701 11281 7704
rect 11223 7695 11281 7701
rect 24836 7692 24842 7704
rect 24894 7692 24900 7744
rect 25020 7692 25026 7744
rect 25078 7732 25084 7744
rect 25848 7732 25854 7744
rect 25078 7704 25854 7732
rect 25078 7692 25084 7704
rect 25848 7692 25854 7704
rect 25906 7692 25912 7744
rect 26492 7692 26498 7744
rect 26550 7732 26556 7744
rect 27320 7732 27326 7744
rect 26550 7704 27326 7732
rect 26550 7692 26556 7704
rect 27320 7692 27326 7704
rect 27378 7692 27384 7744
rect 28332 7692 28338 7744
rect 28390 7732 28396 7744
rect 28792 7732 28798 7744
rect 28390 7704 28798 7732
rect 28390 7692 28396 7704
rect 28792 7692 28798 7704
rect 28850 7692 28856 7744
rect 41580 7732 41586 7744
rect 41541 7704 41586 7732
rect 41580 7692 41586 7704
rect 41638 7692 41644 7744
rect 57882 7732 57910 7772
rect 58419 7735 58477 7741
rect 58419 7732 58431 7735
rect 57882 7704 58431 7732
rect 58419 7701 58431 7704
rect 58465 7701 58477 7735
rect 58419 7695 58477 7701
rect 1086 7642 58862 7664
rect 1086 7590 4228 7642
rect 4280 7590 4292 7642
rect 4344 7590 4356 7642
rect 4408 7590 4420 7642
rect 4472 7590 34948 7642
rect 35000 7590 35012 7642
rect 35064 7590 35076 7642
rect 35128 7590 35140 7642
rect 35192 7590 58862 7642
rect 1086 7568 58862 7590
rect 12600 7488 12606 7540
rect 12658 7528 12664 7540
rect 13336 7528 13342 7540
rect 12658 7500 13342 7528
rect 12658 7488 12664 7500
rect 13336 7488 13342 7500
rect 13394 7488 13400 7540
rect 15544 7488 15550 7540
rect 15602 7528 15608 7540
rect 16188 7528 16194 7540
rect 15602 7500 16194 7528
rect 15602 7488 15608 7500
rect 16188 7488 16194 7500
rect 16246 7488 16252 7540
rect 17568 7528 17574 7540
rect 17529 7500 17574 7528
rect 17568 7488 17574 7500
rect 17626 7488 17632 7540
rect 19960 7488 19966 7540
rect 20018 7528 20024 7540
rect 20420 7528 20426 7540
rect 20018 7500 20426 7528
rect 20018 7488 20024 7500
rect 20420 7488 20426 7500
rect 20478 7488 20484 7540
rect 20880 7488 20886 7540
rect 20938 7528 20944 7540
rect 41580 7528 41586 7540
rect 20938 7500 41586 7528
rect 20938 7488 20944 7500
rect 41580 7488 41586 7500
rect 41638 7488 41644 7540
rect 49679 7531 49737 7537
rect 49679 7497 49691 7531
rect 49725 7528 49737 7531
rect 49768 7528 49774 7540
rect 49725 7500 49774 7528
rect 49725 7497 49737 7500
rect 49679 7491 49737 7497
rect 49768 7488 49774 7500
rect 49826 7488 49832 7540
rect 12784 7420 12790 7472
rect 12842 7460 12848 7472
rect 13704 7460 13710 7472
rect 12842 7432 13710 7460
rect 12842 7420 12848 7432
rect 13704 7420 13710 7432
rect 13762 7420 13768 7472
rect 15268 7420 15274 7472
rect 15326 7460 15332 7472
rect 15912 7460 15918 7472
rect 15326 7432 15918 7460
rect 15326 7420 15332 7432
rect 15912 7420 15918 7432
rect 15970 7420 15976 7472
rect 12692 7352 12698 7404
rect 12750 7392 12756 7404
rect 23456 7392 23462 7404
rect 12750 7364 23462 7392
rect 12750 7352 12756 7364
rect 23456 7352 23462 7364
rect 23514 7352 23520 7404
rect 8230 7250 8236 7302
rect 8288 7250 8294 7302
rect 9104 7284 9110 7336
rect 9162 7324 9168 7336
rect 9843 7327 9901 7333
rect 9843 7324 9855 7327
rect 9162 7296 9855 7324
rect 9162 7284 9168 7296
rect 9843 7293 9855 7296
rect 9889 7293 9901 7327
rect 9843 7287 9901 7293
rect 22079 7327 22137 7333
rect 22079 7293 22091 7327
rect 22125 7324 22137 7327
rect 28884 7324 28890 7336
rect 22125 7296 28890 7324
rect 22125 7293 22137 7296
rect 22079 7287 22137 7293
rect 28884 7284 28890 7296
rect 28942 7284 28948 7336
rect 44987 7327 45045 7333
rect 44987 7293 44999 7327
rect 45033 7324 45045 7327
rect 53172 7324 53178 7336
rect 45033 7296 53178 7324
rect 45033 7293 45045 7296
rect 44987 7287 45045 7293
rect 53172 7284 53178 7296
rect 53230 7284 53236 7336
rect 28976 7216 28982 7268
rect 29034 7256 29040 7268
rect 45996 7256 46002 7268
rect 29034 7228 46002 7256
rect 29034 7216 29040 7228
rect 45996 7216 46002 7228
rect 46054 7216 46060 7268
rect 24100 7188 24106 7200
rect 8538 7160 24106 7188
rect 24100 7148 24106 7160
rect 24158 7148 24164 7200
rect 1086 7098 58862 7120
rect 1086 7046 19588 7098
rect 19640 7046 19652 7098
rect 19704 7046 19716 7098
rect 19768 7046 19780 7098
rect 19832 7046 50308 7098
rect 50360 7046 50372 7098
rect 50424 7046 50436 7098
rect 50488 7046 50500 7098
rect 50552 7046 58862 7098
rect 1086 7024 58862 7046
rect 39648 6984 39654 6996
rect 39574 6956 39654 6984
rect 39574 6928 39602 6956
rect 39648 6944 39654 6956
rect 39706 6944 39712 6996
rect 39556 6876 39562 6928
rect 39614 6876 39620 6928
rect 8092 6808 8098 6860
rect 8150 6848 8156 6860
rect 15176 6848 15182 6860
rect 8150 6820 15182 6848
rect 8150 6808 8156 6820
rect 15176 6808 15182 6820
rect 15234 6808 15240 6860
rect 8000 6740 8006 6792
rect 8058 6780 8064 6792
rect 8058 6752 17338 6780
rect 8058 6740 8064 6752
rect 8371 6715 8429 6721
rect 8371 6681 8383 6715
rect 8417 6712 8429 6715
rect 17200 6712 17206 6724
rect 8417 6684 17206 6712
rect 8417 6681 8429 6684
rect 8371 6675 8429 6681
rect 17200 6672 17206 6684
rect 17258 6672 17264 6724
rect 8460 6604 8466 6656
rect 8518 6644 8524 6656
rect 16556 6644 16562 6656
rect 8518 6616 16562 6644
rect 8518 6604 8524 6616
rect 16556 6604 16562 6616
rect 16614 6604 16620 6656
rect 17310 6644 17338 6752
rect 46916 6740 46922 6792
rect 46974 6780 46980 6792
rect 51795 6783 51853 6789
rect 51795 6780 51807 6783
rect 46974 6752 51807 6780
rect 46974 6740 46980 6752
rect 51795 6749 51807 6752
rect 51841 6749 51853 6783
rect 51795 6743 51853 6749
rect 27688 6644 27694 6656
rect 17310 6616 27694 6644
rect 27688 6604 27694 6616
rect 27746 6604 27752 6656
rect 38820 6604 38826 6656
rect 38878 6644 38884 6656
rect 46916 6644 46922 6656
rect 38878 6616 46922 6644
rect 38878 6604 38884 6616
rect 46916 6604 46922 6616
rect 46974 6604 46980 6656
rect 52436 6644 52442 6656
rect 52397 6616 52442 6644
rect 52436 6604 52442 6616
rect 52494 6604 52500 6656
rect 1086 6554 58862 6576
rect 1086 6502 4228 6554
rect 4280 6502 4292 6554
rect 4344 6502 4356 6554
rect 4408 6502 4420 6554
rect 4472 6502 34948 6554
rect 35000 6502 35012 6554
rect 35064 6502 35076 6554
rect 35128 6502 35140 6554
rect 35192 6502 58862 6554
rect 1086 6480 58862 6502
rect 8460 6440 8466 6452
rect 8432 6400 8466 6440
rect 8518 6400 8524 6452
rect 8616 6412 14486 6440
rect 8432 6324 8460 6400
rect 8616 6324 8644 6412
rect 14458 6372 14486 6412
rect 17476 6400 17482 6452
rect 17534 6440 17540 6452
rect 36980 6440 36986 6452
rect 17534 6412 36986 6440
rect 17534 6400 17540 6412
rect 36980 6400 36986 6412
rect 37038 6400 37044 6452
rect 38636 6400 38642 6452
rect 38694 6440 38700 6452
rect 52436 6440 52442 6452
rect 38694 6412 52442 6440
rect 38694 6400 38700 6412
rect 52436 6400 52442 6412
rect 52494 6400 52500 6452
rect 21340 6372 21346 6384
rect 14458 6344 21346 6372
rect 21340 6332 21346 6344
rect 21398 6332 21404 6384
rect 27688 6332 27694 6384
rect 27746 6372 27752 6384
rect 38820 6372 38826 6384
rect 27746 6344 38826 6372
rect 27746 6332 27752 6344
rect 38820 6332 38826 6344
rect 38878 6332 38884 6384
rect 8092 6264 8098 6316
rect 8150 6304 8156 6316
rect 18304 6304 18310 6316
rect 8150 6276 8262 6304
rect 8814 6276 18310 6304
rect 8150 6264 8156 6276
rect 18304 6264 18310 6276
rect 18362 6264 18368 6316
rect 36980 6264 36986 6316
rect 37038 6304 37044 6316
rect 38636 6304 38642 6316
rect 37038 6276 38642 6304
rect 37038 6264 37044 6276
rect 38636 6264 38642 6276
rect 38694 6264 38700 6316
rect 38728 6264 38734 6316
rect 38786 6304 38792 6316
rect 43147 6307 43205 6313
rect 43147 6304 43159 6307
rect 38786 6276 43159 6304
rect 38786 6264 38792 6276
rect 43147 6273 43159 6276
rect 43193 6273 43205 6307
rect 43147 6267 43205 6273
rect 14532 6196 14538 6248
rect 14590 6236 14596 6248
rect 34499 6239 34557 6245
rect 34499 6236 34511 6239
rect 14590 6208 34511 6236
rect 14590 6196 14596 6208
rect 34499 6205 34511 6208
rect 34545 6205 34557 6239
rect 34499 6199 34557 6205
rect 35787 6239 35845 6245
rect 35787 6205 35799 6239
rect 35833 6205 35845 6239
rect 35787 6199 35845 6205
rect 35802 6168 35830 6199
rect 40108 6196 40114 6248
rect 40166 6236 40172 6248
rect 42779 6239 42837 6245
rect 42779 6236 42791 6239
rect 40166 6208 42791 6236
rect 40166 6196 40172 6208
rect 42779 6205 42791 6208
rect 42825 6205 42837 6239
rect 42779 6199 42837 6205
rect 51056 6168 51062 6180
rect 35802 6140 51062 6168
rect 51056 6128 51062 6140
rect 51114 6128 51120 6180
rect 14440 6100 14446 6112
rect 8906 6072 14446 6100
rect 14440 6060 14446 6072
rect 14498 6060 14504 6112
rect 1086 6010 58862 6032
rect 1086 5958 19588 6010
rect 19640 5958 19652 6010
rect 19704 5958 19716 6010
rect 19768 5958 19780 6010
rect 19832 5958 50308 6010
rect 50360 5958 50372 6010
rect 50424 5958 50436 6010
rect 50488 5958 50500 6010
rect 50552 5958 58862 6010
rect 1086 5936 58862 5958
rect 17200 5856 17206 5908
rect 17258 5896 17264 5908
rect 40016 5896 40022 5908
rect 17258 5868 40022 5896
rect 17258 5856 17264 5868
rect 40016 5856 40022 5868
rect 40074 5856 40080 5908
rect 5424 5788 5430 5840
rect 5482 5828 5488 5840
rect 21895 5831 21953 5837
rect 21895 5828 21907 5831
rect 5482 5800 21907 5828
rect 5482 5788 5488 5800
rect 21895 5797 21907 5800
rect 21941 5797 21953 5831
rect 21895 5791 21953 5797
rect 26311 5831 26369 5837
rect 26311 5797 26323 5831
rect 26357 5828 26369 5831
rect 28976 5828 28982 5840
rect 26357 5800 28982 5828
rect 26357 5797 26369 5800
rect 26311 5791 26369 5797
rect 28976 5788 28982 5800
rect 29034 5788 29040 5840
rect 10944 5720 10950 5772
rect 11002 5760 11008 5772
rect 28151 5763 28209 5769
rect 28151 5760 28163 5763
rect 11002 5732 28163 5760
rect 11002 5720 11008 5732
rect 28151 5729 28163 5732
rect 28197 5729 28209 5763
rect 28151 5723 28209 5729
rect 32472 5720 32478 5772
rect 32530 5720 32536 5772
rect 10303 5695 10361 5701
rect 10303 5661 10315 5695
rect 10349 5692 10361 5695
rect 32490 5692 32518 5720
rect 10349 5664 32518 5692
rect 10349 5661 10361 5664
rect 10303 5655 10361 5661
rect 5703 5627 5761 5633
rect 5703 5593 5715 5627
rect 5749 5624 5761 5627
rect 26311 5627 26369 5633
rect 26311 5624 26323 5627
rect 5749 5596 26323 5624
rect 5749 5593 5761 5596
rect 5703 5587 5761 5593
rect 26311 5593 26323 5596
rect 26357 5593 26369 5627
rect 26311 5587 26369 5593
rect 1192 5516 1198 5568
rect 1250 5556 1256 5568
rect 35695 5559 35753 5565
rect 35695 5556 35707 5559
rect 1250 5528 35707 5556
rect 1250 5516 1256 5528
rect 35695 5525 35707 5528
rect 35741 5525 35753 5559
rect 35695 5519 35753 5525
rect 1086 5466 58862 5488
rect 1086 5414 4228 5466
rect 4280 5414 4292 5466
rect 4344 5414 4356 5466
rect 4408 5414 4420 5466
rect 4472 5414 34948 5466
rect 35000 5414 35012 5466
rect 35064 5414 35076 5466
rect 35128 5414 35140 5466
rect 35192 5414 58862 5466
rect 1086 5392 58862 5414
rect 8368 5352 8374 5364
rect 8248 5324 8374 5352
rect 8248 5236 8276 5324
rect 8368 5312 8374 5324
rect 8426 5312 8432 5364
rect 10300 5352 10306 5364
rect 8524 5324 10306 5352
rect 8524 5216 8552 5324
rect 10300 5312 10306 5324
rect 10358 5312 10364 5364
rect 11036 5216 11042 5228
rect 8446 5188 8552 5216
rect 8630 5188 11042 5216
rect 11036 5176 11042 5188
rect 11094 5176 11100 5228
rect 46180 5216 46186 5228
rect 46141 5188 46186 5216
rect 46180 5176 46186 5188
rect 46238 5176 46244 5228
rect 8736 5108 8742 5160
rect 8794 5148 8800 5160
rect 15636 5148 15642 5160
rect 8794 5120 15642 5148
rect 8794 5108 8800 5120
rect 15636 5108 15642 5120
rect 15694 5108 15700 5160
rect 32380 5108 32386 5160
rect 32438 5148 32444 5160
rect 33763 5151 33821 5157
rect 33763 5148 33775 5151
rect 32438 5120 33775 5148
rect 32438 5108 32444 5120
rect 33763 5117 33775 5120
rect 33809 5117 33821 5151
rect 33763 5111 33821 5117
rect 52436 5108 52442 5160
rect 52494 5148 52500 5160
rect 55107 5151 55165 5157
rect 55107 5148 55119 5151
rect 52494 5120 55119 5148
rect 52494 5108 52500 5120
rect 55107 5117 55119 5120
rect 55153 5117 55165 5151
rect 55107 5111 55165 5117
rect 8644 4972 8650 5024
rect 8702 4972 8708 5024
rect 20052 4972 20058 5024
rect 20110 5012 20116 5024
rect 22628 5012 22634 5024
rect 20110 4984 22634 5012
rect 20110 4972 20116 4984
rect 22628 4972 22634 4984
rect 22686 4972 22692 5024
rect 50136 4972 50142 5024
rect 50194 5012 50200 5024
rect 55288 5012 55294 5024
rect 50194 4984 55294 5012
rect 50194 4972 50200 4984
rect 55288 4972 55294 4984
rect 55346 4972 55352 5024
rect 1086 4922 58862 4944
rect 1086 4870 19588 4922
rect 19640 4870 19652 4922
rect 19704 4870 19716 4922
rect 19768 4870 19780 4922
rect 19832 4870 50308 4922
rect 50360 4870 50372 4922
rect 50424 4870 50436 4922
rect 50488 4870 50500 4922
rect 50552 4870 58862 4922
rect 1086 4848 58862 4870
rect 20052 4768 20058 4820
rect 20110 4808 20116 4820
rect 20328 4808 20334 4820
rect 20110 4780 20334 4808
rect 20110 4768 20116 4780
rect 20328 4768 20334 4780
rect 20386 4768 20392 4820
rect 32840 4768 32846 4820
rect 32898 4808 32904 4820
rect 33116 4808 33122 4820
rect 32898 4780 33122 4808
rect 32898 4768 32904 4780
rect 33116 4768 33122 4780
rect 33174 4768 33180 4820
rect 48940 4768 48946 4820
rect 48998 4808 49004 4820
rect 52712 4808 52718 4820
rect 48998 4780 52718 4808
rect 48998 4768 49004 4780
rect 52712 4768 52718 4780
rect 52770 4768 52776 4820
rect 17108 4700 17114 4752
rect 17166 4740 17172 4752
rect 18580 4740 18586 4752
rect 17166 4712 18586 4740
rect 17166 4700 17172 4712
rect 18580 4700 18586 4712
rect 18638 4700 18644 4752
rect 6896 4632 6902 4684
rect 6954 4672 6960 4684
rect 9012 4672 9018 4684
rect 6954 4644 9018 4672
rect 6954 4632 6960 4644
rect 9012 4632 9018 4644
rect 9070 4632 9076 4684
rect 13060 4564 13066 4616
rect 13118 4604 13124 4616
rect 14808 4604 14814 4616
rect 13118 4576 14814 4604
rect 13118 4564 13124 4576
rect 14808 4564 14814 4576
rect 14866 4564 14872 4616
rect 1086 4378 58862 4400
rect 1086 4326 4228 4378
rect 4280 4326 4292 4378
rect 4344 4326 4356 4378
rect 4408 4326 4420 4378
rect 4472 4326 34948 4378
rect 35000 4326 35012 4378
rect 35064 4326 35076 4378
rect 35128 4326 35140 4378
rect 35192 4326 58862 4378
rect 1086 4304 58862 4326
rect 16740 4224 16746 4276
rect 16798 4264 16804 4276
rect 17016 4264 17022 4276
rect 16798 4236 17022 4264
rect 16798 4224 16804 4236
rect 17016 4224 17022 4236
rect 17074 4224 17080 4276
rect 20420 4224 20426 4276
rect 20478 4264 20484 4276
rect 23827 4267 23885 4273
rect 23827 4264 23839 4267
rect 20478 4236 23839 4264
rect 20478 4224 20484 4236
rect 23827 4233 23839 4236
rect 23873 4233 23885 4267
rect 23827 4227 23885 4233
rect 32564 4224 32570 4276
rect 32622 4264 32628 4276
rect 32622 4236 34542 4264
rect 32622 4224 32628 4236
rect 22922 4168 23410 4196
rect 3676 4088 3682 4140
rect 3734 4128 3740 4140
rect 3952 4128 3958 4140
rect 3734 4100 3958 4128
rect 3734 4088 3740 4100
rect 3952 4088 3958 4100
rect 4010 4088 4016 4140
rect 6160 4088 6166 4140
rect 6218 4128 6224 4140
rect 6712 4128 6718 4140
rect 6218 4100 6718 4128
rect 6218 4088 6224 4100
rect 6712 4088 6718 4100
rect 6770 4088 6776 4140
rect 7264 4088 7270 4140
rect 7322 4128 7328 4140
rect 7724 4128 7730 4140
rect 7322 4100 7730 4128
rect 7322 4088 7328 4100
rect 7724 4088 7730 4100
rect 7782 4088 7788 4140
rect 8920 4128 8926 4140
rect 8722 4100 8926 4128
rect 8920 4088 8926 4100
rect 8978 4088 8984 4140
rect 10208 4088 10214 4140
rect 10266 4128 10272 4140
rect 10760 4128 10766 4140
rect 10266 4100 10766 4128
rect 10266 4088 10272 4100
rect 10760 4088 10766 4100
rect 10818 4088 10824 4140
rect 11680 4088 11686 4140
rect 11738 4128 11744 4140
rect 12324 4128 12330 4140
rect 11738 4100 12330 4128
rect 11738 4088 11744 4100
rect 12324 4088 12330 4100
rect 12382 4088 12388 4140
rect 12968 4088 12974 4140
rect 13026 4128 13032 4140
rect 13428 4128 13434 4140
rect 13026 4100 13434 4128
rect 13026 4088 13032 4100
rect 13428 4088 13434 4100
rect 13486 4088 13492 4140
rect 14624 4088 14630 4140
rect 14682 4128 14688 4140
rect 15452 4128 15458 4140
rect 14682 4100 15458 4128
rect 14682 4088 14688 4100
rect 15452 4088 15458 4100
rect 15510 4088 15516 4140
rect 16004 4088 16010 4140
rect 16062 4128 16068 4140
rect 16464 4128 16470 4140
rect 16062 4100 16470 4128
rect 16062 4088 16068 4100
rect 16464 4088 16470 4100
rect 16522 4088 16528 4140
rect 17108 4088 17114 4140
rect 17166 4128 17172 4140
rect 17844 4128 17850 4140
rect 17166 4100 17850 4128
rect 17166 4088 17172 4100
rect 17844 4088 17850 4100
rect 17902 4088 17908 4140
rect 18672 4088 18678 4140
rect 18730 4128 18736 4140
rect 19316 4128 19322 4140
rect 18730 4100 19322 4128
rect 18730 4088 18736 4100
rect 19316 4088 19322 4100
rect 19374 4088 19380 4140
rect 21432 4088 21438 4140
rect 21490 4128 21496 4140
rect 22168 4128 22174 4140
rect 21490 4100 22174 4128
rect 21490 4088 21496 4100
rect 22168 4088 22174 4100
rect 22226 4088 22232 4140
rect 22260 4088 22266 4140
rect 22318 4128 22324 4140
rect 22922 4128 22950 4168
rect 23382 4140 23410 4168
rect 30926 4168 31598 4196
rect 22318 4100 22950 4128
rect 22318 4088 22324 4100
rect 22996 4088 23002 4140
rect 23054 4128 23060 4140
rect 23272 4128 23278 4140
rect 23054 4100 23278 4128
rect 23054 4088 23060 4100
rect 23272 4088 23278 4100
rect 23330 4088 23336 4140
rect 23364 4088 23370 4140
rect 23422 4088 23428 4140
rect 24100 4088 24106 4140
rect 24158 4128 24164 4140
rect 24744 4128 24750 4140
rect 24158 4100 24750 4128
rect 24158 4088 24164 4100
rect 24744 4088 24750 4100
rect 24802 4088 24808 4140
rect 25572 4088 25578 4140
rect 25630 4128 25636 4140
rect 26124 4128 26130 4140
rect 25630 4100 26130 4128
rect 25630 4088 25636 4100
rect 26124 4088 26130 4100
rect 26182 4088 26188 4140
rect 27136 4088 27142 4140
rect 27194 4128 27200 4140
rect 27780 4128 27786 4140
rect 27194 4100 27786 4128
rect 27194 4088 27200 4100
rect 27780 4088 27786 4100
rect 27838 4088 27844 4140
rect 29712 4088 29718 4140
rect 29770 4128 29776 4140
rect 30926 4128 30954 4168
rect 29770 4100 30954 4128
rect 29770 4088 29776 4100
rect 31000 4088 31006 4140
rect 31058 4128 31064 4140
rect 31460 4128 31466 4140
rect 31058 4100 31466 4128
rect 31058 4088 31064 4100
rect 31460 4088 31466 4100
rect 31518 4088 31524 4140
rect 31570 4128 31598 4168
rect 32030 4168 33070 4196
rect 32030 4128 32058 4168
rect 31570 4100 32058 4128
rect 32104 4088 32110 4140
rect 32162 4128 32168 4140
rect 32932 4128 32938 4140
rect 32162 4100 32938 4128
rect 32162 4088 32168 4100
rect 32932 4088 32938 4100
rect 32990 4088 32996 4140
rect 33042 4128 33070 4168
rect 33042 4100 33530 4128
rect 2848 4020 2854 4072
rect 2906 4060 2912 4072
rect 3860 4060 3866 4072
rect 2906 4032 3866 4060
rect 2906 4020 2912 4032
rect 3860 4020 3866 4032
rect 3918 4020 3924 4072
rect 4596 4020 4602 4072
rect 4654 4060 4660 4072
rect 5056 4060 5062 4072
rect 4654 4032 5062 4060
rect 4654 4020 4660 4032
rect 5056 4020 5062 4032
rect 5114 4020 5120 4072
rect 6804 4020 6810 4072
rect 6862 4060 6868 4072
rect 6862 4032 8262 4060
rect 6862 4020 6868 4032
rect 9840 4020 9846 4072
rect 9898 4060 9904 4072
rect 10852 4060 10858 4072
rect 9898 4032 10858 4060
rect 9898 4020 9904 4032
rect 10852 4020 10858 4032
rect 10910 4020 10916 4072
rect 11312 4020 11318 4072
rect 11370 4060 11376 4072
rect 12140 4060 12146 4072
rect 11370 4032 12146 4060
rect 11370 4020 11376 4032
rect 12140 4020 12146 4032
rect 12198 4020 12204 4072
rect 13060 4020 13066 4072
rect 13118 4060 13124 4072
rect 13612 4060 13618 4072
rect 13118 4032 13618 4060
rect 13118 4020 13124 4032
rect 13612 4020 13618 4032
rect 13670 4020 13676 4072
rect 13796 4020 13802 4072
rect 13854 4060 13860 4072
rect 14992 4060 14998 4072
rect 13854 4032 14998 4060
rect 13854 4020 13860 4032
rect 14992 4020 14998 4032
rect 15050 4020 15056 4072
rect 15636 4020 15642 4072
rect 15694 4060 15700 4072
rect 16372 4060 16378 4072
rect 15694 4032 16378 4060
rect 15694 4020 15700 4032
rect 16372 4020 16378 4032
rect 16430 4020 16436 4072
rect 24836 4020 24842 4072
rect 24894 4060 24900 4072
rect 26308 4060 26314 4072
rect 24894 4032 26314 4060
rect 24894 4020 24900 4032
rect 26308 4020 26314 4032
rect 26366 4020 26372 4072
rect 27044 4020 27050 4072
rect 27102 4060 27108 4072
rect 30080 4060 30086 4072
rect 27102 4032 30086 4060
rect 27102 4020 27108 4032
rect 30080 4020 30086 4032
rect 30138 4020 30144 4072
rect 30632 4020 30638 4072
rect 30690 4060 30696 4072
rect 31552 4060 31558 4072
rect 30690 4032 31558 4060
rect 30690 4020 30696 4032
rect 31552 4020 31558 4032
rect 31610 4020 31616 4072
rect 31736 4020 31742 4072
rect 31794 4060 31800 4072
rect 33024 4060 33030 4072
rect 31794 4032 33030 4060
rect 31794 4020 31800 4032
rect 33024 4020 33030 4032
rect 33082 4020 33088 4072
rect 33502 4060 33530 4100
rect 33576 4088 33582 4140
rect 33634 4128 33640 4140
rect 34404 4128 34410 4140
rect 33634 4100 34410 4128
rect 33634 4088 33640 4100
rect 34404 4088 34410 4100
rect 34462 4088 34468 4140
rect 34514 4128 34542 4236
rect 50596 4224 50602 4276
rect 50654 4264 50660 4276
rect 56392 4264 56398 4276
rect 50654 4236 56398 4264
rect 50654 4224 50660 4236
rect 56392 4224 56398 4236
rect 56450 4224 56456 4276
rect 37550 4168 38682 4196
rect 37550 4128 37578 4168
rect 34514 4100 37578 4128
rect 37624 4088 37630 4140
rect 37682 4128 37688 4140
rect 38544 4128 38550 4140
rect 37682 4100 38550 4128
rect 37682 4088 37688 4100
rect 38544 4088 38550 4100
rect 38602 4088 38608 4140
rect 33502 4032 35554 4060
rect 5056 3884 5062 3936
rect 5114 3924 5120 3936
rect 5240 3924 5246 3936
rect 5114 3896 5246 3924
rect 5114 3884 5120 3896
rect 5240 3884 5246 3896
rect 5298 3884 5304 3936
rect 7540 3884 7546 3936
rect 7598 3924 7604 3936
rect 8432 3924 8460 4012
rect 12784 3952 12790 4004
rect 12842 3992 12848 4004
rect 13244 3992 13250 4004
rect 12842 3964 13250 3992
rect 12842 3952 12848 3964
rect 13244 3952 13250 3964
rect 13302 3952 13308 4004
rect 18488 3952 18494 4004
rect 18546 3992 18552 4004
rect 20696 3992 20702 4004
rect 18546 3964 20702 3992
rect 18546 3952 18552 3964
rect 20696 3952 20702 3964
rect 20754 3952 20760 4004
rect 21156 3952 21162 4004
rect 21214 3992 21220 4004
rect 21800 3992 21806 4004
rect 21214 3964 21806 3992
rect 21214 3952 21220 3964
rect 21800 3952 21806 3964
rect 21858 3952 21864 4004
rect 25112 3952 25118 4004
rect 25170 3992 25176 4004
rect 26124 3992 26130 4004
rect 25170 3964 26130 3992
rect 25170 3952 25176 3964
rect 26124 3952 26130 3964
rect 26182 3952 26188 4004
rect 7598 3896 8460 3924
rect 7598 3884 7604 3896
rect 13152 3884 13158 3936
rect 13210 3924 13216 3936
rect 14440 3924 14446 3936
rect 13210 3896 14446 3924
rect 13210 3884 13216 3896
rect 14440 3884 14446 3896
rect 14498 3884 14504 3936
rect 18120 3884 18126 3936
rect 18178 3924 18184 3936
rect 20420 3924 20426 3936
rect 18178 3896 20426 3924
rect 18178 3884 18184 3896
rect 20420 3884 20426 3896
rect 20478 3884 20484 3936
rect 25664 3884 25670 3936
rect 25722 3924 25728 3936
rect 29252 3924 29258 3936
rect 25722 3896 29258 3924
rect 25722 3884 25728 3896
rect 29252 3884 29258 3896
rect 29310 3884 29316 3936
rect 29344 3884 29350 3936
rect 29402 3924 29408 3936
rect 32840 3924 32846 3936
rect 29402 3896 32846 3924
rect 29402 3884 29408 3896
rect 32840 3884 32846 3896
rect 32898 3884 32904 3936
rect 35526 3924 35554 4032
rect 37256 4020 37262 4072
rect 37314 4060 37320 4072
rect 38452 4060 38458 4072
rect 37314 4032 38458 4060
rect 37314 4020 37320 4032
rect 38452 4020 38458 4032
rect 38510 4020 38516 4072
rect 38654 4060 38682 4168
rect 41304 4156 41310 4208
rect 41362 4196 41368 4208
rect 41362 4168 41534 4196
rect 41362 4156 41368 4168
rect 40752 4088 40758 4140
rect 40810 4128 40816 4140
rect 40810 4100 41074 4128
rect 40810 4088 40816 4100
rect 40936 4060 40942 4072
rect 38654 4032 40942 4060
rect 40936 4020 40942 4032
rect 40994 4020 41000 4072
rect 41046 4060 41074 4100
rect 41322 4100 41442 4128
rect 41322 4060 41350 4100
rect 41046 4032 41350 4060
rect 36704 3952 36710 4004
rect 36762 3992 36768 4004
rect 41304 3992 41310 4004
rect 36762 3964 41310 3992
rect 36762 3952 36768 3964
rect 41304 3952 41310 3964
rect 41362 3952 41368 4004
rect 41414 3992 41442 4100
rect 41506 4060 41534 4168
rect 41580 4156 41586 4208
rect 41638 4196 41644 4208
rect 41638 4168 41718 4196
rect 41638 4156 41644 4168
rect 41690 4128 41718 4168
rect 42224 4156 42230 4208
rect 42282 4196 42288 4208
rect 42282 4168 43282 4196
rect 42282 4156 42288 4168
rect 43144 4128 43150 4140
rect 41690 4100 43150 4128
rect 43144 4088 43150 4100
rect 43202 4088 43208 4140
rect 43254 4128 43282 4168
rect 45646 4168 46870 4196
rect 43254 4100 43650 4128
rect 43512 4060 43518 4072
rect 41506 4032 43518 4060
rect 43512 4020 43518 4032
rect 43570 4020 43576 4072
rect 43622 4060 43650 4100
rect 43696 4088 43702 4140
rect 43754 4128 43760 4140
rect 45646 4128 45674 4168
rect 43754 4100 45674 4128
rect 43754 4088 43760 4100
rect 45720 4088 45726 4140
rect 45778 4128 45784 4140
rect 46732 4128 46738 4140
rect 45778 4100 46738 4128
rect 45778 4088 45784 4100
rect 46732 4088 46738 4100
rect 46790 4088 46796 4140
rect 46842 4128 46870 4168
rect 47468 4156 47474 4208
rect 47526 4196 47532 4208
rect 47836 4196 47842 4208
rect 47526 4168 47842 4196
rect 47526 4156 47532 4168
rect 47836 4156 47842 4168
rect 47894 4156 47900 4208
rect 48756 4128 48762 4140
rect 46842 4100 48762 4128
rect 48756 4088 48762 4100
rect 48814 4088 48820 4140
rect 45904 4060 45910 4072
rect 43622 4032 45910 4060
rect 45904 4020 45910 4032
rect 45962 4020 45968 4072
rect 46088 4020 46094 4072
rect 46146 4060 46152 4072
rect 46824 4060 46830 4072
rect 46146 4032 46830 4060
rect 46146 4020 46152 4032
rect 46824 4020 46830 4032
rect 46882 4020 46888 4072
rect 47560 4020 47566 4072
rect 47618 4060 47624 4072
rect 49400 4060 49406 4072
rect 47618 4032 49406 4060
rect 47618 4020 47624 4032
rect 49400 4020 49406 4032
rect 49458 4020 49464 4072
rect 45536 3992 45542 4004
rect 41414 3964 45542 3992
rect 45536 3952 45542 3964
rect 45594 3952 45600 4004
rect 45996 3952 46002 4004
rect 46054 3992 46060 4004
rect 49952 3992 49958 4004
rect 46054 3964 49958 3992
rect 46054 3952 46060 3964
rect 49952 3952 49958 3964
rect 50010 3952 50016 4004
rect 37716 3924 37722 3936
rect 35526 3896 37722 3924
rect 37716 3884 37722 3896
rect 37774 3884 37780 3936
rect 39280 3884 39286 3936
rect 39338 3924 39344 3936
rect 46456 3924 46462 3936
rect 39338 3896 46462 3924
rect 39338 3884 39344 3896
rect 46456 3884 46462 3896
rect 46514 3884 46520 3936
rect 49768 3884 49774 3936
rect 49826 3924 49832 3936
rect 50964 3924 50970 3936
rect 49826 3896 50970 3924
rect 49826 3884 49832 3896
rect 50964 3884 50970 3896
rect 51022 3884 51028 3936
rect 51056 3884 51062 3936
rect 51114 3924 51120 3936
rect 58968 3924 58974 3936
rect 51114 3896 58974 3924
rect 51114 3884 51120 3896
rect 58968 3884 58974 3896
rect 59026 3884 59032 3936
rect 1086 3834 58862 3856
rect 1086 3782 19588 3834
rect 19640 3782 19652 3834
rect 19704 3782 19716 3834
rect 19768 3782 19780 3834
rect 19832 3782 50308 3834
rect 50360 3782 50372 3834
rect 50424 3782 50436 3834
rect 50488 3782 50500 3834
rect 50552 3782 58862 3834
rect 1086 3760 58862 3782
rect 8368 3680 8374 3732
rect 8426 3720 8432 3732
rect 9196 3720 9202 3732
rect 8426 3692 9202 3720
rect 8426 3680 8432 3692
rect 9196 3680 9202 3692
rect 9254 3680 9260 3732
rect 22168 3680 22174 3732
rect 22226 3720 22232 3732
rect 25940 3720 25946 3732
rect 22226 3692 25946 3720
rect 22226 3680 22232 3692
rect 25940 3680 25946 3692
rect 25998 3680 26004 3732
rect 28976 3680 28982 3732
rect 29034 3720 29040 3732
rect 29034 3692 32702 3720
rect 29034 3680 29040 3692
rect 21524 3612 21530 3664
rect 21582 3652 21588 3664
rect 24836 3652 24842 3664
rect 21582 3624 24842 3652
rect 21582 3612 21588 3624
rect 24836 3612 24842 3624
rect 24894 3612 24900 3664
rect 26860 3612 26866 3664
rect 26918 3652 26924 3664
rect 29344 3652 29350 3664
rect 26918 3624 29350 3652
rect 26918 3612 26924 3624
rect 29344 3612 29350 3624
rect 29402 3612 29408 3664
rect 32674 3652 32702 3692
rect 32748 3680 32754 3732
rect 32806 3720 32812 3732
rect 33944 3720 33950 3732
rect 32806 3692 33950 3720
rect 32806 3680 32812 3692
rect 33944 3680 33950 3692
rect 34002 3680 34008 3732
rect 34680 3680 34686 3732
rect 34738 3720 34744 3732
rect 35784 3720 35790 3732
rect 34738 3692 35790 3720
rect 34738 3680 34744 3692
rect 35784 3680 35790 3692
rect 35842 3680 35848 3732
rect 35876 3680 35882 3732
rect 35934 3720 35940 3732
rect 40200 3720 40206 3732
rect 35934 3692 40206 3720
rect 35934 3680 35940 3692
rect 40200 3680 40206 3692
rect 40258 3680 40264 3732
rect 41120 3680 41126 3732
rect 41178 3720 41184 3732
rect 41178 3692 42914 3720
rect 41178 3680 41184 3692
rect 32674 3624 37302 3652
rect 2112 3584 2118 3596
rect 2073 3556 2118 3584
rect 2112 3544 2118 3556
rect 2170 3544 2176 3596
rect 7356 3544 7362 3596
rect 7414 3584 7420 3596
rect 10944 3584 10950 3596
rect 7414 3556 10950 3584
rect 7414 3544 7420 3556
rect 10944 3544 10950 3556
rect 11002 3544 11008 3596
rect 24284 3544 24290 3596
rect 24342 3584 24348 3596
rect 28148 3584 28154 3596
rect 24342 3556 28154 3584
rect 24342 3544 24348 3556
rect 28148 3544 28154 3556
rect 28206 3544 28212 3596
rect 32472 3544 32478 3596
rect 32530 3584 32536 3596
rect 35876 3584 35882 3596
rect 32530 3556 35882 3584
rect 32530 3544 32536 3556
rect 35876 3544 35882 3556
rect 35934 3544 35940 3596
rect 36520 3544 36526 3596
rect 36578 3584 36584 3596
rect 37164 3584 37170 3596
rect 36578 3556 37170 3584
rect 36578 3544 36584 3556
rect 37164 3544 37170 3556
rect 37222 3544 37228 3596
rect 37274 3584 37302 3624
rect 39096 3612 39102 3664
rect 39154 3652 39160 3664
rect 39556 3652 39562 3664
rect 39154 3624 39562 3652
rect 39154 3612 39160 3624
rect 39556 3612 39562 3624
rect 39614 3612 39620 3664
rect 40016 3612 40022 3664
rect 40074 3652 40080 3664
rect 42776 3652 42782 3664
rect 40074 3624 42782 3652
rect 40074 3612 40080 3624
rect 42776 3612 42782 3624
rect 42834 3612 42840 3664
rect 40568 3584 40574 3596
rect 37274 3556 40574 3584
rect 40568 3544 40574 3556
rect 40626 3544 40632 3596
rect 40660 3544 40666 3596
rect 40718 3584 40724 3596
rect 42319 3587 42377 3593
rect 42319 3584 42331 3587
rect 40718 3556 42331 3584
rect 40718 3544 40724 3556
rect 42319 3553 42331 3556
rect 42365 3553 42377 3587
rect 42886 3584 42914 3692
rect 43604 3680 43610 3732
rect 43662 3720 43668 3732
rect 49032 3720 49038 3732
rect 43662 3692 49038 3720
rect 43662 3680 43668 3692
rect 49032 3680 49038 3692
rect 49090 3680 49096 3732
rect 50688 3680 50694 3732
rect 50746 3720 50752 3732
rect 51332 3720 51338 3732
rect 50746 3692 51338 3720
rect 50746 3680 50752 3692
rect 51332 3680 51338 3692
rect 51390 3680 51396 3732
rect 52068 3680 52074 3732
rect 52126 3720 52132 3732
rect 59336 3720 59342 3732
rect 52126 3692 59342 3720
rect 52126 3680 52132 3692
rect 59336 3680 59342 3692
rect 59394 3680 59400 3732
rect 43420 3612 43426 3664
rect 43478 3652 43484 3664
rect 45444 3652 45450 3664
rect 43478 3624 45450 3652
rect 43478 3612 43484 3624
rect 45444 3612 45450 3624
rect 45502 3612 45508 3664
rect 45536 3612 45542 3664
rect 45594 3652 45600 3664
rect 46824 3652 46830 3664
rect 45594 3624 46830 3652
rect 45594 3612 45600 3624
rect 46824 3612 46830 3624
rect 46882 3612 46888 3664
rect 46916 3612 46922 3664
rect 46974 3652 46980 3664
rect 50872 3652 50878 3664
rect 46974 3624 50878 3652
rect 46974 3612 46980 3624
rect 50872 3612 50878 3624
rect 50930 3612 50936 3664
rect 51976 3612 51982 3664
rect 52034 3652 52040 3664
rect 58232 3652 58238 3664
rect 52034 3624 58238 3652
rect 52034 3612 52040 3624
rect 58232 3612 58238 3624
rect 58290 3612 58296 3664
rect 48296 3584 48302 3596
rect 42886 3556 48302 3584
rect 42319 3547 42377 3553
rect 48296 3544 48302 3556
rect 48354 3544 48360 3596
rect 50136 3544 50142 3596
rect 50194 3584 50200 3596
rect 50964 3584 50970 3596
rect 50194 3556 50970 3584
rect 50194 3544 50200 3556
rect 50964 3544 50970 3556
rect 51022 3544 51028 3596
rect 51792 3544 51798 3596
rect 51850 3584 51856 3596
rect 59704 3584 59710 3596
rect 51850 3556 59710 3584
rect 51850 3544 51856 3556
rect 59704 3544 59710 3556
rect 59762 3544 59768 3596
rect 180 3476 186 3528
rect 238 3516 244 3528
rect 1100 3516 1106 3528
rect 238 3488 1106 3516
rect 238 3476 244 3488
rect 1100 3476 1106 3488
rect 1158 3476 1164 3528
rect 1928 3476 1934 3528
rect 1986 3516 1992 3528
rect 2480 3516 2486 3528
rect 1986 3488 2486 3516
rect 1986 3476 1992 3488
rect 2480 3476 2486 3488
rect 2538 3476 2544 3528
rect 8736 3476 8742 3528
rect 8794 3516 8800 3528
rect 9472 3516 9478 3528
rect 8794 3488 9478 3516
rect 8794 3476 8800 3488
rect 9472 3476 9478 3488
rect 9530 3476 9536 3528
rect 14716 3476 14722 3528
rect 14774 3516 14780 3528
rect 26860 3516 26866 3528
rect 14774 3488 26866 3516
rect 14774 3476 14780 3488
rect 26860 3476 26866 3488
rect 26918 3476 26924 3528
rect 31184 3476 31190 3528
rect 31242 3516 31248 3528
rect 36428 3516 36434 3528
rect 31242 3488 36434 3516
rect 31242 3476 31248 3488
rect 36428 3476 36434 3488
rect 36486 3476 36492 3528
rect 37900 3476 37906 3528
rect 37958 3516 37964 3528
rect 41304 3516 41310 3528
rect 37958 3488 41310 3516
rect 37958 3476 37964 3488
rect 41304 3476 41310 3488
rect 41362 3476 41368 3528
rect 41396 3476 41402 3528
rect 41454 3516 41460 3528
rect 47192 3516 47198 3528
rect 41454 3488 47198 3516
rect 41454 3476 41460 3488
rect 47192 3476 47198 3488
rect 47250 3476 47256 3528
rect 50044 3476 50050 3528
rect 50102 3516 50108 3528
rect 52528 3516 52534 3528
rect 50102 3488 52534 3516
rect 50102 3476 50108 3488
rect 52528 3476 52534 3488
rect 52586 3476 52592 3528
rect 53080 3476 53086 3528
rect 53138 3516 53144 3528
rect 53816 3516 53822 3528
rect 53138 3488 53822 3516
rect 53138 3476 53144 3488
rect 53816 3476 53822 3488
rect 53874 3476 53880 3528
rect 53926 3488 55518 3516
rect 916 3408 922 3460
rect 974 3448 980 3460
rect 974 3420 16326 3448
rect 974 3408 980 3420
rect 12508 3380 12514 3392
rect 12469 3352 12514 3380
rect 12508 3340 12514 3352
rect 12566 3340 12572 3392
rect 16298 3380 16326 3420
rect 22812 3408 22818 3460
rect 22870 3448 22876 3460
rect 27044 3448 27050 3460
rect 22870 3420 27050 3448
rect 22870 3408 22876 3420
rect 27044 3408 27050 3420
rect 27102 3408 27108 3460
rect 28516 3408 28522 3460
rect 28574 3448 28580 3460
rect 40108 3448 40114 3460
rect 28574 3420 40114 3448
rect 28574 3408 28580 3420
rect 40108 3408 40114 3420
rect 40166 3408 40172 3460
rect 40200 3408 40206 3460
rect 40258 3448 40264 3460
rect 41672 3448 41678 3460
rect 40258 3420 41678 3448
rect 40258 3408 40264 3420
rect 41672 3408 41678 3420
rect 41730 3408 41736 3460
rect 42702 3420 51654 3448
rect 42702 3380 42730 3420
rect 16298 3352 42730 3380
rect 42776 3340 42782 3392
rect 42834 3380 42840 3392
rect 50596 3380 50602 3392
rect 42834 3352 50602 3380
rect 42834 3340 42840 3352
rect 50596 3340 50602 3352
rect 50654 3340 50660 3392
rect 51626 3380 51654 3420
rect 51700 3408 51706 3460
rect 51758 3448 51764 3460
rect 53926 3448 53954 3488
rect 51758 3420 53954 3448
rect 51758 3408 51764 3420
rect 55291 3383 55349 3389
rect 55291 3380 55303 3383
rect 51626 3352 55303 3380
rect 55291 3349 55303 3352
rect 55337 3349 55349 3383
rect 55490 3380 55518 3488
rect 55840 3476 55846 3528
rect 55898 3516 55904 3528
rect 57864 3516 57870 3528
rect 55898 3488 57870 3516
rect 55898 3476 55904 3488
rect 57864 3476 57870 3488
rect 57922 3476 57928 3528
rect 58600 3380 58606 3392
rect 55490 3352 58606 3380
rect 55291 3343 55349 3349
rect 58600 3340 58606 3352
rect 58658 3340 58664 3392
rect 1086 3290 58862 3312
rect 1086 3238 4228 3290
rect 4280 3238 4292 3290
rect 4344 3238 4356 3290
rect 4408 3238 4420 3290
rect 4472 3238 34948 3290
rect 35000 3238 35012 3290
rect 35064 3238 35076 3290
rect 35128 3238 35140 3290
rect 35192 3238 58862 3290
rect 1086 3216 58862 3238
rect 5332 3136 5338 3188
rect 5390 3176 5396 3188
rect 5390 3148 8722 3176
rect 5390 3136 5396 3148
rect 12508 3136 12514 3188
rect 12566 3176 12572 3188
rect 51608 3176 51614 3188
rect 12566 3148 51614 3176
rect 12566 3136 12572 3148
rect 51608 3136 51614 3148
rect 51666 3136 51672 3188
rect 51884 3136 51890 3188
rect 51942 3176 51948 3188
rect 57496 3176 57502 3188
rect 51942 3148 57502 3176
rect 51942 3136 51948 3148
rect 57496 3136 57502 3148
rect 57554 3136 57560 3188
rect 1376 3068 1382 3120
rect 1434 3108 1440 3120
rect 2572 3108 2578 3120
rect 1434 3080 2578 3108
rect 1434 3068 1440 3080
rect 2572 3068 2578 3080
rect 2630 3068 2636 3120
rect 26860 3068 26866 3120
rect 26918 3108 26924 3120
rect 32472 3108 32478 3120
rect 26918 3080 32478 3108
rect 26918 3068 26924 3080
rect 32472 3068 32478 3080
rect 32530 3068 32536 3120
rect 35232 3068 35238 3120
rect 35290 3108 35296 3120
rect 38084 3108 38090 3120
rect 35290 3080 38090 3108
rect 35290 3068 35296 3080
rect 38084 3068 38090 3080
rect 38142 3068 38148 3120
rect 39372 3068 39378 3120
rect 39430 3108 39436 3120
rect 45352 3108 45358 3120
rect 39430 3080 45358 3108
rect 39430 3068 39436 3080
rect 45352 3068 45358 3080
rect 45410 3068 45416 3120
rect 45444 3068 45450 3120
rect 45502 3108 45508 3120
rect 51240 3108 51246 3120
rect 45502 3080 51246 3108
rect 45502 3068 45508 3080
rect 51240 3068 51246 3080
rect 51298 3068 51304 3120
rect 51332 3068 51338 3120
rect 51390 3108 51396 3120
rect 55656 3108 55662 3120
rect 51390 3080 55662 3108
rect 51390 3068 51396 3080
rect 55656 3068 55662 3080
rect 55714 3068 55720 3120
rect 2664 3000 2670 3052
rect 2722 3040 2728 3052
rect 2722 3012 8262 3040
rect 2722 3000 2728 3012
rect 20512 3000 20518 3052
rect 20570 3040 20576 3052
rect 24468 3040 24474 3052
rect 20570 3012 24474 3040
rect 20570 3000 20576 3012
rect 24468 3000 24474 3012
rect 24526 3000 24532 3052
rect 28424 3000 28430 3052
rect 28482 3040 28488 3052
rect 36152 3040 36158 3052
rect 28482 3012 36158 3040
rect 28482 3000 28488 3012
rect 36152 3000 36158 3012
rect 36210 3000 36216 3052
rect 37992 3000 37998 3052
rect 38050 3040 38056 3052
rect 44616 3040 44622 3052
rect 38050 3012 44622 3040
rect 38050 3000 38056 3012
rect 44616 3000 44622 3012
rect 44674 3000 44680 3052
rect 44800 3000 44806 3052
rect 44858 3040 44864 3052
rect 52344 3040 52350 3052
rect 44858 3012 52350 3040
rect 44858 3000 44864 3012
rect 52344 3000 52350 3012
rect 52402 3000 52408 3052
rect 56024 3040 56030 3052
rect 52454 3012 56030 3040
rect 12416 2932 12422 2984
rect 12474 2972 12480 2984
rect 13520 2972 13526 2984
rect 12474 2944 13526 2972
rect 12474 2932 12480 2944
rect 13520 2932 13526 2944
rect 13578 2932 13584 2984
rect 24192 2932 24198 2984
rect 24250 2972 24256 2984
rect 28884 2972 28890 2984
rect 24250 2944 28890 2972
rect 24250 2932 24256 2944
rect 28884 2932 28890 2944
rect 28942 2932 28948 2984
rect 29620 2932 29626 2984
rect 29678 2972 29684 2984
rect 30264 2972 30270 2984
rect 29678 2944 30270 2972
rect 29678 2932 29684 2944
rect 30264 2932 30270 2944
rect 30322 2932 30328 2984
rect 31092 2932 31098 2984
rect 31150 2972 31156 2984
rect 40200 2972 40206 2984
rect 31150 2944 40206 2972
rect 31150 2932 31156 2944
rect 40200 2932 40206 2944
rect 40258 2932 40264 2984
rect 40844 2932 40850 2984
rect 40902 2972 40908 2984
rect 41396 2972 41402 2984
rect 40902 2944 41402 2972
rect 40902 2932 40908 2944
rect 41396 2932 41402 2944
rect 41454 2932 41460 2984
rect 41488 2932 41494 2984
rect 41546 2972 41552 2984
rect 44984 2972 44990 2984
rect 41546 2944 44990 2972
rect 41546 2932 41552 2944
rect 44984 2932 44990 2944
rect 45042 2932 45048 2984
rect 49676 2972 49682 2984
rect 45094 2944 49682 2972
rect 1284 2796 1290 2848
rect 1342 2836 1348 2848
rect 8432 2836 8460 2924
rect 28608 2864 28614 2916
rect 28666 2904 28672 2916
rect 37992 2904 37998 2916
rect 28666 2876 37998 2904
rect 28666 2864 28672 2876
rect 37992 2864 37998 2876
rect 38050 2864 38056 2916
rect 38084 2864 38090 2916
rect 38142 2904 38148 2916
rect 42040 2904 42046 2916
rect 38142 2876 42046 2904
rect 38142 2864 38148 2876
rect 42040 2864 42046 2876
rect 42098 2864 42104 2916
rect 42132 2864 42138 2916
rect 42190 2904 42196 2916
rect 42190 2876 42914 2904
rect 42190 2864 42196 2876
rect 1342 2808 8460 2836
rect 1342 2796 1348 2808
rect 27412 2796 27418 2848
rect 27470 2836 27476 2848
rect 32380 2836 32386 2848
rect 27470 2808 32386 2836
rect 27470 2796 27476 2808
rect 32380 2796 32386 2808
rect 32438 2796 32444 2848
rect 32656 2796 32662 2848
rect 32714 2836 32720 2848
rect 36336 2836 36342 2848
rect 32714 2808 36342 2836
rect 32714 2796 32720 2808
rect 36336 2796 36342 2808
rect 36394 2796 36400 2848
rect 36428 2796 36434 2848
rect 36486 2836 36492 2848
rect 42776 2836 42782 2848
rect 36486 2808 42782 2836
rect 36486 2796 36492 2808
rect 42776 2796 42782 2808
rect 42834 2796 42840 2848
rect 42886 2836 42914 2876
rect 43880 2864 43886 2916
rect 43938 2904 43944 2916
rect 45094 2904 45122 2944
rect 49676 2932 49682 2944
rect 49734 2932 49740 2984
rect 50780 2932 50786 2984
rect 50838 2972 50844 2984
rect 52454 2972 52482 3012
rect 56024 3000 56030 3012
rect 56082 3000 56088 3052
rect 50838 2944 52482 2972
rect 50838 2932 50844 2944
rect 52528 2932 52534 2984
rect 52586 2972 52592 2984
rect 56760 2972 56766 2984
rect 52586 2944 56766 2972
rect 52586 2932 52592 2944
rect 56760 2932 56766 2944
rect 56818 2932 56824 2984
rect 43938 2876 45122 2904
rect 43938 2864 43944 2876
rect 47928 2864 47934 2916
rect 47986 2904 47992 2916
rect 52436 2904 52442 2916
rect 47986 2876 52442 2904
rect 47986 2864 47992 2876
rect 52436 2864 52442 2876
rect 52494 2864 52500 2916
rect 53172 2864 53178 2916
rect 53230 2904 53236 2916
rect 57128 2904 57134 2916
rect 53230 2876 57134 2904
rect 53230 2864 53236 2876
rect 57128 2864 57134 2876
rect 57186 2864 57192 2916
rect 48664 2836 48670 2848
rect 42886 2808 48670 2836
rect 48664 2796 48670 2808
rect 48722 2796 48728 2848
rect 48756 2796 48762 2848
rect 48814 2836 48820 2848
rect 51976 2836 51982 2848
rect 48814 2808 51982 2836
rect 48814 2796 48820 2808
rect 51976 2796 51982 2808
rect 52034 2796 52040 2848
rect 1086 2746 58862 2768
rect 1086 2694 19588 2746
rect 19640 2694 19652 2746
rect 19704 2694 19716 2746
rect 19768 2694 19780 2746
rect 19832 2694 50308 2746
rect 50360 2694 50372 2746
rect 50424 2694 50436 2746
rect 50488 2694 50500 2746
rect 50552 2694 58862 2746
rect 1086 2672 58862 2694
rect 17384 2592 17390 2644
rect 17442 2632 17448 2644
rect 17844 2632 17850 2644
rect 17442 2604 17850 2632
rect 17442 2592 17448 2604
rect 17844 2592 17850 2604
rect 17902 2592 17908 2644
rect 17936 2592 17942 2644
rect 17994 2632 18000 2644
rect 18396 2632 18402 2644
rect 17994 2604 18402 2632
rect 17994 2592 18000 2604
rect 18396 2592 18402 2604
rect 18454 2592 18460 2644
rect 36612 2592 36618 2644
rect 36670 2632 36676 2644
rect 44248 2632 44254 2644
rect 36670 2604 44254 2632
rect 36670 2592 36676 2604
rect 44248 2592 44254 2604
rect 44306 2592 44312 2644
rect 46272 2592 46278 2644
rect 46330 2632 46336 2644
rect 53448 2632 53454 2644
rect 46330 2604 53454 2632
rect 46330 2592 46336 2604
rect 53448 2592 53454 2604
rect 53506 2592 53512 2644
rect 37716 2524 37722 2576
rect 37774 2564 37780 2576
rect 39372 2564 39378 2576
rect 37774 2536 39378 2564
rect 37774 2524 37780 2536
rect 39372 2524 39378 2536
rect 39430 2524 39436 2576
rect 49400 2524 49406 2576
rect 49458 2564 49464 2576
rect 54184 2564 54190 2576
rect 49458 2536 54190 2564
rect 49458 2524 49464 2536
rect 54184 2524 54190 2536
rect 54242 2524 54248 2576
rect 14903 2295 14961 2301
rect 14903 2261 14915 2295
rect 14949 2292 14961 2295
rect 29988 2292 29994 2304
rect 14949 2264 29994 2292
rect 14949 2261 14961 2264
rect 14903 2255 14961 2261
rect 29988 2252 29994 2264
rect 30046 2252 30052 2304
rect 1086 2202 58862 2224
rect 1086 2150 4228 2202
rect 4280 2150 4292 2202
rect 4344 2150 4356 2202
rect 4408 2150 4420 2202
rect 4472 2150 34948 2202
rect 35000 2150 35012 2202
rect 35064 2150 35076 2202
rect 35128 2150 35140 2202
rect 35192 2150 58862 2202
rect 1086 2128 58862 2150
rect 49952 1980 49958 2032
rect 50010 2020 50016 2032
rect 53080 2020 53086 2032
rect 50010 1992 53086 2020
rect 50010 1980 50016 1992
rect 53080 1980 53086 1992
rect 53138 1980 53144 2032
rect 20788 1504 20794 1556
rect 20846 1544 20852 1556
rect 21340 1544 21346 1556
rect 20846 1516 21346 1544
rect 20846 1504 20852 1516
rect 21340 1504 21346 1516
rect 21398 1504 21404 1556
rect 19684 1096 19690 1148
rect 19742 1136 19748 1148
rect 20880 1136 20886 1148
rect 19742 1108 20886 1136
rect 19742 1096 19748 1108
rect 20880 1096 20886 1108
rect 20938 1096 20944 1148
<< via1 >>
rect 15090 59100 15142 59152
rect 15366 59100 15418 59152
rect 23830 59143 23882 59152
rect 23830 59109 23839 59143
rect 23839 59109 23873 59143
rect 23873 59109 23882 59143
rect 23830 59100 23882 59109
rect 23830 57919 23882 57928
rect 23830 57885 23839 57919
rect 23839 57885 23873 57919
rect 23873 57885 23882 57919
rect 23830 57876 23882 57885
rect 4228 57638 4280 57690
rect 4292 57638 4344 57690
rect 4356 57638 4408 57690
rect 4420 57638 4472 57690
rect 34948 57638 35000 57690
rect 35012 57638 35064 57690
rect 35076 57638 35128 57690
rect 35140 57638 35192 57690
rect 19588 57094 19640 57146
rect 19652 57094 19704 57146
rect 19716 57094 19768 57146
rect 19780 57094 19832 57146
rect 50308 57094 50360 57146
rect 50372 57094 50424 57146
rect 50436 57094 50488 57146
rect 50500 57094 50552 57146
rect 4970 56720 5022 56772
rect 32662 56720 32714 56772
rect 15090 56652 15142 56704
rect 15274 56652 15326 56704
rect 17850 56652 17902 56704
rect 29994 56652 30046 56704
rect 32202 56652 32254 56704
rect 4228 56550 4280 56602
rect 4292 56550 4344 56602
rect 4356 56550 4408 56602
rect 4420 56550 4472 56602
rect 34948 56550 35000 56602
rect 35012 56550 35064 56602
rect 35076 56550 35128 56602
rect 35140 56550 35192 56602
rect 646 56448 698 56500
rect 1106 56448 1158 56500
rect 1750 56448 1802 56500
rect 2670 56448 2722 56500
rect 10306 56448 10358 56500
rect 12790 56448 12842 56500
rect 186 56380 238 56432
rect 1290 56380 1342 56432
rect 1382 56380 1434 56432
rect 2210 56380 2262 56432
rect 2578 56380 2630 56432
rect 21714 56448 21766 56500
rect 24290 56448 24342 56500
rect 29994 56448 30046 56500
rect 1566 56312 1618 56364
rect 17298 56380 17350 56432
rect 21162 56380 21214 56432
rect 21990 56380 22042 56432
rect 22818 56380 22870 56432
rect 28062 56380 28114 56432
rect 28154 56380 28206 56432
rect 30638 56380 30690 56432
rect 31006 56380 31058 56432
rect 33858 56448 33910 56500
rect 16930 56312 16982 56364
rect 24842 56312 24894 56364
rect 24934 56312 24986 56364
rect 29074 56312 29126 56364
rect 29718 56312 29770 56364
rect 32754 56380 32806 56432
rect 33766 56380 33818 56432
rect 35238 56380 35290 56432
rect 40022 56380 40074 56432
rect 40206 56448 40258 56500
rect 41678 56448 41730 56500
rect 44714 56448 44766 56500
rect 48026 56448 48078 56500
rect 48302 56448 48354 56500
rect 49590 56448 49642 56500
rect 40758 56380 40810 56432
rect 40850 56380 40902 56432
rect 45542 56380 45594 56432
rect 46186 56380 46238 56432
rect 51706 56380 51758 56432
rect 31650 56312 31702 56364
rect 38642 56312 38694 56364
rect 49590 56312 49642 56364
rect 53270 56312 53322 56364
rect 3682 56244 3734 56296
rect 35882 56244 35934 56296
rect 35974 56244 36026 56296
rect 40850 56244 40902 56296
rect 40942 56244 40994 56296
rect 46002 56244 46054 56296
rect 57502 56244 57554 56296
rect 10122 56176 10174 56228
rect 13158 56176 13210 56228
rect 14446 56176 14498 56228
rect 20794 56176 20846 56228
rect 20886 56176 20938 56228
rect 11686 56108 11738 56160
rect 16838 56108 16890 56160
rect 17114 56108 17166 56160
rect 41310 56108 41362 56160
rect 41402 56108 41454 56160
rect 45358 56108 45410 56160
rect 45542 56176 45594 56228
rect 48578 56108 48630 56160
rect 49130 56176 49182 56228
rect 52718 56176 52770 56228
rect 54834 56108 54886 56160
rect 19588 56006 19640 56058
rect 19652 56006 19704 56058
rect 19716 56006 19768 56058
rect 19780 56006 19832 56058
rect 50308 56006 50360 56058
rect 50372 56006 50424 56058
rect 50436 56006 50488 56058
rect 50500 56006 50552 56058
rect 4050 55904 4102 55956
rect 17758 55904 17810 55956
rect 41218 55904 41270 55956
rect 41310 55904 41362 55956
rect 44714 55904 44766 55956
rect 46002 55904 46054 55956
rect 59066 55904 59118 55956
rect 31742 55836 31794 55888
rect 31834 55836 31886 55888
rect 35422 55836 35474 55888
rect 36158 55836 36210 55888
rect 40666 55836 40718 55888
rect 40758 55836 40810 55888
rect 42230 55836 42282 55888
rect 42322 55836 42374 55888
rect 46094 55836 46146 55888
rect 46186 55836 46238 55888
rect 55938 55836 55990 55888
rect 6350 55768 6402 55820
rect 16930 55768 16982 55820
rect 11410 55700 11462 55752
rect 17114 55700 17166 55752
rect 1842 55632 1894 55684
rect 2578 55632 2630 55684
rect 8190 55632 8242 55684
rect 17574 55768 17626 55820
rect 17666 55768 17718 55820
rect 22726 55768 22778 55820
rect 22910 55768 22962 55820
rect 24934 55768 24986 55820
rect 25670 55768 25722 55820
rect 17298 55700 17350 55752
rect 24382 55700 24434 55752
rect 17390 55632 17442 55684
rect 20886 55632 20938 55684
rect 21346 55632 21398 55684
rect 25946 55700 25998 55752
rect 26130 55768 26182 55820
rect 28154 55768 28206 55820
rect 28338 55768 28390 55820
rect 51154 55768 51206 55820
rect 41402 55700 41454 55752
rect 41494 55700 41546 55752
rect 49130 55700 49182 55752
rect 25210 55632 25262 55684
rect 34318 55632 34370 55684
rect 35330 55632 35382 55684
rect 59618 55632 59670 55684
rect 30454 55564 30506 55616
rect 31742 55564 31794 55616
rect 36158 55564 36210 55616
rect 39654 55564 39706 55616
rect 42046 55564 42098 55616
rect 42138 55564 42190 55616
rect 43794 55564 43846 55616
rect 43886 55564 43938 55616
rect 48302 55564 48354 55616
rect 4228 55462 4280 55514
rect 4292 55462 4344 55514
rect 4356 55462 4408 55514
rect 4420 55462 4472 55514
rect 34948 55462 35000 55514
rect 35012 55462 35064 55514
rect 35076 55462 35128 55514
rect 35140 55462 35192 55514
rect 4878 55360 4930 55412
rect 7454 55360 7506 55412
rect 9846 55360 9898 55412
rect 6994 55292 7046 55344
rect 7914 55292 7966 55344
rect 8282 55292 8334 55344
rect 9570 55292 9622 55344
rect 13066 55292 13118 55344
rect 17114 55292 17166 55344
rect 2762 55224 2814 55276
rect 3774 55224 3826 55276
rect 4602 55224 4654 55276
rect 7546 55224 7598 55276
rect 8098 55224 8150 55276
rect 13250 55224 13302 55276
rect 13710 55224 13762 55276
rect 17574 55360 17626 55412
rect 18034 55292 18086 55344
rect 19230 55292 19282 55344
rect 19874 55292 19926 55344
rect 20610 55292 20662 55344
rect 20794 55360 20846 55412
rect 23278 55360 23330 55412
rect 31282 55360 31334 55412
rect 24106 55292 24158 55344
rect 26406 55292 26458 55344
rect 27050 55292 27102 55344
rect 35238 55360 35290 55412
rect 35422 55360 35474 55412
rect 40758 55360 40810 55412
rect 41678 55360 41730 55412
rect 54374 55360 54426 55412
rect 38550 55292 38602 55344
rect 40666 55292 40718 55344
rect 41034 55292 41086 55344
rect 56398 55292 56450 55344
rect 25210 55224 25262 55276
rect 25578 55224 25630 55276
rect 24198 55156 24250 55208
rect 26130 55156 26182 55208
rect 32202 55156 32254 55208
rect 41678 55156 41730 55208
rect 43242 55224 43294 55276
rect 44070 55224 44122 55276
rect 44898 55156 44950 55208
rect 5338 55020 5390 55072
rect 19588 54918 19640 54970
rect 19652 54918 19704 54970
rect 19716 54918 19768 54970
rect 19780 54918 19832 54970
rect 50308 54918 50360 54970
rect 50372 54918 50424 54970
rect 50436 54918 50488 54970
rect 50500 54918 50552 54970
rect 16838 54816 16890 54868
rect 8558 54748 8610 54800
rect 21438 54680 21490 54732
rect 27602 54680 27654 54732
rect 38642 54680 38694 54732
rect 19138 54612 19190 54664
rect 17390 54519 17442 54528
rect 17390 54485 17399 54519
rect 17399 54485 17433 54519
rect 17433 54485 17442 54519
rect 17390 54476 17442 54485
rect 19138 54476 19190 54528
rect 21438 54476 21490 54528
rect 21622 54519 21674 54528
rect 21622 54485 21631 54519
rect 21631 54485 21665 54519
rect 21665 54485 21674 54519
rect 21622 54476 21674 54485
rect 27602 54476 27654 54528
rect 38642 54476 38694 54528
rect 42414 54519 42466 54528
rect 42414 54485 42423 54519
rect 42423 54485 42457 54519
rect 42457 54485 42466 54519
rect 42414 54476 42466 54485
rect 4228 54374 4280 54426
rect 4292 54374 4344 54426
rect 4356 54374 4408 54426
rect 4420 54374 4472 54426
rect 34948 54374 35000 54426
rect 35012 54374 35064 54426
rect 35076 54374 35128 54426
rect 35140 54374 35192 54426
rect 17390 54272 17442 54324
rect 50602 54272 50654 54324
rect 14814 54204 14866 54256
rect 42414 54204 42466 54256
rect 21622 54136 21674 54188
rect 43426 54136 43478 54188
rect 47566 54068 47618 54120
rect 19588 53830 19640 53882
rect 19652 53830 19704 53882
rect 19716 53830 19768 53882
rect 19780 53830 19832 53882
rect 50308 53830 50360 53882
rect 50372 53830 50424 53882
rect 50436 53830 50488 53882
rect 50500 53830 50552 53882
rect 58054 53592 58106 53644
rect 4228 53286 4280 53338
rect 4292 53286 4344 53338
rect 4356 53286 4408 53338
rect 4420 53286 4472 53338
rect 34948 53286 35000 53338
rect 35012 53286 35064 53338
rect 35076 53286 35128 53338
rect 35140 53286 35192 53338
rect 17022 53227 17074 53236
rect 17022 53193 17031 53227
rect 17031 53193 17065 53227
rect 17065 53193 17074 53227
rect 17022 53184 17074 53193
rect 15274 53116 15326 53168
rect 15734 53116 15786 53168
rect 26498 53116 26550 53168
rect 26958 53116 27010 53168
rect 15274 52980 15326 53032
rect 15918 52980 15970 53032
rect 18586 52980 18638 53032
rect 33030 52912 33082 52964
rect 19588 52742 19640 52794
rect 19652 52742 19704 52794
rect 19716 52742 19768 52794
rect 19780 52742 19832 52794
rect 50308 52742 50360 52794
rect 50372 52742 50424 52794
rect 50436 52742 50488 52794
rect 50500 52742 50552 52794
rect 20334 52300 20386 52352
rect 4228 52198 4280 52250
rect 4292 52198 4344 52250
rect 4356 52198 4408 52250
rect 4420 52198 4472 52250
rect 34948 52198 35000 52250
rect 35012 52198 35064 52250
rect 35076 52198 35128 52250
rect 35140 52198 35192 52250
rect 30454 51892 30506 51944
rect 32386 51892 32438 51944
rect 38550 51892 38602 51944
rect 19588 51654 19640 51706
rect 19652 51654 19704 51706
rect 19716 51654 19768 51706
rect 19780 51654 19832 51706
rect 50308 51654 50360 51706
rect 50372 51654 50424 51706
rect 50436 51654 50488 51706
rect 50500 51654 50552 51706
rect 48394 51484 48446 51536
rect 49038 51484 49090 51536
rect 35238 51212 35290 51264
rect 4228 51110 4280 51162
rect 4292 51110 4344 51162
rect 4356 51110 4408 51162
rect 4420 51110 4472 51162
rect 34948 51110 35000 51162
rect 35012 51110 35064 51162
rect 35076 51110 35128 51162
rect 35140 51110 35192 51162
rect 1382 50668 1434 50720
rect 19588 50566 19640 50618
rect 19652 50566 19704 50618
rect 19716 50566 19768 50618
rect 19780 50566 19832 50618
rect 50308 50566 50360 50618
rect 50372 50566 50424 50618
rect 50436 50566 50488 50618
rect 50500 50566 50552 50618
rect 42046 50124 42098 50176
rect 4228 50022 4280 50074
rect 4292 50022 4344 50074
rect 4356 50022 4408 50074
rect 4420 50022 4472 50074
rect 34948 50022 35000 50074
rect 35012 50022 35064 50074
rect 35076 50022 35128 50074
rect 35140 50022 35192 50074
rect 19588 49478 19640 49530
rect 19652 49478 19704 49530
rect 19716 49478 19768 49530
rect 19780 49478 19832 49530
rect 50308 49478 50360 49530
rect 50372 49478 50424 49530
rect 50436 49478 50488 49530
rect 50500 49478 50552 49530
rect 18310 49308 18362 49360
rect 19046 49308 19098 49360
rect 12330 49036 12382 49088
rect 39286 49036 39338 49088
rect 4228 48934 4280 48986
rect 4292 48934 4344 48986
rect 4356 48934 4408 48986
rect 4420 48934 4472 48986
rect 34948 48934 35000 48986
rect 35012 48934 35064 48986
rect 35076 48934 35128 48986
rect 35140 48934 35192 48986
rect 8006 48628 8058 48680
rect 53086 48628 53138 48680
rect 19588 48390 19640 48442
rect 19652 48390 19704 48442
rect 19716 48390 19768 48442
rect 19780 48390 19832 48442
rect 50308 48390 50360 48442
rect 50372 48390 50424 48442
rect 50436 48390 50488 48442
rect 50500 48390 50552 48442
rect 29350 48288 29402 48340
rect 30178 48288 30230 48340
rect 31650 48288 31702 48340
rect 32662 48288 32714 48340
rect 39102 48288 39154 48340
rect 39470 48288 39522 48340
rect 6718 47948 6770 48000
rect 4228 47846 4280 47898
rect 4292 47846 4344 47898
rect 4356 47846 4408 47898
rect 4420 47846 4472 47898
rect 34948 47846 35000 47898
rect 35012 47846 35064 47898
rect 35076 47846 35128 47898
rect 35140 47846 35192 47898
rect 19414 47608 19466 47660
rect 3866 47540 3918 47592
rect 24198 47404 24250 47456
rect 44070 47404 44122 47456
rect 19588 47302 19640 47354
rect 19652 47302 19704 47354
rect 19716 47302 19768 47354
rect 19780 47302 19832 47354
rect 50308 47302 50360 47354
rect 50372 47302 50424 47354
rect 50436 47302 50488 47354
rect 50500 47302 50552 47354
rect 8650 47132 8702 47184
rect 9110 47132 9162 47184
rect 24750 46928 24802 46980
rect 26406 46860 26458 46912
rect 26498 46860 26550 46912
rect 29350 46860 29402 46912
rect 29534 46860 29586 46912
rect 48302 46860 48354 46912
rect 48394 46860 48446 46912
rect 4228 46758 4280 46810
rect 4292 46758 4344 46810
rect 4356 46758 4408 46810
rect 4420 46758 4472 46810
rect 34948 46758 35000 46810
rect 35012 46758 35064 46810
rect 35076 46758 35128 46810
rect 35140 46758 35192 46810
rect 46830 46452 46882 46504
rect 50694 46384 50746 46436
rect 19588 46214 19640 46266
rect 19652 46214 19704 46266
rect 19716 46214 19768 46266
rect 19780 46214 19832 46266
rect 50308 46214 50360 46266
rect 50372 46214 50424 46266
rect 50436 46214 50488 46266
rect 50500 46214 50552 46266
rect 4228 45670 4280 45722
rect 4292 45670 4344 45722
rect 4356 45670 4408 45722
rect 4420 45670 4472 45722
rect 34948 45670 35000 45722
rect 35012 45670 35064 45722
rect 35076 45670 35128 45722
rect 35140 45670 35192 45722
rect 34318 45568 34370 45620
rect 34778 45568 34830 45620
rect 8926 45500 8978 45552
rect 9110 45500 9162 45552
rect 14170 45500 14222 45552
rect 14446 45500 14498 45552
rect 39838 45364 39890 45416
rect 19588 45126 19640 45178
rect 19652 45126 19704 45178
rect 19716 45126 19768 45178
rect 19780 45126 19832 45178
rect 50308 45126 50360 45178
rect 50372 45126 50424 45178
rect 50436 45126 50488 45178
rect 50500 45126 50552 45178
rect 16838 45067 16890 45076
rect 16838 45033 16847 45067
rect 16847 45033 16881 45067
rect 16881 45033 16890 45067
rect 16838 45024 16890 45033
rect 2302 44727 2354 44736
rect 2302 44693 2311 44727
rect 2311 44693 2345 44727
rect 2345 44693 2354 44727
rect 2302 44684 2354 44693
rect 26866 44684 26918 44736
rect 37170 44684 37222 44736
rect 50970 44684 51022 44736
rect 56950 44727 57002 44736
rect 56950 44693 56959 44727
rect 56959 44693 56993 44727
rect 56993 44693 57002 44727
rect 56950 44684 57002 44693
rect 4228 44582 4280 44634
rect 4292 44582 4344 44634
rect 4356 44582 4408 44634
rect 4420 44582 4472 44634
rect 34948 44582 35000 44634
rect 35012 44582 35064 44634
rect 35076 44582 35128 44634
rect 35140 44582 35192 44634
rect 23370 44480 23422 44532
rect 56950 44480 57002 44532
rect 2302 44412 2354 44464
rect 39378 44412 39430 44464
rect 19588 44038 19640 44090
rect 19652 44038 19704 44090
rect 19716 44038 19768 44090
rect 19780 44038 19832 44090
rect 50308 44038 50360 44090
rect 50372 44038 50424 44090
rect 50436 44038 50488 44090
rect 50500 44038 50552 44090
rect 4228 43494 4280 43546
rect 4292 43494 4344 43546
rect 4356 43494 4408 43546
rect 4420 43494 4472 43546
rect 34948 43494 35000 43546
rect 35012 43494 35064 43546
rect 35076 43494 35128 43546
rect 35140 43494 35192 43546
rect 40114 43435 40166 43444
rect 40114 43401 40123 43435
rect 40123 43401 40157 43435
rect 40157 43401 40166 43435
rect 40114 43392 40166 43401
rect 2578 43188 2630 43240
rect 40758 43120 40810 43172
rect 19588 42950 19640 43002
rect 19652 42950 19704 43002
rect 19716 42950 19768 43002
rect 19780 42950 19832 43002
rect 50308 42950 50360 43002
rect 50372 42950 50424 43002
rect 50436 42950 50488 43002
rect 50500 42950 50552 43002
rect 16470 42644 16522 42696
rect 4228 42406 4280 42458
rect 4292 42406 4344 42458
rect 4356 42406 4408 42458
rect 4420 42406 4472 42458
rect 34948 42406 35000 42458
rect 35012 42406 35064 42458
rect 35076 42406 35128 42458
rect 35140 42406 35192 42458
rect 42138 42304 42190 42356
rect 13618 42236 13670 42288
rect 17206 42100 17258 42152
rect 31006 42168 31058 42220
rect 37906 42032 37958 42084
rect 3866 41964 3918 42016
rect 19588 41862 19640 41914
rect 19652 41862 19704 41914
rect 19716 41862 19768 41914
rect 19780 41862 19832 41914
rect 50308 41862 50360 41914
rect 50372 41862 50424 41914
rect 50436 41862 50488 41914
rect 50500 41862 50552 41914
rect 17206 41760 17258 41812
rect 27050 41760 27102 41812
rect 13802 41624 13854 41676
rect 43518 41420 43570 41472
rect 4228 41318 4280 41370
rect 4292 41318 4344 41370
rect 4356 41318 4408 41370
rect 4420 41318 4472 41370
rect 34948 41318 35000 41370
rect 35012 41318 35064 41370
rect 35076 41318 35128 41370
rect 35140 41318 35192 41370
rect 38826 41080 38878 41132
rect 39102 41080 39154 41132
rect 43150 41012 43202 41064
rect 50878 41012 50930 41064
rect 19588 40774 19640 40826
rect 19652 40774 19704 40826
rect 19716 40774 19768 40826
rect 19780 40774 19832 40826
rect 50308 40774 50360 40826
rect 50372 40774 50424 40826
rect 50436 40774 50488 40826
rect 50500 40774 50552 40826
rect 3682 40400 3734 40452
rect 11870 40375 11922 40384
rect 11870 40341 11879 40375
rect 11879 40341 11913 40375
rect 11913 40341 11922 40375
rect 11870 40332 11922 40341
rect 4228 40230 4280 40282
rect 4292 40230 4344 40282
rect 4356 40230 4408 40282
rect 4420 40230 4472 40282
rect 34948 40230 35000 40282
rect 35012 40230 35064 40282
rect 35076 40230 35128 40282
rect 35140 40230 35192 40282
rect 11870 40128 11922 40180
rect 24198 40128 24250 40180
rect 38458 40128 38510 40180
rect 23278 40060 23330 40112
rect 26958 40035 27010 40044
rect 26958 40001 26967 40035
rect 26967 40001 27001 40035
rect 27001 40001 27010 40035
rect 26958 39992 27010 40001
rect 19588 39686 19640 39738
rect 19652 39686 19704 39738
rect 19716 39686 19768 39738
rect 19780 39686 19832 39738
rect 50308 39686 50360 39738
rect 50372 39686 50424 39738
rect 50436 39686 50488 39738
rect 50500 39686 50552 39738
rect 42138 39244 42190 39296
rect 4228 39142 4280 39194
rect 4292 39142 4344 39194
rect 4356 39142 4408 39194
rect 4420 39142 4472 39194
rect 34948 39142 35000 39194
rect 35012 39142 35064 39194
rect 35076 39142 35128 39194
rect 35140 39142 35192 39194
rect 1842 39083 1894 39092
rect 1842 39049 1851 39083
rect 1851 39049 1885 39083
rect 1885 39049 1894 39083
rect 1842 39040 1894 39049
rect 4786 38904 4838 38956
rect 16286 38836 16338 38888
rect 19588 38598 19640 38650
rect 19652 38598 19704 38650
rect 19716 38598 19768 38650
rect 19780 38598 19832 38650
rect 50308 38598 50360 38650
rect 50372 38598 50424 38650
rect 50436 38598 50488 38650
rect 50500 38598 50552 38650
rect 28246 38156 28298 38208
rect 47842 38199 47894 38208
rect 47842 38165 47851 38199
rect 47851 38165 47885 38199
rect 47885 38165 47894 38199
rect 47842 38156 47894 38165
rect 4228 38054 4280 38106
rect 4292 38054 4344 38106
rect 4356 38054 4408 38106
rect 4420 38054 4472 38106
rect 34948 38054 35000 38106
rect 35012 38054 35064 38106
rect 35076 38054 35128 38106
rect 35140 38054 35192 38106
rect 49498 37748 49550 37800
rect 21898 37680 21950 37732
rect 8558 37612 8610 37664
rect 19588 37510 19640 37562
rect 19652 37510 19704 37562
rect 19716 37510 19768 37562
rect 19780 37510 19832 37562
rect 50308 37510 50360 37562
rect 50372 37510 50424 37562
rect 50436 37510 50488 37562
rect 50500 37510 50552 37562
rect 3498 37272 3550 37324
rect 4786 37272 4838 37324
rect 12054 37272 12106 37324
rect 19138 37272 19190 37324
rect 26406 37272 26458 37324
rect 26498 37272 26550 37324
rect 27510 37272 27562 37324
rect 48302 37272 48354 37324
rect 48394 37272 48446 37324
rect 49774 37272 49826 37324
rect 49866 37272 49918 37324
rect 27786 37204 27838 37256
rect 12974 37111 13026 37120
rect 12974 37077 12983 37111
rect 12983 37077 13017 37111
rect 13017 37077 13026 37111
rect 12974 37068 13026 37077
rect 26682 37111 26734 37120
rect 26682 37077 26691 37111
rect 26691 37077 26725 37111
rect 26725 37077 26734 37111
rect 26682 37068 26734 37077
rect 29258 37111 29310 37120
rect 29258 37077 29267 37111
rect 29267 37077 29301 37111
rect 29301 37077 29310 37111
rect 29258 37068 29310 37077
rect 31098 37111 31150 37120
rect 31098 37077 31107 37111
rect 31107 37077 31141 37111
rect 31141 37077 31150 37111
rect 31098 37068 31150 37077
rect 47842 37204 47894 37256
rect 48026 37204 48078 37256
rect 42782 37136 42834 37188
rect 43150 37136 43202 37188
rect 4228 36966 4280 37018
rect 4292 36966 4344 37018
rect 4356 36966 4408 37018
rect 4420 36966 4472 37018
rect 34948 36966 35000 37018
rect 35012 36966 35064 37018
rect 35076 36966 35128 37018
rect 35140 36966 35192 37018
rect 14998 36864 15050 36916
rect 26682 36864 26734 36916
rect 29258 36864 29310 36916
rect 46278 36864 46330 36916
rect 37078 36660 37130 36712
rect 50786 36592 50838 36644
rect 19588 36422 19640 36474
rect 19652 36422 19704 36474
rect 19716 36422 19768 36474
rect 19780 36422 19832 36474
rect 50308 36422 50360 36474
rect 50372 36422 50424 36474
rect 50436 36422 50488 36474
rect 50500 36422 50552 36474
rect 13526 35980 13578 36032
rect 4228 35878 4280 35930
rect 4292 35878 4344 35930
rect 4356 35878 4408 35930
rect 4420 35878 4472 35930
rect 34948 35878 35000 35930
rect 35012 35878 35064 35930
rect 35076 35878 35128 35930
rect 35140 35878 35192 35930
rect 12238 35572 12290 35624
rect 19588 35334 19640 35386
rect 19652 35334 19704 35386
rect 19716 35334 19768 35386
rect 19780 35334 19832 35386
rect 50308 35334 50360 35386
rect 50372 35334 50424 35386
rect 50436 35334 50488 35386
rect 50500 35334 50552 35386
rect 32570 35096 32622 35148
rect 52902 34935 52954 34944
rect 52902 34901 52911 34935
rect 52911 34901 52945 34935
rect 52945 34901 52954 34935
rect 52902 34892 52954 34901
rect 4228 34790 4280 34842
rect 4292 34790 4344 34842
rect 4356 34790 4408 34842
rect 4420 34790 4472 34842
rect 34948 34790 35000 34842
rect 35012 34790 35064 34842
rect 35076 34790 35128 34842
rect 35140 34790 35192 34842
rect 2486 34688 2538 34740
rect 52902 34688 52954 34740
rect 25578 34620 25630 34672
rect 10858 34552 10910 34604
rect 19588 34246 19640 34298
rect 19652 34246 19704 34298
rect 19716 34246 19768 34298
rect 19780 34246 19832 34298
rect 50308 34246 50360 34298
rect 50372 34246 50424 34298
rect 50436 34246 50488 34298
rect 50500 34246 50552 34298
rect 21806 33804 21858 33856
rect 43610 33847 43662 33856
rect 43610 33813 43619 33847
rect 43619 33813 43653 33847
rect 43653 33813 43662 33847
rect 43610 33804 43662 33813
rect 58422 33847 58474 33856
rect 58422 33813 58431 33847
rect 58431 33813 58465 33847
rect 58465 33813 58474 33847
rect 58422 33804 58474 33813
rect 4228 33702 4280 33754
rect 4292 33702 4344 33754
rect 4356 33702 4408 33754
rect 4420 33702 4472 33754
rect 34948 33702 35000 33754
rect 35012 33702 35064 33754
rect 35076 33702 35128 33754
rect 35140 33702 35192 33754
rect 35790 33600 35842 33652
rect 43610 33600 43662 33652
rect 32938 33532 32990 33584
rect 58422 33532 58474 33584
rect 22818 33464 22870 33516
rect 2394 33396 2446 33448
rect 19588 33158 19640 33210
rect 19652 33158 19704 33210
rect 19716 33158 19768 33210
rect 19780 33158 19832 33210
rect 50308 33158 50360 33210
rect 50372 33158 50424 33210
rect 50436 33158 50488 33210
rect 50500 33158 50552 33210
rect 50142 32716 50194 32768
rect 4228 32614 4280 32666
rect 4292 32614 4344 32666
rect 4356 32614 4408 32666
rect 4420 32614 4472 32666
rect 34948 32614 35000 32666
rect 35012 32614 35064 32666
rect 35076 32614 35128 32666
rect 35140 32614 35192 32666
rect 39838 32376 39890 32428
rect 14538 32308 14590 32360
rect 54006 32308 54058 32360
rect 19588 32070 19640 32122
rect 19652 32070 19704 32122
rect 19716 32070 19768 32122
rect 19780 32070 19832 32122
rect 50308 32070 50360 32122
rect 50372 32070 50424 32122
rect 50436 32070 50488 32122
rect 50500 32070 50552 32122
rect 37998 31968 38050 32020
rect 10766 31900 10818 31952
rect 31558 31900 31610 31952
rect 9294 31832 9346 31884
rect 24290 31764 24342 31816
rect 40850 31764 40902 31816
rect 23462 31696 23514 31748
rect 23646 31696 23698 31748
rect 4228 31526 4280 31578
rect 4292 31526 4344 31578
rect 4356 31526 4408 31578
rect 4420 31526 4472 31578
rect 34948 31526 35000 31578
rect 35012 31526 35064 31578
rect 35076 31526 35128 31578
rect 35140 31526 35192 31578
rect 8742 31220 8794 31272
rect 36526 31220 36578 31272
rect 17206 31152 17258 31204
rect 5246 31084 5298 31136
rect 5430 31084 5482 31136
rect 8834 31084 8886 31136
rect 9018 31084 9070 31136
rect 25578 31084 25630 31136
rect 19588 30982 19640 31034
rect 19652 30982 19704 31034
rect 19716 30982 19768 31034
rect 19780 30982 19832 31034
rect 50308 30982 50360 31034
rect 50372 30982 50424 31034
rect 50436 30982 50488 31034
rect 50500 30982 50552 31034
rect 17206 30880 17258 30932
rect 28798 30880 28850 30932
rect 8742 30812 8794 30864
rect 28706 30812 28758 30864
rect 22726 30744 22778 30796
rect 7362 30583 7414 30592
rect 7362 30549 7371 30583
rect 7371 30549 7405 30583
rect 7405 30549 7414 30583
rect 7362 30540 7414 30549
rect 21162 30540 21214 30592
rect 4228 30438 4280 30490
rect 4292 30438 4344 30490
rect 4356 30438 4408 30490
rect 4420 30438 4472 30490
rect 34948 30438 35000 30490
rect 35012 30438 35064 30490
rect 35076 30438 35128 30490
rect 35140 30438 35192 30490
rect 25670 30268 25722 30320
rect 14906 30200 14958 30252
rect 8466 30132 8518 30184
rect 12146 30132 12198 30184
rect 12882 30064 12934 30116
rect 8834 29996 8886 30048
rect 9018 29996 9070 30048
rect 16010 30039 16062 30048
rect 16010 30005 16019 30039
rect 16019 30005 16053 30039
rect 16053 30005 16062 30039
rect 16010 29996 16062 30005
rect 26130 30064 26182 30116
rect 24290 29996 24342 30048
rect 19588 29894 19640 29946
rect 19652 29894 19704 29946
rect 19716 29894 19768 29946
rect 19780 29894 19832 29946
rect 50308 29894 50360 29946
rect 50372 29894 50424 29946
rect 50436 29894 50488 29946
rect 50500 29894 50552 29946
rect 12882 29792 12934 29844
rect 27234 29792 27286 29844
rect 1106 29724 1158 29776
rect 16010 29724 16062 29776
rect 8466 29656 8518 29708
rect 27602 29656 27654 29708
rect 26682 29495 26734 29504
rect 26682 29461 26691 29495
rect 26691 29461 26725 29495
rect 26725 29461 26734 29495
rect 26682 29452 26734 29461
rect 48946 29452 48998 29504
rect 4228 29350 4280 29402
rect 4292 29350 4344 29402
rect 4356 29350 4408 29402
rect 4420 29350 4472 29402
rect 34948 29350 35000 29402
rect 35012 29350 35064 29402
rect 35076 29350 35128 29402
rect 35140 29350 35192 29402
rect 3498 29044 3550 29096
rect 3590 29010 3642 29062
rect 8558 29112 8610 29164
rect 25118 29248 25170 29300
rect 26682 29248 26734 29300
rect 51706 29248 51758 29300
rect 34318 29112 34370 29164
rect 27326 29044 27378 29096
rect 7822 28976 7874 29028
rect 15550 28976 15602 29028
rect 15642 28976 15694 29028
rect 34410 28976 34462 29028
rect 22726 28908 22778 28960
rect 19588 28806 19640 28858
rect 19652 28806 19704 28858
rect 19716 28806 19768 28858
rect 19780 28806 19832 28858
rect 50308 28806 50360 28858
rect 50372 28806 50424 28858
rect 50436 28806 50488 28858
rect 50500 28806 50552 28858
rect 3774 28611 3826 28620
rect 3774 28577 3783 28611
rect 3783 28577 3817 28611
rect 3817 28577 3826 28611
rect 3774 28568 3826 28577
rect 36802 28364 36854 28416
rect 4228 28262 4280 28314
rect 4292 28262 4344 28314
rect 4356 28262 4408 28314
rect 4420 28262 4472 28314
rect 34948 28262 35000 28314
rect 35012 28262 35064 28314
rect 35076 28262 35128 28314
rect 35140 28262 35192 28314
rect 28062 28160 28114 28212
rect 28246 28160 28298 28212
rect 8558 28024 8610 28076
rect 8926 28024 8978 28076
rect 25394 28024 25446 28076
rect 8834 27956 8886 28008
rect 25854 27956 25906 28008
rect 8558 27820 8610 27872
rect 21438 27820 21490 27872
rect 19588 27718 19640 27770
rect 19652 27718 19704 27770
rect 19716 27718 19768 27770
rect 19780 27718 19832 27770
rect 50308 27718 50360 27770
rect 50372 27718 50424 27770
rect 50436 27718 50488 27770
rect 50500 27718 50552 27770
rect 5338 27616 5390 27668
rect 28062 27616 28114 27668
rect 28154 27616 28206 27668
rect 34502 27616 34554 27668
rect 34778 27616 34830 27668
rect 38734 27616 38786 27668
rect 38826 27616 38878 27668
rect 47842 27616 47894 27668
rect 48026 27616 48078 27668
rect 3406 27548 3458 27600
rect 3590 27548 3642 27600
rect 14814 27548 14866 27600
rect 14906 27548 14958 27600
rect 18218 27548 18270 27600
rect 18310 27548 18362 27600
rect 26498 27548 26550 27600
rect 26590 27548 26642 27600
rect 5338 27412 5390 27464
rect 17206 27276 17258 27328
rect 4228 27174 4280 27226
rect 4292 27174 4344 27226
rect 4356 27174 4408 27226
rect 4420 27174 4472 27226
rect 34948 27174 35000 27226
rect 35012 27174 35064 27226
rect 35076 27174 35128 27226
rect 35140 27174 35192 27226
rect 7638 26936 7690 26988
rect 7914 26936 7966 26988
rect 8558 26936 8610 26988
rect 8834 26936 8886 26988
rect 23646 26936 23698 26988
rect 8466 26868 8518 26920
rect 8926 26868 8978 26920
rect 24382 26868 24434 26920
rect 46738 26868 46790 26920
rect 55846 26868 55898 26920
rect 21530 26732 21582 26784
rect 19588 26630 19640 26682
rect 19652 26630 19704 26682
rect 19716 26630 19768 26682
rect 19780 26630 19832 26682
rect 50308 26630 50360 26682
rect 50372 26630 50424 26682
rect 50436 26630 50488 26682
rect 50500 26630 50552 26682
rect 5522 26392 5574 26444
rect 36986 26392 37038 26444
rect 50050 26392 50102 26444
rect 20610 26324 20662 26376
rect 6626 26256 6678 26308
rect 25670 26188 25722 26240
rect 25762 26188 25814 26240
rect 39746 26188 39798 26240
rect 39930 26188 39982 26240
rect 4228 26086 4280 26138
rect 4292 26086 4344 26138
rect 4356 26086 4408 26138
rect 4420 26086 4472 26138
rect 34948 26086 35000 26138
rect 35012 26086 35064 26138
rect 35076 26086 35128 26138
rect 35140 26086 35192 26138
rect 8558 25984 8610 26036
rect 11410 26027 11462 26036
rect 11410 25993 11419 26027
rect 11419 25993 11453 26027
rect 11453 25993 11462 26027
rect 11410 25984 11462 25993
rect 8558 25848 8610 25900
rect 7730 25780 7782 25832
rect 35698 25780 35750 25832
rect 8926 25712 8978 25764
rect 22910 25712 22962 25764
rect 8696 25644 8748 25696
rect 8834 25644 8886 25696
rect 22542 25644 22594 25696
rect 19588 25542 19640 25594
rect 19652 25542 19704 25594
rect 19716 25542 19768 25594
rect 19780 25542 19832 25594
rect 50308 25542 50360 25594
rect 50372 25542 50424 25594
rect 50436 25542 50488 25594
rect 50500 25542 50552 25594
rect 8696 25440 8748 25492
rect 20058 25440 20110 25492
rect 7730 25372 7782 25424
rect 32570 25372 32622 25424
rect 8282 25100 8334 25152
rect 12422 25100 12474 25152
rect 4228 24998 4280 25050
rect 4292 24998 4344 25050
rect 4356 24998 4408 25050
rect 4420 24998 4472 25050
rect 34948 24998 35000 25050
rect 35012 24998 35064 25050
rect 35076 24998 35128 25050
rect 35140 24998 35192 25050
rect 8282 24896 8334 24948
rect 12422 24896 12474 24948
rect 19966 24896 20018 24948
rect 1566 24760 1618 24812
rect 8604 24760 8656 24812
rect 8926 24760 8978 24812
rect 10214 24760 10266 24812
rect 21070 24760 21122 24812
rect 8466 24624 8518 24676
rect 22082 24692 22134 24744
rect 21714 24624 21766 24676
rect 10214 24556 10266 24608
rect 19588 24454 19640 24506
rect 19652 24454 19704 24506
rect 19716 24454 19768 24506
rect 19780 24454 19832 24506
rect 50308 24454 50360 24506
rect 50372 24454 50424 24506
rect 50436 24454 50488 24506
rect 50500 24454 50552 24506
rect 8466 24352 8518 24404
rect 20794 24352 20846 24404
rect 9846 24259 9898 24268
rect 9846 24225 9855 24259
rect 9855 24225 9889 24259
rect 9889 24225 9898 24259
rect 9846 24216 9898 24225
rect 51062 24148 51114 24200
rect 3774 24080 3826 24132
rect 34226 24080 34278 24132
rect 16470 24012 16522 24064
rect 31558 24012 31610 24064
rect 51062 24012 51114 24064
rect 4228 23910 4280 23962
rect 4292 23910 4344 23962
rect 4356 23910 4408 23962
rect 4420 23910 4472 23962
rect 34948 23910 35000 23962
rect 35012 23910 35064 23962
rect 35076 23910 35128 23962
rect 35140 23910 35192 23962
rect 8650 23808 8702 23860
rect 8834 23808 8886 23860
rect 18586 23808 18638 23860
rect 34226 23808 34278 23860
rect 8604 23706 8656 23758
rect 9478 23740 9530 23792
rect 8742 23672 8794 23724
rect 20426 23672 20478 23724
rect 8466 23604 8518 23656
rect 8834 23604 8886 23656
rect 19874 23604 19926 23656
rect 8466 23468 8518 23520
rect 11778 23468 11830 23520
rect 20242 23468 20294 23520
rect 30270 23536 30322 23588
rect 19588 23366 19640 23418
rect 19652 23366 19704 23418
rect 19716 23366 19768 23418
rect 19780 23366 19832 23418
rect 50308 23366 50360 23418
rect 50372 23366 50424 23418
rect 50436 23366 50488 23418
rect 50500 23366 50552 23418
rect 9662 22924 9714 22976
rect 20610 22924 20662 22976
rect 4228 22822 4280 22874
rect 4292 22822 4344 22874
rect 4356 22822 4408 22874
rect 4420 22822 4472 22874
rect 34948 22822 35000 22874
rect 35012 22822 35064 22874
rect 35076 22822 35128 22874
rect 35140 22822 35192 22874
rect 18678 22720 18730 22772
rect 18034 22584 18086 22636
rect 18770 22516 18822 22568
rect 41494 22559 41546 22568
rect 41494 22525 41503 22559
rect 41503 22525 41537 22559
rect 41537 22525 41546 22559
rect 41494 22516 41546 22525
rect 18126 22380 18178 22432
rect 19588 22278 19640 22330
rect 19652 22278 19704 22330
rect 19716 22278 19768 22330
rect 19780 22278 19832 22330
rect 50308 22278 50360 22330
rect 50372 22278 50424 22330
rect 50436 22278 50488 22330
rect 50500 22278 50552 22330
rect 9662 22176 9714 22228
rect 28430 22176 28482 22228
rect 35422 22040 35474 22092
rect 9386 21836 9438 21888
rect 4228 21734 4280 21786
rect 4292 21734 4344 21786
rect 4356 21734 4408 21786
rect 4420 21734 4472 21786
rect 34948 21734 35000 21786
rect 35012 21734 35064 21786
rect 35076 21734 35128 21786
rect 35140 21734 35192 21786
rect 17298 21496 17350 21548
rect 16930 21428 16982 21480
rect 8466 21292 8518 21344
rect 8650 21292 8702 21344
rect 17390 21292 17442 21344
rect 19588 21190 19640 21242
rect 19652 21190 19704 21242
rect 19716 21190 19768 21242
rect 19780 21190 19832 21242
rect 50308 21190 50360 21242
rect 50372 21190 50424 21242
rect 50436 21190 50488 21242
rect 50500 21190 50552 21242
rect 28338 20952 28390 21004
rect 7730 20884 7782 20936
rect 43610 20816 43662 20868
rect 4228 20646 4280 20698
rect 4292 20646 4344 20698
rect 4356 20646 4408 20698
rect 4420 20646 4472 20698
rect 34948 20646 35000 20698
rect 35012 20646 35064 20698
rect 35076 20646 35128 20698
rect 35140 20646 35192 20698
rect 4050 20587 4102 20596
rect 4050 20553 4059 20587
rect 4059 20553 4093 20587
rect 4093 20553 4102 20587
rect 4050 20544 4102 20553
rect 8466 20544 8518 20596
rect 8650 20544 8702 20596
rect 16838 20544 16890 20596
rect 51798 20408 51850 20460
rect 15550 20340 15602 20392
rect 28614 20383 28666 20392
rect 28614 20349 28623 20383
rect 28623 20349 28657 20383
rect 28657 20349 28666 20383
rect 28614 20340 28666 20349
rect 8282 20204 8334 20256
rect 15826 20272 15878 20324
rect 38366 20272 38418 20324
rect 11410 20204 11462 20256
rect 14630 20204 14682 20256
rect 19588 20102 19640 20154
rect 19652 20102 19704 20154
rect 19716 20102 19768 20154
rect 19780 20102 19832 20154
rect 50308 20102 50360 20154
rect 50372 20102 50424 20154
rect 50436 20102 50488 20154
rect 50500 20102 50552 20154
rect 8282 20000 8334 20052
rect 11410 20000 11462 20052
rect 5154 19932 5206 19984
rect 28614 20000 28666 20052
rect 39562 20043 39614 20052
rect 39562 20009 39571 20043
rect 39571 20009 39605 20043
rect 39605 20009 39614 20043
rect 39562 20000 39614 20009
rect 49590 19907 49642 19916
rect 49590 19873 49599 19907
rect 49599 19873 49633 19907
rect 49633 19873 49642 19907
rect 49590 19864 49642 19873
rect 8466 19660 8518 19712
rect 15918 19660 15970 19712
rect 16378 19660 16430 19712
rect 4228 19558 4280 19610
rect 4292 19558 4344 19610
rect 4356 19558 4408 19610
rect 4420 19558 4472 19610
rect 34948 19558 35000 19610
rect 35012 19558 35064 19610
rect 35076 19558 35128 19610
rect 35140 19558 35192 19610
rect 8466 19456 8518 19508
rect 34778 19388 34830 19440
rect 7454 19252 7506 19304
rect 7822 19286 7874 19338
rect 21346 19320 21398 19372
rect 29258 19320 29310 19372
rect 29350 19320 29402 19372
rect 32662 19320 32714 19372
rect 34594 19320 34646 19372
rect 8006 19252 8058 19304
rect 13158 19295 13210 19304
rect 8420 19218 8472 19270
rect 13158 19261 13167 19295
rect 13167 19261 13201 19295
rect 13201 19261 13210 19295
rect 13158 19252 13210 19261
rect 20978 19252 21030 19304
rect 21070 19252 21122 19304
rect 22910 19252 22962 19304
rect 23094 19252 23146 19304
rect 23646 19252 23698 19304
rect 23922 19252 23974 19304
rect 36894 19252 36946 19304
rect 37078 19252 37130 19304
rect 48394 19252 48446 19304
rect 52074 19252 52126 19304
rect 56674 19252 56726 19304
rect 8926 19116 8978 19168
rect 13158 19116 13210 19168
rect 48394 19116 48446 19168
rect 19588 19014 19640 19066
rect 19652 19014 19704 19066
rect 19716 19014 19768 19066
rect 19780 19014 19832 19066
rect 50308 19014 50360 19066
rect 50372 19014 50424 19066
rect 50436 19014 50488 19066
rect 50500 19014 50552 19066
rect 8466 18912 8518 18964
rect 13342 18912 13394 18964
rect 7638 18640 7690 18692
rect 26774 18640 26826 18692
rect 8650 18572 8702 18624
rect 12790 18572 12842 18624
rect 28338 18572 28390 18624
rect 4228 18470 4280 18522
rect 4292 18470 4344 18522
rect 4356 18470 4408 18522
rect 4420 18470 4472 18522
rect 34948 18470 35000 18522
rect 35012 18470 35064 18522
rect 35076 18470 35128 18522
rect 35140 18470 35192 18522
rect 8834 18368 8886 18420
rect 9018 18368 9070 18420
rect 14170 18368 14222 18420
rect 8650 18232 8702 18284
rect 26774 18232 26826 18284
rect 12606 18164 12658 18216
rect 23186 18164 23238 18216
rect 12882 18028 12934 18080
rect 23462 18028 23514 18080
rect 23554 18028 23606 18080
rect 19588 17926 19640 17978
rect 19652 17926 19704 17978
rect 19716 17926 19768 17978
rect 19780 17926 19832 17978
rect 50308 17926 50360 17978
rect 50372 17926 50424 17978
rect 50436 17926 50488 17978
rect 50500 17926 50552 17978
rect 8834 17620 8886 17672
rect 52074 17620 52126 17672
rect 8742 17552 8794 17604
rect 55386 17552 55438 17604
rect 5062 17484 5114 17536
rect 4228 17382 4280 17434
rect 4292 17382 4344 17434
rect 4356 17382 4408 17434
rect 4420 17382 4472 17434
rect 34948 17382 35000 17434
rect 35012 17382 35064 17434
rect 35076 17382 35128 17434
rect 35140 17382 35192 17434
rect 8834 17280 8886 17332
rect 9110 17246 9162 17298
rect 9570 17212 9622 17264
rect 35330 17212 35382 17264
rect 8006 17076 8058 17128
rect 8742 17076 8794 17128
rect 19588 16838 19640 16890
rect 19652 16838 19704 16890
rect 19716 16838 19768 16890
rect 19780 16838 19832 16890
rect 50308 16838 50360 16890
rect 50372 16838 50424 16890
rect 50436 16838 50488 16890
rect 50500 16838 50552 16890
rect 8006 16736 8058 16788
rect 51890 16736 51942 16788
rect 25762 16600 25814 16652
rect 25946 16600 25998 16652
rect 39654 16600 39706 16652
rect 39930 16600 39982 16652
rect 8650 16396 8702 16448
rect 51062 16396 51114 16448
rect 4228 16294 4280 16346
rect 4292 16294 4344 16346
rect 4356 16294 4408 16346
rect 4420 16294 4472 16346
rect 34948 16294 35000 16346
rect 35012 16294 35064 16346
rect 35076 16294 35128 16346
rect 35140 16294 35192 16346
rect 8742 16192 8794 16244
rect 8650 16074 8702 16126
rect 16654 16031 16706 16040
rect 16654 15997 16663 16031
rect 16663 15997 16697 16031
rect 16697 15997 16706 16031
rect 16654 15988 16706 15997
rect 8742 15852 8794 15904
rect 33858 15852 33910 15904
rect 19588 15750 19640 15802
rect 19652 15750 19704 15802
rect 19716 15750 19768 15802
rect 19780 15750 19832 15802
rect 50308 15750 50360 15802
rect 50372 15750 50424 15802
rect 50436 15750 50488 15802
rect 50500 15750 50552 15802
rect 1106 15648 1158 15700
rect 16654 15648 16706 15700
rect 44806 15308 44858 15360
rect 4228 15206 4280 15258
rect 4292 15206 4344 15258
rect 4356 15206 4408 15258
rect 4420 15206 4472 15258
rect 34948 15206 35000 15258
rect 35012 15206 35064 15258
rect 35076 15206 35128 15258
rect 35140 15206 35192 15258
rect 8466 15104 8518 15156
rect 8650 15104 8702 15156
rect 25486 15104 25538 15156
rect 8650 14968 8702 15020
rect 8282 14866 8334 14918
rect 27142 14943 27194 14952
rect 27142 14909 27151 14943
rect 27151 14909 27185 14943
rect 27185 14909 27194 14943
rect 27142 14900 27194 14909
rect 48394 14900 48446 14952
rect 29718 14832 29770 14884
rect 31466 14832 31518 14884
rect 19588 14662 19640 14714
rect 19652 14662 19704 14714
rect 19716 14662 19768 14714
rect 19780 14662 19832 14714
rect 50308 14662 50360 14714
rect 50372 14662 50424 14714
rect 50436 14662 50488 14714
rect 50500 14662 50552 14714
rect 5246 14492 5298 14544
rect 5430 14492 5482 14544
rect 16838 14492 16890 14544
rect 17022 14492 17074 14544
rect 4228 14118 4280 14170
rect 4292 14118 4344 14170
rect 4356 14118 4408 14170
rect 4420 14118 4472 14170
rect 34948 14118 35000 14170
rect 35012 14118 35064 14170
rect 35076 14118 35128 14170
rect 35140 14118 35192 14170
rect 8834 14016 8886 14068
rect 32202 14059 32254 14068
rect 32202 14025 32211 14059
rect 32211 14025 32245 14059
rect 32245 14025 32254 14059
rect 32202 14016 32254 14025
rect 45726 13948 45778 14000
rect 8006 13880 8058 13932
rect 13066 13880 13118 13932
rect 13434 13880 13486 13932
rect 20150 13812 20202 13864
rect 19588 13574 19640 13626
rect 19652 13574 19704 13626
rect 19716 13574 19768 13626
rect 19780 13574 19832 13626
rect 50308 13574 50360 13626
rect 50372 13574 50424 13626
rect 50436 13574 50488 13626
rect 50500 13574 50552 13626
rect 6534 13379 6586 13388
rect 6534 13345 6543 13379
rect 6543 13345 6577 13379
rect 6577 13345 6586 13379
rect 6534 13336 6586 13345
rect 4228 13030 4280 13082
rect 4292 13030 4344 13082
rect 4356 13030 4408 13082
rect 4420 13030 4472 13082
rect 34948 13030 35000 13082
rect 35012 13030 35064 13082
rect 35076 13030 35128 13082
rect 35140 13030 35192 13082
rect 8144 12928 8196 12980
rect 18954 12860 19006 12912
rect 42966 12792 43018 12844
rect 8926 12724 8978 12776
rect 51982 12724 52034 12776
rect 21990 12588 22042 12640
rect 19588 12486 19640 12538
rect 19652 12486 19704 12538
rect 19716 12486 19768 12538
rect 19780 12486 19832 12538
rect 50308 12486 50360 12538
rect 50372 12486 50424 12538
rect 50436 12486 50488 12538
rect 50500 12486 50552 12538
rect 5798 12044 5850 12096
rect 47198 12087 47250 12096
rect 47198 12053 47207 12087
rect 47207 12053 47241 12087
rect 47241 12053 47250 12087
rect 47198 12044 47250 12053
rect 4228 11942 4280 11994
rect 4292 11942 4344 11994
rect 4356 11942 4408 11994
rect 4420 11942 4472 11994
rect 34948 11942 35000 11994
rect 35012 11942 35064 11994
rect 35076 11942 35128 11994
rect 35140 11942 35192 11994
rect 35330 11840 35382 11892
rect 47198 11840 47250 11892
rect 8236 11602 8288 11654
rect 8466 11636 8518 11688
rect 38734 11636 38786 11688
rect 33766 11500 33818 11552
rect 19588 11398 19640 11450
rect 19652 11398 19704 11450
rect 19716 11398 19768 11450
rect 19780 11398 19832 11450
rect 50308 11398 50360 11450
rect 50372 11398 50424 11450
rect 50436 11398 50488 11450
rect 50500 11398 50552 11450
rect 9202 11160 9254 11212
rect 9386 11160 9438 11212
rect 31190 11135 31242 11144
rect 31190 11101 31199 11135
rect 31199 11101 31233 11135
rect 31233 11101 31242 11135
rect 31190 11092 31242 11101
rect 9294 10956 9346 11008
rect 33306 10956 33358 11008
rect 4228 10854 4280 10906
rect 4292 10854 4344 10906
rect 4356 10854 4408 10906
rect 4420 10854 4472 10906
rect 34948 10854 35000 10906
rect 35012 10854 35064 10906
rect 35076 10854 35128 10906
rect 35140 10854 35192 10906
rect 38642 10752 38694 10804
rect 13250 10548 13302 10600
rect 52074 10548 52126 10600
rect 9294 10480 9346 10532
rect 37262 10412 37314 10464
rect 19588 10310 19640 10362
rect 19652 10310 19704 10362
rect 19716 10310 19768 10362
rect 19780 10310 19832 10362
rect 50308 10310 50360 10362
rect 50372 10310 50424 10362
rect 50436 10310 50488 10362
rect 50500 10310 50552 10362
rect 13250 10208 13302 10260
rect 34594 10208 34646 10260
rect 32846 9936 32898 9988
rect 32754 9868 32806 9920
rect 4228 9766 4280 9818
rect 4292 9766 4344 9818
rect 4356 9766 4408 9818
rect 4420 9766 4472 9818
rect 34948 9766 35000 9818
rect 35012 9766 35064 9818
rect 35076 9766 35128 9818
rect 35140 9766 35192 9818
rect 3222 9664 3274 9716
rect 3498 9664 3550 9716
rect 7454 9664 7506 9716
rect 7822 9664 7874 9716
rect 36894 9664 36946 9716
rect 37078 9664 37130 9716
rect 8374 9426 8426 9478
rect 41126 9460 41178 9512
rect 43518 9503 43570 9512
rect 43518 9469 43527 9503
rect 43527 9469 43561 9503
rect 43561 9469 43570 9503
rect 43518 9460 43570 9469
rect 47474 9503 47526 9512
rect 47474 9469 47483 9503
rect 47483 9469 47517 9503
rect 47517 9469 47526 9503
rect 47474 9460 47526 9469
rect 54926 9460 54978 9512
rect 29626 9392 29678 9444
rect 13710 9324 13762 9376
rect 19588 9222 19640 9274
rect 19652 9222 19704 9274
rect 19716 9222 19768 9274
rect 19780 9222 19832 9274
rect 50308 9222 50360 9274
rect 50372 9222 50424 9274
rect 50436 9222 50488 9274
rect 50500 9222 50552 9274
rect 19230 9120 19282 9172
rect 25210 9120 25262 9172
rect 43518 9120 43570 9172
rect 3958 9052 4010 9104
rect 47474 9052 47526 9104
rect 8374 8984 8426 9036
rect 29258 8984 29310 9036
rect 5246 8780 5298 8832
rect 39746 8780 39798 8832
rect 49682 8780 49734 8832
rect 4228 8678 4280 8730
rect 4292 8678 4344 8730
rect 4356 8678 4408 8730
rect 4420 8678 4472 8730
rect 34948 8678 35000 8730
rect 35012 8678 35064 8730
rect 35076 8678 35128 8730
rect 35140 8678 35192 8730
rect 39746 8619 39798 8628
rect 8834 8508 8886 8560
rect 39746 8585 39755 8619
rect 39755 8585 39789 8619
rect 39789 8585 39798 8619
rect 39746 8576 39798 8585
rect 26590 8508 26642 8560
rect 48302 8508 48354 8560
rect 27418 8440 27470 8492
rect 27510 8440 27562 8492
rect 29074 8440 29126 8492
rect 8558 8372 8610 8424
rect 10582 8372 10634 8424
rect 48210 8372 48262 8424
rect 20150 8304 20202 8356
rect 20518 8304 20570 8356
rect 25670 8304 25722 8356
rect 25946 8304 25998 8356
rect 20058 8236 20110 8288
rect 23738 8236 23790 8288
rect 28154 8236 28206 8288
rect 35422 8236 35474 8288
rect 19588 8134 19640 8186
rect 19652 8134 19704 8186
rect 19716 8134 19768 8186
rect 19780 8134 19832 8186
rect 50308 8134 50360 8186
rect 50372 8134 50424 8186
rect 50436 8134 50488 8186
rect 50500 8134 50552 8186
rect 14538 7896 14590 7948
rect 14722 7896 14774 7948
rect 17942 7760 17994 7812
rect 18126 7760 18178 7812
rect 26682 7760 26734 7812
rect 24842 7692 24894 7744
rect 25026 7692 25078 7744
rect 25854 7692 25906 7744
rect 26498 7692 26550 7744
rect 27326 7692 27378 7744
rect 28338 7692 28390 7744
rect 28798 7692 28850 7744
rect 41586 7735 41638 7744
rect 41586 7701 41595 7735
rect 41595 7701 41629 7735
rect 41629 7701 41638 7735
rect 41586 7692 41638 7701
rect 4228 7590 4280 7642
rect 4292 7590 4344 7642
rect 4356 7590 4408 7642
rect 4420 7590 4472 7642
rect 34948 7590 35000 7642
rect 35012 7590 35064 7642
rect 35076 7590 35128 7642
rect 35140 7590 35192 7642
rect 12606 7488 12658 7540
rect 13342 7488 13394 7540
rect 15550 7488 15602 7540
rect 16194 7488 16246 7540
rect 17574 7531 17626 7540
rect 17574 7497 17583 7531
rect 17583 7497 17617 7531
rect 17617 7497 17626 7531
rect 17574 7488 17626 7497
rect 19966 7488 20018 7540
rect 20426 7488 20478 7540
rect 20886 7488 20938 7540
rect 41586 7488 41638 7540
rect 49774 7488 49826 7540
rect 12790 7420 12842 7472
rect 13710 7420 13762 7472
rect 15274 7420 15326 7472
rect 15918 7420 15970 7472
rect 12698 7352 12750 7404
rect 23462 7352 23514 7404
rect 8236 7250 8288 7302
rect 9110 7284 9162 7336
rect 28890 7284 28942 7336
rect 53178 7284 53230 7336
rect 28982 7216 29034 7268
rect 46002 7216 46054 7268
rect 24106 7148 24158 7200
rect 19588 7046 19640 7098
rect 19652 7046 19704 7098
rect 19716 7046 19768 7098
rect 19780 7046 19832 7098
rect 50308 7046 50360 7098
rect 50372 7046 50424 7098
rect 50436 7046 50488 7098
rect 50500 7046 50552 7098
rect 39654 6944 39706 6996
rect 39562 6876 39614 6928
rect 8098 6808 8150 6860
rect 15182 6808 15234 6860
rect 8006 6740 8058 6792
rect 17206 6672 17258 6724
rect 8466 6604 8518 6656
rect 16562 6604 16614 6656
rect 46922 6740 46974 6792
rect 27694 6604 27746 6656
rect 38826 6604 38878 6656
rect 46922 6604 46974 6656
rect 52442 6647 52494 6656
rect 52442 6613 52451 6647
rect 52451 6613 52485 6647
rect 52485 6613 52494 6647
rect 52442 6604 52494 6613
rect 4228 6502 4280 6554
rect 4292 6502 4344 6554
rect 4356 6502 4408 6554
rect 4420 6502 4472 6554
rect 34948 6502 35000 6554
rect 35012 6502 35064 6554
rect 35076 6502 35128 6554
rect 35140 6502 35192 6554
rect 8466 6400 8518 6452
rect 17482 6400 17534 6452
rect 36986 6400 37038 6452
rect 38642 6400 38694 6452
rect 52442 6400 52494 6452
rect 21346 6332 21398 6384
rect 27694 6332 27746 6384
rect 38826 6332 38878 6384
rect 8098 6264 8150 6316
rect 18310 6264 18362 6316
rect 36986 6264 37038 6316
rect 38642 6264 38694 6316
rect 38734 6264 38786 6316
rect 14538 6196 14590 6248
rect 40114 6196 40166 6248
rect 51062 6128 51114 6180
rect 14446 6060 14498 6112
rect 19588 5958 19640 6010
rect 19652 5958 19704 6010
rect 19716 5958 19768 6010
rect 19780 5958 19832 6010
rect 50308 5958 50360 6010
rect 50372 5958 50424 6010
rect 50436 5958 50488 6010
rect 50500 5958 50552 6010
rect 17206 5856 17258 5908
rect 40022 5856 40074 5908
rect 5430 5788 5482 5840
rect 28982 5788 29034 5840
rect 10950 5720 11002 5772
rect 32478 5720 32530 5772
rect 1198 5516 1250 5568
rect 4228 5414 4280 5466
rect 4292 5414 4344 5466
rect 4356 5414 4408 5466
rect 4420 5414 4472 5466
rect 34948 5414 35000 5466
rect 35012 5414 35064 5466
rect 35076 5414 35128 5466
rect 35140 5414 35192 5466
rect 8374 5312 8426 5364
rect 10306 5312 10358 5364
rect 11042 5176 11094 5228
rect 46186 5219 46238 5228
rect 46186 5185 46195 5219
rect 46195 5185 46229 5219
rect 46229 5185 46238 5219
rect 46186 5176 46238 5185
rect 8742 5108 8794 5160
rect 15642 5108 15694 5160
rect 32386 5108 32438 5160
rect 52442 5108 52494 5160
rect 8650 4972 8702 5024
rect 20058 4972 20110 5024
rect 22634 4972 22686 5024
rect 50142 4972 50194 5024
rect 55294 4972 55346 5024
rect 19588 4870 19640 4922
rect 19652 4870 19704 4922
rect 19716 4870 19768 4922
rect 19780 4870 19832 4922
rect 50308 4870 50360 4922
rect 50372 4870 50424 4922
rect 50436 4870 50488 4922
rect 50500 4870 50552 4922
rect 20058 4768 20110 4820
rect 20334 4768 20386 4820
rect 32846 4768 32898 4820
rect 33122 4768 33174 4820
rect 48946 4768 48998 4820
rect 52718 4768 52770 4820
rect 17114 4700 17166 4752
rect 18586 4700 18638 4752
rect 6902 4632 6954 4684
rect 9018 4632 9070 4684
rect 13066 4564 13118 4616
rect 14814 4564 14866 4616
rect 4228 4326 4280 4378
rect 4292 4326 4344 4378
rect 4356 4326 4408 4378
rect 4420 4326 4472 4378
rect 34948 4326 35000 4378
rect 35012 4326 35064 4378
rect 35076 4326 35128 4378
rect 35140 4326 35192 4378
rect 16746 4224 16798 4276
rect 17022 4224 17074 4276
rect 20426 4224 20478 4276
rect 32570 4224 32622 4276
rect 3682 4088 3734 4140
rect 3958 4088 4010 4140
rect 6166 4088 6218 4140
rect 6718 4088 6770 4140
rect 7270 4088 7322 4140
rect 7730 4088 7782 4140
rect 8926 4088 8978 4140
rect 10214 4088 10266 4140
rect 10766 4088 10818 4140
rect 11686 4088 11738 4140
rect 12330 4088 12382 4140
rect 12974 4088 13026 4140
rect 13434 4088 13486 4140
rect 14630 4088 14682 4140
rect 15458 4088 15510 4140
rect 16010 4088 16062 4140
rect 16470 4088 16522 4140
rect 17114 4088 17166 4140
rect 17850 4088 17902 4140
rect 18678 4088 18730 4140
rect 19322 4088 19374 4140
rect 21438 4088 21490 4140
rect 22174 4088 22226 4140
rect 22266 4088 22318 4140
rect 23002 4088 23054 4140
rect 23278 4088 23330 4140
rect 23370 4088 23422 4140
rect 24106 4088 24158 4140
rect 24750 4088 24802 4140
rect 25578 4088 25630 4140
rect 26130 4088 26182 4140
rect 27142 4088 27194 4140
rect 27786 4088 27838 4140
rect 29718 4088 29770 4140
rect 31006 4088 31058 4140
rect 31466 4088 31518 4140
rect 32110 4088 32162 4140
rect 32938 4088 32990 4140
rect 2854 4020 2906 4072
rect 3866 4020 3918 4072
rect 4602 4020 4654 4072
rect 5062 4020 5114 4072
rect 6810 4020 6862 4072
rect 9846 4020 9898 4072
rect 10858 4020 10910 4072
rect 11318 4020 11370 4072
rect 12146 4020 12198 4072
rect 13066 4020 13118 4072
rect 13618 4020 13670 4072
rect 13802 4020 13854 4072
rect 14998 4020 15050 4072
rect 15642 4020 15694 4072
rect 16378 4020 16430 4072
rect 24842 4020 24894 4072
rect 26314 4020 26366 4072
rect 27050 4020 27102 4072
rect 30086 4020 30138 4072
rect 30638 4020 30690 4072
rect 31558 4020 31610 4072
rect 31742 4020 31794 4072
rect 33030 4020 33082 4072
rect 33582 4088 33634 4140
rect 34410 4088 34462 4140
rect 50602 4224 50654 4276
rect 56398 4224 56450 4276
rect 37630 4088 37682 4140
rect 38550 4088 38602 4140
rect 5062 3884 5114 3936
rect 5246 3884 5298 3936
rect 7546 3884 7598 3936
rect 12790 3952 12842 4004
rect 13250 3952 13302 4004
rect 18494 3952 18546 4004
rect 20702 3952 20754 4004
rect 21162 3952 21214 4004
rect 21806 3952 21858 4004
rect 25118 3952 25170 4004
rect 26130 3952 26182 4004
rect 13158 3884 13210 3936
rect 14446 3884 14498 3936
rect 18126 3884 18178 3936
rect 20426 3884 20478 3936
rect 25670 3884 25722 3936
rect 29258 3884 29310 3936
rect 29350 3884 29402 3936
rect 32846 3884 32898 3936
rect 37262 4020 37314 4072
rect 38458 4020 38510 4072
rect 41310 4156 41362 4208
rect 40758 4088 40810 4140
rect 40942 4020 40994 4072
rect 36710 3952 36762 4004
rect 41310 3952 41362 4004
rect 41586 4156 41638 4208
rect 42230 4156 42282 4208
rect 43150 4088 43202 4140
rect 43518 4020 43570 4072
rect 43702 4088 43754 4140
rect 45726 4088 45778 4140
rect 46738 4088 46790 4140
rect 47474 4156 47526 4208
rect 47842 4156 47894 4208
rect 48762 4088 48814 4140
rect 45910 4020 45962 4072
rect 46094 4020 46146 4072
rect 46830 4020 46882 4072
rect 47566 4020 47618 4072
rect 49406 4020 49458 4072
rect 45542 3952 45594 4004
rect 46002 3952 46054 4004
rect 49958 3952 50010 4004
rect 37722 3884 37774 3936
rect 39286 3884 39338 3936
rect 46462 3884 46514 3936
rect 49774 3884 49826 3936
rect 50970 3884 51022 3936
rect 51062 3884 51114 3936
rect 58974 3884 59026 3936
rect 19588 3782 19640 3834
rect 19652 3782 19704 3834
rect 19716 3782 19768 3834
rect 19780 3782 19832 3834
rect 50308 3782 50360 3834
rect 50372 3782 50424 3834
rect 50436 3782 50488 3834
rect 50500 3782 50552 3834
rect 8374 3680 8426 3732
rect 9202 3680 9254 3732
rect 22174 3680 22226 3732
rect 25946 3680 25998 3732
rect 28982 3680 29034 3732
rect 21530 3612 21582 3664
rect 24842 3612 24894 3664
rect 26866 3612 26918 3664
rect 29350 3612 29402 3664
rect 32754 3680 32806 3732
rect 33950 3680 34002 3732
rect 34686 3680 34738 3732
rect 35790 3680 35842 3732
rect 35882 3680 35934 3732
rect 40206 3680 40258 3732
rect 41126 3680 41178 3732
rect 2118 3587 2170 3596
rect 2118 3553 2127 3587
rect 2127 3553 2161 3587
rect 2161 3553 2170 3587
rect 2118 3544 2170 3553
rect 7362 3544 7414 3596
rect 10950 3544 11002 3596
rect 24290 3544 24342 3596
rect 28154 3544 28206 3596
rect 32478 3544 32530 3596
rect 35882 3544 35934 3596
rect 36526 3544 36578 3596
rect 37170 3544 37222 3596
rect 39102 3612 39154 3664
rect 39562 3612 39614 3664
rect 40022 3612 40074 3664
rect 42782 3612 42834 3664
rect 40574 3544 40626 3596
rect 40666 3544 40718 3596
rect 43610 3680 43662 3732
rect 49038 3680 49090 3732
rect 50694 3680 50746 3732
rect 51338 3680 51390 3732
rect 52074 3680 52126 3732
rect 59342 3680 59394 3732
rect 43426 3612 43478 3664
rect 45450 3612 45502 3664
rect 45542 3612 45594 3664
rect 46830 3612 46882 3664
rect 46922 3612 46974 3664
rect 50878 3612 50930 3664
rect 51982 3612 52034 3664
rect 58238 3612 58290 3664
rect 48302 3544 48354 3596
rect 50142 3544 50194 3596
rect 50970 3544 51022 3596
rect 51798 3544 51850 3596
rect 59710 3544 59762 3596
rect 186 3476 238 3528
rect 1106 3476 1158 3528
rect 1934 3476 1986 3528
rect 2486 3476 2538 3528
rect 8742 3476 8794 3528
rect 9478 3476 9530 3528
rect 14722 3476 14774 3528
rect 26866 3476 26918 3528
rect 31190 3476 31242 3528
rect 36434 3476 36486 3528
rect 37906 3476 37958 3528
rect 41310 3476 41362 3528
rect 41402 3476 41454 3528
rect 47198 3476 47250 3528
rect 50050 3476 50102 3528
rect 52534 3476 52586 3528
rect 53086 3476 53138 3528
rect 53822 3476 53874 3528
rect 922 3408 974 3460
rect 12514 3383 12566 3392
rect 12514 3349 12523 3383
rect 12523 3349 12557 3383
rect 12557 3349 12566 3383
rect 12514 3340 12566 3349
rect 22818 3408 22870 3460
rect 27050 3408 27102 3460
rect 28522 3408 28574 3460
rect 40114 3408 40166 3460
rect 40206 3408 40258 3460
rect 41678 3408 41730 3460
rect 42782 3340 42834 3392
rect 50602 3340 50654 3392
rect 51706 3408 51758 3460
rect 55846 3476 55898 3528
rect 57870 3476 57922 3528
rect 58606 3340 58658 3392
rect 4228 3238 4280 3290
rect 4292 3238 4344 3290
rect 4356 3238 4408 3290
rect 4420 3238 4472 3290
rect 34948 3238 35000 3290
rect 35012 3238 35064 3290
rect 35076 3238 35128 3290
rect 35140 3238 35192 3290
rect 5338 3136 5390 3188
rect 12514 3136 12566 3188
rect 51614 3136 51666 3188
rect 51890 3136 51942 3188
rect 57502 3136 57554 3188
rect 1382 3068 1434 3120
rect 2578 3068 2630 3120
rect 26866 3068 26918 3120
rect 32478 3068 32530 3120
rect 35238 3068 35290 3120
rect 38090 3068 38142 3120
rect 39378 3068 39430 3120
rect 45358 3068 45410 3120
rect 45450 3068 45502 3120
rect 51246 3068 51298 3120
rect 51338 3068 51390 3120
rect 55662 3068 55714 3120
rect 2670 3000 2722 3052
rect 20518 3000 20570 3052
rect 24474 3000 24526 3052
rect 28430 3000 28482 3052
rect 36158 3000 36210 3052
rect 37998 3000 38050 3052
rect 44622 3000 44674 3052
rect 44806 3000 44858 3052
rect 52350 3000 52402 3052
rect 12422 2932 12474 2984
rect 13526 2932 13578 2984
rect 24198 2932 24250 2984
rect 28890 2932 28942 2984
rect 29626 2932 29678 2984
rect 30270 2932 30322 2984
rect 31098 2932 31150 2984
rect 40206 2932 40258 2984
rect 40850 2932 40902 2984
rect 41402 2932 41454 2984
rect 41494 2932 41546 2984
rect 44990 2932 45042 2984
rect 1290 2796 1342 2848
rect 28614 2864 28666 2916
rect 37998 2864 38050 2916
rect 38090 2864 38142 2916
rect 42046 2864 42098 2916
rect 42138 2864 42190 2916
rect 27418 2796 27470 2848
rect 32386 2796 32438 2848
rect 32662 2796 32714 2848
rect 36342 2796 36394 2848
rect 36434 2796 36486 2848
rect 42782 2796 42834 2848
rect 43886 2864 43938 2916
rect 49682 2932 49734 2984
rect 50786 2932 50838 2984
rect 56030 3000 56082 3052
rect 52534 2932 52586 2984
rect 56766 2932 56818 2984
rect 47934 2864 47986 2916
rect 52442 2864 52494 2916
rect 53178 2864 53230 2916
rect 57134 2864 57186 2916
rect 48670 2796 48722 2848
rect 48762 2796 48814 2848
rect 51982 2796 52034 2848
rect 19588 2694 19640 2746
rect 19652 2694 19704 2746
rect 19716 2694 19768 2746
rect 19780 2694 19832 2746
rect 50308 2694 50360 2746
rect 50372 2694 50424 2746
rect 50436 2694 50488 2746
rect 50500 2694 50552 2746
rect 17390 2592 17442 2644
rect 17850 2592 17902 2644
rect 17942 2592 17994 2644
rect 18402 2592 18454 2644
rect 36618 2592 36670 2644
rect 44254 2592 44306 2644
rect 46278 2592 46330 2644
rect 53454 2592 53506 2644
rect 37722 2524 37774 2576
rect 39378 2524 39430 2576
rect 49406 2524 49458 2576
rect 54190 2524 54242 2576
rect 29994 2252 30046 2304
rect 4228 2150 4280 2202
rect 4292 2150 4344 2202
rect 4356 2150 4408 2202
rect 4420 2150 4472 2202
rect 34948 2150 35000 2202
rect 35012 2150 35064 2202
rect 35076 2150 35128 2202
rect 35140 2150 35192 2202
rect 49958 1980 50010 2032
rect 53086 1980 53138 2032
rect 20794 1504 20846 1556
rect 21346 1504 21398 1556
rect 19690 1096 19742 1148
rect 20886 1096 20938 1148
<< metal2 >>
rect 184 59200 240 60000
rect 644 59200 700 60000
rect 1196 59200 1252 60000
rect 1748 59200 1804 60000
rect 2208 59200 2264 60000
rect 2760 59200 2816 60000
rect 3312 59200 3368 60000
rect 3864 59200 3920 60000
rect 4324 59200 4380 60000
rect 4876 59200 4932 60000
rect 5428 59200 5484 60000
rect 5888 59200 5944 60000
rect 6440 59200 6496 60000
rect 6992 59200 7048 60000
rect 7544 59200 7600 60000
rect 8004 59200 8060 60000
rect 8556 59200 8612 60000
rect 9108 59200 9164 60000
rect 9568 59200 9624 60000
rect 10120 59200 10176 60000
rect 10672 59200 10728 60000
rect 11224 59200 11280 60000
rect 11684 59200 11740 60000
rect 12236 59200 12292 60000
rect 12788 59200 12844 60000
rect 13248 59200 13304 60000
rect 13800 59200 13856 60000
rect 14352 59200 14408 60000
rect 14904 59200 14960 60000
rect 15364 59200 15420 60000
rect 15916 59200 15972 60000
rect 16468 59200 16524 60000
rect 17020 59200 17076 60000
rect 17480 59200 17536 60000
rect 18032 59200 18088 60000
rect 18584 59200 18640 60000
rect 19044 59200 19100 60000
rect 19596 59200 19652 60000
rect 20148 59200 20204 60000
rect 20700 59200 20756 60000
rect 21160 59200 21216 60000
rect 21712 59200 21768 60000
rect 22264 59200 22320 60000
rect 22724 59200 22780 60000
rect 23276 59200 23332 60000
rect 23828 59200 23884 60000
rect 24380 59200 24436 60000
rect 24840 59200 24896 60000
rect 25392 59200 25448 60000
rect 25944 59200 26000 60000
rect 26404 59200 26460 60000
rect 26956 59200 27012 60000
rect 27508 59200 27564 60000
rect 28060 59200 28116 60000
rect 28520 59200 28576 60000
rect 29072 59200 29128 60000
rect 29624 59200 29680 60000
rect 30176 59200 30232 60000
rect 30636 59200 30692 60000
rect 31188 59200 31244 60000
rect 31740 59200 31796 60000
rect 32200 59200 32256 60000
rect 32752 59200 32808 60000
rect 33304 59200 33360 60000
rect 33856 59200 33912 60000
rect 34316 59200 34372 60000
rect 34868 59200 34924 60000
rect 35420 59200 35476 60000
rect 35880 59200 35936 60000
rect 36432 59200 36488 60000
rect 36984 59200 37040 60000
rect 37536 59200 37592 60000
rect 37996 59200 38052 60000
rect 38548 59200 38604 60000
rect 39100 59200 39156 60000
rect 39560 59200 39616 60000
rect 40112 59200 40168 60000
rect 40664 59200 40720 60000
rect 41216 59200 41272 60000
rect 41676 59200 41732 60000
rect 42228 59200 42284 60000
rect 42780 59200 42836 60000
rect 43240 59200 43296 60000
rect 43792 59200 43848 60000
rect 44344 59200 44400 60000
rect 44896 59200 44952 60000
rect 45356 59200 45412 60000
rect 45908 59200 45964 60000
rect 46460 59200 46516 60000
rect 47012 59200 47068 60000
rect 47472 59200 47528 60000
rect 48024 59200 48080 60000
rect 48576 59200 48632 60000
rect 49036 59200 49092 60000
rect 49588 59200 49644 60000
rect 50140 59200 50196 60000
rect 50692 59200 50748 60000
rect 51152 59200 51208 60000
rect 51704 59200 51760 60000
rect 52256 59200 52312 60000
rect 52716 59200 52772 60000
rect 53268 59200 53324 60000
rect 53820 59200 53876 60000
rect 54372 59200 54428 60000
rect 54832 59200 54888 60000
rect 55384 59200 55440 60000
rect 55936 59200 55992 60000
rect 56396 59200 56452 60000
rect 56948 59200 57004 60000
rect 57500 59200 57556 60000
rect 58052 59200 58108 60000
rect 58512 59200 58568 60000
rect 59064 59200 59120 60000
rect 59616 59200 59672 60000
rect 198 56438 226 59200
rect 658 56506 686 59200
rect 646 56500 698 56506
rect 646 56442 698 56448
rect 1106 56500 1158 56506
rect 1106 56442 1158 56448
rect 186 56432 238 56438
rect 186 56374 238 56380
rect 1118 29782 1146 56442
rect 1106 29776 1158 29782
rect 1106 29718 1158 29724
rect 1106 15700 1158 15706
rect 1106 15642 1158 15648
rect 1118 3534 1146 15642
rect 1210 5574 1238 59200
rect 1762 56506 1790 59200
rect 1750 56500 1802 56506
rect 1750 56442 1802 56448
rect 2222 56438 2250 59200
rect 2670 56500 2722 56506
rect 2670 56442 2722 56448
rect 1290 56432 1342 56438
rect 1290 56374 1342 56380
rect 1382 56432 1434 56438
rect 1382 56374 1434 56380
rect 2210 56432 2262 56438
rect 2210 56374 2262 56380
rect 2578 56432 2630 56438
rect 2578 56374 2630 56380
rect 1198 5568 1250 5574
rect 1198 5510 1250 5516
rect 186 3528 238 3534
rect 186 3470 238 3476
rect 1106 3528 1158 3534
rect 1106 3470 1158 3476
rect 198 800 226 3470
rect 922 3460 974 3466
rect 922 3402 974 3408
rect 934 800 962 3402
rect 1302 2854 1330 56374
rect 1394 50726 1422 56374
rect 1566 56364 1618 56370
rect 1566 56306 1618 56312
rect 1382 50720 1434 50726
rect 1382 50662 1434 50668
rect 1578 24818 1606 56306
rect 2116 55856 2172 55865
rect 2116 55791 2172 55800
rect 1842 55684 1894 55690
rect 1842 55626 1894 55632
rect 1854 39098 1882 55626
rect 1842 39092 1894 39098
rect 1842 39034 1894 39040
rect 1566 24812 1618 24818
rect 1566 24754 1618 24760
rect 2130 3602 2158 55791
rect 2590 55690 2618 56374
rect 2578 55684 2630 55690
rect 2578 55626 2630 55632
rect 2302 44736 2354 44742
rect 2302 44678 2354 44684
rect 2314 44470 2342 44678
rect 2302 44464 2354 44470
rect 2302 44406 2354 44412
rect 2578 43240 2630 43246
rect 2578 43182 2630 43188
rect 2486 34740 2538 34746
rect 2486 34682 2538 34688
rect 2394 33448 2446 33454
rect 2394 33390 2446 33396
rect 2118 3596 2170 3602
rect 2118 3538 2170 3544
rect 1934 3528 1986 3534
rect 1934 3470 1986 3476
rect 1382 3120 1434 3126
rect 1382 3062 1434 3068
rect 1290 2848 1342 2854
rect 1290 2790 1342 2796
rect 1394 800 1422 3062
rect 1946 800 1974 3470
rect 2406 800 2434 33390
rect 2498 3534 2526 34682
rect 2486 3528 2538 3534
rect 2486 3470 2538 3476
rect 2590 3126 2618 43182
rect 2578 3120 2630 3126
rect 2578 3062 2630 3068
rect 2682 3058 2710 56442
rect 2774 55282 2802 59200
rect 3682 56296 3734 56302
rect 3682 56238 3734 56244
rect 2762 55276 2814 55282
rect 2762 55218 2814 55224
rect 3694 53666 3722 56238
rect 3774 55276 3826 55282
rect 3774 55218 3826 55224
rect 3786 54210 3814 55218
rect 3878 54346 3906 59200
rect 4338 57882 4366 59200
rect 4338 57854 4642 57882
rect 4202 57692 4498 57712
rect 4258 57690 4282 57692
rect 4338 57690 4362 57692
rect 4418 57690 4442 57692
rect 4280 57638 4282 57690
rect 4344 57638 4356 57690
rect 4418 57638 4420 57690
rect 4258 57636 4282 57638
rect 4338 57636 4362 57638
rect 4418 57636 4442 57638
rect 4202 57616 4498 57636
rect 4202 56604 4498 56624
rect 4258 56602 4282 56604
rect 4338 56602 4362 56604
rect 4418 56602 4442 56604
rect 4280 56550 4282 56602
rect 4344 56550 4356 56602
rect 4418 56550 4420 56602
rect 4258 56548 4282 56550
rect 4338 56548 4362 56550
rect 4418 56548 4442 56550
rect 4202 56528 4498 56548
rect 4050 55956 4102 55962
rect 4050 55898 4102 55904
rect 3878 54318 3998 54346
rect 3786 54182 3906 54210
rect 3694 53638 3814 53666
rect 3682 40452 3734 40458
rect 3682 40394 3734 40400
rect 3498 37324 3550 37330
rect 3498 37266 3550 37272
rect 3510 29102 3538 37266
rect 3498 29096 3550 29102
rect 3498 29038 3550 29044
rect 3590 29062 3642 29068
rect 3590 29004 3642 29010
rect 3602 27606 3630 29004
rect 3406 27600 3458 27606
rect 3406 27542 3458 27548
rect 3590 27600 3642 27606
rect 3590 27542 3642 27548
rect 3418 18193 3446 27542
rect 3404 18184 3460 18193
rect 3404 18119 3460 18128
rect 3588 18048 3644 18057
rect 3588 17983 3644 17992
rect 3602 9738 3630 17983
rect 3510 9722 3630 9738
rect 3222 9716 3274 9722
rect 3222 9658 3274 9664
rect 3498 9716 3630 9722
rect 3550 9710 3630 9716
rect 3498 9658 3550 9664
rect 2854 4072 2906 4078
rect 2854 4014 2906 4020
rect 2670 3052 2722 3058
rect 2670 2994 2722 3000
rect 2866 800 2894 4014
rect 3234 800 3262 9658
rect 3694 4146 3722 40394
rect 3786 28626 3814 53638
rect 3878 47598 3906 54182
rect 3866 47592 3918 47598
rect 3866 47534 3918 47540
rect 3866 42016 3918 42022
rect 3866 41958 3918 41964
rect 3774 28620 3826 28626
rect 3774 28562 3826 28568
rect 3774 24132 3826 24138
rect 3774 24074 3826 24080
rect 3682 4140 3734 4146
rect 3682 4082 3734 4088
rect 3786 2802 3814 24074
rect 3878 4078 3906 41958
rect 3970 9110 3998 54318
rect 4062 20602 4090 55898
rect 4202 55516 4498 55536
rect 4258 55514 4282 55516
rect 4338 55514 4362 55516
rect 4418 55514 4442 55516
rect 4280 55462 4282 55514
rect 4344 55462 4356 55514
rect 4418 55462 4420 55514
rect 4258 55460 4282 55462
rect 4338 55460 4362 55462
rect 4418 55460 4442 55462
rect 4202 55440 4498 55460
rect 4614 55282 4642 57854
rect 4890 55418 4918 59200
rect 4970 56772 5022 56778
rect 4970 56714 5022 56720
rect 4878 55412 4930 55418
rect 4878 55354 4930 55360
rect 4602 55276 4654 55282
rect 4602 55218 4654 55224
rect 4202 54428 4498 54448
rect 4258 54426 4282 54428
rect 4338 54426 4362 54428
rect 4418 54426 4442 54428
rect 4280 54374 4282 54426
rect 4344 54374 4356 54426
rect 4418 54374 4420 54426
rect 4258 54372 4282 54374
rect 4338 54372 4362 54374
rect 4418 54372 4442 54374
rect 4202 54352 4498 54372
rect 4202 53340 4498 53360
rect 4258 53338 4282 53340
rect 4338 53338 4362 53340
rect 4418 53338 4442 53340
rect 4280 53286 4282 53338
rect 4344 53286 4356 53338
rect 4418 53286 4420 53338
rect 4258 53284 4282 53286
rect 4338 53284 4362 53286
rect 4418 53284 4442 53286
rect 4202 53264 4498 53284
rect 4202 52252 4498 52272
rect 4258 52250 4282 52252
rect 4338 52250 4362 52252
rect 4418 52250 4442 52252
rect 4280 52198 4282 52250
rect 4344 52198 4356 52250
rect 4418 52198 4420 52250
rect 4258 52196 4282 52198
rect 4338 52196 4362 52198
rect 4418 52196 4442 52198
rect 4202 52176 4498 52196
rect 4202 51164 4498 51184
rect 4258 51162 4282 51164
rect 4338 51162 4362 51164
rect 4418 51162 4442 51164
rect 4280 51110 4282 51162
rect 4344 51110 4356 51162
rect 4418 51110 4420 51162
rect 4258 51108 4282 51110
rect 4338 51108 4362 51110
rect 4418 51108 4442 51110
rect 4202 51088 4498 51108
rect 4202 50076 4498 50096
rect 4258 50074 4282 50076
rect 4338 50074 4362 50076
rect 4418 50074 4442 50076
rect 4280 50022 4282 50074
rect 4344 50022 4356 50074
rect 4418 50022 4420 50074
rect 4258 50020 4282 50022
rect 4338 50020 4362 50022
rect 4418 50020 4442 50022
rect 4202 50000 4498 50020
rect 4202 48988 4498 49008
rect 4258 48986 4282 48988
rect 4338 48986 4362 48988
rect 4418 48986 4442 48988
rect 4280 48934 4282 48986
rect 4344 48934 4356 48986
rect 4418 48934 4420 48986
rect 4258 48932 4282 48934
rect 4338 48932 4362 48934
rect 4418 48932 4442 48934
rect 4202 48912 4498 48932
rect 4202 47900 4498 47920
rect 4258 47898 4282 47900
rect 4338 47898 4362 47900
rect 4418 47898 4442 47900
rect 4280 47846 4282 47898
rect 4344 47846 4356 47898
rect 4418 47846 4420 47898
rect 4258 47844 4282 47846
rect 4338 47844 4362 47846
rect 4418 47844 4442 47846
rect 4202 47824 4498 47844
rect 4202 46812 4498 46832
rect 4258 46810 4282 46812
rect 4338 46810 4362 46812
rect 4418 46810 4442 46812
rect 4280 46758 4282 46810
rect 4344 46758 4356 46810
rect 4418 46758 4420 46810
rect 4258 46756 4282 46758
rect 4338 46756 4362 46758
rect 4418 46756 4442 46758
rect 4202 46736 4498 46756
rect 4202 45724 4498 45744
rect 4258 45722 4282 45724
rect 4338 45722 4362 45724
rect 4418 45722 4442 45724
rect 4280 45670 4282 45722
rect 4344 45670 4356 45722
rect 4418 45670 4420 45722
rect 4258 45668 4282 45670
rect 4338 45668 4362 45670
rect 4418 45668 4442 45670
rect 4202 45648 4498 45668
rect 4202 44636 4498 44656
rect 4258 44634 4282 44636
rect 4338 44634 4362 44636
rect 4418 44634 4442 44636
rect 4280 44582 4282 44634
rect 4344 44582 4356 44634
rect 4418 44582 4420 44634
rect 4258 44580 4282 44582
rect 4338 44580 4362 44582
rect 4418 44580 4442 44582
rect 4202 44560 4498 44580
rect 4202 43548 4498 43568
rect 4258 43546 4282 43548
rect 4338 43546 4362 43548
rect 4418 43546 4442 43548
rect 4280 43494 4282 43546
rect 4344 43494 4356 43546
rect 4418 43494 4420 43546
rect 4258 43492 4282 43494
rect 4338 43492 4362 43494
rect 4418 43492 4442 43494
rect 4202 43472 4498 43492
rect 4202 42460 4498 42480
rect 4258 42458 4282 42460
rect 4338 42458 4362 42460
rect 4418 42458 4442 42460
rect 4280 42406 4282 42458
rect 4344 42406 4356 42458
rect 4418 42406 4420 42458
rect 4258 42404 4282 42406
rect 4338 42404 4362 42406
rect 4418 42404 4442 42406
rect 4202 42384 4498 42404
rect 4202 41372 4498 41392
rect 4258 41370 4282 41372
rect 4338 41370 4362 41372
rect 4418 41370 4442 41372
rect 4280 41318 4282 41370
rect 4344 41318 4356 41370
rect 4418 41318 4420 41370
rect 4258 41316 4282 41318
rect 4338 41316 4362 41318
rect 4418 41316 4442 41318
rect 4202 41296 4498 41316
rect 4202 40284 4498 40304
rect 4258 40282 4282 40284
rect 4338 40282 4362 40284
rect 4418 40282 4442 40284
rect 4280 40230 4282 40282
rect 4344 40230 4356 40282
rect 4418 40230 4420 40282
rect 4258 40228 4282 40230
rect 4338 40228 4362 40230
rect 4418 40228 4442 40230
rect 4202 40208 4498 40228
rect 4202 39196 4498 39216
rect 4258 39194 4282 39196
rect 4338 39194 4362 39196
rect 4418 39194 4442 39196
rect 4280 39142 4282 39194
rect 4344 39142 4356 39194
rect 4418 39142 4420 39194
rect 4258 39140 4282 39142
rect 4338 39140 4362 39142
rect 4418 39140 4442 39142
rect 4202 39120 4498 39140
rect 4786 38956 4838 38962
rect 4786 38898 4838 38904
rect 4202 38108 4498 38128
rect 4258 38106 4282 38108
rect 4338 38106 4362 38108
rect 4418 38106 4442 38108
rect 4280 38054 4282 38106
rect 4344 38054 4356 38106
rect 4418 38054 4420 38106
rect 4258 38052 4282 38054
rect 4338 38052 4362 38054
rect 4418 38052 4442 38054
rect 4202 38032 4498 38052
rect 4798 37330 4826 38898
rect 4786 37324 4838 37330
rect 4786 37266 4838 37272
rect 4202 37020 4498 37040
rect 4258 37018 4282 37020
rect 4338 37018 4362 37020
rect 4418 37018 4442 37020
rect 4280 36966 4282 37018
rect 4344 36966 4356 37018
rect 4418 36966 4420 37018
rect 4258 36964 4282 36966
rect 4338 36964 4362 36966
rect 4418 36964 4442 36966
rect 4202 36944 4498 36964
rect 4202 35932 4498 35952
rect 4258 35930 4282 35932
rect 4338 35930 4362 35932
rect 4418 35930 4442 35932
rect 4280 35878 4282 35930
rect 4344 35878 4356 35930
rect 4418 35878 4420 35930
rect 4258 35876 4282 35878
rect 4338 35876 4362 35878
rect 4418 35876 4442 35878
rect 4202 35856 4498 35876
rect 4202 34844 4498 34864
rect 4258 34842 4282 34844
rect 4338 34842 4362 34844
rect 4418 34842 4442 34844
rect 4280 34790 4282 34842
rect 4344 34790 4356 34842
rect 4418 34790 4420 34842
rect 4258 34788 4282 34790
rect 4338 34788 4362 34790
rect 4418 34788 4442 34790
rect 4202 34768 4498 34788
rect 4202 33756 4498 33776
rect 4258 33754 4282 33756
rect 4338 33754 4362 33756
rect 4418 33754 4442 33756
rect 4280 33702 4282 33754
rect 4344 33702 4356 33754
rect 4418 33702 4420 33754
rect 4258 33700 4282 33702
rect 4338 33700 4362 33702
rect 4418 33700 4442 33702
rect 4202 33680 4498 33700
rect 4202 32668 4498 32688
rect 4258 32666 4282 32668
rect 4338 32666 4362 32668
rect 4418 32666 4442 32668
rect 4280 32614 4282 32666
rect 4344 32614 4356 32666
rect 4418 32614 4420 32666
rect 4258 32612 4282 32614
rect 4338 32612 4362 32614
rect 4418 32612 4442 32614
rect 4202 32592 4498 32612
rect 4202 31580 4498 31600
rect 4258 31578 4282 31580
rect 4338 31578 4362 31580
rect 4418 31578 4442 31580
rect 4280 31526 4282 31578
rect 4344 31526 4356 31578
rect 4418 31526 4420 31578
rect 4258 31524 4282 31526
rect 4338 31524 4362 31526
rect 4418 31524 4442 31526
rect 4202 31504 4498 31524
rect 4202 30492 4498 30512
rect 4258 30490 4282 30492
rect 4338 30490 4362 30492
rect 4418 30490 4442 30492
rect 4280 30438 4282 30490
rect 4344 30438 4356 30490
rect 4418 30438 4420 30490
rect 4258 30436 4282 30438
rect 4338 30436 4362 30438
rect 4418 30436 4442 30438
rect 4202 30416 4498 30436
rect 4202 29404 4498 29424
rect 4258 29402 4282 29404
rect 4338 29402 4362 29404
rect 4418 29402 4442 29404
rect 4280 29350 4282 29402
rect 4344 29350 4356 29402
rect 4418 29350 4420 29402
rect 4258 29348 4282 29350
rect 4338 29348 4362 29350
rect 4418 29348 4442 29350
rect 4202 29328 4498 29348
rect 4202 28316 4498 28336
rect 4258 28314 4282 28316
rect 4338 28314 4362 28316
rect 4418 28314 4442 28316
rect 4280 28262 4282 28314
rect 4344 28262 4356 28314
rect 4418 28262 4420 28314
rect 4258 28260 4282 28262
rect 4338 28260 4362 28262
rect 4418 28260 4442 28262
rect 4202 28240 4498 28260
rect 4202 27228 4498 27248
rect 4258 27226 4282 27228
rect 4338 27226 4362 27228
rect 4418 27226 4442 27228
rect 4280 27174 4282 27226
rect 4344 27174 4356 27226
rect 4418 27174 4420 27226
rect 4258 27172 4282 27174
rect 4338 27172 4362 27174
rect 4418 27172 4442 27174
rect 4202 27152 4498 27172
rect 4202 26140 4498 26160
rect 4258 26138 4282 26140
rect 4338 26138 4362 26140
rect 4418 26138 4442 26140
rect 4280 26086 4282 26138
rect 4344 26086 4356 26138
rect 4418 26086 4420 26138
rect 4258 26084 4282 26086
rect 4338 26084 4362 26086
rect 4418 26084 4442 26086
rect 4202 26064 4498 26084
rect 4202 25052 4498 25072
rect 4258 25050 4282 25052
rect 4338 25050 4362 25052
rect 4418 25050 4442 25052
rect 4280 24998 4282 25050
rect 4344 24998 4356 25050
rect 4418 24998 4420 25050
rect 4258 24996 4282 24998
rect 4338 24996 4362 24998
rect 4418 24996 4442 24998
rect 4202 24976 4498 24996
rect 4202 23964 4498 23984
rect 4258 23962 4282 23964
rect 4338 23962 4362 23964
rect 4418 23962 4442 23964
rect 4280 23910 4282 23962
rect 4344 23910 4356 23962
rect 4418 23910 4420 23962
rect 4258 23908 4282 23910
rect 4338 23908 4362 23910
rect 4418 23908 4442 23910
rect 4202 23888 4498 23908
rect 4202 22876 4498 22896
rect 4258 22874 4282 22876
rect 4338 22874 4362 22876
rect 4418 22874 4442 22876
rect 4280 22822 4282 22874
rect 4344 22822 4356 22874
rect 4418 22822 4420 22874
rect 4258 22820 4282 22822
rect 4338 22820 4362 22822
rect 4418 22820 4442 22822
rect 4202 22800 4498 22820
rect 4202 21788 4498 21808
rect 4258 21786 4282 21788
rect 4338 21786 4362 21788
rect 4418 21786 4442 21788
rect 4280 21734 4282 21786
rect 4344 21734 4356 21786
rect 4418 21734 4420 21786
rect 4258 21732 4282 21734
rect 4338 21732 4362 21734
rect 4418 21732 4442 21734
rect 4202 21712 4498 21732
rect 4202 20700 4498 20720
rect 4258 20698 4282 20700
rect 4338 20698 4362 20700
rect 4418 20698 4442 20700
rect 4280 20646 4282 20698
rect 4344 20646 4356 20698
rect 4418 20646 4420 20698
rect 4258 20644 4282 20646
rect 4338 20644 4362 20646
rect 4418 20644 4442 20646
rect 4202 20624 4498 20644
rect 4050 20596 4102 20602
rect 4050 20538 4102 20544
rect 4202 19612 4498 19632
rect 4258 19610 4282 19612
rect 4338 19610 4362 19612
rect 4418 19610 4442 19612
rect 4280 19558 4282 19610
rect 4344 19558 4356 19610
rect 4418 19558 4420 19610
rect 4258 19556 4282 19558
rect 4338 19556 4362 19558
rect 4418 19556 4442 19558
rect 4202 19536 4498 19556
rect 4202 18524 4498 18544
rect 4258 18522 4282 18524
rect 4338 18522 4362 18524
rect 4418 18522 4442 18524
rect 4280 18470 4282 18522
rect 4344 18470 4356 18522
rect 4418 18470 4420 18522
rect 4258 18468 4282 18470
rect 4338 18468 4362 18470
rect 4418 18468 4442 18470
rect 4202 18448 4498 18468
rect 4202 17436 4498 17456
rect 4258 17434 4282 17436
rect 4338 17434 4362 17436
rect 4418 17434 4442 17436
rect 4280 17382 4282 17434
rect 4344 17382 4356 17434
rect 4418 17382 4420 17434
rect 4258 17380 4282 17382
rect 4338 17380 4362 17382
rect 4418 17380 4442 17382
rect 4202 17360 4498 17380
rect 4202 16348 4498 16368
rect 4258 16346 4282 16348
rect 4338 16346 4362 16348
rect 4418 16346 4442 16348
rect 4280 16294 4282 16346
rect 4344 16294 4356 16346
rect 4418 16294 4420 16346
rect 4258 16292 4282 16294
rect 4338 16292 4362 16294
rect 4418 16292 4442 16294
rect 4202 16272 4498 16292
rect 4202 15260 4498 15280
rect 4258 15258 4282 15260
rect 4338 15258 4362 15260
rect 4418 15258 4442 15260
rect 4280 15206 4282 15258
rect 4344 15206 4356 15258
rect 4418 15206 4420 15258
rect 4258 15204 4282 15206
rect 4338 15204 4362 15206
rect 4418 15204 4442 15206
rect 4202 15184 4498 15204
rect 4202 14172 4498 14192
rect 4258 14170 4282 14172
rect 4338 14170 4362 14172
rect 4418 14170 4442 14172
rect 4280 14118 4282 14170
rect 4344 14118 4356 14170
rect 4418 14118 4420 14170
rect 4258 14116 4282 14118
rect 4338 14116 4362 14118
rect 4418 14116 4442 14118
rect 4202 14096 4498 14116
rect 4202 13084 4498 13104
rect 4258 13082 4282 13084
rect 4338 13082 4362 13084
rect 4418 13082 4442 13084
rect 4280 13030 4282 13082
rect 4344 13030 4356 13082
rect 4418 13030 4420 13082
rect 4258 13028 4282 13030
rect 4338 13028 4362 13030
rect 4418 13028 4442 13030
rect 4202 13008 4498 13028
rect 4202 11996 4498 12016
rect 4258 11994 4282 11996
rect 4338 11994 4362 11996
rect 4418 11994 4442 11996
rect 4280 11942 4282 11994
rect 4344 11942 4356 11994
rect 4418 11942 4420 11994
rect 4258 11940 4282 11942
rect 4338 11940 4362 11942
rect 4418 11940 4442 11942
rect 4202 11920 4498 11940
rect 4202 10908 4498 10928
rect 4258 10906 4282 10908
rect 4338 10906 4362 10908
rect 4418 10906 4442 10908
rect 4280 10854 4282 10906
rect 4344 10854 4356 10906
rect 4418 10854 4420 10906
rect 4258 10852 4282 10854
rect 4338 10852 4362 10854
rect 4418 10852 4442 10854
rect 4202 10832 4498 10852
rect 4202 9820 4498 9840
rect 4258 9818 4282 9820
rect 4338 9818 4362 9820
rect 4418 9818 4442 9820
rect 4280 9766 4282 9818
rect 4344 9766 4356 9818
rect 4418 9766 4420 9818
rect 4258 9764 4282 9766
rect 4338 9764 4362 9766
rect 4418 9764 4442 9766
rect 4202 9744 4498 9764
rect 3958 9104 4010 9110
rect 3958 9046 4010 9052
rect 4202 8732 4498 8752
rect 4258 8730 4282 8732
rect 4338 8730 4362 8732
rect 4418 8730 4442 8732
rect 4280 8678 4282 8730
rect 4344 8678 4356 8730
rect 4418 8678 4420 8730
rect 4258 8676 4282 8678
rect 4338 8676 4362 8678
rect 4418 8676 4442 8678
rect 4202 8656 4498 8676
rect 4202 7644 4498 7664
rect 4258 7642 4282 7644
rect 4338 7642 4362 7644
rect 4418 7642 4442 7644
rect 4280 7590 4282 7642
rect 4344 7590 4356 7642
rect 4418 7590 4420 7642
rect 4258 7588 4282 7590
rect 4338 7588 4362 7590
rect 4418 7588 4442 7590
rect 4202 7568 4498 7588
rect 4202 6556 4498 6576
rect 4258 6554 4282 6556
rect 4338 6554 4362 6556
rect 4418 6554 4442 6556
rect 4280 6502 4282 6554
rect 4344 6502 4356 6554
rect 4418 6502 4420 6554
rect 4258 6500 4282 6502
rect 4338 6500 4362 6502
rect 4418 6500 4442 6502
rect 4202 6480 4498 6500
rect 4202 5468 4498 5488
rect 4258 5466 4282 5468
rect 4338 5466 4362 5468
rect 4418 5466 4442 5468
rect 4280 5414 4282 5466
rect 4344 5414 4356 5466
rect 4418 5414 4420 5466
rect 4258 5412 4282 5414
rect 4338 5412 4362 5414
rect 4418 5412 4442 5414
rect 4202 5392 4498 5412
rect 4982 4842 5010 56714
rect 5442 55162 5470 59200
rect 5902 55162 5930 59200
rect 6350 55820 6402 55826
rect 6350 55762 6402 55768
rect 5258 55134 5470 55162
rect 5534 55134 5930 55162
rect 5258 37346 5286 55134
rect 5338 55072 5390 55078
rect 5338 55014 5390 55020
rect 5166 37318 5286 37346
rect 5166 36258 5194 37318
rect 5166 36230 5286 36258
rect 5258 31142 5286 36230
rect 5246 31136 5298 31142
rect 5246 31078 5298 31084
rect 5350 27674 5378 55014
rect 5430 31136 5482 31142
rect 5430 31078 5482 31084
rect 5338 27668 5390 27674
rect 5338 27610 5390 27616
rect 5338 27464 5390 27470
rect 5338 27406 5390 27412
rect 5154 19984 5206 19990
rect 5154 19926 5206 19932
rect 5062 17536 5114 17542
rect 5062 17478 5114 17484
rect 4706 4814 5010 4842
rect 4202 4380 4498 4400
rect 4258 4378 4282 4380
rect 4338 4378 4362 4380
rect 4418 4378 4442 4380
rect 4280 4326 4282 4378
rect 4344 4326 4356 4378
rect 4418 4326 4420 4378
rect 4258 4324 4282 4326
rect 4338 4324 4362 4326
rect 4418 4324 4442 4326
rect 4202 4304 4498 4324
rect 3958 4140 4010 4146
rect 3958 4082 4010 4088
rect 3866 4072 3918 4078
rect 3866 4014 3918 4020
rect 3510 2774 3814 2802
rect 3510 2666 3538 2774
rect 3510 2638 3630 2666
rect 3602 800 3630 2638
rect 3970 800 3998 4082
rect 4602 4072 4654 4078
rect 4602 4014 4654 4020
rect 4202 3292 4498 3312
rect 4258 3290 4282 3292
rect 4338 3290 4362 3292
rect 4418 3290 4442 3292
rect 4280 3238 4282 3290
rect 4344 3238 4356 3290
rect 4418 3238 4420 3290
rect 4258 3236 4282 3238
rect 4338 3236 4362 3238
rect 4418 3236 4442 3238
rect 4202 3216 4498 3236
rect 4202 2204 4498 2224
rect 4258 2202 4282 2204
rect 4338 2202 4362 2204
rect 4418 2202 4442 2204
rect 4280 2150 4282 2202
rect 4344 2150 4356 2202
rect 4418 2150 4420 2202
rect 4258 2148 4282 2150
rect 4338 2148 4362 2150
rect 4418 2148 4442 2150
rect 4202 2128 4498 2148
rect 4614 1442 4642 4014
rect 4338 1414 4642 1442
rect 4338 800 4366 1414
rect 4706 800 4734 4814
rect 5074 4078 5102 17478
rect 5062 4072 5114 4078
rect 5062 4014 5114 4020
rect 5062 3936 5114 3942
rect 5062 3878 5114 3884
rect 5074 800 5102 3878
rect 5166 2836 5194 19926
rect 5244 18048 5300 18057
rect 5244 17983 5300 17992
rect 5258 14550 5286 17983
rect 5246 14544 5298 14550
rect 5246 14486 5298 14492
rect 5246 8832 5298 8838
rect 5246 8774 5298 8780
rect 5258 3942 5286 8774
rect 5246 3936 5298 3942
rect 5246 3878 5298 3884
rect 5350 3194 5378 27406
rect 5442 18057 5470 31078
rect 5534 26450 5562 55134
rect 6362 53394 6390 55762
rect 6454 55162 6482 59200
rect 7006 55350 7034 59200
rect 7454 55412 7506 55418
rect 7454 55354 7506 55360
rect 6994 55344 7046 55350
rect 6994 55286 7046 55292
rect 7466 55162 7494 55354
rect 7558 55282 7586 59200
rect 8190 55684 8242 55690
rect 8190 55626 8242 55632
rect 7914 55344 7966 55350
rect 7914 55286 7966 55292
rect 7546 55276 7598 55282
rect 7546 55218 7598 55224
rect 6454 55134 6850 55162
rect 7466 55134 7586 55162
rect 6362 53366 6574 53394
rect 5522 26444 5574 26450
rect 5522 26386 5574 26392
rect 5428 18048 5484 18057
rect 5428 17983 5484 17992
rect 5430 14544 5482 14550
rect 5430 14486 5482 14492
rect 5442 5846 5470 14486
rect 6546 13394 6574 53366
rect 6718 48000 6770 48006
rect 6718 47942 6770 47948
rect 6626 26308 6678 26314
rect 6626 26250 6678 26256
rect 6534 13388 6586 13394
rect 6534 13330 6586 13336
rect 5798 12096 5850 12102
rect 5798 12038 5850 12044
rect 5430 5840 5482 5846
rect 5430 5782 5482 5788
rect 5338 3188 5390 3194
rect 5338 3130 5390 3136
rect 5166 2808 5378 2836
rect 5350 2666 5378 2808
rect 5350 2638 5470 2666
rect 5442 800 5470 2638
rect 5810 800 5838 12038
rect 6638 4842 6666 26250
rect 6546 4814 6666 4842
rect 6166 4140 6218 4146
rect 6166 4082 6218 4088
rect 6178 800 6206 4082
rect 6546 800 6574 4814
rect 6730 4146 6758 47942
rect 6718 4140 6770 4146
rect 6718 4082 6770 4088
rect 6822 4078 6850 55134
rect 7362 30592 7414 30598
rect 7362 30534 7414 30540
rect 6902 4684 6954 4690
rect 6902 4626 6954 4632
rect 6810 4072 6862 4078
rect 6810 4014 6862 4020
rect 6914 800 6942 4626
rect 7270 4140 7322 4146
rect 7270 4082 7322 4088
rect 7282 800 7310 4082
rect 7374 3602 7402 30534
rect 7454 19304 7506 19310
rect 7454 19246 7506 19252
rect 7466 9722 7494 19246
rect 7454 9716 7506 9722
rect 7454 9658 7506 9664
rect 7558 3942 7586 55134
rect 7822 29028 7874 29034
rect 7822 28970 7874 28976
rect 7638 26988 7690 26994
rect 7638 26930 7690 26936
rect 7650 18698 7678 26930
rect 7730 25832 7782 25838
rect 7730 25774 7782 25780
rect 7742 25430 7770 25774
rect 7730 25424 7782 25430
rect 7730 25366 7782 25372
rect 7730 20936 7782 20942
rect 7730 20878 7782 20884
rect 7638 18692 7690 18698
rect 7638 18634 7690 18640
rect 7742 4146 7770 20878
rect 7834 19344 7862 28970
rect 7926 26994 7954 55286
rect 8098 55276 8150 55282
rect 8098 55218 8150 55224
rect 8006 48680 8058 48686
rect 8006 48622 8058 48628
rect 7914 26988 7966 26994
rect 7914 26930 7966 26936
rect 8018 24154 8046 48622
rect 7926 24126 8046 24154
rect 7822 19338 7874 19344
rect 7822 19280 7874 19286
rect 7822 9716 7874 9722
rect 7822 9658 7874 9664
rect 7730 4140 7782 4146
rect 7730 4082 7782 4088
rect 7834 4026 7862 9658
rect 7650 3998 7862 4026
rect 7546 3936 7598 3942
rect 7546 3878 7598 3884
rect 7362 3596 7414 3602
rect 7362 3538 7414 3544
rect 7650 800 7678 3998
rect 7926 3176 7954 24126
rect 8006 19304 8058 19310
rect 8004 19272 8006 19281
rect 8058 19272 8060 19281
rect 8004 19207 8060 19216
rect 8006 17128 8058 17134
rect 8006 17070 8058 17076
rect 8018 16794 8046 17070
rect 8006 16788 8058 16794
rect 8006 16730 8058 16736
rect 8004 13968 8060 13977
rect 8004 13903 8006 13912
rect 8058 13903 8060 13912
rect 8006 13874 8058 13880
rect 8110 13410 8138 55218
rect 8018 13382 8138 13410
rect 8018 6798 8046 13382
rect 8202 13274 8230 55626
rect 8282 55344 8334 55350
rect 8282 55286 8334 55292
rect 8294 31770 8322 55286
rect 8570 54806 8598 59200
rect 8558 54800 8610 54806
rect 8558 54742 8610 54748
rect 9122 47190 9150 59200
rect 9582 55350 9610 59200
rect 10134 56234 10162 59200
rect 10306 56500 10358 56506
rect 10306 56442 10358 56448
rect 10122 56228 10174 56234
rect 10122 56170 10174 56176
rect 9846 55412 9898 55418
rect 9846 55354 9898 55360
rect 9570 55344 9622 55350
rect 9570 55286 9622 55292
rect 8650 47184 8702 47190
rect 8650 47126 8702 47132
rect 9110 47184 9162 47190
rect 9110 47126 9162 47132
rect 8662 46866 8690 47126
rect 8662 46838 8966 46866
rect 8938 45558 8966 46838
rect 8926 45552 8978 45558
rect 8926 45494 8978 45500
rect 9110 45552 9162 45558
rect 9110 45494 9162 45500
rect 8558 37664 8610 37670
rect 8558 37606 8610 37612
rect 8294 31742 8460 31770
rect 8432 31634 8460 31742
rect 8386 31606 8460 31634
rect 8282 25152 8334 25158
rect 8282 25094 8334 25100
rect 8294 24954 8322 25094
rect 8282 24948 8334 24954
rect 8282 24890 8334 24896
rect 8282 20256 8334 20262
rect 8282 20198 8334 20204
rect 8294 20058 8322 20198
rect 8282 20052 8334 20058
rect 8282 19994 8334 20000
rect 8386 19938 8414 31606
rect 8466 30184 8518 30190
rect 8466 30126 8518 30132
rect 8478 29714 8506 30126
rect 8466 29708 8518 29714
rect 8466 29650 8518 29656
rect 8570 29170 8598 37606
rect 9122 37108 9150 45494
rect 8938 37080 9150 37108
rect 8938 32450 8966 37080
rect 8938 32422 9150 32450
rect 8742 31272 8794 31278
rect 8742 31214 8794 31220
rect 8754 30870 8782 31214
rect 8834 31136 8886 31142
rect 9018 31136 9070 31142
rect 8886 31084 9018 31090
rect 8834 31078 9070 31084
rect 8846 31062 9058 31078
rect 8742 30864 8794 30870
rect 8742 30806 8794 30812
rect 8834 30048 8886 30054
rect 9018 30048 9070 30054
rect 8886 29996 9018 30002
rect 8834 29990 9070 29996
rect 8846 29974 9058 29990
rect 8558 29164 8610 29170
rect 8558 29106 8610 29112
rect 8570 28082 8966 28098
rect 8558 28076 8978 28082
rect 8610 28070 8926 28076
rect 8558 28018 8610 28024
rect 8926 28018 8978 28024
rect 8834 28008 8886 28014
rect 8570 27956 8834 27962
rect 8570 27950 8886 27956
rect 8570 27934 8874 27950
rect 8570 27878 8598 27934
rect 8558 27872 8610 27878
rect 8558 27814 8610 27820
rect 8558 26988 8610 26994
rect 8834 26988 8886 26994
rect 8610 26948 8834 26976
rect 8558 26930 8610 26936
rect 8834 26930 8886 26936
rect 8466 26920 8518 26926
rect 8926 26920 8978 26926
rect 8518 26868 8926 26874
rect 8466 26862 8978 26868
rect 8478 26846 8966 26862
rect 8558 26036 8610 26042
rect 8610 25996 8966 26024
rect 8558 25978 8610 25984
rect 8558 25900 8610 25906
rect 8558 25842 8610 25848
rect 8570 25786 8598 25842
rect 8570 25758 8874 25786
rect 8938 25770 8966 25996
rect 8846 25702 8874 25758
rect 8926 25764 8978 25770
rect 8926 25706 8978 25712
rect 8696 25696 8748 25702
rect 8696 25638 8748 25644
rect 8834 25696 8886 25702
rect 8834 25638 8886 25644
rect 8708 25498 8736 25638
rect 8696 25492 8748 25498
rect 8696 25434 8748 25440
rect 8604 24812 8656 24818
rect 8926 24812 8978 24818
rect 8656 24772 8926 24800
rect 8604 24754 8656 24760
rect 8926 24754 8978 24760
rect 8466 24676 8518 24682
rect 8466 24618 8518 24624
rect 8478 24410 8506 24618
rect 8466 24404 8518 24410
rect 8466 24346 8518 24352
rect 8650 23860 8702 23866
rect 8834 23860 8886 23866
rect 8702 23820 8834 23848
rect 8650 23802 8702 23808
rect 8834 23802 8886 23808
rect 8604 23758 8656 23764
rect 8656 23730 8782 23746
rect 8656 23724 8794 23730
rect 8656 23718 8742 23724
rect 8604 23700 8656 23706
rect 8742 23666 8794 23672
rect 8466 23656 8518 23662
rect 8464 23624 8466 23633
rect 8834 23656 8886 23662
rect 8518 23624 8520 23633
rect 8834 23598 8886 23604
rect 8464 23559 8520 23568
rect 8466 23520 8518 23526
rect 8846 23508 8874 23598
rect 8518 23480 8874 23508
rect 8466 23462 8518 23468
rect 8466 21344 8518 21350
rect 8650 21344 8702 21350
rect 8518 21292 8650 21298
rect 8466 21286 8702 21292
rect 8478 21270 8690 21286
rect 8478 20602 8690 20618
rect 8466 20596 8702 20602
rect 8518 20590 8650 20596
rect 8466 20538 8518 20544
rect 8650 20538 8702 20544
rect 8294 19910 8414 19938
rect 8294 15042 8322 19910
rect 8466 19712 8518 19718
rect 8466 19654 8518 19660
rect 8478 19514 8506 19654
rect 8466 19508 8518 19514
rect 8466 19450 8518 19456
rect 8420 19270 8472 19276
rect 8420 19212 8472 19218
rect 8924 19272 8980 19281
rect 8432 18986 8460 19212
rect 8924 19207 8980 19216
rect 8938 19174 8966 19207
rect 8926 19168 8978 19174
rect 8926 19110 8978 19116
rect 8432 18970 8506 18986
rect 8432 18964 8518 18970
rect 8432 18958 8466 18964
rect 8466 18906 8518 18912
rect 8650 18624 8702 18630
rect 8650 18566 8702 18572
rect 8662 18290 8690 18566
rect 8832 18456 8888 18465
rect 8832 18391 8834 18400
rect 8886 18391 8888 18400
rect 9016 18456 9072 18465
rect 9016 18391 9018 18400
rect 8834 18362 8886 18368
rect 9070 18391 9072 18400
rect 9018 18362 9070 18368
rect 9122 18306 9150 32422
rect 9294 31884 9346 31890
rect 9294 31826 9346 31832
rect 8650 18284 8702 18290
rect 8650 18226 8702 18232
rect 9030 18278 9150 18306
rect 8834 17672 8886 17678
rect 8834 17614 8886 17620
rect 8742 17604 8794 17610
rect 8742 17546 8794 17552
rect 8754 17134 8782 17546
rect 8846 17338 8874 17614
rect 8834 17332 8886 17338
rect 8834 17274 8886 17280
rect 8742 17128 8794 17134
rect 8742 17070 8794 17076
rect 8650 16448 8702 16454
rect 8650 16390 8702 16396
rect 8662 16132 8690 16390
rect 8742 16244 8794 16250
rect 8742 16186 8794 16192
rect 8650 16126 8702 16132
rect 8650 16068 8702 16074
rect 8754 15910 8782 16186
rect 8742 15904 8794 15910
rect 8742 15846 8794 15852
rect 8466 15156 8518 15162
rect 8650 15156 8702 15162
rect 8518 15116 8650 15144
rect 8466 15098 8518 15104
rect 8650 15098 8702 15104
rect 8294 15014 8414 15042
rect 8280 14920 8336 14929
rect 8386 14906 8414 15014
rect 8650 15020 8702 15026
rect 8650 14962 8702 14968
rect 8662 14929 8690 14962
rect 8648 14920 8704 14929
rect 8386 14878 8598 14906
rect 8280 14855 8336 14864
rect 8156 13246 8230 13274
rect 8156 12986 8184 13246
rect 8144 12980 8196 12986
rect 8144 12922 8196 12928
rect 8466 11688 8518 11694
rect 8236 11654 8288 11660
rect 8288 11636 8466 11642
rect 8288 11630 8518 11636
rect 8288 11614 8506 11630
rect 8236 11596 8288 11602
rect 8374 9478 8426 9484
rect 8374 9420 8426 9426
rect 8386 9042 8414 9420
rect 8374 9036 8426 9042
rect 8374 8978 8426 8984
rect 8570 8650 8598 14878
rect 8648 14855 8704 14864
rect 8834 14068 8886 14074
rect 8834 14010 8886 14016
rect 8846 13977 8874 14010
rect 8832 13968 8888 13977
rect 8832 13903 8888 13912
rect 9030 12866 9058 18278
rect 9110 17298 9162 17304
rect 9110 17241 9162 17246
rect 9108 17232 9164 17241
rect 9108 17167 9164 17176
rect 8846 12838 9058 12866
rect 8846 10418 8874 12838
rect 8926 12776 8978 12782
rect 8926 12718 8978 12724
rect 8938 10520 8966 12718
rect 9202 11212 9254 11218
rect 9202 11154 9254 11160
rect 8938 10492 9058 10520
rect 8846 10390 8966 10418
rect 8386 8622 8598 8650
rect 8234 7304 8290 7313
rect 8234 7239 8290 7248
rect 8098 6860 8150 6866
rect 8098 6802 8150 6808
rect 8006 6792 8058 6798
rect 8006 6734 8058 6740
rect 8110 6322 8138 6802
rect 8098 6316 8150 6322
rect 8098 6258 8150 6264
rect 8386 5370 8414 8622
rect 8834 8560 8886 8566
rect 8834 8502 8886 8508
rect 8558 8424 8610 8430
rect 8846 8412 8874 8502
rect 8610 8384 8874 8412
rect 8558 8366 8610 8372
rect 8466 6656 8518 6662
rect 8466 6598 8518 6604
rect 8478 6458 8506 6598
rect 8466 6452 8518 6458
rect 8466 6394 8518 6400
rect 8374 5364 8426 5370
rect 8374 5306 8426 5312
rect 8742 5160 8794 5166
rect 8742 5102 8794 5108
rect 8650 5024 8702 5030
rect 8754 4978 8782 5102
rect 8702 4972 8782 4978
rect 8650 4966 8782 4972
rect 8662 4950 8782 4966
rect 8938 4146 8966 10390
rect 9030 4690 9058 10492
rect 9110 7336 9162 7342
rect 9110 7278 9162 7284
rect 9018 4684 9070 4690
rect 9018 4626 9070 4632
rect 8926 4140 8978 4146
rect 8926 4082 8978 4088
rect 8374 3732 8426 3738
rect 8374 3674 8426 3680
rect 7926 3148 8046 3176
rect 8018 800 8046 3148
rect 8386 800 8414 3674
rect 8742 3528 8794 3534
rect 8742 3470 8794 3476
rect 8754 800 8782 3470
rect 9122 800 9150 7278
rect 9214 3738 9242 11154
rect 9306 11098 9334 31826
rect 9858 24274 9886 55354
rect 10214 24812 10266 24818
rect 10214 24754 10266 24760
rect 10226 24614 10254 24754
rect 10214 24608 10266 24614
rect 10214 24550 10266 24556
rect 9846 24268 9898 24274
rect 9846 24210 9898 24216
rect 9478 23792 9530 23798
rect 9478 23734 9530 23740
rect 9386 21888 9438 21894
rect 9386 21830 9438 21836
rect 9398 11218 9426 21830
rect 9386 11212 9438 11218
rect 9386 11154 9438 11160
rect 9306 11070 9426 11098
rect 9294 11008 9346 11014
rect 9294 10950 9346 10956
rect 9306 10538 9334 10950
rect 9294 10532 9346 10538
rect 9294 10474 9346 10480
rect 9202 3732 9254 3738
rect 9202 3674 9254 3680
rect 9398 3380 9426 11070
rect 9490 3534 9518 23734
rect 9662 22976 9714 22982
rect 9662 22918 9714 22924
rect 9674 22234 9702 22918
rect 9662 22228 9714 22234
rect 9662 22170 9714 22176
rect 9570 17264 9622 17270
rect 9568 17232 9570 17241
rect 9622 17232 9624 17241
rect 9568 17167 9624 17176
rect 10318 5370 10346 56442
rect 10686 55162 10714 59200
rect 11238 55162 11266 59200
rect 11698 56166 11726 59200
rect 11686 56160 11738 56166
rect 11686 56102 11738 56108
rect 11410 55752 11462 55758
rect 11410 55694 11462 55700
rect 10686 55134 10990 55162
rect 10858 34604 10910 34610
rect 10858 34546 10910 34552
rect 10766 31952 10818 31958
rect 10766 31894 10818 31900
rect 10582 8424 10634 8430
rect 10582 8366 10634 8372
rect 10306 5364 10358 5370
rect 10306 5306 10358 5312
rect 10214 4140 10266 4146
rect 10214 4082 10266 4088
rect 9846 4072 9898 4078
rect 9846 4014 9898 4020
rect 9478 3528 9530 3534
rect 9478 3470 9530 3476
rect 9398 3352 9518 3380
rect 9490 800 9518 3352
rect 9858 800 9886 4014
rect 10226 800 10254 4082
rect 10594 800 10622 8366
rect 10778 4146 10806 31894
rect 10766 4140 10818 4146
rect 10766 4082 10818 4088
rect 10870 4078 10898 34546
rect 10962 5778 10990 55134
rect 11054 55134 11266 55162
rect 10950 5772 11002 5778
rect 10950 5714 11002 5720
rect 11054 5234 11082 55134
rect 11422 26042 11450 55694
rect 11870 40384 11922 40390
rect 11870 40326 11922 40332
rect 11882 40186 11910 40326
rect 11870 40180 11922 40186
rect 11870 40122 11922 40128
rect 12054 37324 12106 37330
rect 12054 37266 12106 37272
rect 11410 26036 11462 26042
rect 11410 25978 11462 25984
rect 11776 23624 11832 23633
rect 11776 23559 11832 23568
rect 11790 23526 11818 23559
rect 11778 23520 11830 23526
rect 11778 23462 11830 23468
rect 11410 20256 11462 20262
rect 11410 20198 11462 20204
rect 11422 20058 11450 20198
rect 11410 20052 11462 20058
rect 11410 19994 11462 20000
rect 11042 5228 11094 5234
rect 11042 5170 11094 5176
rect 11686 4140 11738 4146
rect 11686 4082 11738 4088
rect 10858 4072 10910 4078
rect 10858 4014 10910 4020
rect 11318 4072 11370 4078
rect 11318 4014 11370 4020
rect 10950 3596 11002 3602
rect 10950 3538 11002 3544
rect 10962 800 10990 3538
rect 11330 800 11358 4014
rect 11698 800 11726 4082
rect 12066 800 12094 37266
rect 12250 35630 12278 59200
rect 12802 56506 12830 59200
rect 12790 56500 12842 56506
rect 12790 56442 12842 56448
rect 13158 56228 13210 56234
rect 13158 56170 13210 56176
rect 13066 55344 13118 55350
rect 13066 55286 13118 55292
rect 12330 49088 12382 49094
rect 12330 49030 12382 49036
rect 12238 35624 12290 35630
rect 12238 35566 12290 35572
rect 12146 30184 12198 30190
rect 12146 30126 12198 30132
rect 12158 4078 12186 30126
rect 12342 4146 12370 49030
rect 12974 37120 13026 37126
rect 12974 37062 13026 37068
rect 12882 30116 12934 30122
rect 12882 30058 12934 30064
rect 12894 29850 12922 30058
rect 12882 29844 12934 29850
rect 12882 29786 12934 29792
rect 12422 25152 12474 25158
rect 12422 25094 12474 25100
rect 12434 24954 12462 25094
rect 12422 24948 12474 24954
rect 12422 24890 12474 24896
rect 12790 18624 12842 18630
rect 12790 18566 12842 18572
rect 12606 18216 12658 18222
rect 12606 18158 12658 18164
rect 12618 7546 12646 18158
rect 12606 7540 12658 7546
rect 12606 7482 12658 7488
rect 12802 7478 12830 18566
rect 12882 18080 12934 18086
rect 12882 18022 12934 18028
rect 12790 7472 12842 7478
rect 12790 7414 12842 7420
rect 12698 7404 12750 7410
rect 12698 7346 12750 7352
rect 12710 7313 12738 7346
rect 12696 7304 12752 7313
rect 12696 7239 12752 7248
rect 12330 4140 12382 4146
rect 12330 4082 12382 4088
rect 12146 4072 12198 4078
rect 12146 4014 12198 4020
rect 12790 4004 12842 4010
rect 12790 3946 12842 3952
rect 12514 3392 12566 3398
rect 12514 3334 12566 3340
rect 12526 3194 12554 3334
rect 12514 3188 12566 3194
rect 12514 3130 12566 3136
rect 12422 2984 12474 2990
rect 12422 2926 12474 2932
rect 12434 800 12462 2926
rect 12802 800 12830 3946
rect 12894 2802 12922 18022
rect 12986 4146 13014 37062
rect 13078 13938 13106 55286
rect 13170 19310 13198 56170
rect 13262 55282 13290 59200
rect 13250 55276 13302 55282
rect 13250 55218 13302 55224
rect 13710 55276 13762 55282
rect 13710 55218 13762 55224
rect 13618 42288 13670 42294
rect 13618 42230 13670 42236
rect 13526 36032 13578 36038
rect 13526 35974 13578 35980
rect 13158 19304 13210 19310
rect 13158 19246 13210 19252
rect 13158 19168 13210 19174
rect 13158 19110 13210 19116
rect 13066 13932 13118 13938
rect 13066 13874 13118 13880
rect 13170 13818 13198 19110
rect 13342 18964 13394 18970
rect 13342 18906 13394 18912
rect 13078 13790 13198 13818
rect 13078 4622 13106 13790
rect 13250 10600 13302 10606
rect 13250 10542 13302 10548
rect 13262 10266 13290 10542
rect 13250 10260 13302 10266
rect 13250 10202 13302 10208
rect 13354 7834 13382 18906
rect 13434 13932 13486 13938
rect 13434 13874 13486 13880
rect 13170 7806 13382 7834
rect 13066 4616 13118 4622
rect 13066 4558 13118 4564
rect 12974 4140 13026 4146
rect 12974 4082 13026 4088
rect 13066 4072 13118 4078
rect 13066 4014 13118 4020
rect 12894 2774 13014 2802
rect 12986 800 13014 2774
rect 13078 800 13106 4014
rect 13170 3942 13198 7806
rect 13446 7698 13474 13874
rect 13262 7670 13474 7698
rect 13262 4010 13290 7670
rect 13342 7540 13394 7546
rect 13342 7482 13394 7488
rect 13250 4004 13302 4010
rect 13250 3946 13302 3952
rect 13158 3936 13210 3942
rect 13158 3878 13210 3884
rect 13354 800 13382 7482
rect 13434 4140 13486 4146
rect 13434 4082 13486 4088
rect 13446 800 13474 4082
rect 13538 2990 13566 35974
rect 13630 4078 13658 42230
rect 13722 9382 13750 55218
rect 13814 41682 13842 59200
rect 14446 56228 14498 56234
rect 14446 56170 14498 56176
rect 14458 45558 14486 56170
rect 14814 54256 14866 54262
rect 14814 54198 14866 54204
rect 14170 45552 14222 45558
rect 14170 45494 14222 45500
rect 14446 45552 14498 45558
rect 14446 45494 14498 45500
rect 13802 41676 13854 41682
rect 13802 41618 13854 41624
rect 14182 36009 14210 45494
rect 14168 36000 14224 36009
rect 14168 35935 14224 35944
rect 14352 36000 14408 36009
rect 14352 35935 14408 35944
rect 14170 18420 14222 18426
rect 14170 18362 14222 18368
rect 13710 9376 13762 9382
rect 13710 9318 13762 9324
rect 13710 7472 13762 7478
rect 13710 7414 13762 7420
rect 13618 4072 13670 4078
rect 13618 4014 13670 4020
rect 13526 2984 13578 2990
rect 13526 2926 13578 2932
rect 13722 800 13750 7414
rect 13802 4072 13854 4078
rect 13802 4014 13854 4020
rect 13814 800 13842 4014
rect 14182 800 14210 18362
rect 14366 13138 14394 35935
rect 14538 32360 14590 32366
rect 14538 32302 14590 32308
rect 14366 13110 14486 13138
rect 14458 6118 14486 13110
rect 14550 7954 14578 32302
rect 14826 27606 14854 54198
rect 14918 30258 14946 59200
rect 15378 59158 15406 59200
rect 15090 59152 15142 59158
rect 15090 59094 15142 59100
rect 15366 59152 15418 59158
rect 15366 59094 15418 59100
rect 15102 56710 15130 59094
rect 15090 56704 15142 56710
rect 15090 56646 15142 56652
rect 15274 56704 15326 56710
rect 15274 56646 15326 56652
rect 15286 53174 15314 56646
rect 15274 53168 15326 53174
rect 15274 53110 15326 53116
rect 15734 53168 15786 53174
rect 15734 53110 15786 53116
rect 15274 53032 15326 53038
rect 15274 52974 15326 52980
rect 14998 36916 15050 36922
rect 14998 36858 15050 36864
rect 14906 30252 14958 30258
rect 14906 30194 14958 30200
rect 14814 27600 14866 27606
rect 14814 27542 14866 27548
rect 14906 27600 14958 27606
rect 14906 27542 14958 27548
rect 14630 20256 14682 20262
rect 14630 20198 14682 20204
rect 14538 7948 14590 7954
rect 14538 7890 14590 7896
rect 14538 6248 14590 6254
rect 14538 6190 14590 6196
rect 14446 6112 14498 6118
rect 14446 6054 14498 6060
rect 14446 3936 14498 3942
rect 14446 3878 14498 3884
rect 14458 800 14486 3878
rect 14550 800 14578 6190
rect 14642 4146 14670 20198
rect 14722 7948 14774 7954
rect 14722 7890 14774 7896
rect 14630 4140 14682 4146
rect 14630 4082 14682 4088
rect 14734 3534 14762 7890
rect 14814 4616 14866 4622
rect 14814 4558 14866 4564
rect 14722 3528 14774 3534
rect 14722 3470 14774 3476
rect 14826 800 14854 4558
rect 14918 800 14946 27542
rect 15010 4078 15038 36858
rect 15286 14498 15314 52974
rect 15746 37312 15774 53110
rect 15930 53038 15958 59200
rect 15918 53032 15970 53038
rect 15918 52974 15970 52980
rect 16482 42702 16510 59200
rect 16930 56364 16982 56370
rect 16930 56306 16982 56312
rect 16838 56160 16890 56166
rect 16838 56102 16890 56108
rect 16850 54874 16878 56102
rect 16942 55826 16970 56306
rect 16930 55820 16982 55826
rect 16930 55762 16982 55768
rect 16838 54868 16890 54874
rect 16838 54810 16890 54816
rect 17034 53242 17062 59200
rect 17298 56432 17350 56438
rect 17298 56374 17350 56380
rect 17114 56160 17166 56166
rect 17114 56102 17166 56108
rect 17126 55758 17154 56102
rect 17310 55758 17338 56374
rect 17114 55752 17166 55758
rect 17114 55694 17166 55700
rect 17298 55752 17350 55758
rect 17298 55694 17350 55700
rect 17390 55684 17442 55690
rect 17390 55626 17442 55632
rect 17402 55434 17430 55626
rect 17126 55406 17430 55434
rect 17126 55350 17154 55406
rect 17114 55344 17166 55350
rect 17114 55286 17166 55292
rect 17390 54528 17442 54534
rect 17390 54470 17442 54476
rect 17402 54330 17430 54470
rect 17390 54324 17442 54330
rect 17390 54266 17442 54272
rect 17022 53236 17074 53242
rect 17022 53178 17074 53184
rect 17494 51490 17522 59200
rect 17850 56704 17902 56710
rect 17850 56646 17902 56652
rect 17586 55962 17798 55978
rect 17586 55956 17810 55962
rect 17586 55950 17758 55956
rect 17586 55826 17614 55950
rect 17758 55898 17810 55904
rect 17574 55820 17626 55826
rect 17574 55762 17626 55768
rect 17666 55820 17718 55826
rect 17666 55762 17718 55768
rect 17574 55412 17626 55418
rect 17574 55354 17626 55360
rect 16574 51462 17522 51490
rect 16470 42696 16522 42702
rect 16470 42638 16522 42644
rect 16286 38888 16338 38894
rect 16286 38830 16338 38836
rect 15562 37284 15774 37312
rect 15562 29034 15590 37284
rect 16010 30048 16062 30054
rect 16010 29990 16062 29996
rect 16022 29782 16050 29990
rect 16010 29776 16062 29782
rect 16010 29718 16062 29724
rect 15550 29028 15602 29034
rect 15550 28970 15602 28976
rect 15642 29028 15694 29034
rect 15642 28970 15694 28976
rect 15550 20392 15602 20398
rect 15550 20334 15602 20340
rect 15194 14470 15314 14498
rect 15194 6866 15222 14470
rect 15562 7546 15590 20334
rect 15550 7540 15602 7546
rect 15550 7482 15602 7488
rect 15274 7472 15326 7478
rect 15274 7414 15326 7420
rect 15182 6860 15234 6866
rect 15182 6802 15234 6808
rect 14998 4072 15050 4078
rect 14998 4014 15050 4020
rect 15286 800 15314 7414
rect 15654 5166 15682 28970
rect 15826 20324 15878 20330
rect 15826 20266 15878 20272
rect 15642 5160 15694 5166
rect 15642 5102 15694 5108
rect 15458 4140 15510 4146
rect 15458 4082 15510 4088
rect 15470 800 15498 4082
rect 15642 4072 15694 4078
rect 15642 4014 15694 4020
rect 15654 800 15682 4014
rect 15838 800 15866 20266
rect 15918 19712 15970 19718
rect 15918 19654 15970 19660
rect 15930 7478 15958 19654
rect 16194 7540 16246 7546
rect 16194 7482 16246 7488
rect 15918 7472 15970 7478
rect 15918 7414 15970 7420
rect 16010 4140 16062 4146
rect 16010 4082 16062 4088
rect 16022 800 16050 4082
rect 16206 800 16234 7482
rect 16298 3924 16326 38830
rect 16470 24064 16522 24070
rect 16470 24006 16522 24012
rect 16378 19712 16430 19718
rect 16378 19654 16430 19660
rect 16390 4078 16418 19654
rect 16482 4146 16510 24006
rect 16574 6662 16602 51462
rect 17586 51354 17614 55354
rect 16850 51326 17614 51354
rect 16850 45082 16878 51326
rect 17678 51218 17706 55762
rect 17586 51190 17706 51218
rect 16838 45076 16890 45082
rect 16838 45018 16890 45024
rect 17206 42152 17258 42158
rect 17206 42094 17258 42100
rect 17218 41818 17246 42094
rect 17206 41812 17258 41818
rect 17206 41754 17258 41760
rect 17206 31204 17258 31210
rect 17206 31146 17258 31152
rect 17218 30938 17246 31146
rect 17206 30932 17258 30938
rect 17206 30874 17258 30880
rect 17206 27328 17258 27334
rect 17206 27270 17258 27276
rect 16930 21480 16982 21486
rect 16930 21422 16982 21428
rect 16838 20596 16890 20602
rect 16838 20538 16890 20544
rect 16654 16040 16706 16046
rect 16654 15982 16706 15988
rect 16666 15706 16694 15982
rect 16654 15700 16706 15706
rect 16654 15642 16706 15648
rect 16850 14550 16878 20538
rect 16838 14544 16890 14550
rect 16838 14486 16890 14492
rect 16562 6656 16614 6662
rect 16562 6598 16614 6604
rect 16746 4276 16798 4282
rect 16746 4218 16798 4224
rect 16470 4140 16522 4146
rect 16470 4082 16522 4088
rect 16378 4072 16430 4078
rect 16378 4014 16430 4020
rect 16298 3896 16418 3924
rect 16390 800 16418 3896
rect 16758 800 16786 4218
rect 16942 800 16970 21422
rect 17022 14544 17074 14550
rect 17218 14498 17246 27270
rect 17298 21548 17350 21554
rect 17298 21490 17350 21496
rect 17022 14486 17074 14492
rect 17034 4282 17062 14486
rect 17126 14470 17246 14498
rect 17126 4758 17154 14470
rect 17206 6724 17258 6730
rect 17206 6666 17258 6672
rect 17218 5914 17246 6666
rect 17206 5908 17258 5914
rect 17206 5850 17258 5856
rect 17114 4752 17166 4758
rect 17114 4694 17166 4700
rect 17022 4276 17074 4282
rect 17022 4218 17074 4224
rect 17114 4140 17166 4146
rect 17114 4082 17166 4088
rect 17126 800 17154 4082
rect 17310 800 17338 21490
rect 17390 21344 17442 21350
rect 17390 21286 17442 21292
rect 17402 2650 17430 21286
rect 17586 7546 17614 51190
rect 17574 7540 17626 7546
rect 17574 7482 17626 7488
rect 17482 6452 17534 6458
rect 17482 6394 17534 6400
rect 17390 2644 17442 2650
rect 17390 2586 17442 2592
rect 17494 800 17522 6394
rect 17862 4146 17890 56646
rect 18046 55350 18074 59200
rect 18034 55344 18086 55350
rect 18034 55286 18086 55292
rect 18598 53038 18626 59200
rect 18586 53032 18638 53038
rect 18586 52974 18638 52980
rect 19058 49366 19086 59200
rect 19610 57338 19638 59200
rect 19610 57310 19914 57338
rect 19562 57148 19858 57168
rect 19618 57146 19642 57148
rect 19698 57146 19722 57148
rect 19778 57146 19802 57148
rect 19640 57094 19642 57146
rect 19704 57094 19716 57146
rect 19778 57094 19780 57146
rect 19618 57092 19642 57094
rect 19698 57092 19722 57094
rect 19778 57092 19802 57094
rect 19562 57072 19858 57092
rect 19562 56060 19858 56080
rect 19618 56058 19642 56060
rect 19698 56058 19722 56060
rect 19778 56058 19802 56060
rect 19640 56006 19642 56058
rect 19704 56006 19716 56058
rect 19778 56006 19780 56058
rect 19618 56004 19642 56006
rect 19698 56004 19722 56006
rect 19778 56004 19802 56006
rect 19562 55984 19858 56004
rect 19886 55350 19914 57310
rect 19230 55344 19282 55350
rect 19230 55286 19282 55292
rect 19874 55344 19926 55350
rect 19874 55286 19926 55292
rect 19138 54664 19190 54670
rect 19138 54606 19190 54612
rect 19150 54534 19178 54606
rect 19138 54528 19190 54534
rect 19138 54470 19190 54476
rect 18310 49360 18362 49366
rect 18310 49302 18362 49308
rect 19046 49360 19098 49366
rect 19046 49302 19098 49308
rect 18322 37346 18350 49302
rect 18230 37318 18350 37346
rect 19138 37324 19190 37330
rect 18230 27606 18258 37318
rect 19138 37266 19190 37272
rect 19150 37233 19178 37266
rect 19136 37224 19192 37233
rect 19136 37159 19192 37168
rect 18218 27600 18270 27606
rect 18218 27542 18270 27548
rect 18310 27600 18362 27606
rect 18310 27542 18362 27548
rect 18034 22636 18086 22642
rect 18034 22578 18086 22584
rect 17942 7812 17994 7818
rect 17942 7754 17994 7760
rect 17850 4140 17902 4146
rect 17850 4082 17902 4088
rect 17954 2650 17982 7754
rect 17850 2644 17902 2650
rect 17850 2586 17902 2592
rect 17942 2644 17994 2650
rect 17942 2586 17994 2592
rect 17862 800 17890 2586
rect 18046 800 18074 22578
rect 18126 22432 18178 22438
rect 18126 22374 18178 22380
rect 18138 7818 18166 22374
rect 18322 18034 18350 27542
rect 18586 23860 18638 23866
rect 18586 23802 18638 23808
rect 18230 18006 18350 18034
rect 18230 9602 18258 18006
rect 18598 14498 18626 23802
rect 18678 22772 18730 22778
rect 18678 22714 18730 22720
rect 18506 14470 18626 14498
rect 18230 9574 18350 9602
rect 18126 7812 18178 7818
rect 18126 7754 18178 7760
rect 18322 6322 18350 9574
rect 18310 6316 18362 6322
rect 18310 6258 18362 6264
rect 18506 4010 18534 14470
rect 18586 4752 18638 4758
rect 18586 4694 18638 4700
rect 18494 4004 18546 4010
rect 18494 3946 18546 3952
rect 18126 3936 18178 3942
rect 18126 3878 18178 3884
rect 18138 1442 18166 3878
rect 18402 2644 18454 2650
rect 18402 2586 18454 2592
rect 18138 1414 18258 1442
rect 18230 800 18258 1414
rect 18414 800 18442 2586
rect 18598 800 18626 4694
rect 18690 4146 18718 22714
rect 18770 22568 18822 22574
rect 18770 22510 18822 22516
rect 18678 4140 18730 4146
rect 18678 4082 18730 4088
rect 18782 800 18810 22510
rect 18954 12912 19006 12918
rect 18954 12854 19006 12860
rect 18966 800 18994 12854
rect 19242 9178 19270 55286
rect 20162 55162 20190 59200
rect 20610 55344 20662 55350
rect 20610 55286 20662 55292
rect 19426 55134 20190 55162
rect 19426 47666 19454 55134
rect 19562 54972 19858 54992
rect 19618 54970 19642 54972
rect 19698 54970 19722 54972
rect 19778 54970 19802 54972
rect 19640 54918 19642 54970
rect 19704 54918 19716 54970
rect 19778 54918 19780 54970
rect 19618 54916 19642 54918
rect 19698 54916 19722 54918
rect 19778 54916 19802 54918
rect 19562 54896 19858 54916
rect 19562 53884 19858 53904
rect 19618 53882 19642 53884
rect 19698 53882 19722 53884
rect 19778 53882 19802 53884
rect 19640 53830 19642 53882
rect 19704 53830 19716 53882
rect 19778 53830 19780 53882
rect 19618 53828 19642 53830
rect 19698 53828 19722 53830
rect 19778 53828 19802 53830
rect 19562 53808 19858 53828
rect 19562 52796 19858 52816
rect 19618 52794 19642 52796
rect 19698 52794 19722 52796
rect 19778 52794 19802 52796
rect 19640 52742 19642 52794
rect 19704 52742 19716 52794
rect 19778 52742 19780 52794
rect 19618 52740 19642 52742
rect 19698 52740 19722 52742
rect 19778 52740 19802 52742
rect 19562 52720 19858 52740
rect 20334 52352 20386 52358
rect 20334 52294 20386 52300
rect 19562 51708 19858 51728
rect 19618 51706 19642 51708
rect 19698 51706 19722 51708
rect 19778 51706 19802 51708
rect 19640 51654 19642 51706
rect 19704 51654 19716 51706
rect 19778 51654 19780 51706
rect 19618 51652 19642 51654
rect 19698 51652 19722 51654
rect 19778 51652 19802 51654
rect 19562 51632 19858 51652
rect 19562 50620 19858 50640
rect 19618 50618 19642 50620
rect 19698 50618 19722 50620
rect 19778 50618 19802 50620
rect 19640 50566 19642 50618
rect 19704 50566 19716 50618
rect 19778 50566 19780 50618
rect 19618 50564 19642 50566
rect 19698 50564 19722 50566
rect 19778 50564 19802 50566
rect 19562 50544 19858 50564
rect 19562 49532 19858 49552
rect 19618 49530 19642 49532
rect 19698 49530 19722 49532
rect 19778 49530 19802 49532
rect 19640 49478 19642 49530
rect 19704 49478 19716 49530
rect 19778 49478 19780 49530
rect 19618 49476 19642 49478
rect 19698 49476 19722 49478
rect 19778 49476 19802 49478
rect 19562 49456 19858 49476
rect 19562 48444 19858 48464
rect 19618 48442 19642 48444
rect 19698 48442 19722 48444
rect 19778 48442 19802 48444
rect 19640 48390 19642 48442
rect 19704 48390 19716 48442
rect 19778 48390 19780 48442
rect 19618 48388 19642 48390
rect 19698 48388 19722 48390
rect 19778 48388 19802 48390
rect 19562 48368 19858 48388
rect 19414 47660 19466 47666
rect 19414 47602 19466 47608
rect 19562 47356 19858 47376
rect 19618 47354 19642 47356
rect 19698 47354 19722 47356
rect 19778 47354 19802 47356
rect 19640 47302 19642 47354
rect 19704 47302 19716 47354
rect 19778 47302 19780 47354
rect 19618 47300 19642 47302
rect 19698 47300 19722 47302
rect 19778 47300 19802 47302
rect 19562 47280 19858 47300
rect 19562 46268 19858 46288
rect 19618 46266 19642 46268
rect 19698 46266 19722 46268
rect 19778 46266 19802 46268
rect 19640 46214 19642 46266
rect 19704 46214 19716 46266
rect 19778 46214 19780 46266
rect 19618 46212 19642 46214
rect 19698 46212 19722 46214
rect 19778 46212 19802 46214
rect 19562 46192 19858 46212
rect 19562 45180 19858 45200
rect 19618 45178 19642 45180
rect 19698 45178 19722 45180
rect 19778 45178 19802 45180
rect 19640 45126 19642 45178
rect 19704 45126 19716 45178
rect 19778 45126 19780 45178
rect 19618 45124 19642 45126
rect 19698 45124 19722 45126
rect 19778 45124 19802 45126
rect 19562 45104 19858 45124
rect 19562 44092 19858 44112
rect 19618 44090 19642 44092
rect 19698 44090 19722 44092
rect 19778 44090 19802 44092
rect 19640 44038 19642 44090
rect 19704 44038 19716 44090
rect 19778 44038 19780 44090
rect 19618 44036 19642 44038
rect 19698 44036 19722 44038
rect 19778 44036 19802 44038
rect 19562 44016 19858 44036
rect 19562 43004 19858 43024
rect 19618 43002 19642 43004
rect 19698 43002 19722 43004
rect 19778 43002 19802 43004
rect 19640 42950 19642 43002
rect 19704 42950 19716 43002
rect 19778 42950 19780 43002
rect 19618 42948 19642 42950
rect 19698 42948 19722 42950
rect 19778 42948 19802 42950
rect 19562 42928 19858 42948
rect 19562 41916 19858 41936
rect 19618 41914 19642 41916
rect 19698 41914 19722 41916
rect 19778 41914 19802 41916
rect 19640 41862 19642 41914
rect 19704 41862 19716 41914
rect 19778 41862 19780 41914
rect 19618 41860 19642 41862
rect 19698 41860 19722 41862
rect 19778 41860 19802 41862
rect 19562 41840 19858 41860
rect 19562 40828 19858 40848
rect 19618 40826 19642 40828
rect 19698 40826 19722 40828
rect 19778 40826 19802 40828
rect 19640 40774 19642 40826
rect 19704 40774 19716 40826
rect 19778 40774 19780 40826
rect 19618 40772 19642 40774
rect 19698 40772 19722 40774
rect 19778 40772 19802 40774
rect 19562 40752 19858 40772
rect 19562 39740 19858 39760
rect 19618 39738 19642 39740
rect 19698 39738 19722 39740
rect 19778 39738 19802 39740
rect 19640 39686 19642 39738
rect 19704 39686 19716 39738
rect 19778 39686 19780 39738
rect 19618 39684 19642 39686
rect 19698 39684 19722 39686
rect 19778 39684 19802 39686
rect 19562 39664 19858 39684
rect 19562 38652 19858 38672
rect 19618 38650 19642 38652
rect 19698 38650 19722 38652
rect 19778 38650 19802 38652
rect 19640 38598 19642 38650
rect 19704 38598 19716 38650
rect 19778 38598 19780 38650
rect 19618 38596 19642 38598
rect 19698 38596 19722 38598
rect 19778 38596 19802 38598
rect 19562 38576 19858 38596
rect 19562 37564 19858 37584
rect 19618 37562 19642 37564
rect 19698 37562 19722 37564
rect 19778 37562 19802 37564
rect 19640 37510 19642 37562
rect 19704 37510 19716 37562
rect 19778 37510 19780 37562
rect 19618 37508 19642 37510
rect 19698 37508 19722 37510
rect 19778 37508 19802 37510
rect 19562 37488 19858 37508
rect 19562 36476 19858 36496
rect 19618 36474 19642 36476
rect 19698 36474 19722 36476
rect 19778 36474 19802 36476
rect 19640 36422 19642 36474
rect 19704 36422 19716 36474
rect 19778 36422 19780 36474
rect 19618 36420 19642 36422
rect 19698 36420 19722 36422
rect 19778 36420 19802 36422
rect 19562 36400 19858 36420
rect 19562 35388 19858 35408
rect 19618 35386 19642 35388
rect 19698 35386 19722 35388
rect 19778 35386 19802 35388
rect 19640 35334 19642 35386
rect 19704 35334 19716 35386
rect 19778 35334 19780 35386
rect 19618 35332 19642 35334
rect 19698 35332 19722 35334
rect 19778 35332 19802 35334
rect 19562 35312 19858 35332
rect 19562 34300 19858 34320
rect 19618 34298 19642 34300
rect 19698 34298 19722 34300
rect 19778 34298 19802 34300
rect 19640 34246 19642 34298
rect 19704 34246 19716 34298
rect 19778 34246 19780 34298
rect 19618 34244 19642 34246
rect 19698 34244 19722 34246
rect 19778 34244 19802 34246
rect 19562 34224 19858 34244
rect 19562 33212 19858 33232
rect 19618 33210 19642 33212
rect 19698 33210 19722 33212
rect 19778 33210 19802 33212
rect 19640 33158 19642 33210
rect 19704 33158 19716 33210
rect 19778 33158 19780 33210
rect 19618 33156 19642 33158
rect 19698 33156 19722 33158
rect 19778 33156 19802 33158
rect 19562 33136 19858 33156
rect 19562 32124 19858 32144
rect 19618 32122 19642 32124
rect 19698 32122 19722 32124
rect 19778 32122 19802 32124
rect 19640 32070 19642 32122
rect 19704 32070 19716 32122
rect 19778 32070 19780 32122
rect 19618 32068 19642 32070
rect 19698 32068 19722 32070
rect 19778 32068 19802 32070
rect 19562 32048 19858 32068
rect 19562 31036 19858 31056
rect 19618 31034 19642 31036
rect 19698 31034 19722 31036
rect 19778 31034 19802 31036
rect 19640 30982 19642 31034
rect 19704 30982 19716 31034
rect 19778 30982 19780 31034
rect 19618 30980 19642 30982
rect 19698 30980 19722 30982
rect 19778 30980 19802 30982
rect 19562 30960 19858 30980
rect 19562 29948 19858 29968
rect 19618 29946 19642 29948
rect 19698 29946 19722 29948
rect 19778 29946 19802 29948
rect 19640 29894 19642 29946
rect 19704 29894 19716 29946
rect 19778 29894 19780 29946
rect 19618 29892 19642 29894
rect 19698 29892 19722 29894
rect 19778 29892 19802 29894
rect 19562 29872 19858 29892
rect 19562 28860 19858 28880
rect 19618 28858 19642 28860
rect 19698 28858 19722 28860
rect 19778 28858 19802 28860
rect 19640 28806 19642 28858
rect 19704 28806 19716 28858
rect 19778 28806 19780 28858
rect 19618 28804 19642 28806
rect 19698 28804 19722 28806
rect 19778 28804 19802 28806
rect 19562 28784 19858 28804
rect 19562 27772 19858 27792
rect 19618 27770 19642 27772
rect 19698 27770 19722 27772
rect 19778 27770 19802 27772
rect 19640 27718 19642 27770
rect 19704 27718 19716 27770
rect 19778 27718 19780 27770
rect 19618 27716 19642 27718
rect 19698 27716 19722 27718
rect 19778 27716 19802 27718
rect 19562 27696 19858 27716
rect 19562 26684 19858 26704
rect 19618 26682 19642 26684
rect 19698 26682 19722 26684
rect 19778 26682 19802 26684
rect 19640 26630 19642 26682
rect 19704 26630 19716 26682
rect 19778 26630 19780 26682
rect 19618 26628 19642 26630
rect 19698 26628 19722 26630
rect 19778 26628 19802 26630
rect 19562 26608 19858 26628
rect 19562 25596 19858 25616
rect 19618 25594 19642 25596
rect 19698 25594 19722 25596
rect 19778 25594 19802 25596
rect 19640 25542 19642 25594
rect 19704 25542 19716 25594
rect 19778 25542 19780 25594
rect 19618 25540 19642 25542
rect 19698 25540 19722 25542
rect 19778 25540 19802 25542
rect 19562 25520 19858 25540
rect 20058 25492 20110 25498
rect 20058 25434 20110 25440
rect 19966 24948 20018 24954
rect 19966 24890 20018 24896
rect 19562 24508 19858 24528
rect 19618 24506 19642 24508
rect 19698 24506 19722 24508
rect 19778 24506 19802 24508
rect 19640 24454 19642 24506
rect 19704 24454 19716 24506
rect 19778 24454 19780 24506
rect 19618 24452 19642 24454
rect 19698 24452 19722 24454
rect 19778 24452 19802 24454
rect 19562 24432 19858 24452
rect 19874 23656 19926 23662
rect 19874 23598 19926 23604
rect 19562 23420 19858 23440
rect 19618 23418 19642 23420
rect 19698 23418 19722 23420
rect 19778 23418 19802 23420
rect 19640 23366 19642 23418
rect 19704 23366 19716 23418
rect 19778 23366 19780 23418
rect 19618 23364 19642 23366
rect 19698 23364 19722 23366
rect 19778 23364 19802 23366
rect 19562 23344 19858 23364
rect 19562 22332 19858 22352
rect 19618 22330 19642 22332
rect 19698 22330 19722 22332
rect 19778 22330 19802 22332
rect 19640 22278 19642 22330
rect 19704 22278 19716 22330
rect 19778 22278 19780 22330
rect 19618 22276 19642 22278
rect 19698 22276 19722 22278
rect 19778 22276 19802 22278
rect 19562 22256 19858 22276
rect 19562 21244 19858 21264
rect 19618 21242 19642 21244
rect 19698 21242 19722 21244
rect 19778 21242 19802 21244
rect 19640 21190 19642 21242
rect 19704 21190 19716 21242
rect 19778 21190 19780 21242
rect 19618 21188 19642 21190
rect 19698 21188 19722 21190
rect 19778 21188 19802 21190
rect 19562 21168 19858 21188
rect 19562 20156 19858 20176
rect 19618 20154 19642 20156
rect 19698 20154 19722 20156
rect 19778 20154 19802 20156
rect 19640 20102 19642 20154
rect 19704 20102 19716 20154
rect 19778 20102 19780 20154
rect 19618 20100 19642 20102
rect 19698 20100 19722 20102
rect 19778 20100 19802 20102
rect 19562 20080 19858 20100
rect 19562 19068 19858 19088
rect 19618 19066 19642 19068
rect 19698 19066 19722 19068
rect 19778 19066 19802 19068
rect 19640 19014 19642 19066
rect 19704 19014 19716 19066
rect 19778 19014 19780 19066
rect 19618 19012 19642 19014
rect 19698 19012 19722 19014
rect 19778 19012 19802 19014
rect 19562 18992 19858 19012
rect 19562 17980 19858 18000
rect 19618 17978 19642 17980
rect 19698 17978 19722 17980
rect 19778 17978 19802 17980
rect 19640 17926 19642 17978
rect 19704 17926 19716 17978
rect 19778 17926 19780 17978
rect 19618 17924 19642 17926
rect 19698 17924 19722 17926
rect 19778 17924 19802 17926
rect 19562 17904 19858 17924
rect 19562 16892 19858 16912
rect 19618 16890 19642 16892
rect 19698 16890 19722 16892
rect 19778 16890 19802 16892
rect 19640 16838 19642 16890
rect 19704 16838 19716 16890
rect 19778 16838 19780 16890
rect 19618 16836 19642 16838
rect 19698 16836 19722 16838
rect 19778 16836 19802 16838
rect 19562 16816 19858 16836
rect 19562 15804 19858 15824
rect 19618 15802 19642 15804
rect 19698 15802 19722 15804
rect 19778 15802 19802 15804
rect 19640 15750 19642 15802
rect 19704 15750 19716 15802
rect 19778 15750 19780 15802
rect 19618 15748 19642 15750
rect 19698 15748 19722 15750
rect 19778 15748 19802 15750
rect 19562 15728 19858 15748
rect 19562 14716 19858 14736
rect 19618 14714 19642 14716
rect 19698 14714 19722 14716
rect 19778 14714 19802 14716
rect 19640 14662 19642 14714
rect 19704 14662 19716 14714
rect 19778 14662 19780 14714
rect 19618 14660 19642 14662
rect 19698 14660 19722 14662
rect 19778 14660 19802 14662
rect 19562 14640 19858 14660
rect 19562 13628 19858 13648
rect 19618 13626 19642 13628
rect 19698 13626 19722 13628
rect 19778 13626 19802 13628
rect 19640 13574 19642 13626
rect 19704 13574 19716 13626
rect 19778 13574 19780 13626
rect 19618 13572 19642 13574
rect 19698 13572 19722 13574
rect 19778 13572 19802 13574
rect 19562 13552 19858 13572
rect 19562 12540 19858 12560
rect 19618 12538 19642 12540
rect 19698 12538 19722 12540
rect 19778 12538 19802 12540
rect 19640 12486 19642 12538
rect 19704 12486 19716 12538
rect 19778 12486 19780 12538
rect 19618 12484 19642 12486
rect 19698 12484 19722 12486
rect 19778 12484 19802 12486
rect 19562 12464 19858 12484
rect 19562 11452 19858 11472
rect 19618 11450 19642 11452
rect 19698 11450 19722 11452
rect 19778 11450 19802 11452
rect 19640 11398 19642 11450
rect 19704 11398 19716 11450
rect 19778 11398 19780 11450
rect 19618 11396 19642 11398
rect 19698 11396 19722 11398
rect 19778 11396 19802 11398
rect 19562 11376 19858 11396
rect 19562 10364 19858 10384
rect 19618 10362 19642 10364
rect 19698 10362 19722 10364
rect 19778 10362 19802 10364
rect 19640 10310 19642 10362
rect 19704 10310 19716 10362
rect 19778 10310 19780 10362
rect 19618 10308 19642 10310
rect 19698 10308 19722 10310
rect 19778 10308 19802 10310
rect 19562 10288 19858 10308
rect 19562 9276 19858 9296
rect 19618 9274 19642 9276
rect 19698 9274 19722 9276
rect 19778 9274 19802 9276
rect 19640 9222 19642 9274
rect 19704 9222 19716 9274
rect 19778 9222 19780 9274
rect 19618 9220 19642 9222
rect 19698 9220 19722 9222
rect 19778 9220 19802 9222
rect 19562 9200 19858 9220
rect 19230 9172 19282 9178
rect 19230 9114 19282 9120
rect 19562 8188 19858 8208
rect 19618 8186 19642 8188
rect 19698 8186 19722 8188
rect 19778 8186 19802 8188
rect 19640 8134 19642 8186
rect 19704 8134 19716 8186
rect 19778 8134 19780 8186
rect 19618 8132 19642 8134
rect 19698 8132 19722 8134
rect 19778 8132 19802 8134
rect 19562 8112 19858 8132
rect 19562 7100 19858 7120
rect 19618 7098 19642 7100
rect 19698 7098 19722 7100
rect 19778 7098 19802 7100
rect 19640 7046 19642 7098
rect 19704 7046 19716 7098
rect 19778 7046 19780 7098
rect 19618 7044 19642 7046
rect 19698 7044 19722 7046
rect 19778 7044 19802 7046
rect 19562 7024 19858 7044
rect 19562 6012 19858 6032
rect 19618 6010 19642 6012
rect 19698 6010 19722 6012
rect 19778 6010 19802 6012
rect 19640 5958 19642 6010
rect 19704 5958 19716 6010
rect 19778 5958 19780 6010
rect 19618 5956 19642 5958
rect 19698 5956 19722 5958
rect 19778 5956 19802 5958
rect 19562 5936 19858 5956
rect 19562 4924 19858 4944
rect 19618 4922 19642 4924
rect 19698 4922 19722 4924
rect 19778 4922 19802 4924
rect 19640 4870 19642 4922
rect 19704 4870 19716 4922
rect 19778 4870 19780 4922
rect 19618 4868 19642 4870
rect 19698 4868 19722 4870
rect 19778 4868 19802 4870
rect 19562 4848 19858 4868
rect 19322 4140 19374 4146
rect 19322 4082 19374 4088
rect 19334 800 19362 4082
rect 19562 3836 19858 3856
rect 19618 3834 19642 3836
rect 19698 3834 19722 3836
rect 19778 3834 19802 3836
rect 19640 3782 19642 3834
rect 19704 3782 19716 3834
rect 19778 3782 19780 3834
rect 19618 3780 19642 3782
rect 19698 3780 19722 3782
rect 19778 3780 19802 3782
rect 19562 3760 19858 3780
rect 19562 2748 19858 2768
rect 19618 2746 19642 2748
rect 19698 2746 19722 2748
rect 19778 2746 19802 2748
rect 19640 2694 19642 2746
rect 19704 2694 19716 2746
rect 19778 2694 19780 2746
rect 19618 2692 19642 2694
rect 19698 2692 19722 2694
rect 19778 2692 19802 2694
rect 19562 2672 19858 2692
rect 19886 1306 19914 23598
rect 19978 7698 20006 24890
rect 20070 8294 20098 25434
rect 20242 23520 20294 23526
rect 20242 23462 20294 23468
rect 20150 13864 20202 13870
rect 20150 13806 20202 13812
rect 20162 8362 20190 13806
rect 20150 8356 20202 8362
rect 20150 8298 20202 8304
rect 20058 8288 20110 8294
rect 20058 8230 20110 8236
rect 19978 7670 20098 7698
rect 19966 7540 20018 7546
rect 19966 7482 20018 7488
rect 19518 1278 19914 1306
rect 19518 800 19546 1278
rect 19690 1148 19742 1154
rect 19690 1090 19742 1096
rect 19702 800 19730 1090
rect 19978 898 20006 7482
rect 20070 5030 20098 7670
rect 20058 5024 20110 5030
rect 20058 4966 20110 4972
rect 20058 4820 20110 4826
rect 20058 4762 20110 4768
rect 19886 870 20006 898
rect 19886 800 19914 870
rect 20070 800 20098 4762
rect 20254 800 20282 23462
rect 20346 4826 20374 52294
rect 20622 26382 20650 55286
rect 20714 55162 20742 59200
rect 21174 56438 21202 59200
rect 21726 56506 21754 59200
rect 21714 56500 21766 56506
rect 21714 56442 21766 56448
rect 21162 56432 21214 56438
rect 21162 56374 21214 56380
rect 21990 56432 22042 56438
rect 21990 56374 22042 56380
rect 20794 56228 20846 56234
rect 20794 56170 20846 56176
rect 20886 56228 20938 56234
rect 20886 56170 20938 56176
rect 20806 55418 20834 56170
rect 20898 55690 20926 56170
rect 20886 55684 20938 55690
rect 20886 55626 20938 55632
rect 21346 55684 21398 55690
rect 21346 55626 21398 55632
rect 20794 55412 20846 55418
rect 20794 55354 20846 55360
rect 20714 55134 21294 55162
rect 21162 30592 21214 30598
rect 21162 30534 21214 30540
rect 20610 26376 20662 26382
rect 20610 26318 20662 26324
rect 21070 24812 21122 24818
rect 21070 24754 21122 24760
rect 20794 24404 20846 24410
rect 20794 24346 20846 24352
rect 20426 23724 20478 23730
rect 20426 23666 20478 23672
rect 20438 7546 20466 23666
rect 20610 22976 20662 22982
rect 20610 22918 20662 22924
rect 20518 8356 20570 8362
rect 20518 8298 20570 8304
rect 20426 7540 20478 7546
rect 20426 7482 20478 7488
rect 20334 4820 20386 4826
rect 20334 4762 20386 4768
rect 20426 4276 20478 4282
rect 20426 4218 20478 4224
rect 20438 3942 20466 4218
rect 20426 3936 20478 3942
rect 20426 3878 20478 3884
rect 20530 3058 20558 8298
rect 20518 3052 20570 3058
rect 20518 2994 20570 3000
rect 20622 2938 20650 22918
rect 20702 4004 20754 4010
rect 20702 3946 20754 3952
rect 20438 2910 20650 2938
rect 20438 800 20466 2910
rect 20714 1442 20742 3946
rect 20806 1562 20834 24346
rect 21082 19310 21110 24754
rect 20978 19304 21030 19310
rect 20978 19246 21030 19252
rect 21070 19304 21122 19310
rect 21070 19246 21122 19252
rect 20886 7540 20938 7546
rect 20886 7482 20938 7488
rect 20794 1556 20846 1562
rect 20794 1498 20846 1504
rect 20714 1414 20834 1442
rect 20806 800 20834 1414
rect 20898 1154 20926 7482
rect 20886 1148 20938 1154
rect 20886 1090 20938 1096
rect 20990 800 21018 19246
rect 21174 4842 21202 30534
rect 21266 14498 21294 55134
rect 21358 19378 21386 55626
rect 21438 54732 21490 54738
rect 21438 54674 21490 54680
rect 21450 54534 21478 54674
rect 21438 54528 21490 54534
rect 21438 54470 21490 54476
rect 21622 54528 21674 54534
rect 21622 54470 21674 54476
rect 21634 54194 21662 54470
rect 21622 54188 21674 54194
rect 21622 54130 21674 54136
rect 21898 37732 21950 37738
rect 21898 37674 21950 37680
rect 21806 33856 21858 33862
rect 21806 33798 21858 33804
rect 21438 27872 21490 27878
rect 21438 27814 21490 27820
rect 21346 19372 21398 19378
rect 21346 19314 21398 19320
rect 21266 14470 21386 14498
rect 21358 6390 21386 14470
rect 21346 6384 21398 6390
rect 21346 6326 21398 6332
rect 21174 4814 21386 4842
rect 21162 4004 21214 4010
rect 21162 3946 21214 3952
rect 21174 800 21202 3946
rect 21358 3516 21386 4814
rect 21450 4146 21478 27814
rect 21530 26784 21582 26790
rect 21530 26726 21582 26732
rect 21438 4140 21490 4146
rect 21438 4082 21490 4088
rect 21542 3670 21570 26726
rect 21714 24676 21766 24682
rect 21714 24618 21766 24624
rect 21530 3664 21582 3670
rect 21530 3606 21582 3612
rect 21358 3488 21570 3516
rect 21346 1556 21398 1562
rect 21346 1498 21398 1504
rect 21358 800 21386 1498
rect 21542 800 21570 3488
rect 21726 800 21754 24618
rect 21818 4010 21846 33798
rect 21806 4004 21858 4010
rect 21806 3946 21858 3952
rect 21910 800 21938 37674
rect 22002 12646 22030 56374
rect 22738 55826 22766 59200
rect 22818 56432 22870 56438
rect 22818 56374 22870 56380
rect 22726 55820 22778 55826
rect 22726 55762 22778 55768
rect 22830 55162 22858 56374
rect 22910 55820 22962 55826
rect 22910 55762 22962 55768
rect 22738 55134 22858 55162
rect 22738 30802 22766 55134
rect 22922 55026 22950 55762
rect 23290 55418 23318 59200
rect 23842 59158 23870 59200
rect 23830 59152 23882 59158
rect 23830 59094 23882 59100
rect 23830 57928 23882 57934
rect 23830 57870 23882 57876
rect 23842 56658 23870 57870
rect 23750 56630 23870 56658
rect 23278 55412 23330 55418
rect 23278 55354 23330 55360
rect 22830 54998 22950 55026
rect 22830 33522 22858 54998
rect 23750 48362 23778 56630
rect 24290 56500 24342 56506
rect 24290 56442 24342 56448
rect 24106 55344 24158 55350
rect 24106 55286 24158 55292
rect 23658 48334 23778 48362
rect 23370 44532 23422 44538
rect 23370 44474 23422 44480
rect 23278 40112 23330 40118
rect 23278 40054 23330 40060
rect 22818 33516 22870 33522
rect 22818 33458 22870 33464
rect 22726 30796 22778 30802
rect 22726 30738 22778 30744
rect 22726 28960 22778 28966
rect 22726 28902 22778 28908
rect 22542 25696 22594 25702
rect 22542 25638 22594 25644
rect 22082 24744 22134 24750
rect 22082 24686 22134 24692
rect 21990 12640 22042 12646
rect 21990 12582 22042 12588
rect 22094 800 22122 24686
rect 22554 14362 22582 25638
rect 22738 14498 22766 28902
rect 22910 25764 22962 25770
rect 22910 25706 22962 25712
rect 22922 19310 22950 25706
rect 22910 19304 22962 19310
rect 22910 19246 22962 19252
rect 23094 19304 23146 19310
rect 23094 19246 23146 19252
rect 22738 14470 22858 14498
rect 22554 14334 22766 14362
rect 22634 5024 22686 5030
rect 22634 4966 22686 4972
rect 22174 4140 22226 4146
rect 22174 4082 22226 4088
rect 22266 4140 22318 4146
rect 22266 4082 22318 4088
rect 22186 3738 22214 4082
rect 22174 3732 22226 3738
rect 22174 3674 22226 3680
rect 22278 800 22306 4082
rect 22646 800 22674 4966
rect 22738 3346 22766 14334
rect 22830 3466 22858 14470
rect 23002 4140 23054 4146
rect 23002 4082 23054 4088
rect 22818 3460 22870 3466
rect 22818 3402 22870 3408
rect 22738 3318 22858 3346
rect 22830 800 22858 3318
rect 23014 800 23042 4082
rect 23106 3924 23134 19246
rect 23186 18216 23238 18222
rect 23186 18158 23238 18164
rect 23198 4026 23226 18158
rect 23290 4146 23318 40054
rect 23382 4146 23410 44474
rect 23658 37312 23686 48334
rect 23566 37284 23686 37312
rect 23566 37210 23594 37284
rect 23566 37182 23686 37210
rect 23658 31754 23686 37182
rect 23462 31748 23514 31754
rect 23462 31690 23514 31696
rect 23646 31748 23698 31754
rect 23646 31690 23698 31696
rect 23474 27554 23502 31690
rect 23474 27526 23594 27554
rect 23566 18086 23594 27526
rect 23646 26988 23698 26994
rect 23646 26930 23698 26936
rect 23658 19310 23686 26930
rect 23646 19304 23698 19310
rect 23646 19246 23698 19252
rect 23922 19304 23974 19310
rect 23922 19246 23974 19252
rect 23462 18080 23514 18086
rect 23462 18022 23514 18028
rect 23554 18080 23606 18086
rect 23554 18022 23606 18028
rect 23474 7410 23502 18022
rect 23738 8288 23790 8294
rect 23738 8230 23790 8236
rect 23462 7404 23514 7410
rect 23462 7346 23514 7352
rect 23278 4140 23330 4146
rect 23278 4082 23330 4088
rect 23370 4140 23422 4146
rect 23370 4082 23422 4088
rect 23198 3998 23410 4026
rect 23106 3896 23226 3924
rect 23198 800 23226 3896
rect 23382 800 23410 3998
rect 23750 800 23778 8230
rect 23934 800 23962 19246
rect 24118 7206 24146 55286
rect 24198 55208 24250 55214
rect 24198 55150 24250 55156
rect 24210 47462 24238 55150
rect 24198 47456 24250 47462
rect 24198 47398 24250 47404
rect 24198 40180 24250 40186
rect 24198 40122 24250 40128
rect 24106 7200 24158 7206
rect 24106 7142 24158 7148
rect 24106 4140 24158 4146
rect 24106 4082 24158 4088
rect 24118 800 24146 4082
rect 24210 2990 24238 40122
rect 24302 31822 24330 56442
rect 24394 55758 24422 59200
rect 24854 56370 24882 59200
rect 24842 56364 24894 56370
rect 24842 56306 24894 56312
rect 24934 56364 24986 56370
rect 24934 56306 24986 56312
rect 24946 55826 24974 56306
rect 25484 56264 25540 56273
rect 25484 56199 25540 56208
rect 24934 55820 24986 55826
rect 24934 55762 24986 55768
rect 24382 55752 24434 55758
rect 24382 55694 24434 55700
rect 25210 55684 25262 55690
rect 25210 55626 25262 55632
rect 25222 55282 25250 55626
rect 25210 55276 25262 55282
rect 25210 55218 25262 55224
rect 24750 46980 24802 46986
rect 24750 46922 24802 46928
rect 24290 31816 24342 31822
rect 24290 31758 24342 31764
rect 24290 30048 24342 30054
rect 24290 29990 24342 29996
rect 24302 3602 24330 29990
rect 24382 26920 24434 26926
rect 24382 26862 24434 26868
rect 24290 3596 24342 3602
rect 24290 3538 24342 3544
rect 24394 3482 24422 26862
rect 24762 4146 24790 46922
rect 25118 29300 25170 29306
rect 25118 29242 25170 29248
rect 24842 7744 24894 7750
rect 24842 7686 24894 7692
rect 25026 7744 25078 7750
rect 25026 7686 25078 7692
rect 24750 4140 24802 4146
rect 24750 4082 24802 4088
rect 24854 4078 24882 7686
rect 24842 4072 24894 4078
rect 24842 4014 24894 4020
rect 24842 3664 24894 3670
rect 24842 3606 24894 3612
rect 24302 3454 24422 3482
rect 24198 2984 24250 2990
rect 24198 2926 24250 2932
rect 24302 800 24330 3454
rect 24474 3052 24526 3058
rect 24474 2994 24526 3000
rect 24486 800 24514 2994
rect 24854 800 24882 3606
rect 25038 800 25066 7686
rect 25130 4010 25158 29242
rect 25394 28076 25446 28082
rect 25394 28018 25446 28024
rect 25210 9172 25262 9178
rect 25210 9114 25262 9120
rect 25118 4004 25170 4010
rect 25118 3946 25170 3952
rect 25222 800 25250 9114
rect 25406 800 25434 28018
rect 25498 15162 25526 56199
rect 25670 55820 25722 55826
rect 25670 55762 25722 55768
rect 25578 55276 25630 55282
rect 25578 55218 25630 55224
rect 25590 34678 25618 55218
rect 25578 34672 25630 34678
rect 25578 34614 25630 34620
rect 25578 31136 25630 31142
rect 25578 31078 25630 31084
rect 25590 27690 25618 31078
rect 25682 30326 25710 55762
rect 25958 55758 25986 59200
rect 26130 55820 26182 55826
rect 26130 55762 26182 55768
rect 25946 55752 25998 55758
rect 25946 55694 25998 55700
rect 26142 55214 26170 55762
rect 26418 55350 26446 59200
rect 26406 55344 26458 55350
rect 26406 55286 26458 55292
rect 26130 55208 26182 55214
rect 26130 55150 26182 55156
rect 26970 53174 26998 59200
rect 27050 55344 27102 55350
rect 27050 55286 27102 55292
rect 26498 53168 26550 53174
rect 26498 53110 26550 53116
rect 26958 53168 27010 53174
rect 26958 53110 27010 53116
rect 26510 46918 26538 53110
rect 27062 52714 27090 55286
rect 26970 52686 27090 52714
rect 26406 46912 26458 46918
rect 26406 46854 26458 46860
rect 26498 46912 26550 46918
rect 26498 46854 26550 46860
rect 26418 37330 26446 46854
rect 26866 44736 26918 44742
rect 26866 44678 26918 44684
rect 26406 37324 26458 37330
rect 26406 37266 26458 37272
rect 26498 37324 26550 37330
rect 26498 37266 26550 37272
rect 25670 30320 25722 30326
rect 25670 30262 25722 30268
rect 26130 30116 26182 30122
rect 26130 30058 26182 30064
rect 25854 28008 25906 28014
rect 25854 27950 25906 27956
rect 25590 27662 25710 27690
rect 25682 26246 25710 27662
rect 25670 26240 25722 26246
rect 25670 26182 25722 26188
rect 25762 26240 25814 26246
rect 25762 26182 25814 26188
rect 25774 16658 25802 26182
rect 25866 18057 25894 27950
rect 25852 18048 25908 18057
rect 25852 17983 25908 17992
rect 25852 17912 25908 17921
rect 25852 17847 25908 17856
rect 25762 16652 25814 16658
rect 25762 16594 25814 16600
rect 25486 15156 25538 15162
rect 25486 15098 25538 15104
rect 25670 8356 25722 8362
rect 25670 8298 25722 8304
rect 25578 4140 25630 4146
rect 25578 4082 25630 4088
rect 25590 800 25618 4082
rect 25682 3942 25710 8298
rect 25866 7750 25894 17847
rect 25946 16652 25998 16658
rect 25946 16594 25998 16600
rect 25958 8362 25986 16594
rect 25946 8356 25998 8362
rect 25946 8298 25998 8304
rect 25854 7744 25906 7750
rect 25854 7686 25906 7692
rect 26142 4146 26170 30058
rect 26510 27606 26538 37266
rect 26682 37120 26734 37126
rect 26682 37062 26734 37068
rect 26694 36922 26722 37062
rect 26682 36916 26734 36922
rect 26682 36858 26734 36864
rect 26682 29504 26734 29510
rect 26682 29446 26734 29452
rect 26694 29306 26722 29446
rect 26682 29300 26734 29306
rect 26682 29242 26734 29248
rect 26498 27600 26550 27606
rect 26498 27542 26550 27548
rect 26590 27600 26642 27606
rect 26590 27542 26642 27548
rect 26602 8566 26630 27542
rect 26774 18692 26826 18698
rect 26774 18634 26826 18640
rect 26786 18290 26814 18634
rect 26774 18284 26826 18290
rect 26774 18226 26826 18232
rect 26590 8560 26642 8566
rect 26590 8502 26642 8508
rect 26682 7812 26734 7818
rect 26682 7754 26734 7760
rect 26498 7744 26550 7750
rect 26498 7686 26550 7692
rect 26130 4140 26182 4146
rect 26130 4082 26182 4088
rect 26314 4072 26366 4078
rect 26314 4014 26366 4020
rect 26130 4004 26182 4010
rect 26130 3946 26182 3952
rect 25670 3936 25722 3942
rect 25670 3878 25722 3884
rect 25946 3732 25998 3738
rect 25946 3674 25998 3680
rect 25958 800 25986 3674
rect 26142 800 26170 3946
rect 26326 800 26354 4014
rect 26510 800 26538 7686
rect 26694 800 26722 7754
rect 26878 3670 26906 44678
rect 26970 40050 26998 52686
rect 27050 41812 27102 41818
rect 27050 41754 27102 41760
rect 26958 40044 27010 40050
rect 26958 39986 27010 39992
rect 27062 4078 27090 41754
rect 27522 37330 27550 59200
rect 28074 56438 28102 59200
rect 28062 56432 28114 56438
rect 28062 56374 28114 56380
rect 28154 56432 28206 56438
rect 28154 56374 28206 56380
rect 28166 55826 28194 56374
rect 29086 56370 29114 59200
rect 29074 56364 29126 56370
rect 29074 56306 29126 56312
rect 28154 55820 28206 55826
rect 28154 55762 28206 55768
rect 28338 55820 28390 55826
rect 28338 55762 28390 55768
rect 27602 54732 27654 54738
rect 27602 54674 27654 54680
rect 27614 54534 27642 54674
rect 27602 54528 27654 54534
rect 27602 54470 27654 54476
rect 28246 38208 28298 38214
rect 28246 38150 28298 38156
rect 27510 37324 27562 37330
rect 27510 37266 27562 37272
rect 27786 37256 27838 37262
rect 27784 37224 27786 37233
rect 27838 37224 27840 37233
rect 27784 37159 27840 37168
rect 27234 29844 27286 29850
rect 27234 29786 27286 29792
rect 27142 14952 27194 14958
rect 27142 14894 27194 14900
rect 27154 4146 27182 14894
rect 27142 4140 27194 4146
rect 27142 4082 27194 4088
rect 27050 4072 27102 4078
rect 27050 4014 27102 4020
rect 26866 3664 26918 3670
rect 26866 3606 26918 3612
rect 26866 3528 26918 3534
rect 26866 3470 26918 3476
rect 26878 3126 26906 3470
rect 27050 3460 27102 3466
rect 27050 3402 27102 3408
rect 26866 3120 26918 3126
rect 26866 3062 26918 3068
rect 27062 800 27090 3402
rect 27246 800 27274 29786
rect 27602 29708 27654 29714
rect 27602 29650 27654 29656
rect 27326 29096 27378 29102
rect 27326 29038 27378 29044
rect 27338 7750 27366 29038
rect 27430 8498 27550 8514
rect 27418 8492 27562 8498
rect 27470 8486 27510 8492
rect 27418 8434 27470 8440
rect 27510 8434 27562 8440
rect 27326 7744 27378 7750
rect 27326 7686 27378 7692
rect 27418 2848 27470 2854
rect 27418 2790 27470 2796
rect 27430 800 27458 2790
rect 27614 800 27642 29650
rect 28258 28218 28286 38150
rect 28062 28212 28114 28218
rect 28062 28154 28114 28160
rect 28246 28212 28298 28218
rect 28246 28154 28298 28160
rect 28074 27674 28102 28154
rect 28062 27668 28114 27674
rect 28062 27610 28114 27616
rect 28154 27668 28206 27674
rect 28154 27610 28206 27616
rect 28166 8294 28194 27610
rect 28350 21010 28378 55762
rect 29638 55298 29666 59200
rect 29994 56704 30046 56710
rect 29994 56646 30046 56652
rect 30006 56506 30034 56646
rect 29994 56500 30046 56506
rect 29994 56442 30046 56448
rect 29718 56364 29770 56370
rect 29718 56306 29770 56312
rect 29086 55270 29666 55298
rect 28798 30932 28850 30938
rect 28798 30874 28850 30880
rect 28706 30864 28758 30870
rect 28706 30806 28758 30812
rect 28430 22228 28482 22234
rect 28430 22170 28482 22176
rect 28338 21004 28390 21010
rect 28338 20946 28390 20952
rect 28338 18624 28390 18630
rect 28338 18566 28390 18572
rect 28154 8288 28206 8294
rect 28154 8230 28206 8236
rect 28350 7834 28378 18566
rect 28442 12322 28470 22170
rect 28614 20392 28666 20398
rect 28614 20334 28666 20340
rect 28626 20058 28654 20334
rect 28614 20052 28666 20058
rect 28614 19994 28666 20000
rect 28442 12294 28654 12322
rect 28350 7806 28470 7834
rect 28338 7744 28390 7750
rect 28338 7686 28390 7692
rect 27694 6656 27746 6662
rect 27694 6598 27746 6604
rect 27706 6390 27734 6598
rect 27694 6384 27746 6390
rect 27694 6326 27746 6332
rect 27786 4140 27838 4146
rect 27786 4082 27838 4088
rect 27798 800 27826 4082
rect 28154 3596 28206 3602
rect 28154 3538 28206 3544
rect 28166 800 28194 3538
rect 28350 800 28378 7686
rect 28442 3058 28470 7806
rect 28522 3460 28574 3466
rect 28522 3402 28574 3408
rect 28430 3052 28482 3058
rect 28430 2994 28482 3000
rect 28534 800 28562 3402
rect 28626 2922 28654 12294
rect 28614 2916 28666 2922
rect 28614 2858 28666 2864
rect 28718 800 28746 30806
rect 28810 7750 28838 30874
rect 29086 8498 29114 55270
rect 29730 53802 29758 56306
rect 29638 53774 29758 53802
rect 29350 48340 29402 48346
rect 29350 48282 29402 48288
rect 29362 46918 29390 48282
rect 29350 46912 29402 46918
rect 29350 46854 29402 46860
rect 29534 46912 29586 46918
rect 29534 46854 29586 46860
rect 29546 37312 29574 46854
rect 29454 37284 29574 37312
rect 29454 37210 29482 37284
rect 29362 37182 29482 37210
rect 29258 37120 29310 37126
rect 29258 37062 29310 37068
rect 29270 36922 29298 37062
rect 29258 36916 29310 36922
rect 29258 36858 29310 36864
rect 29362 19378 29390 37182
rect 29258 19372 29310 19378
rect 29258 19314 29310 19320
rect 29350 19372 29402 19378
rect 29350 19314 29402 19320
rect 29270 9042 29298 19314
rect 29638 9450 29666 53774
rect 30190 48346 30218 59200
rect 30650 56438 30678 59200
rect 30638 56432 30690 56438
rect 30638 56374 30690 56380
rect 31006 56432 31058 56438
rect 31006 56374 31058 56380
rect 30454 55616 30506 55622
rect 30454 55558 30506 55564
rect 30466 51950 30494 55558
rect 30454 51944 30506 51950
rect 30454 51886 30506 51892
rect 30178 48340 30230 48346
rect 30178 48282 30230 48288
rect 31018 42226 31046 56374
rect 31202 53802 31230 59200
rect 32214 56710 32242 59200
rect 32662 56772 32714 56778
rect 32662 56714 32714 56720
rect 32202 56704 32254 56710
rect 32202 56646 32254 56652
rect 31650 56364 31702 56370
rect 31650 56306 31702 56312
rect 31662 56273 31690 56306
rect 31648 56264 31704 56273
rect 31648 56199 31704 56208
rect 32568 56128 32624 56137
rect 32568 56063 32624 56072
rect 31280 55992 31336 56001
rect 31280 55927 31336 55936
rect 31832 55992 31888 56001
rect 31832 55927 31888 55936
rect 32476 55992 32532 56001
rect 32476 55927 32532 55936
rect 31294 55418 31322 55927
rect 31846 55894 31874 55927
rect 31742 55888 31794 55894
rect 31742 55830 31794 55836
rect 31834 55888 31886 55894
rect 31834 55830 31886 55836
rect 31754 55622 31782 55830
rect 31742 55616 31794 55622
rect 31742 55558 31794 55564
rect 31282 55412 31334 55418
rect 31282 55354 31334 55360
rect 32202 55208 32254 55214
rect 32202 55150 32254 55156
rect 31202 53774 31598 53802
rect 31006 42220 31058 42226
rect 31006 42162 31058 42168
rect 31098 37120 31150 37126
rect 31098 37062 31150 37068
rect 30270 23588 30322 23594
rect 30270 23530 30322 23536
rect 29718 14884 29770 14890
rect 29718 14826 29770 14832
rect 29626 9444 29678 9450
rect 29626 9386 29678 9392
rect 29258 9036 29310 9042
rect 29258 8978 29310 8984
rect 29074 8492 29126 8498
rect 29074 8434 29126 8440
rect 28798 7744 28850 7750
rect 28798 7686 28850 7692
rect 28890 7336 28942 7342
rect 28942 7284 29022 7290
rect 28890 7278 29022 7284
rect 28902 7274 29022 7278
rect 28902 7268 29034 7274
rect 28902 7262 28982 7268
rect 28982 7210 29034 7216
rect 28982 5840 29034 5846
rect 28982 5782 29034 5788
rect 28994 3738 29022 5782
rect 29730 4146 29758 14826
rect 29718 4140 29770 4146
rect 29718 4082 29770 4088
rect 30086 4072 30138 4078
rect 30086 4014 30138 4020
rect 29258 3936 29310 3942
rect 29258 3878 29310 3884
rect 29350 3936 29402 3942
rect 29350 3878 29402 3884
rect 28982 3732 29034 3738
rect 28982 3674 29034 3680
rect 28890 2984 28942 2990
rect 28890 2926 28942 2932
rect 28902 800 28930 2926
rect 29270 800 29298 3878
rect 29362 3670 29390 3878
rect 29350 3664 29402 3670
rect 29350 3606 29402 3612
rect 29626 2984 29678 2990
rect 29626 2926 29678 2932
rect 29638 800 29666 2926
rect 29994 2304 30046 2310
rect 30098 2292 30126 4014
rect 30282 2990 30310 23530
rect 31006 4140 31058 4146
rect 31006 4082 31058 4088
rect 30638 4072 30690 4078
rect 30638 4014 30690 4020
rect 30270 2984 30322 2990
rect 30270 2926 30322 2932
rect 30098 2264 30310 2292
rect 29994 2246 30046 2252
rect 30006 800 30034 2246
rect 30282 800 30310 2264
rect 30650 800 30678 4014
rect 31018 800 31046 4082
rect 31110 2990 31138 37062
rect 31570 31958 31598 53774
rect 31650 48340 31702 48346
rect 31650 48282 31702 48288
rect 31558 31952 31610 31958
rect 31558 31894 31610 31900
rect 31558 24064 31610 24070
rect 31558 24006 31610 24012
rect 31466 14884 31518 14890
rect 31466 14826 31518 14832
rect 31190 11144 31242 11150
rect 31190 11086 31242 11092
rect 31202 3534 31230 11086
rect 31478 4146 31506 14826
rect 31466 4140 31518 4146
rect 31466 4082 31518 4088
rect 31570 4078 31598 24006
rect 31558 4072 31610 4078
rect 31558 4014 31610 4020
rect 31190 3528 31242 3534
rect 31190 3470 31242 3476
rect 31098 2984 31150 2990
rect 31098 2926 31150 2932
rect 31662 2666 31690 48282
rect 32214 14074 32242 55150
rect 32386 51944 32438 51950
rect 32386 51886 32438 51892
rect 32202 14068 32254 14074
rect 32202 14010 32254 14016
rect 32398 5658 32426 51886
rect 32490 5778 32518 55927
rect 32582 35154 32610 56063
rect 32674 48346 32702 56714
rect 32766 56438 32794 59200
rect 32754 56432 32806 56438
rect 32754 56374 32806 56380
rect 33030 52964 33082 52970
rect 33030 52906 33082 52912
rect 32662 48340 32714 48346
rect 32662 48282 32714 48288
rect 32570 35148 32622 35154
rect 32570 35090 32622 35096
rect 32938 33584 32990 33590
rect 32938 33526 32990 33532
rect 32570 25424 32622 25430
rect 32570 25366 32622 25372
rect 32478 5772 32530 5778
rect 32478 5714 32530 5720
rect 32398 5630 32518 5658
rect 32386 5160 32438 5166
rect 32386 5102 32438 5108
rect 32110 4140 32162 4146
rect 32110 4082 32162 4088
rect 31742 4072 31794 4078
rect 31742 4014 31794 4020
rect 31386 2638 31690 2666
rect 31386 800 31414 2638
rect 31754 800 31782 4014
rect 32122 800 32150 4082
rect 32398 2854 32426 5102
rect 32490 3602 32518 5630
rect 32582 4282 32610 25366
rect 32662 19372 32714 19378
rect 32662 19314 32714 19320
rect 32570 4276 32622 4282
rect 32570 4218 32622 4224
rect 32478 3596 32530 3602
rect 32478 3538 32530 3544
rect 32478 3120 32530 3126
rect 32478 3062 32530 3068
rect 32386 2848 32438 2854
rect 32386 2790 32438 2796
rect 32490 800 32518 3062
rect 32674 2854 32702 19314
rect 32846 9988 32898 9994
rect 32846 9930 32898 9936
rect 32754 9920 32806 9926
rect 32754 9862 32806 9868
rect 32766 3738 32794 9862
rect 32858 4826 32886 9930
rect 32846 4820 32898 4826
rect 32846 4762 32898 4768
rect 32950 4146 32978 33526
rect 32938 4140 32990 4146
rect 32938 4082 32990 4088
rect 33042 4078 33070 52906
rect 33318 11014 33346 59200
rect 33870 56506 33898 59200
rect 33858 56500 33910 56506
rect 33858 56442 33910 56448
rect 33766 56432 33818 56438
rect 33766 56374 33818 56380
rect 33778 11558 33806 56374
rect 33856 56264 33912 56273
rect 33856 56199 33912 56208
rect 33870 15910 33898 56199
rect 34330 55690 34358 59200
rect 34882 57882 34910 59200
rect 34790 57854 34910 57882
rect 34318 55684 34370 55690
rect 34318 55626 34370 55632
rect 34790 45626 34818 57854
rect 34922 57692 35218 57712
rect 34978 57690 35002 57692
rect 35058 57690 35082 57692
rect 35138 57690 35162 57692
rect 35000 57638 35002 57690
rect 35064 57638 35076 57690
rect 35138 57638 35140 57690
rect 34978 57636 35002 57638
rect 35058 57636 35082 57638
rect 35138 57636 35162 57638
rect 34922 57616 35218 57636
rect 34922 56604 35218 56624
rect 34978 56602 35002 56604
rect 35058 56602 35082 56604
rect 35138 56602 35162 56604
rect 35000 56550 35002 56602
rect 35064 56550 35076 56602
rect 35138 56550 35140 56602
rect 34978 56548 35002 56550
rect 35058 56548 35082 56550
rect 35138 56548 35162 56550
rect 34922 56528 35218 56548
rect 35238 56432 35290 56438
rect 35238 56374 35290 56380
rect 34922 55516 35218 55536
rect 34978 55514 35002 55516
rect 35058 55514 35082 55516
rect 35138 55514 35162 55516
rect 35000 55462 35002 55514
rect 35064 55462 35076 55514
rect 35138 55462 35140 55514
rect 34978 55460 35002 55462
rect 35058 55460 35082 55462
rect 35138 55460 35162 55462
rect 34922 55440 35218 55460
rect 35250 55418 35278 56374
rect 35434 55894 35462 59200
rect 35894 56302 35922 59200
rect 35882 56296 35934 56302
rect 35974 56296 36026 56302
rect 35882 56238 35934 56244
rect 35972 56264 35974 56273
rect 36026 56264 36028 56273
rect 35972 56199 36028 56208
rect 35422 55888 35474 55894
rect 35422 55830 35474 55836
rect 36158 55888 36210 55894
rect 36158 55830 36210 55836
rect 35330 55684 35382 55690
rect 35330 55626 35382 55632
rect 35238 55412 35290 55418
rect 35238 55354 35290 55360
rect 34922 54428 35218 54448
rect 34978 54426 35002 54428
rect 35058 54426 35082 54428
rect 35138 54426 35162 54428
rect 35000 54374 35002 54426
rect 35064 54374 35076 54426
rect 35138 54374 35140 54426
rect 34978 54372 35002 54374
rect 35058 54372 35082 54374
rect 35138 54372 35162 54374
rect 34922 54352 35218 54372
rect 34922 53340 35218 53360
rect 34978 53338 35002 53340
rect 35058 53338 35082 53340
rect 35138 53338 35162 53340
rect 35000 53286 35002 53338
rect 35064 53286 35076 53338
rect 35138 53286 35140 53338
rect 34978 53284 35002 53286
rect 35058 53284 35082 53286
rect 35138 53284 35162 53286
rect 34922 53264 35218 53284
rect 34922 52252 35218 52272
rect 34978 52250 35002 52252
rect 35058 52250 35082 52252
rect 35138 52250 35162 52252
rect 35000 52198 35002 52250
rect 35064 52198 35076 52250
rect 35138 52198 35140 52250
rect 34978 52196 35002 52198
rect 35058 52196 35082 52198
rect 35138 52196 35162 52198
rect 34922 52176 35218 52196
rect 35238 51264 35290 51270
rect 35238 51206 35290 51212
rect 34922 51164 35218 51184
rect 34978 51162 35002 51164
rect 35058 51162 35082 51164
rect 35138 51162 35162 51164
rect 35000 51110 35002 51162
rect 35064 51110 35076 51162
rect 35138 51110 35140 51162
rect 34978 51108 35002 51110
rect 35058 51108 35082 51110
rect 35138 51108 35162 51110
rect 34922 51088 35218 51108
rect 34922 50076 35218 50096
rect 34978 50074 35002 50076
rect 35058 50074 35082 50076
rect 35138 50074 35162 50076
rect 35000 50022 35002 50074
rect 35064 50022 35076 50074
rect 35138 50022 35140 50074
rect 34978 50020 35002 50022
rect 35058 50020 35082 50022
rect 35138 50020 35162 50022
rect 34922 50000 35218 50020
rect 34922 48988 35218 49008
rect 34978 48986 35002 48988
rect 35058 48986 35082 48988
rect 35138 48986 35162 48988
rect 35000 48934 35002 48986
rect 35064 48934 35076 48986
rect 35138 48934 35140 48986
rect 34978 48932 35002 48934
rect 35058 48932 35082 48934
rect 35138 48932 35162 48934
rect 34922 48912 35218 48932
rect 34922 47900 35218 47920
rect 34978 47898 35002 47900
rect 35058 47898 35082 47900
rect 35138 47898 35162 47900
rect 35000 47846 35002 47898
rect 35064 47846 35076 47898
rect 35138 47846 35140 47898
rect 34978 47844 35002 47846
rect 35058 47844 35082 47846
rect 35138 47844 35162 47846
rect 34922 47824 35218 47844
rect 34922 46812 35218 46832
rect 34978 46810 35002 46812
rect 35058 46810 35082 46812
rect 35138 46810 35162 46812
rect 35000 46758 35002 46810
rect 35064 46758 35076 46810
rect 35138 46758 35140 46810
rect 34978 46756 35002 46758
rect 35058 46756 35082 46758
rect 35138 46756 35162 46758
rect 34922 46736 35218 46756
rect 34922 45724 35218 45744
rect 34978 45722 35002 45724
rect 35058 45722 35082 45724
rect 35138 45722 35162 45724
rect 35000 45670 35002 45722
rect 35064 45670 35076 45722
rect 35138 45670 35140 45722
rect 34978 45668 35002 45670
rect 35058 45668 35082 45670
rect 35138 45668 35162 45670
rect 34922 45648 35218 45668
rect 34318 45620 34370 45626
rect 34318 45562 34370 45568
rect 34778 45620 34830 45626
rect 34778 45562 34830 45568
rect 34330 36145 34358 45562
rect 34922 44636 35218 44656
rect 34978 44634 35002 44636
rect 35058 44634 35082 44636
rect 35138 44634 35162 44636
rect 35000 44582 35002 44634
rect 35064 44582 35076 44634
rect 35138 44582 35140 44634
rect 34978 44580 35002 44582
rect 35058 44580 35082 44582
rect 35138 44580 35162 44582
rect 34922 44560 35218 44580
rect 34922 43548 35218 43568
rect 34978 43546 35002 43548
rect 35058 43546 35082 43548
rect 35138 43546 35162 43548
rect 35000 43494 35002 43546
rect 35064 43494 35076 43546
rect 35138 43494 35140 43546
rect 34978 43492 35002 43494
rect 35058 43492 35082 43494
rect 35138 43492 35162 43494
rect 34922 43472 35218 43492
rect 34922 42460 35218 42480
rect 34978 42458 35002 42460
rect 35058 42458 35082 42460
rect 35138 42458 35162 42460
rect 35000 42406 35002 42458
rect 35064 42406 35076 42458
rect 35138 42406 35140 42458
rect 34978 42404 35002 42406
rect 35058 42404 35082 42406
rect 35138 42404 35162 42406
rect 34922 42384 35218 42404
rect 34922 41372 35218 41392
rect 34978 41370 35002 41372
rect 35058 41370 35082 41372
rect 35138 41370 35162 41372
rect 35000 41318 35002 41370
rect 35064 41318 35076 41370
rect 35138 41318 35140 41370
rect 34978 41316 35002 41318
rect 35058 41316 35082 41318
rect 35138 41316 35162 41318
rect 34922 41296 35218 41316
rect 34922 40284 35218 40304
rect 34978 40282 35002 40284
rect 35058 40282 35082 40284
rect 35138 40282 35162 40284
rect 35000 40230 35002 40282
rect 35064 40230 35076 40282
rect 35138 40230 35140 40282
rect 34978 40228 35002 40230
rect 35058 40228 35082 40230
rect 35138 40228 35162 40230
rect 34922 40208 35218 40228
rect 34922 39196 35218 39216
rect 34978 39194 35002 39196
rect 35058 39194 35082 39196
rect 35138 39194 35162 39196
rect 35000 39142 35002 39194
rect 35064 39142 35076 39194
rect 35138 39142 35140 39194
rect 34978 39140 35002 39142
rect 35058 39140 35082 39142
rect 35138 39140 35162 39142
rect 34922 39120 35218 39140
rect 34922 38108 35218 38128
rect 34978 38106 35002 38108
rect 35058 38106 35082 38108
rect 35138 38106 35162 38108
rect 35000 38054 35002 38106
rect 35064 38054 35076 38106
rect 35138 38054 35140 38106
rect 34978 38052 35002 38054
rect 35058 38052 35082 38054
rect 35138 38052 35162 38054
rect 34922 38032 35218 38052
rect 34922 37020 35218 37040
rect 34978 37018 35002 37020
rect 35058 37018 35082 37020
rect 35138 37018 35162 37020
rect 35000 36966 35002 37018
rect 35064 36966 35076 37018
rect 35138 36966 35140 37018
rect 34978 36964 35002 36966
rect 35058 36964 35082 36966
rect 35138 36964 35162 36966
rect 34922 36944 35218 36964
rect 34316 36136 34372 36145
rect 34316 36071 34372 36080
rect 34500 36000 34556 36009
rect 34500 35935 34556 35944
rect 34318 29164 34370 29170
rect 34318 29106 34370 29112
rect 34226 24132 34278 24138
rect 34226 24074 34278 24080
rect 34238 23866 34266 24074
rect 34226 23860 34278 23866
rect 34226 23802 34278 23808
rect 33858 15904 33910 15910
rect 33858 15846 33910 15852
rect 33766 11552 33818 11558
rect 33766 11494 33818 11500
rect 33306 11008 33358 11014
rect 33306 10950 33358 10956
rect 33122 4820 33174 4826
rect 33122 4762 33174 4768
rect 33030 4072 33082 4078
rect 33030 4014 33082 4020
rect 32846 3936 32898 3942
rect 32846 3878 32898 3884
rect 32754 3732 32806 3738
rect 32754 3674 32806 3680
rect 32662 2848 32714 2854
rect 32662 2790 32714 2796
rect 32858 800 32886 3878
rect 33134 2666 33162 4762
rect 33582 4140 33634 4146
rect 33582 4082 33634 4088
rect 33134 2638 33254 2666
rect 33226 800 33254 2638
rect 33594 800 33622 4082
rect 33950 3732 34002 3738
rect 33950 3674 34002 3680
rect 33962 800 33990 3674
rect 34330 800 34358 29106
rect 34410 29028 34462 29034
rect 34410 28970 34462 28976
rect 34422 4146 34450 28970
rect 34514 27674 34542 35935
rect 34922 35932 35218 35952
rect 34978 35930 35002 35932
rect 35058 35930 35082 35932
rect 35138 35930 35162 35932
rect 35000 35878 35002 35930
rect 35064 35878 35076 35930
rect 35138 35878 35140 35930
rect 34978 35876 35002 35878
rect 35058 35876 35082 35878
rect 35138 35876 35162 35878
rect 34922 35856 35218 35876
rect 34922 34844 35218 34864
rect 34978 34842 35002 34844
rect 35058 34842 35082 34844
rect 35138 34842 35162 34844
rect 35000 34790 35002 34842
rect 35064 34790 35076 34842
rect 35138 34790 35140 34842
rect 34978 34788 35002 34790
rect 35058 34788 35082 34790
rect 35138 34788 35162 34790
rect 34922 34768 35218 34788
rect 34922 33756 35218 33776
rect 34978 33754 35002 33756
rect 35058 33754 35082 33756
rect 35138 33754 35162 33756
rect 35000 33702 35002 33754
rect 35064 33702 35076 33754
rect 35138 33702 35140 33754
rect 34978 33700 35002 33702
rect 35058 33700 35082 33702
rect 35138 33700 35162 33702
rect 34922 33680 35218 33700
rect 34922 32668 35218 32688
rect 34978 32666 35002 32668
rect 35058 32666 35082 32668
rect 35138 32666 35162 32668
rect 35000 32614 35002 32666
rect 35064 32614 35076 32666
rect 35138 32614 35140 32666
rect 34978 32612 35002 32614
rect 35058 32612 35082 32614
rect 35138 32612 35162 32614
rect 34922 32592 35218 32612
rect 34922 31580 35218 31600
rect 34978 31578 35002 31580
rect 35058 31578 35082 31580
rect 35138 31578 35162 31580
rect 35000 31526 35002 31578
rect 35064 31526 35076 31578
rect 35138 31526 35140 31578
rect 34978 31524 35002 31526
rect 35058 31524 35082 31526
rect 35138 31524 35162 31526
rect 34922 31504 35218 31524
rect 34922 30492 35218 30512
rect 34978 30490 35002 30492
rect 35058 30490 35082 30492
rect 35138 30490 35162 30492
rect 35000 30438 35002 30490
rect 35064 30438 35076 30490
rect 35138 30438 35140 30490
rect 34978 30436 35002 30438
rect 35058 30436 35082 30438
rect 35138 30436 35162 30438
rect 34922 30416 35218 30436
rect 34922 29404 35218 29424
rect 34978 29402 35002 29404
rect 35058 29402 35082 29404
rect 35138 29402 35162 29404
rect 35000 29350 35002 29402
rect 35064 29350 35076 29402
rect 35138 29350 35140 29402
rect 34978 29348 35002 29350
rect 35058 29348 35082 29350
rect 35138 29348 35162 29350
rect 34922 29328 35218 29348
rect 34922 28316 35218 28336
rect 34978 28314 35002 28316
rect 35058 28314 35082 28316
rect 35138 28314 35162 28316
rect 35000 28262 35002 28314
rect 35064 28262 35076 28314
rect 35138 28262 35140 28314
rect 34978 28260 35002 28262
rect 35058 28260 35082 28262
rect 35138 28260 35162 28262
rect 34922 28240 35218 28260
rect 34502 27668 34554 27674
rect 34502 27610 34554 27616
rect 34778 27668 34830 27674
rect 34778 27610 34830 27616
rect 34790 22250 34818 27610
rect 34922 27228 35218 27248
rect 34978 27226 35002 27228
rect 35058 27226 35082 27228
rect 35138 27226 35162 27228
rect 35000 27174 35002 27226
rect 35064 27174 35076 27226
rect 35138 27174 35140 27226
rect 34978 27172 35002 27174
rect 35058 27172 35082 27174
rect 35138 27172 35162 27174
rect 34922 27152 35218 27172
rect 34922 26140 35218 26160
rect 34978 26138 35002 26140
rect 35058 26138 35082 26140
rect 35138 26138 35162 26140
rect 35000 26086 35002 26138
rect 35064 26086 35076 26138
rect 35138 26086 35140 26138
rect 34978 26084 35002 26086
rect 35058 26084 35082 26086
rect 35138 26084 35162 26086
rect 34922 26064 35218 26084
rect 34922 25052 35218 25072
rect 34978 25050 35002 25052
rect 35058 25050 35082 25052
rect 35138 25050 35162 25052
rect 35000 24998 35002 25050
rect 35064 24998 35076 25050
rect 35138 24998 35140 25050
rect 34978 24996 35002 24998
rect 35058 24996 35082 24998
rect 35138 24996 35162 24998
rect 34922 24976 35218 24996
rect 34922 23964 35218 23984
rect 34978 23962 35002 23964
rect 35058 23962 35082 23964
rect 35138 23962 35162 23964
rect 35000 23910 35002 23962
rect 35064 23910 35076 23962
rect 35138 23910 35140 23962
rect 34978 23908 35002 23910
rect 35058 23908 35082 23910
rect 35138 23908 35162 23910
rect 34922 23888 35218 23908
rect 34922 22876 35218 22896
rect 34978 22874 35002 22876
rect 35058 22874 35082 22876
rect 35138 22874 35162 22876
rect 35000 22822 35002 22874
rect 35064 22822 35076 22874
rect 35138 22822 35140 22874
rect 34978 22820 35002 22822
rect 35058 22820 35082 22822
rect 35138 22820 35162 22822
rect 34922 22800 35218 22820
rect 34790 22222 34910 22250
rect 34882 21978 34910 22222
rect 34790 21950 34910 21978
rect 34790 19446 34818 21950
rect 34922 21788 35218 21808
rect 34978 21786 35002 21788
rect 35058 21786 35082 21788
rect 35138 21786 35162 21788
rect 35000 21734 35002 21786
rect 35064 21734 35076 21786
rect 35138 21734 35140 21786
rect 34978 21732 35002 21734
rect 35058 21732 35082 21734
rect 35138 21732 35162 21734
rect 34922 21712 35218 21732
rect 34922 20700 35218 20720
rect 34978 20698 35002 20700
rect 35058 20698 35082 20700
rect 35138 20698 35162 20700
rect 35000 20646 35002 20698
rect 35064 20646 35076 20698
rect 35138 20646 35140 20698
rect 34978 20644 35002 20646
rect 35058 20644 35082 20646
rect 35138 20644 35162 20646
rect 34922 20624 35218 20644
rect 34922 19612 35218 19632
rect 34978 19610 35002 19612
rect 35058 19610 35082 19612
rect 35138 19610 35162 19612
rect 35000 19558 35002 19610
rect 35064 19558 35076 19610
rect 35138 19558 35140 19610
rect 34978 19556 35002 19558
rect 35058 19556 35082 19558
rect 35138 19556 35162 19558
rect 34922 19536 35218 19556
rect 34778 19440 34830 19446
rect 34778 19382 34830 19388
rect 34594 19372 34646 19378
rect 34594 19314 34646 19320
rect 34606 10266 34634 19314
rect 34922 18524 35218 18544
rect 34978 18522 35002 18524
rect 35058 18522 35082 18524
rect 35138 18522 35162 18524
rect 35000 18470 35002 18522
rect 35064 18470 35076 18522
rect 35138 18470 35140 18522
rect 34978 18468 35002 18470
rect 35058 18468 35082 18470
rect 35138 18468 35162 18470
rect 34922 18448 35218 18468
rect 34922 17436 35218 17456
rect 34978 17434 35002 17436
rect 35058 17434 35082 17436
rect 35138 17434 35162 17436
rect 35000 17382 35002 17434
rect 35064 17382 35076 17434
rect 35138 17382 35140 17434
rect 34978 17380 35002 17382
rect 35058 17380 35082 17382
rect 35138 17380 35162 17382
rect 34922 17360 35218 17380
rect 34922 16348 35218 16368
rect 34978 16346 35002 16348
rect 35058 16346 35082 16348
rect 35138 16346 35162 16348
rect 35000 16294 35002 16346
rect 35064 16294 35076 16346
rect 35138 16294 35140 16346
rect 34978 16292 35002 16294
rect 35058 16292 35082 16294
rect 35138 16292 35162 16294
rect 34922 16272 35218 16292
rect 34922 15260 35218 15280
rect 34978 15258 35002 15260
rect 35058 15258 35082 15260
rect 35138 15258 35162 15260
rect 35000 15206 35002 15258
rect 35064 15206 35076 15258
rect 35138 15206 35140 15258
rect 34978 15204 35002 15206
rect 35058 15204 35082 15206
rect 35138 15204 35162 15206
rect 34922 15184 35218 15204
rect 34922 14172 35218 14192
rect 34978 14170 35002 14172
rect 35058 14170 35082 14172
rect 35138 14170 35162 14172
rect 35000 14118 35002 14170
rect 35064 14118 35076 14170
rect 35138 14118 35140 14170
rect 34978 14116 35002 14118
rect 35058 14116 35082 14118
rect 35138 14116 35162 14118
rect 34922 14096 35218 14116
rect 34922 13084 35218 13104
rect 34978 13082 35002 13084
rect 35058 13082 35082 13084
rect 35138 13082 35162 13084
rect 35000 13030 35002 13082
rect 35064 13030 35076 13082
rect 35138 13030 35140 13082
rect 34978 13028 35002 13030
rect 35058 13028 35082 13030
rect 35138 13028 35162 13030
rect 34922 13008 35218 13028
rect 34922 11996 35218 12016
rect 34978 11994 35002 11996
rect 35058 11994 35082 11996
rect 35138 11994 35162 11996
rect 35000 11942 35002 11994
rect 35064 11942 35076 11994
rect 35138 11942 35140 11994
rect 34978 11940 35002 11942
rect 35058 11940 35082 11942
rect 35138 11940 35162 11942
rect 34922 11920 35218 11940
rect 34922 10908 35218 10928
rect 34978 10906 35002 10908
rect 35058 10906 35082 10908
rect 35138 10906 35162 10908
rect 35000 10854 35002 10906
rect 35064 10854 35076 10906
rect 35138 10854 35140 10906
rect 34978 10852 35002 10854
rect 35058 10852 35082 10854
rect 35138 10852 35162 10854
rect 34922 10832 35218 10852
rect 34594 10260 34646 10266
rect 34594 10202 34646 10208
rect 34922 9820 35218 9840
rect 34978 9818 35002 9820
rect 35058 9818 35082 9820
rect 35138 9818 35162 9820
rect 35000 9766 35002 9818
rect 35064 9766 35076 9818
rect 35138 9766 35140 9818
rect 34978 9764 35002 9766
rect 35058 9764 35082 9766
rect 35138 9764 35162 9766
rect 34922 9744 35218 9764
rect 34922 8732 35218 8752
rect 34978 8730 35002 8732
rect 35058 8730 35082 8732
rect 35138 8730 35162 8732
rect 35000 8678 35002 8730
rect 35064 8678 35076 8730
rect 35138 8678 35140 8730
rect 34978 8676 35002 8678
rect 35058 8676 35082 8678
rect 35138 8676 35162 8678
rect 34922 8656 35218 8676
rect 34922 7644 35218 7664
rect 34978 7642 35002 7644
rect 35058 7642 35082 7644
rect 35138 7642 35162 7644
rect 35000 7590 35002 7642
rect 35064 7590 35076 7642
rect 35138 7590 35140 7642
rect 34978 7588 35002 7590
rect 35058 7588 35082 7590
rect 35138 7588 35162 7590
rect 34922 7568 35218 7588
rect 34922 6556 35218 6576
rect 34978 6554 35002 6556
rect 35058 6554 35082 6556
rect 35138 6554 35162 6556
rect 35000 6502 35002 6554
rect 35064 6502 35076 6554
rect 35138 6502 35140 6554
rect 34978 6500 35002 6502
rect 35058 6500 35082 6502
rect 35138 6500 35162 6502
rect 34922 6480 35218 6500
rect 34922 5468 35218 5488
rect 34978 5466 35002 5468
rect 35058 5466 35082 5468
rect 35138 5466 35162 5468
rect 35000 5414 35002 5466
rect 35064 5414 35076 5466
rect 35138 5414 35140 5466
rect 34978 5412 35002 5414
rect 35058 5412 35082 5414
rect 35138 5412 35162 5414
rect 34922 5392 35218 5412
rect 34922 4380 35218 4400
rect 34978 4378 35002 4380
rect 35058 4378 35082 4380
rect 35138 4378 35162 4380
rect 35000 4326 35002 4378
rect 35064 4326 35076 4378
rect 35138 4326 35140 4378
rect 34978 4324 35002 4326
rect 35058 4324 35082 4326
rect 35138 4324 35162 4326
rect 34922 4304 35218 4324
rect 34410 4140 34462 4146
rect 34410 4082 34462 4088
rect 34686 3732 34738 3738
rect 34686 3674 34738 3680
rect 34698 800 34726 3674
rect 34922 3292 35218 3312
rect 34978 3290 35002 3292
rect 35058 3290 35082 3292
rect 35138 3290 35162 3292
rect 35000 3238 35002 3290
rect 35064 3238 35076 3290
rect 35138 3238 35140 3290
rect 34978 3236 35002 3238
rect 35058 3236 35082 3238
rect 35138 3236 35162 3238
rect 34922 3216 35218 3236
rect 35250 3126 35278 51206
rect 35342 17270 35370 55626
rect 36170 55622 36198 55830
rect 36158 55616 36210 55622
rect 36158 55558 36210 55564
rect 35422 55412 35474 55418
rect 35422 55354 35474 55360
rect 35434 22098 35462 55354
rect 35790 33652 35842 33658
rect 35790 33594 35842 33600
rect 35698 25832 35750 25838
rect 35698 25774 35750 25780
rect 35422 22092 35474 22098
rect 35422 22034 35474 22040
rect 35330 17264 35382 17270
rect 35330 17206 35382 17212
rect 35330 11892 35382 11898
rect 35330 11834 35382 11840
rect 35238 3120 35290 3126
rect 35238 3062 35290 3068
rect 34922 2204 35218 2224
rect 34978 2202 35002 2204
rect 35058 2202 35082 2204
rect 35138 2202 35162 2204
rect 35000 2150 35002 2202
rect 35064 2150 35076 2202
rect 35138 2150 35140 2202
rect 34978 2148 35002 2150
rect 35058 2148 35082 2150
rect 35138 2148 35162 2150
rect 34922 2128 35218 2148
rect 35342 2122 35370 11834
rect 35422 8288 35474 8294
rect 35422 8230 35474 8236
rect 35250 2094 35370 2122
rect 35250 1986 35278 2094
rect 35066 1958 35278 1986
rect 35066 800 35094 1958
rect 35434 800 35462 8230
rect 35710 3618 35738 25774
rect 35802 3738 35830 33594
rect 36526 31272 36578 31278
rect 36526 31214 36578 31220
rect 36538 7562 36566 31214
rect 36802 28416 36854 28422
rect 36802 28358 36854 28364
rect 36814 21978 36842 28358
rect 36998 26450 37026 59200
rect 37550 55162 37578 59200
rect 38562 56828 38590 59200
rect 38470 56800 38590 56828
rect 38470 55332 38498 56800
rect 38640 56400 38696 56409
rect 38640 56335 38642 56344
rect 38694 56335 38696 56344
rect 38642 56306 38694 56312
rect 38550 55344 38602 55350
rect 38470 55304 38550 55332
rect 38550 55286 38602 55292
rect 37274 55134 37578 55162
rect 37170 44736 37222 44742
rect 37170 44678 37222 44684
rect 37078 36712 37130 36718
rect 37078 36654 37130 36660
rect 36986 26444 37038 26450
rect 36986 26386 37038 26392
rect 36722 21950 36842 21978
rect 36538 7534 36658 7562
rect 35790 3732 35842 3738
rect 35790 3674 35842 3680
rect 35882 3732 35934 3738
rect 35882 3674 35934 3680
rect 35710 3590 35830 3618
rect 35894 3602 35922 3674
rect 35802 800 35830 3590
rect 35882 3596 35934 3602
rect 35882 3538 35934 3544
rect 36526 3596 36578 3602
rect 36526 3538 36578 3544
rect 36434 3528 36486 3534
rect 36434 3470 36486 3476
rect 36158 3052 36210 3058
rect 36158 2994 36210 3000
rect 36170 800 36198 2994
rect 36446 2854 36474 3470
rect 36342 2848 36394 2854
rect 36340 2816 36342 2825
rect 36434 2848 36486 2854
rect 36394 2816 36396 2825
rect 36434 2790 36486 2796
rect 36340 2751 36396 2760
rect 36538 800 36566 3538
rect 36630 2650 36658 7534
rect 36722 4010 36750 21950
rect 37090 19310 37118 36654
rect 36894 19304 36946 19310
rect 36894 19246 36946 19252
rect 37078 19304 37130 19310
rect 37078 19246 37130 19252
rect 36906 9722 36934 19246
rect 36894 9716 36946 9722
rect 36894 9658 36946 9664
rect 37078 9716 37130 9722
rect 37078 9658 37130 9664
rect 36986 6452 37038 6458
rect 36986 6394 37038 6400
rect 36998 6322 37026 6394
rect 36986 6316 37038 6322
rect 36986 6258 37038 6264
rect 36710 4004 36762 4010
rect 36710 3946 36762 3952
rect 37090 2836 37118 9658
rect 37182 3602 37210 44678
rect 37274 10470 37302 55134
rect 38642 54732 38694 54738
rect 38642 54674 38694 54680
rect 38654 54534 38682 54674
rect 38642 54528 38694 54534
rect 38642 54470 38694 54476
rect 39114 52850 39142 59200
rect 38654 52822 39142 52850
rect 38550 51944 38602 51950
rect 38550 51886 38602 51892
rect 37906 42084 37958 42090
rect 37906 42026 37958 42032
rect 37262 10464 37314 10470
rect 37262 10406 37314 10412
rect 37630 4140 37682 4146
rect 37630 4082 37682 4088
rect 37262 4072 37314 4078
rect 37262 4014 37314 4020
rect 37170 3596 37222 3602
rect 37170 3538 37222 3544
rect 37090 2808 37210 2836
rect 36618 2644 36670 2650
rect 36618 2586 36670 2592
rect 37182 921 37210 2808
rect 36892 912 36948 921
rect 36892 847 36948 856
rect 37168 912 37224 921
rect 37168 847 37224 856
rect 36906 800 36934 847
rect 37274 800 37302 4014
rect 37642 800 37670 4082
rect 37722 3936 37774 3942
rect 37722 3878 37774 3884
rect 37734 2582 37762 3878
rect 37918 3534 37946 42026
rect 38458 40180 38510 40186
rect 38458 40122 38510 40128
rect 37998 32020 38050 32026
rect 37998 31962 38050 31968
rect 37906 3528 37958 3534
rect 37906 3470 37958 3476
rect 38010 3058 38038 31962
rect 38366 20324 38418 20330
rect 38366 20266 38418 20272
rect 38090 3120 38142 3126
rect 38090 3062 38142 3068
rect 37998 3052 38050 3058
rect 37998 2994 38050 3000
rect 38102 2922 38130 3062
rect 37998 2916 38050 2922
rect 37998 2858 38050 2864
rect 38090 2916 38142 2922
rect 38090 2858 38142 2864
rect 37722 2576 37774 2582
rect 37722 2518 37774 2524
rect 38010 800 38038 2858
rect 38378 800 38406 20266
rect 38470 4078 38498 40122
rect 38562 4146 38590 51886
rect 38654 10810 38682 52822
rect 39574 51218 39602 59200
rect 40126 56828 40154 59200
rect 40034 56800 40154 56828
rect 40034 56438 40062 56800
rect 40206 56500 40258 56506
rect 40126 56460 40206 56488
rect 40022 56432 40074 56438
rect 40022 56374 40074 56380
rect 39654 55616 39706 55622
rect 39654 55558 39706 55564
rect 39482 51190 39602 51218
rect 39286 49088 39338 49094
rect 39286 49030 39338 49036
rect 39102 48340 39154 48346
rect 39102 48282 39154 48288
rect 39114 41138 39142 48282
rect 38826 41132 38878 41138
rect 38826 41074 38878 41080
rect 39102 41132 39154 41138
rect 39102 41074 39154 41080
rect 38838 27674 38866 41074
rect 38734 27668 38786 27674
rect 38734 27610 38786 27616
rect 38826 27668 38878 27674
rect 38826 27610 38878 27616
rect 38746 11694 38774 27610
rect 38734 11688 38786 11694
rect 38734 11630 38786 11636
rect 38642 10804 38694 10810
rect 38642 10746 38694 10752
rect 38826 6656 38878 6662
rect 38826 6598 38878 6604
rect 38642 6452 38694 6458
rect 38642 6394 38694 6400
rect 38654 6322 38682 6394
rect 38838 6390 38866 6598
rect 38826 6384 38878 6390
rect 38826 6326 38878 6332
rect 38642 6316 38694 6322
rect 38642 6258 38694 6264
rect 38734 6316 38786 6322
rect 38734 6258 38786 6264
rect 38550 4140 38602 4146
rect 38550 4082 38602 4088
rect 38458 4072 38510 4078
rect 38458 4014 38510 4020
rect 38746 800 38774 6258
rect 39298 3942 39326 49030
rect 39482 48346 39510 51190
rect 39666 51082 39694 55558
rect 39574 51054 39694 51082
rect 39470 48340 39522 48346
rect 39470 48282 39522 48288
rect 39378 44464 39430 44470
rect 39378 44406 39430 44412
rect 39286 3936 39338 3942
rect 39286 3878 39338 3884
rect 39102 3664 39154 3670
rect 39102 3606 39154 3612
rect 39114 800 39142 3606
rect 39390 3126 39418 44406
rect 39574 20058 39602 51054
rect 39838 45416 39890 45422
rect 39838 45358 39890 45364
rect 39850 38865 39878 45358
rect 40126 43450 40154 56460
rect 40206 56442 40258 56448
rect 40678 55894 40706 59200
rect 41690 56506 41718 59200
rect 41678 56500 41730 56506
rect 41678 56442 41730 56448
rect 40758 56432 40810 56438
rect 40758 56374 40810 56380
rect 40850 56432 40902 56438
rect 40850 56374 40902 56380
rect 40770 55894 40798 56374
rect 40862 56302 40890 56374
rect 40850 56296 40902 56302
rect 40850 56238 40902 56244
rect 40942 56296 40994 56302
rect 40942 56238 40994 56244
rect 40954 56137 40982 56238
rect 41310 56160 41362 56166
rect 40940 56128 40996 56137
rect 40940 56063 40996 56072
rect 41216 56128 41272 56137
rect 41402 56160 41454 56166
rect 41310 56102 41362 56108
rect 41400 56128 41402 56137
rect 41454 56128 41456 56137
rect 41216 56063 41272 56072
rect 41230 55962 41258 56063
rect 41322 55962 41350 56102
rect 41400 56063 41456 56072
rect 41492 55992 41548 56001
rect 41218 55956 41270 55962
rect 41218 55898 41270 55904
rect 41310 55956 41362 55962
rect 41492 55927 41548 55936
rect 41310 55898 41362 55904
rect 40666 55888 40718 55894
rect 40666 55830 40718 55836
rect 40758 55888 40810 55894
rect 40758 55830 40810 55836
rect 41506 55758 41534 55927
rect 42242 55894 42270 59200
rect 42230 55888 42282 55894
rect 42230 55830 42282 55836
rect 42322 55888 42374 55894
rect 42322 55830 42374 55836
rect 41402 55752 41454 55758
rect 41400 55720 41402 55729
rect 41494 55752 41546 55758
rect 41454 55720 41456 55729
rect 42334 55706 42362 55830
rect 41494 55694 41546 55700
rect 41400 55655 41456 55664
rect 42058 55678 42362 55706
rect 42058 55622 42086 55678
rect 42046 55616 42098 55622
rect 42046 55558 42098 55564
rect 42138 55616 42190 55622
rect 42138 55558 42190 55564
rect 40758 55412 40810 55418
rect 40758 55354 40810 55360
rect 41678 55412 41730 55418
rect 41678 55354 41730 55360
rect 40666 55344 40718 55350
rect 40666 55286 40718 55292
rect 40770 55298 40798 55354
rect 41034 55344 41086 55350
rect 40770 55292 41034 55298
rect 40770 55286 41086 55292
rect 40114 43444 40166 43450
rect 40114 43386 40166 43392
rect 39836 38856 39892 38865
rect 39836 38791 39892 38800
rect 39652 38720 39708 38729
rect 39652 38655 39708 38664
rect 39666 32450 39694 38655
rect 39666 32422 39786 32450
rect 39758 26246 39786 32422
rect 39838 32428 39890 32434
rect 39838 32370 39890 32376
rect 39746 26240 39798 26246
rect 39746 26182 39798 26188
rect 39562 20052 39614 20058
rect 39562 19994 39614 20000
rect 39654 16652 39706 16658
rect 39654 16594 39706 16600
rect 39666 7002 39694 16594
rect 39746 8832 39798 8838
rect 39746 8774 39798 8780
rect 39758 8634 39786 8774
rect 39746 8628 39798 8634
rect 39746 8570 39798 8576
rect 39654 6996 39706 7002
rect 39654 6938 39706 6944
rect 39562 6928 39614 6934
rect 39562 6870 39614 6876
rect 39574 3670 39602 6870
rect 39562 3664 39614 3670
rect 39562 3606 39614 3612
rect 39378 3120 39430 3126
rect 39378 3062 39430 3068
rect 39378 2576 39430 2582
rect 39378 2518 39430 2524
rect 39390 898 39418 2518
rect 39390 870 39510 898
rect 39482 800 39510 870
rect 39850 800 39878 32370
rect 39930 26240 39982 26246
rect 39930 26182 39982 26188
rect 39942 16658 39970 26182
rect 39930 16652 39982 16658
rect 39930 16594 39982 16600
rect 40114 6248 40166 6254
rect 40114 6190 40166 6196
rect 40022 5908 40074 5914
rect 40022 5850 40074 5856
rect 40034 3670 40062 5850
rect 40022 3664 40074 3670
rect 40022 3606 40074 3612
rect 40126 3466 40154 6190
rect 40206 3732 40258 3738
rect 40206 3674 40258 3680
rect 40218 3466 40246 3674
rect 40678 3602 40706 55286
rect 40770 55270 41074 55286
rect 41690 55214 41718 55354
rect 41678 55208 41730 55214
rect 41678 55150 41730 55156
rect 42046 50176 42098 50182
rect 42046 50118 42098 50124
rect 40758 43172 40810 43178
rect 40758 43114 40810 43120
rect 40770 4146 40798 43114
rect 40850 31816 40902 31822
rect 40850 31758 40902 31764
rect 40758 4140 40810 4146
rect 40758 4082 40810 4088
rect 40574 3596 40626 3602
rect 40574 3538 40626 3544
rect 40666 3596 40718 3602
rect 40666 3538 40718 3544
rect 40114 3460 40166 3466
rect 40114 3402 40166 3408
rect 40206 3460 40258 3466
rect 40206 3402 40258 3408
rect 40206 2984 40258 2990
rect 40206 2926 40258 2932
rect 40218 800 40246 2926
rect 40586 800 40614 3538
rect 40862 2990 40890 31758
rect 41494 22568 41546 22574
rect 41494 22510 41546 22516
rect 41126 9512 41178 9518
rect 41126 9454 41178 9460
rect 40942 4072 40994 4078
rect 40942 4014 40994 4020
rect 40850 2984 40902 2990
rect 40850 2926 40902 2932
rect 40954 800 40982 4014
rect 41138 3738 41166 9454
rect 41310 4208 41362 4214
rect 41506 4196 41534 22510
rect 41586 7744 41638 7750
rect 41586 7686 41638 7692
rect 41598 7546 41626 7686
rect 42058 7562 42086 50118
rect 42150 42362 42178 55558
rect 42794 55162 42822 59200
rect 43254 55282 43282 59200
rect 43806 55622 43834 59200
rect 44714 56500 44766 56506
rect 44714 56442 44766 56448
rect 44726 55962 44754 56442
rect 44714 55956 44766 55962
rect 44714 55898 44766 55904
rect 43884 55720 43940 55729
rect 43884 55655 43940 55664
rect 43898 55622 43926 55655
rect 43794 55616 43846 55622
rect 43794 55558 43846 55564
rect 43886 55616 43938 55622
rect 43886 55558 43938 55564
rect 43242 55276 43294 55282
rect 43242 55218 43294 55224
rect 44070 55276 44122 55282
rect 44070 55218 44122 55224
rect 42794 55134 43006 55162
rect 42414 54528 42466 54534
rect 42414 54470 42466 54476
rect 42426 54262 42454 54470
rect 42414 54256 42466 54262
rect 42414 54198 42466 54204
rect 42138 42356 42190 42362
rect 42138 42298 42190 42304
rect 42138 39296 42190 39302
rect 42138 39238 42190 39244
rect 42150 7698 42178 39238
rect 42782 37188 42834 37194
rect 42782 37130 42834 37136
rect 42794 31090 42822 37130
rect 42610 31062 42822 31090
rect 42610 26353 42638 31062
rect 42596 26344 42652 26353
rect 42596 26279 42652 26288
rect 42872 26344 42928 26353
rect 42872 26279 42928 26288
rect 42886 16674 42914 26279
rect 42702 16646 42914 16674
rect 42150 7670 42270 7698
rect 41586 7540 41638 7546
rect 42058 7534 42178 7562
rect 41586 7482 41638 7488
rect 41586 4208 41638 4214
rect 41506 4168 41586 4196
rect 41310 4150 41362 4156
rect 41586 4150 41638 4156
rect 41322 4010 41350 4150
rect 41310 4004 41362 4010
rect 41310 3946 41362 3952
rect 41126 3732 41178 3738
rect 41126 3674 41178 3680
rect 41310 3528 41362 3534
rect 41310 3470 41362 3476
rect 41402 3528 41454 3534
rect 41402 3470 41454 3476
rect 41322 2961 41350 3470
rect 41414 2990 41442 3470
rect 41678 3460 41730 3466
rect 41678 3402 41730 3408
rect 41402 2984 41454 2990
rect 41308 2952 41364 2961
rect 41494 2984 41546 2990
rect 41402 2926 41454 2932
rect 41492 2952 41494 2961
rect 41546 2952 41548 2961
rect 41308 2887 41364 2896
rect 41492 2887 41548 2896
rect 41308 2816 41364 2825
rect 41308 2751 41364 2760
rect 41322 800 41350 2751
rect 41690 800 41718 3402
rect 42150 2922 42178 7534
rect 42242 4214 42270 7670
rect 42702 6882 42730 16646
rect 42978 12850 43006 55134
rect 43426 54188 43478 54194
rect 43426 54130 43478 54136
rect 43150 41064 43202 41070
rect 43150 41006 43202 41012
rect 43162 37194 43190 41006
rect 43150 37188 43202 37194
rect 43150 37130 43202 37136
rect 42966 12844 43018 12850
rect 42966 12786 43018 12792
rect 42426 6854 42730 6882
rect 42230 4208 42282 4214
rect 42230 4150 42282 4156
rect 42046 2916 42098 2922
rect 42046 2858 42098 2864
rect 42138 2916 42190 2922
rect 42138 2858 42190 2864
rect 42058 800 42086 2858
rect 42426 800 42454 6854
rect 43150 4140 43202 4146
rect 43150 4082 43202 4088
rect 42782 3664 42834 3670
rect 42782 3606 42834 3612
rect 42794 3398 42822 3606
rect 42782 3392 42834 3398
rect 42782 3334 42834 3340
rect 42782 2848 42834 2854
rect 42782 2790 42834 2796
rect 42794 800 42822 2790
rect 43162 800 43190 4082
rect 43438 3670 43466 54130
rect 44082 47462 44110 55218
rect 44910 55214 44938 59200
rect 45370 56166 45398 59200
rect 45542 56432 45594 56438
rect 45542 56374 45594 56380
rect 45554 56234 45582 56374
rect 45542 56228 45594 56234
rect 45542 56170 45594 56176
rect 45358 56160 45410 56166
rect 45358 56102 45410 56108
rect 44898 55208 44950 55214
rect 45922 55162 45950 59200
rect 46474 57202 46502 59200
rect 46106 57174 46502 57202
rect 46002 56296 46054 56302
rect 46002 56238 46054 56244
rect 46014 55962 46042 56238
rect 46002 55956 46054 55962
rect 46002 55898 46054 55904
rect 46106 55894 46134 57174
rect 46186 56432 46238 56438
rect 46184 56400 46186 56409
rect 46238 56400 46240 56409
rect 46184 56335 46240 56344
rect 46094 55888 46146 55894
rect 46094 55830 46146 55836
rect 46186 55888 46238 55894
rect 47026 55865 47054 59200
rect 48038 56506 48066 59200
rect 48026 56500 48078 56506
rect 48026 56442 48078 56448
rect 48302 56500 48354 56506
rect 48302 56442 48354 56448
rect 46186 55830 46238 55836
rect 47012 55856 47068 55865
rect 44898 55150 44950 55156
rect 45738 55134 45950 55162
rect 44070 47456 44122 47462
rect 44070 47398 44122 47404
rect 45738 43466 45766 55134
rect 45646 43438 45766 43466
rect 43518 41472 43570 41478
rect 43518 41414 43570 41420
rect 43530 9602 43558 41414
rect 43610 33856 43662 33862
rect 43610 33798 43662 33804
rect 43622 33658 43650 33798
rect 43610 33652 43662 33658
rect 43610 33594 43662 33600
rect 45646 32450 45674 43438
rect 45646 32422 45766 32450
rect 43610 20868 43662 20874
rect 43610 20810 43662 20816
rect 43622 9738 43650 20810
rect 44806 15360 44858 15366
rect 44806 15302 44858 15308
rect 43622 9710 43742 9738
rect 43530 9574 43650 9602
rect 43518 9512 43570 9518
rect 43518 9454 43570 9460
rect 43530 9178 43558 9454
rect 43518 9172 43570 9178
rect 43518 9114 43570 9120
rect 43518 4072 43570 4078
rect 43518 4014 43570 4020
rect 43426 3664 43478 3670
rect 43426 3606 43478 3612
rect 43530 800 43558 4014
rect 43622 3738 43650 9574
rect 43714 4146 43742 9710
rect 43702 4140 43754 4146
rect 43702 4082 43754 4088
rect 43610 3732 43662 3738
rect 43610 3674 43662 3680
rect 44818 3058 44846 15302
rect 45738 14006 45766 32422
rect 45726 14000 45778 14006
rect 45726 13942 45778 13948
rect 46002 7268 46054 7274
rect 46002 7210 46054 7216
rect 45726 4140 45778 4146
rect 45726 4082 45778 4088
rect 45542 4004 45594 4010
rect 45542 3946 45594 3952
rect 45554 3670 45582 3946
rect 45450 3664 45502 3670
rect 45450 3606 45502 3612
rect 45542 3664 45594 3670
rect 45542 3606 45594 3612
rect 45462 3126 45490 3606
rect 45358 3120 45410 3126
rect 45358 3062 45410 3068
rect 45450 3120 45502 3126
rect 45450 3062 45502 3068
rect 44622 3052 44674 3058
rect 44622 2994 44674 3000
rect 44806 3052 44858 3058
rect 44806 2994 44858 3000
rect 43886 2916 43938 2922
rect 43886 2858 43938 2864
rect 43898 800 43926 2858
rect 44254 2644 44306 2650
rect 44254 2586 44306 2592
rect 44266 800 44294 2586
rect 44634 800 44662 2994
rect 44990 2984 45042 2990
rect 44990 2926 45042 2932
rect 45002 800 45030 2926
rect 45370 800 45398 3062
rect 45738 800 45766 4082
rect 45910 4072 45962 4078
rect 45910 4014 45962 4020
rect 45922 3777 45950 4014
rect 46014 4010 46042 7210
rect 46198 5234 46226 55830
rect 47012 55791 47068 55800
rect 48314 55622 48342 56442
rect 48590 56166 48618 59200
rect 48578 56160 48630 56166
rect 48578 56102 48630 56108
rect 48302 55616 48354 55622
rect 48302 55558 48354 55564
rect 47566 54120 47618 54126
rect 47566 54062 47618 54068
rect 46830 46504 46882 46510
rect 46830 46446 46882 46452
rect 46278 36916 46330 36922
rect 46278 36858 46330 36864
rect 46186 5228 46238 5234
rect 46186 5170 46238 5176
rect 46094 4072 46146 4078
rect 46094 4014 46146 4020
rect 46002 4004 46054 4010
rect 46002 3946 46054 3952
rect 45908 3768 45964 3777
rect 45908 3703 45964 3712
rect 46106 800 46134 4014
rect 46290 2650 46318 36858
rect 46738 26920 46790 26926
rect 46738 26862 46790 26868
rect 46750 4146 46778 26862
rect 46738 4140 46790 4146
rect 46738 4082 46790 4088
rect 46842 4078 46870 46446
rect 47198 12096 47250 12102
rect 47198 12038 47250 12044
rect 47210 11898 47238 12038
rect 47198 11892 47250 11898
rect 47198 11834 47250 11840
rect 47474 9512 47526 9518
rect 47474 9454 47526 9460
rect 47486 9110 47514 9454
rect 47474 9104 47526 9110
rect 47474 9046 47526 9052
rect 46922 6792 46974 6798
rect 46922 6734 46974 6740
rect 46934 6662 46962 6734
rect 46922 6656 46974 6662
rect 46922 6598 46974 6604
rect 47474 4208 47526 4214
rect 47474 4150 47526 4156
rect 46830 4072 46882 4078
rect 46830 4014 46882 4020
rect 46462 3936 46514 3942
rect 46462 3878 46514 3884
rect 46278 2644 46330 2650
rect 46278 2586 46330 2592
rect 46474 800 46502 3878
rect 46920 3768 46976 3777
rect 46920 3703 46976 3712
rect 46934 3670 46962 3703
rect 46830 3664 46882 3670
rect 46830 3606 46882 3612
rect 46922 3664 46974 3670
rect 46922 3606 46974 3612
rect 46842 800 46870 3606
rect 47198 3528 47250 3534
rect 47198 3470 47250 3476
rect 47210 800 47238 3470
rect 47486 898 47514 4150
rect 47578 4078 47606 54062
rect 49050 51542 49078 59200
rect 49602 56506 49630 59200
rect 49590 56500 49642 56506
rect 49590 56442 49642 56448
rect 49590 56364 49642 56370
rect 49590 56306 49642 56312
rect 49130 56228 49182 56234
rect 49130 56170 49182 56176
rect 49142 55758 49170 56170
rect 49130 55752 49182 55758
rect 49130 55694 49182 55700
rect 48394 51536 48446 51542
rect 48394 51478 48446 51484
rect 49038 51536 49090 51542
rect 49038 51478 49090 51484
rect 48406 46918 48434 51478
rect 48302 46912 48354 46918
rect 48302 46854 48354 46860
rect 48394 46912 48446 46918
rect 48394 46854 48446 46860
rect 47842 38208 47894 38214
rect 47842 38150 47894 38156
rect 47854 37262 47882 38150
rect 48314 37330 48342 46854
rect 49602 41562 49630 56306
rect 50154 51626 50182 59200
rect 50282 57148 50578 57168
rect 50338 57146 50362 57148
rect 50418 57146 50442 57148
rect 50498 57146 50522 57148
rect 50360 57094 50362 57146
rect 50424 57094 50436 57146
rect 50498 57094 50500 57146
rect 50338 57092 50362 57094
rect 50418 57092 50442 57094
rect 50498 57092 50522 57094
rect 50282 57072 50578 57092
rect 50282 56060 50578 56080
rect 50338 56058 50362 56060
rect 50418 56058 50442 56060
rect 50498 56058 50522 56060
rect 50360 56006 50362 56058
rect 50424 56006 50436 56058
rect 50498 56006 50500 56058
rect 50338 56004 50362 56006
rect 50418 56004 50442 56006
rect 50498 56004 50522 56006
rect 50282 55984 50578 56004
rect 51166 55826 51194 59200
rect 51244 56672 51300 56681
rect 51244 56607 51300 56616
rect 51154 55820 51206 55826
rect 51154 55762 51206 55768
rect 50282 54972 50578 54992
rect 50338 54970 50362 54972
rect 50418 54970 50442 54972
rect 50498 54970 50522 54972
rect 50360 54918 50362 54970
rect 50424 54918 50436 54970
rect 50498 54918 50500 54970
rect 50338 54916 50362 54918
rect 50418 54916 50442 54918
rect 50498 54916 50522 54918
rect 50282 54896 50578 54916
rect 50602 54324 50654 54330
rect 50602 54266 50654 54272
rect 50282 53884 50578 53904
rect 50338 53882 50362 53884
rect 50418 53882 50442 53884
rect 50498 53882 50522 53884
rect 50360 53830 50362 53882
rect 50424 53830 50436 53882
rect 50498 53830 50500 53882
rect 50338 53828 50362 53830
rect 50418 53828 50442 53830
rect 50498 53828 50522 53830
rect 50282 53808 50578 53828
rect 50282 52796 50578 52816
rect 50338 52794 50362 52796
rect 50418 52794 50442 52796
rect 50498 52794 50522 52796
rect 50360 52742 50362 52794
rect 50424 52742 50436 52794
rect 50498 52742 50500 52794
rect 50338 52740 50362 52742
rect 50418 52740 50442 52742
rect 50498 52740 50522 52742
rect 50282 52720 50578 52740
rect 50282 51708 50578 51728
rect 50338 51706 50362 51708
rect 50418 51706 50442 51708
rect 50498 51706 50522 51708
rect 50360 51654 50362 51706
rect 50424 51654 50436 51706
rect 50498 51654 50500 51706
rect 50338 51652 50362 51654
rect 50418 51652 50442 51654
rect 50498 51652 50522 51654
rect 50282 51632 50578 51652
rect 49510 41534 49630 41562
rect 49878 51598 50182 51626
rect 49510 38729 49538 41534
rect 49496 38720 49552 38729
rect 49496 38655 49552 38664
rect 49588 38584 49644 38593
rect 49588 38519 49644 38528
rect 49498 37800 49550 37806
rect 49498 37742 49550 37748
rect 48302 37324 48354 37330
rect 48302 37266 48354 37272
rect 48394 37324 48446 37330
rect 48394 37266 48446 37272
rect 47842 37256 47894 37262
rect 47842 37198 47894 37204
rect 48026 37256 48078 37262
rect 48026 37198 48078 37204
rect 48038 27674 48066 37198
rect 47842 27668 47894 27674
rect 47842 27610 47894 27616
rect 48026 27668 48078 27674
rect 48026 27610 48078 27616
rect 47854 4214 47882 27610
rect 48406 19310 48434 37266
rect 48946 29504 48998 29510
rect 48946 29446 48998 29452
rect 48394 19304 48446 19310
rect 48394 19246 48446 19252
rect 48394 19168 48446 19174
rect 48394 19110 48446 19116
rect 48406 14958 48434 19110
rect 48394 14952 48446 14958
rect 48394 14894 48446 14900
rect 48302 8560 48354 8566
rect 48222 8508 48302 8514
rect 48222 8502 48354 8508
rect 48222 8486 48342 8502
rect 48222 8430 48250 8486
rect 48210 8424 48262 8430
rect 48210 8366 48262 8372
rect 48958 4826 48986 29446
rect 48946 4820 48998 4826
rect 48946 4762 48998 4768
rect 47842 4208 47894 4214
rect 47842 4150 47894 4156
rect 48762 4140 48814 4146
rect 48762 4082 48814 4088
rect 47566 4072 47618 4078
rect 47566 4014 47618 4020
rect 48302 3596 48354 3602
rect 48302 3538 48354 3544
rect 47934 2916 47986 2922
rect 47934 2858 47986 2864
rect 47486 870 47606 898
rect 47578 800 47606 870
rect 47946 800 47974 2858
rect 48314 800 48342 3538
rect 48774 2854 48802 4082
rect 49406 4072 49458 4078
rect 49406 4014 49458 4020
rect 49038 3732 49090 3738
rect 49038 3674 49090 3680
rect 48670 2848 48722 2854
rect 48670 2790 48722 2796
rect 48762 2848 48814 2854
rect 48762 2790 48814 2796
rect 48682 800 48710 2790
rect 49050 800 49078 3674
rect 49418 2582 49446 4014
rect 49406 2576 49458 2582
rect 49406 2518 49458 2524
rect 49510 898 49538 37742
rect 49602 19922 49630 38519
rect 49878 37330 49906 51598
rect 50282 50620 50578 50640
rect 50338 50618 50362 50620
rect 50418 50618 50442 50620
rect 50498 50618 50522 50620
rect 50360 50566 50362 50618
rect 50424 50566 50436 50618
rect 50498 50566 50500 50618
rect 50338 50564 50362 50566
rect 50418 50564 50442 50566
rect 50498 50564 50522 50566
rect 50282 50544 50578 50564
rect 50282 49532 50578 49552
rect 50338 49530 50362 49532
rect 50418 49530 50442 49532
rect 50498 49530 50522 49532
rect 50360 49478 50362 49530
rect 50424 49478 50436 49530
rect 50498 49478 50500 49530
rect 50338 49476 50362 49478
rect 50418 49476 50442 49478
rect 50498 49476 50522 49478
rect 50282 49456 50578 49476
rect 50282 48444 50578 48464
rect 50338 48442 50362 48444
rect 50418 48442 50442 48444
rect 50498 48442 50522 48444
rect 50360 48390 50362 48442
rect 50424 48390 50436 48442
rect 50498 48390 50500 48442
rect 50338 48388 50362 48390
rect 50418 48388 50442 48390
rect 50498 48388 50522 48390
rect 50282 48368 50578 48388
rect 50282 47356 50578 47376
rect 50338 47354 50362 47356
rect 50418 47354 50442 47356
rect 50498 47354 50522 47356
rect 50360 47302 50362 47354
rect 50424 47302 50436 47354
rect 50498 47302 50500 47354
rect 50338 47300 50362 47302
rect 50418 47300 50442 47302
rect 50498 47300 50522 47302
rect 50282 47280 50578 47300
rect 50282 46268 50578 46288
rect 50338 46266 50362 46268
rect 50418 46266 50442 46268
rect 50498 46266 50522 46268
rect 50360 46214 50362 46266
rect 50424 46214 50436 46266
rect 50498 46214 50500 46266
rect 50338 46212 50362 46214
rect 50418 46212 50442 46214
rect 50498 46212 50522 46214
rect 50282 46192 50578 46212
rect 50282 45180 50578 45200
rect 50338 45178 50362 45180
rect 50418 45178 50442 45180
rect 50498 45178 50522 45180
rect 50360 45126 50362 45178
rect 50424 45126 50436 45178
rect 50498 45126 50500 45178
rect 50338 45124 50362 45126
rect 50418 45124 50442 45126
rect 50498 45124 50522 45126
rect 50282 45104 50578 45124
rect 50282 44092 50578 44112
rect 50338 44090 50362 44092
rect 50418 44090 50442 44092
rect 50498 44090 50522 44092
rect 50360 44038 50362 44090
rect 50424 44038 50436 44090
rect 50498 44038 50500 44090
rect 50338 44036 50362 44038
rect 50418 44036 50442 44038
rect 50498 44036 50522 44038
rect 50282 44016 50578 44036
rect 50282 43004 50578 43024
rect 50338 43002 50362 43004
rect 50418 43002 50442 43004
rect 50498 43002 50522 43004
rect 50360 42950 50362 43002
rect 50424 42950 50436 43002
rect 50498 42950 50500 43002
rect 50338 42948 50362 42950
rect 50418 42948 50442 42950
rect 50498 42948 50522 42950
rect 50282 42928 50578 42948
rect 50282 41916 50578 41936
rect 50338 41914 50362 41916
rect 50418 41914 50442 41916
rect 50498 41914 50522 41916
rect 50360 41862 50362 41914
rect 50424 41862 50436 41914
rect 50498 41862 50500 41914
rect 50338 41860 50362 41862
rect 50418 41860 50442 41862
rect 50498 41860 50522 41862
rect 50282 41840 50578 41860
rect 50282 40828 50578 40848
rect 50338 40826 50362 40828
rect 50418 40826 50442 40828
rect 50498 40826 50522 40828
rect 50360 40774 50362 40826
rect 50424 40774 50436 40826
rect 50498 40774 50500 40826
rect 50338 40772 50362 40774
rect 50418 40772 50442 40774
rect 50498 40772 50522 40774
rect 50282 40752 50578 40772
rect 50282 39740 50578 39760
rect 50338 39738 50362 39740
rect 50418 39738 50442 39740
rect 50498 39738 50522 39740
rect 50360 39686 50362 39738
rect 50424 39686 50436 39738
rect 50498 39686 50500 39738
rect 50338 39684 50362 39686
rect 50418 39684 50442 39686
rect 50498 39684 50522 39686
rect 50282 39664 50578 39684
rect 50282 38652 50578 38672
rect 50338 38650 50362 38652
rect 50418 38650 50442 38652
rect 50498 38650 50522 38652
rect 50360 38598 50362 38650
rect 50424 38598 50436 38650
rect 50498 38598 50500 38650
rect 50338 38596 50362 38598
rect 50418 38596 50442 38598
rect 50498 38596 50522 38598
rect 50282 38576 50578 38596
rect 50282 37564 50578 37584
rect 50338 37562 50362 37564
rect 50418 37562 50442 37564
rect 50498 37562 50522 37564
rect 50360 37510 50362 37562
rect 50424 37510 50436 37562
rect 50498 37510 50500 37562
rect 50338 37508 50362 37510
rect 50418 37508 50442 37510
rect 50498 37508 50522 37510
rect 50282 37488 50578 37508
rect 49774 37324 49826 37330
rect 49774 37266 49826 37272
rect 49866 37324 49918 37330
rect 49866 37266 49918 37272
rect 49786 29050 49814 37266
rect 50282 36476 50578 36496
rect 50338 36474 50362 36476
rect 50418 36474 50442 36476
rect 50498 36474 50522 36476
rect 50360 36422 50362 36474
rect 50424 36422 50436 36474
rect 50498 36422 50500 36474
rect 50338 36420 50362 36422
rect 50418 36420 50442 36422
rect 50498 36420 50522 36422
rect 50282 36400 50578 36420
rect 50282 35388 50578 35408
rect 50338 35386 50362 35388
rect 50418 35386 50442 35388
rect 50498 35386 50522 35388
rect 50360 35334 50362 35386
rect 50424 35334 50436 35386
rect 50498 35334 50500 35386
rect 50338 35332 50362 35334
rect 50418 35332 50442 35334
rect 50498 35332 50522 35334
rect 50282 35312 50578 35332
rect 50282 34300 50578 34320
rect 50338 34298 50362 34300
rect 50418 34298 50442 34300
rect 50498 34298 50522 34300
rect 50360 34246 50362 34298
rect 50424 34246 50436 34298
rect 50498 34246 50500 34298
rect 50338 34244 50362 34246
rect 50418 34244 50442 34246
rect 50498 34244 50522 34246
rect 50282 34224 50578 34244
rect 50282 33212 50578 33232
rect 50338 33210 50362 33212
rect 50418 33210 50442 33212
rect 50498 33210 50522 33212
rect 50360 33158 50362 33210
rect 50424 33158 50436 33210
rect 50498 33158 50500 33210
rect 50338 33156 50362 33158
rect 50418 33156 50442 33158
rect 50498 33156 50522 33158
rect 50282 33136 50578 33156
rect 50142 32768 50194 32774
rect 50142 32710 50194 32716
rect 49786 29022 49906 29050
rect 49878 28914 49906 29022
rect 49694 28886 49906 28914
rect 49590 19916 49642 19922
rect 49590 19858 49642 19864
rect 49694 14498 49722 28886
rect 50050 26444 50102 26450
rect 50050 26386 50102 26392
rect 49694 14470 49814 14498
rect 49682 8832 49734 8838
rect 49682 8774 49734 8780
rect 49694 2990 49722 8774
rect 49786 7546 49814 14470
rect 49774 7540 49826 7546
rect 49774 7482 49826 7488
rect 49958 4004 50010 4010
rect 49958 3946 50010 3952
rect 49774 3936 49826 3942
rect 49774 3878 49826 3884
rect 49682 2984 49734 2990
rect 49682 2926 49734 2932
rect 49418 870 49538 898
rect 49418 800 49446 870
rect 49786 800 49814 3878
rect 49970 2038 49998 3946
rect 50062 3534 50090 26386
rect 50154 5030 50182 32710
rect 50282 32124 50578 32144
rect 50338 32122 50362 32124
rect 50418 32122 50442 32124
rect 50498 32122 50522 32124
rect 50360 32070 50362 32122
rect 50424 32070 50436 32122
rect 50498 32070 50500 32122
rect 50338 32068 50362 32070
rect 50418 32068 50442 32070
rect 50498 32068 50522 32070
rect 50282 32048 50578 32068
rect 50282 31036 50578 31056
rect 50338 31034 50362 31036
rect 50418 31034 50442 31036
rect 50498 31034 50522 31036
rect 50360 30982 50362 31034
rect 50424 30982 50436 31034
rect 50498 30982 50500 31034
rect 50338 30980 50362 30982
rect 50418 30980 50442 30982
rect 50498 30980 50522 30982
rect 50282 30960 50578 30980
rect 50282 29948 50578 29968
rect 50338 29946 50362 29948
rect 50418 29946 50442 29948
rect 50498 29946 50522 29948
rect 50360 29894 50362 29946
rect 50424 29894 50436 29946
rect 50498 29894 50500 29946
rect 50338 29892 50362 29894
rect 50418 29892 50442 29894
rect 50498 29892 50522 29894
rect 50282 29872 50578 29892
rect 50282 28860 50578 28880
rect 50338 28858 50362 28860
rect 50418 28858 50442 28860
rect 50498 28858 50522 28860
rect 50360 28806 50362 28858
rect 50424 28806 50436 28858
rect 50498 28806 50500 28858
rect 50338 28804 50362 28806
rect 50418 28804 50442 28806
rect 50498 28804 50522 28806
rect 50282 28784 50578 28804
rect 50282 27772 50578 27792
rect 50338 27770 50362 27772
rect 50418 27770 50442 27772
rect 50498 27770 50522 27772
rect 50360 27718 50362 27770
rect 50424 27718 50436 27770
rect 50498 27718 50500 27770
rect 50338 27716 50362 27718
rect 50418 27716 50442 27718
rect 50498 27716 50522 27718
rect 50282 27696 50578 27716
rect 50282 26684 50578 26704
rect 50338 26682 50362 26684
rect 50418 26682 50442 26684
rect 50498 26682 50522 26684
rect 50360 26630 50362 26682
rect 50424 26630 50436 26682
rect 50498 26630 50500 26682
rect 50338 26628 50362 26630
rect 50418 26628 50442 26630
rect 50498 26628 50522 26630
rect 50282 26608 50578 26628
rect 50282 25596 50578 25616
rect 50338 25594 50362 25596
rect 50418 25594 50442 25596
rect 50498 25594 50522 25596
rect 50360 25542 50362 25594
rect 50424 25542 50436 25594
rect 50498 25542 50500 25594
rect 50338 25540 50362 25542
rect 50418 25540 50442 25542
rect 50498 25540 50522 25542
rect 50282 25520 50578 25540
rect 50282 24508 50578 24528
rect 50338 24506 50362 24508
rect 50418 24506 50442 24508
rect 50498 24506 50522 24508
rect 50360 24454 50362 24506
rect 50424 24454 50436 24506
rect 50498 24454 50500 24506
rect 50338 24452 50362 24454
rect 50418 24452 50442 24454
rect 50498 24452 50522 24454
rect 50282 24432 50578 24452
rect 50282 23420 50578 23440
rect 50338 23418 50362 23420
rect 50418 23418 50442 23420
rect 50498 23418 50522 23420
rect 50360 23366 50362 23418
rect 50424 23366 50436 23418
rect 50498 23366 50500 23418
rect 50338 23364 50362 23366
rect 50418 23364 50442 23366
rect 50498 23364 50522 23366
rect 50282 23344 50578 23364
rect 50282 22332 50578 22352
rect 50338 22330 50362 22332
rect 50418 22330 50442 22332
rect 50498 22330 50522 22332
rect 50360 22278 50362 22330
rect 50424 22278 50436 22330
rect 50498 22278 50500 22330
rect 50338 22276 50362 22278
rect 50418 22276 50442 22278
rect 50498 22276 50522 22278
rect 50282 22256 50578 22276
rect 50282 21244 50578 21264
rect 50338 21242 50362 21244
rect 50418 21242 50442 21244
rect 50498 21242 50522 21244
rect 50360 21190 50362 21242
rect 50424 21190 50436 21242
rect 50498 21190 50500 21242
rect 50338 21188 50362 21190
rect 50418 21188 50442 21190
rect 50498 21188 50522 21190
rect 50282 21168 50578 21188
rect 50282 20156 50578 20176
rect 50338 20154 50362 20156
rect 50418 20154 50442 20156
rect 50498 20154 50522 20156
rect 50360 20102 50362 20154
rect 50424 20102 50436 20154
rect 50498 20102 50500 20154
rect 50338 20100 50362 20102
rect 50418 20100 50442 20102
rect 50498 20100 50522 20102
rect 50282 20080 50578 20100
rect 50282 19068 50578 19088
rect 50338 19066 50362 19068
rect 50418 19066 50442 19068
rect 50498 19066 50522 19068
rect 50360 19014 50362 19066
rect 50424 19014 50436 19066
rect 50498 19014 50500 19066
rect 50338 19012 50362 19014
rect 50418 19012 50442 19014
rect 50498 19012 50522 19014
rect 50282 18992 50578 19012
rect 50282 17980 50578 18000
rect 50338 17978 50362 17980
rect 50418 17978 50442 17980
rect 50498 17978 50522 17980
rect 50360 17926 50362 17978
rect 50424 17926 50436 17978
rect 50498 17926 50500 17978
rect 50338 17924 50362 17926
rect 50418 17924 50442 17926
rect 50498 17924 50522 17926
rect 50282 17904 50578 17924
rect 50282 16892 50578 16912
rect 50338 16890 50362 16892
rect 50418 16890 50442 16892
rect 50498 16890 50522 16892
rect 50360 16838 50362 16890
rect 50424 16838 50436 16890
rect 50498 16838 50500 16890
rect 50338 16836 50362 16838
rect 50418 16836 50442 16838
rect 50498 16836 50522 16838
rect 50282 16816 50578 16836
rect 50282 15804 50578 15824
rect 50338 15802 50362 15804
rect 50418 15802 50442 15804
rect 50498 15802 50522 15804
rect 50360 15750 50362 15802
rect 50424 15750 50436 15802
rect 50498 15750 50500 15802
rect 50338 15748 50362 15750
rect 50418 15748 50442 15750
rect 50498 15748 50522 15750
rect 50282 15728 50578 15748
rect 50282 14716 50578 14736
rect 50338 14714 50362 14716
rect 50418 14714 50442 14716
rect 50498 14714 50522 14716
rect 50360 14662 50362 14714
rect 50424 14662 50436 14714
rect 50498 14662 50500 14714
rect 50338 14660 50362 14662
rect 50418 14660 50442 14662
rect 50498 14660 50522 14662
rect 50282 14640 50578 14660
rect 50282 13628 50578 13648
rect 50338 13626 50362 13628
rect 50418 13626 50442 13628
rect 50498 13626 50522 13628
rect 50360 13574 50362 13626
rect 50424 13574 50436 13626
rect 50498 13574 50500 13626
rect 50338 13572 50362 13574
rect 50418 13572 50442 13574
rect 50498 13572 50522 13574
rect 50282 13552 50578 13572
rect 50282 12540 50578 12560
rect 50338 12538 50362 12540
rect 50418 12538 50442 12540
rect 50498 12538 50522 12540
rect 50360 12486 50362 12538
rect 50424 12486 50436 12538
rect 50498 12486 50500 12538
rect 50338 12484 50362 12486
rect 50418 12484 50442 12486
rect 50498 12484 50522 12486
rect 50282 12464 50578 12484
rect 50282 11452 50578 11472
rect 50338 11450 50362 11452
rect 50418 11450 50442 11452
rect 50498 11450 50522 11452
rect 50360 11398 50362 11450
rect 50424 11398 50436 11450
rect 50498 11398 50500 11450
rect 50338 11396 50362 11398
rect 50418 11396 50442 11398
rect 50498 11396 50522 11398
rect 50282 11376 50578 11396
rect 50282 10364 50578 10384
rect 50338 10362 50362 10364
rect 50418 10362 50442 10364
rect 50498 10362 50522 10364
rect 50360 10310 50362 10362
rect 50424 10310 50436 10362
rect 50498 10310 50500 10362
rect 50338 10308 50362 10310
rect 50418 10308 50442 10310
rect 50498 10308 50522 10310
rect 50282 10288 50578 10308
rect 50282 9276 50578 9296
rect 50338 9274 50362 9276
rect 50418 9274 50442 9276
rect 50498 9274 50522 9276
rect 50360 9222 50362 9274
rect 50424 9222 50436 9274
rect 50498 9222 50500 9274
rect 50338 9220 50362 9222
rect 50418 9220 50442 9222
rect 50498 9220 50522 9222
rect 50282 9200 50578 9220
rect 50282 8188 50578 8208
rect 50338 8186 50362 8188
rect 50418 8186 50442 8188
rect 50498 8186 50522 8188
rect 50360 8134 50362 8186
rect 50424 8134 50436 8186
rect 50498 8134 50500 8186
rect 50338 8132 50362 8134
rect 50418 8132 50442 8134
rect 50498 8132 50522 8134
rect 50282 8112 50578 8132
rect 50282 7100 50578 7120
rect 50338 7098 50362 7100
rect 50418 7098 50442 7100
rect 50498 7098 50522 7100
rect 50360 7046 50362 7098
rect 50424 7046 50436 7098
rect 50498 7046 50500 7098
rect 50338 7044 50362 7046
rect 50418 7044 50442 7046
rect 50498 7044 50522 7046
rect 50282 7024 50578 7044
rect 50282 6012 50578 6032
rect 50338 6010 50362 6012
rect 50418 6010 50442 6012
rect 50498 6010 50522 6012
rect 50360 5958 50362 6010
rect 50424 5958 50436 6010
rect 50498 5958 50500 6010
rect 50338 5956 50362 5958
rect 50418 5956 50442 5958
rect 50498 5956 50522 5958
rect 50282 5936 50578 5956
rect 50142 5024 50194 5030
rect 50142 4966 50194 4972
rect 50282 4924 50578 4944
rect 50338 4922 50362 4924
rect 50418 4922 50442 4924
rect 50498 4922 50522 4924
rect 50360 4870 50362 4922
rect 50424 4870 50436 4922
rect 50498 4870 50500 4922
rect 50338 4868 50362 4870
rect 50418 4868 50442 4870
rect 50498 4868 50522 4870
rect 50282 4848 50578 4868
rect 50614 4282 50642 54266
rect 51258 51082 51286 56607
rect 51718 56438 51746 59200
rect 52270 56817 52298 59200
rect 52256 56808 52312 56817
rect 52256 56743 52312 56752
rect 51706 56432 51758 56438
rect 51706 56374 51758 56380
rect 52730 56234 52758 59200
rect 53282 56370 53310 59200
rect 53270 56364 53322 56370
rect 53270 56306 53322 56312
rect 52718 56228 52770 56234
rect 52718 56170 52770 56176
rect 54386 55418 54414 59200
rect 54846 56166 54874 59200
rect 54834 56160 54886 56166
rect 54834 56102 54886 56108
rect 54374 55412 54426 55418
rect 54374 55354 54426 55360
rect 51166 51054 51286 51082
rect 51166 46866 51194 51054
rect 53086 48680 53138 48686
rect 53086 48622 53138 48628
rect 51166 46838 51286 46866
rect 50694 46436 50746 46442
rect 50694 46378 50746 46384
rect 50602 4276 50654 4282
rect 50602 4218 50654 4224
rect 50282 3836 50578 3856
rect 50338 3834 50362 3836
rect 50418 3834 50442 3836
rect 50498 3834 50522 3836
rect 50360 3782 50362 3834
rect 50424 3782 50436 3834
rect 50498 3782 50500 3834
rect 50338 3780 50362 3782
rect 50418 3780 50442 3782
rect 50498 3780 50522 3782
rect 50282 3760 50578 3780
rect 50706 3738 50734 46378
rect 50970 44736 51022 44742
rect 50970 44678 51022 44684
rect 50878 41064 50930 41070
rect 50878 41006 50930 41012
rect 50786 36644 50838 36650
rect 50786 36586 50838 36592
rect 50694 3732 50746 3738
rect 50694 3674 50746 3680
rect 50142 3596 50194 3602
rect 50142 3538 50194 3544
rect 50050 3528 50102 3534
rect 50050 3470 50102 3476
rect 49958 2032 50010 2038
rect 49958 1974 50010 1980
rect 50154 800 50182 3538
rect 50602 3392 50654 3398
rect 50602 3334 50654 3340
rect 50282 2748 50578 2768
rect 50338 2746 50362 2748
rect 50418 2746 50442 2748
rect 50498 2746 50522 2748
rect 50360 2694 50362 2746
rect 50424 2694 50436 2746
rect 50498 2694 50500 2746
rect 50338 2692 50362 2694
rect 50418 2692 50442 2694
rect 50498 2692 50522 2694
rect 50282 2672 50578 2692
rect 50614 2530 50642 3334
rect 50798 2990 50826 36586
rect 50890 3754 50918 41006
rect 50982 3942 51010 44678
rect 51258 29458 51286 46838
rect 52902 34944 52954 34950
rect 52902 34886 52954 34892
rect 52914 34746 52942 34886
rect 52902 34740 52954 34746
rect 52902 34682 52954 34688
rect 51074 29430 51286 29458
rect 51074 24206 51102 29430
rect 51706 29300 51758 29306
rect 51706 29242 51758 29248
rect 51062 24200 51114 24206
rect 51062 24142 51114 24148
rect 51062 24064 51114 24070
rect 51062 24006 51114 24012
rect 51074 16454 51102 24006
rect 51062 16448 51114 16454
rect 51062 16390 51114 16396
rect 51062 6180 51114 6186
rect 51062 6122 51114 6128
rect 51074 3942 51102 6122
rect 50970 3936 51022 3942
rect 50970 3878 51022 3884
rect 51062 3936 51114 3942
rect 51062 3878 51114 3884
rect 50890 3726 51010 3754
rect 50878 3664 50930 3670
rect 50878 3606 50930 3612
rect 50786 2984 50838 2990
rect 50786 2926 50838 2932
rect 50522 2502 50642 2530
rect 50522 800 50550 2502
rect 50890 800 50918 3606
rect 50982 3602 51010 3726
rect 51338 3732 51390 3738
rect 51338 3674 51390 3680
rect 50970 3596 51022 3602
rect 50970 3538 51022 3544
rect 51350 3126 51378 3674
rect 51718 3466 51746 29242
rect 51798 20460 51850 20466
rect 51798 20402 51850 20408
rect 51810 3602 51838 20402
rect 52074 19304 52126 19310
rect 52074 19246 52126 19252
rect 52086 17678 52114 19246
rect 52074 17672 52126 17678
rect 52074 17614 52126 17620
rect 51890 16788 51942 16794
rect 51890 16730 51942 16736
rect 51798 3596 51850 3602
rect 51798 3538 51850 3544
rect 51706 3460 51758 3466
rect 51706 3402 51758 3408
rect 51902 3194 51930 16730
rect 51982 12776 52034 12782
rect 51982 12718 52034 12724
rect 51994 3670 52022 12718
rect 52074 10600 52126 10606
rect 52074 10542 52126 10548
rect 52086 3738 52114 10542
rect 52442 6656 52494 6662
rect 52442 6598 52494 6604
rect 52454 6458 52482 6598
rect 52442 6452 52494 6458
rect 52442 6394 52494 6400
rect 52442 5160 52494 5166
rect 52442 5102 52494 5108
rect 52074 3732 52126 3738
rect 52074 3674 52126 3680
rect 51982 3664 52034 3670
rect 51982 3606 52034 3612
rect 51614 3188 51666 3194
rect 51614 3130 51666 3136
rect 51890 3188 51942 3194
rect 51890 3130 51942 3136
rect 51246 3120 51298 3126
rect 51246 3062 51298 3068
rect 51338 3120 51390 3126
rect 51338 3062 51390 3068
rect 51258 800 51286 3062
rect 51626 800 51654 3130
rect 52350 3052 52402 3058
rect 52350 2994 52402 3000
rect 51982 2848 52034 2854
rect 51982 2790 52034 2796
rect 51994 800 52022 2790
rect 52362 800 52390 2994
rect 52454 2922 52482 5102
rect 52718 4820 52770 4826
rect 52718 4762 52770 4768
rect 52534 3528 52586 3534
rect 52534 3470 52586 3476
rect 52546 2990 52574 3470
rect 52534 2984 52586 2990
rect 52534 2926 52586 2932
rect 52442 2916 52494 2922
rect 52442 2858 52494 2864
rect 52730 800 52758 4762
rect 53098 3534 53126 48622
rect 54006 32360 54058 32366
rect 54006 32302 54058 32308
rect 53178 7336 53230 7342
rect 53178 7278 53230 7284
rect 53086 3528 53138 3534
rect 53086 3470 53138 3476
rect 53190 2922 53218 7278
rect 54018 4298 54046 32302
rect 55398 17610 55426 59200
rect 55950 55894 55978 59200
rect 55938 55888 55990 55894
rect 55938 55830 55990 55836
rect 56410 55350 56438 59200
rect 56962 59106 56990 59200
rect 56778 59078 56990 59106
rect 56398 55344 56450 55350
rect 56398 55286 56450 55292
rect 56778 41426 56806 59078
rect 57514 56302 57542 59200
rect 57502 56296 57554 56302
rect 57502 56238 57554 56244
rect 58066 53650 58094 59200
rect 59078 55962 59106 59200
rect 59066 55956 59118 55962
rect 59066 55898 59118 55904
rect 59630 55690 59658 59200
rect 59618 55684 59670 55690
rect 59618 55626 59670 55632
rect 58054 53644 58106 53650
rect 58054 53586 58106 53592
rect 56950 44736 57002 44742
rect 56950 44678 57002 44684
rect 56962 44538 56990 44678
rect 56950 44532 57002 44538
rect 56950 44474 57002 44480
rect 56686 41398 56806 41426
rect 55846 26920 55898 26926
rect 55846 26862 55898 26868
rect 55386 17604 55438 17610
rect 55386 17546 55438 17552
rect 54926 9512 54978 9518
rect 54926 9454 54978 9460
rect 54018 4270 54506 4298
rect 53822 3528 53874 3534
rect 53822 3470 53874 3476
rect 53178 2916 53230 2922
rect 53178 2858 53230 2864
rect 53454 2644 53506 2650
rect 53454 2586 53506 2592
rect 53086 2032 53138 2038
rect 53086 1974 53138 1980
rect 53098 800 53126 1974
rect 53466 800 53494 2586
rect 53834 800 53862 3470
rect 54190 2576 54242 2582
rect 54190 2518 54242 2524
rect 54202 800 54230 2518
rect 54478 898 54506 4270
rect 54478 870 54598 898
rect 54570 800 54598 870
rect 54938 800 54966 9454
rect 55294 5024 55346 5030
rect 55294 4966 55346 4972
rect 55306 800 55334 4966
rect 55858 3534 55886 26862
rect 56686 19310 56714 41398
rect 58422 33856 58474 33862
rect 58422 33798 58474 33804
rect 58434 33590 58462 33798
rect 58422 33584 58474 33590
rect 58422 33526 58474 33532
rect 56674 19304 56726 19310
rect 56674 19246 56726 19252
rect 56398 4276 56450 4282
rect 56398 4218 56450 4224
rect 55846 3528 55898 3534
rect 55846 3470 55898 3476
rect 55662 3120 55714 3126
rect 55662 3062 55714 3068
rect 55674 800 55702 3062
rect 56030 3052 56082 3058
rect 56030 2994 56082 3000
rect 56042 800 56070 2994
rect 56410 800 56438 4218
rect 58974 3936 59026 3942
rect 58974 3878 59026 3884
rect 58238 3664 58290 3670
rect 58238 3606 58290 3612
rect 57870 3528 57922 3534
rect 57870 3470 57922 3476
rect 57502 3188 57554 3194
rect 57502 3130 57554 3136
rect 56766 2984 56818 2990
rect 56766 2926 56818 2932
rect 56778 800 56806 2926
rect 57134 2916 57186 2922
rect 57134 2858 57186 2864
rect 57146 800 57174 2858
rect 57514 800 57542 3130
rect 57882 800 57910 3470
rect 58250 800 58278 3606
rect 58606 3392 58658 3398
rect 58606 3334 58658 3340
rect 58618 800 58646 3334
rect 58986 800 59014 3878
rect 59342 3732 59394 3738
rect 59342 3674 59394 3680
rect 59354 800 59382 3674
rect 59710 3596 59762 3602
rect 59710 3538 59762 3544
rect 59722 800 59750 3538
rect 0 0 56 800
rect 92 0 148 800
rect 184 0 240 800
rect 276 0 332 800
rect 460 0 516 800
rect 552 0 608 800
rect 644 0 700 800
rect 828 0 884 800
rect 920 0 976 800
rect 1012 0 1068 800
rect 1196 0 1252 800
rect 1288 0 1344 800
rect 1380 0 1436 800
rect 1564 0 1620 800
rect 1656 0 1712 800
rect 1748 0 1804 800
rect 1932 0 1988 800
rect 2024 0 2080 800
rect 2116 0 2172 800
rect 2300 0 2356 800
rect 2392 0 2448 800
rect 2484 0 2540 800
rect 2668 0 2724 800
rect 2760 0 2816 800
rect 2852 0 2908 800
rect 3036 0 3092 800
rect 3128 0 3184 800
rect 3220 0 3276 800
rect 3404 0 3460 800
rect 3496 0 3552 800
rect 3588 0 3644 800
rect 3772 0 3828 800
rect 3864 0 3920 800
rect 3956 0 4012 800
rect 4140 0 4196 800
rect 4232 0 4288 800
rect 4324 0 4380 800
rect 4508 0 4564 800
rect 4600 0 4656 800
rect 4692 0 4748 800
rect 4876 0 4932 800
rect 4968 0 5024 800
rect 5060 0 5116 800
rect 5244 0 5300 800
rect 5336 0 5392 800
rect 5428 0 5484 800
rect 5612 0 5668 800
rect 5704 0 5760 800
rect 5796 0 5852 800
rect 5980 0 6036 800
rect 6072 0 6128 800
rect 6164 0 6220 800
rect 6348 0 6404 800
rect 6440 0 6496 800
rect 6532 0 6588 800
rect 6716 0 6772 800
rect 6808 0 6864 800
rect 6900 0 6956 800
rect 7084 0 7140 800
rect 7176 0 7232 800
rect 7268 0 7324 800
rect 7452 0 7508 800
rect 7544 0 7600 800
rect 7636 0 7692 800
rect 7820 0 7876 800
rect 7912 0 7968 800
rect 8004 0 8060 800
rect 8188 0 8244 800
rect 8280 0 8336 800
rect 8372 0 8428 800
rect 8556 0 8612 800
rect 8648 0 8704 800
rect 8740 0 8796 800
rect 8924 0 8980 800
rect 9016 0 9072 800
rect 9108 0 9164 800
rect 9292 0 9348 800
rect 9384 0 9440 800
rect 9476 0 9532 800
rect 9660 0 9716 800
rect 9752 0 9808 800
rect 9844 0 9900 800
rect 10028 0 10084 800
rect 10120 0 10176 800
rect 10212 0 10268 800
rect 10396 0 10452 800
rect 10488 0 10544 800
rect 10580 0 10636 800
rect 10764 0 10820 800
rect 10856 0 10912 800
rect 10948 0 11004 800
rect 11132 0 11188 800
rect 11224 0 11280 800
rect 11316 0 11372 800
rect 11500 0 11556 800
rect 11592 0 11648 800
rect 11684 0 11740 800
rect 11868 0 11924 800
rect 11960 0 12016 800
rect 12052 0 12108 800
rect 12236 0 12292 800
rect 12328 0 12384 800
rect 12420 0 12476 800
rect 12604 0 12660 800
rect 12696 0 12752 800
rect 12788 0 12844 800
rect 12972 0 13028 800
rect 13064 0 13120 800
rect 13156 0 13212 800
rect 13340 0 13396 800
rect 13432 0 13488 800
rect 13524 0 13580 800
rect 13708 0 13764 800
rect 13800 0 13856 800
rect 13892 0 13948 800
rect 14076 0 14132 800
rect 14168 0 14224 800
rect 14260 0 14316 800
rect 14444 0 14500 800
rect 14536 0 14592 800
rect 14628 0 14684 800
rect 14812 0 14868 800
rect 14904 0 14960 800
rect 14996 0 15052 800
rect 15088 0 15144 800
rect 15272 0 15328 800
rect 15364 0 15420 800
rect 15456 0 15512 800
rect 15640 0 15696 800
rect 15732 0 15788 800
rect 15824 0 15880 800
rect 16008 0 16064 800
rect 16100 0 16156 800
rect 16192 0 16248 800
rect 16376 0 16432 800
rect 16468 0 16524 800
rect 16560 0 16616 800
rect 16744 0 16800 800
rect 16836 0 16892 800
rect 16928 0 16984 800
rect 17112 0 17168 800
rect 17204 0 17260 800
rect 17296 0 17352 800
rect 17480 0 17536 800
rect 17572 0 17628 800
rect 17664 0 17720 800
rect 17848 0 17904 800
rect 17940 0 17996 800
rect 18032 0 18088 800
rect 18216 0 18272 800
rect 18308 0 18364 800
rect 18400 0 18456 800
rect 18584 0 18640 800
rect 18676 0 18732 800
rect 18768 0 18824 800
rect 18952 0 19008 800
rect 19044 0 19100 800
rect 19136 0 19192 800
rect 19320 0 19376 800
rect 19412 0 19468 800
rect 19504 0 19560 800
rect 19688 0 19744 800
rect 19780 0 19836 800
rect 19872 0 19928 800
rect 20056 0 20112 800
rect 20148 0 20204 800
rect 20240 0 20296 800
rect 20424 0 20480 800
rect 20516 0 20572 800
rect 20608 0 20664 800
rect 20792 0 20848 800
rect 20884 0 20940 800
rect 20976 0 21032 800
rect 21160 0 21216 800
rect 21252 0 21308 800
rect 21344 0 21400 800
rect 21528 0 21584 800
rect 21620 0 21676 800
rect 21712 0 21768 800
rect 21896 0 21952 800
rect 21988 0 22044 800
rect 22080 0 22136 800
rect 22264 0 22320 800
rect 22356 0 22412 800
rect 22448 0 22504 800
rect 22632 0 22688 800
rect 22724 0 22780 800
rect 22816 0 22872 800
rect 23000 0 23056 800
rect 23092 0 23148 800
rect 23184 0 23240 800
rect 23368 0 23424 800
rect 23460 0 23516 800
rect 23552 0 23608 800
rect 23736 0 23792 800
rect 23828 0 23884 800
rect 23920 0 23976 800
rect 24104 0 24160 800
rect 24196 0 24252 800
rect 24288 0 24344 800
rect 24472 0 24528 800
rect 24564 0 24620 800
rect 24656 0 24712 800
rect 24840 0 24896 800
rect 24932 0 24988 800
rect 25024 0 25080 800
rect 25208 0 25264 800
rect 25300 0 25356 800
rect 25392 0 25448 800
rect 25576 0 25632 800
rect 25668 0 25724 800
rect 25760 0 25816 800
rect 25944 0 26000 800
rect 26036 0 26092 800
rect 26128 0 26184 800
rect 26312 0 26368 800
rect 26404 0 26460 800
rect 26496 0 26552 800
rect 26680 0 26736 800
rect 26772 0 26828 800
rect 26864 0 26920 800
rect 27048 0 27104 800
rect 27140 0 27196 800
rect 27232 0 27288 800
rect 27416 0 27472 800
rect 27508 0 27564 800
rect 27600 0 27656 800
rect 27784 0 27840 800
rect 27876 0 27932 800
rect 27968 0 28024 800
rect 28152 0 28208 800
rect 28244 0 28300 800
rect 28336 0 28392 800
rect 28520 0 28576 800
rect 28612 0 28668 800
rect 28704 0 28760 800
rect 28888 0 28944 800
rect 28980 0 29036 800
rect 29072 0 29128 800
rect 29256 0 29312 800
rect 29348 0 29404 800
rect 29440 0 29496 800
rect 29624 0 29680 800
rect 29716 0 29772 800
rect 29808 0 29864 800
rect 29992 0 30048 800
rect 30084 0 30140 800
rect 30176 0 30232 800
rect 30268 0 30324 800
rect 30452 0 30508 800
rect 30544 0 30600 800
rect 30636 0 30692 800
rect 30820 0 30876 800
rect 30912 0 30968 800
rect 31004 0 31060 800
rect 31188 0 31244 800
rect 31280 0 31336 800
rect 31372 0 31428 800
rect 31556 0 31612 800
rect 31648 0 31704 800
rect 31740 0 31796 800
rect 31924 0 31980 800
rect 32016 0 32072 800
rect 32108 0 32164 800
rect 32292 0 32348 800
rect 32384 0 32440 800
rect 32476 0 32532 800
rect 32660 0 32716 800
rect 32752 0 32808 800
rect 32844 0 32900 800
rect 33028 0 33084 800
rect 33120 0 33176 800
rect 33212 0 33268 800
rect 33396 0 33452 800
rect 33488 0 33544 800
rect 33580 0 33636 800
rect 33764 0 33820 800
rect 33856 0 33912 800
rect 33948 0 34004 800
rect 34132 0 34188 800
rect 34224 0 34280 800
rect 34316 0 34372 800
rect 34500 0 34556 800
rect 34592 0 34648 800
rect 34684 0 34740 800
rect 34868 0 34924 800
rect 34960 0 35016 800
rect 35052 0 35108 800
rect 35236 0 35292 800
rect 35328 0 35384 800
rect 35420 0 35476 800
rect 35604 0 35660 800
rect 35696 0 35752 800
rect 35788 0 35844 800
rect 35972 0 36028 800
rect 36064 0 36120 800
rect 36156 0 36212 800
rect 36340 0 36396 800
rect 36432 0 36488 800
rect 36524 0 36580 800
rect 36708 0 36764 800
rect 36800 0 36856 800
rect 36892 0 36948 800
rect 37076 0 37132 800
rect 37168 0 37224 800
rect 37260 0 37316 800
rect 37444 0 37500 800
rect 37536 0 37592 800
rect 37628 0 37684 800
rect 37812 0 37868 800
rect 37904 0 37960 800
rect 37996 0 38052 800
rect 38180 0 38236 800
rect 38272 0 38328 800
rect 38364 0 38420 800
rect 38548 0 38604 800
rect 38640 0 38696 800
rect 38732 0 38788 800
rect 38916 0 38972 800
rect 39008 0 39064 800
rect 39100 0 39156 800
rect 39284 0 39340 800
rect 39376 0 39432 800
rect 39468 0 39524 800
rect 39652 0 39708 800
rect 39744 0 39800 800
rect 39836 0 39892 800
rect 40020 0 40076 800
rect 40112 0 40168 800
rect 40204 0 40260 800
rect 40388 0 40444 800
rect 40480 0 40536 800
rect 40572 0 40628 800
rect 40756 0 40812 800
rect 40848 0 40904 800
rect 40940 0 40996 800
rect 41124 0 41180 800
rect 41216 0 41272 800
rect 41308 0 41364 800
rect 41492 0 41548 800
rect 41584 0 41640 800
rect 41676 0 41732 800
rect 41860 0 41916 800
rect 41952 0 42008 800
rect 42044 0 42100 800
rect 42228 0 42284 800
rect 42320 0 42376 800
rect 42412 0 42468 800
rect 42596 0 42652 800
rect 42688 0 42744 800
rect 42780 0 42836 800
rect 42964 0 43020 800
rect 43056 0 43112 800
rect 43148 0 43204 800
rect 43332 0 43388 800
rect 43424 0 43480 800
rect 43516 0 43572 800
rect 43700 0 43756 800
rect 43792 0 43848 800
rect 43884 0 43940 800
rect 44068 0 44124 800
rect 44160 0 44216 800
rect 44252 0 44308 800
rect 44436 0 44492 800
rect 44528 0 44584 800
rect 44620 0 44676 800
rect 44804 0 44860 800
rect 44896 0 44952 800
rect 44988 0 45044 800
rect 45080 0 45136 800
rect 45264 0 45320 800
rect 45356 0 45412 800
rect 45448 0 45504 800
rect 45632 0 45688 800
rect 45724 0 45780 800
rect 45816 0 45872 800
rect 46000 0 46056 800
rect 46092 0 46148 800
rect 46184 0 46240 800
rect 46368 0 46424 800
rect 46460 0 46516 800
rect 46552 0 46608 800
rect 46736 0 46792 800
rect 46828 0 46884 800
rect 46920 0 46976 800
rect 47104 0 47160 800
rect 47196 0 47252 800
rect 47288 0 47344 800
rect 47472 0 47528 800
rect 47564 0 47620 800
rect 47656 0 47712 800
rect 47840 0 47896 800
rect 47932 0 47988 800
rect 48024 0 48080 800
rect 48208 0 48264 800
rect 48300 0 48356 800
rect 48392 0 48448 800
rect 48576 0 48632 800
rect 48668 0 48724 800
rect 48760 0 48816 800
rect 48944 0 49000 800
rect 49036 0 49092 800
rect 49128 0 49184 800
rect 49312 0 49368 800
rect 49404 0 49460 800
rect 49496 0 49552 800
rect 49680 0 49736 800
rect 49772 0 49828 800
rect 49864 0 49920 800
rect 50048 0 50104 800
rect 50140 0 50196 800
rect 50232 0 50288 800
rect 50416 0 50472 800
rect 50508 0 50564 800
rect 50600 0 50656 800
rect 50784 0 50840 800
rect 50876 0 50932 800
rect 50968 0 51024 800
rect 51152 0 51208 800
rect 51244 0 51300 800
rect 51336 0 51392 800
rect 51520 0 51576 800
rect 51612 0 51668 800
rect 51704 0 51760 800
rect 51888 0 51944 800
rect 51980 0 52036 800
rect 52072 0 52128 800
rect 52256 0 52312 800
rect 52348 0 52404 800
rect 52440 0 52496 800
rect 52624 0 52680 800
rect 52716 0 52772 800
rect 52808 0 52864 800
rect 52992 0 53048 800
rect 53084 0 53140 800
rect 53176 0 53232 800
rect 53360 0 53416 800
rect 53452 0 53508 800
rect 53544 0 53600 800
rect 53728 0 53784 800
rect 53820 0 53876 800
rect 53912 0 53968 800
rect 54096 0 54152 800
rect 54188 0 54244 800
rect 54280 0 54336 800
rect 54464 0 54520 800
rect 54556 0 54612 800
rect 54648 0 54704 800
rect 54832 0 54888 800
rect 54924 0 54980 800
rect 55016 0 55072 800
rect 55200 0 55256 800
rect 55292 0 55348 800
rect 55384 0 55440 800
rect 55568 0 55624 800
rect 55660 0 55716 800
rect 55752 0 55808 800
rect 55936 0 55992 800
rect 56028 0 56084 800
rect 56120 0 56176 800
rect 56304 0 56360 800
rect 56396 0 56452 800
rect 56488 0 56544 800
rect 56672 0 56728 800
rect 56764 0 56820 800
rect 56856 0 56912 800
rect 57040 0 57096 800
rect 57132 0 57188 800
rect 57224 0 57280 800
rect 57408 0 57464 800
rect 57500 0 57556 800
rect 57592 0 57648 800
rect 57776 0 57832 800
rect 57868 0 57924 800
rect 57960 0 58016 800
rect 58144 0 58200 800
rect 58236 0 58292 800
rect 58328 0 58384 800
rect 58512 0 58568 800
rect 58604 0 58660 800
rect 58696 0 58752 800
rect 58880 0 58936 800
rect 58972 0 59028 800
rect 59064 0 59120 800
rect 59248 0 59304 800
rect 59340 0 59396 800
rect 59432 0 59488 800
rect 59616 0 59672 800
rect 59708 0 59764 800
rect 59800 0 59856 800
<< via2 >>
rect 2116 55800 2172 55856
rect 4202 57690 4258 57692
rect 4282 57690 4338 57692
rect 4362 57690 4418 57692
rect 4442 57690 4498 57692
rect 4202 57638 4228 57690
rect 4228 57638 4258 57690
rect 4282 57638 4292 57690
rect 4292 57638 4338 57690
rect 4362 57638 4408 57690
rect 4408 57638 4418 57690
rect 4442 57638 4472 57690
rect 4472 57638 4498 57690
rect 4202 57636 4258 57638
rect 4282 57636 4338 57638
rect 4362 57636 4418 57638
rect 4442 57636 4498 57638
rect 4202 56602 4258 56604
rect 4282 56602 4338 56604
rect 4362 56602 4418 56604
rect 4442 56602 4498 56604
rect 4202 56550 4228 56602
rect 4228 56550 4258 56602
rect 4282 56550 4292 56602
rect 4292 56550 4338 56602
rect 4362 56550 4408 56602
rect 4408 56550 4418 56602
rect 4442 56550 4472 56602
rect 4472 56550 4498 56602
rect 4202 56548 4258 56550
rect 4282 56548 4338 56550
rect 4362 56548 4418 56550
rect 4442 56548 4498 56550
rect 3404 18128 3460 18184
rect 3588 17992 3644 18048
rect 4202 55514 4258 55516
rect 4282 55514 4338 55516
rect 4362 55514 4418 55516
rect 4442 55514 4498 55516
rect 4202 55462 4228 55514
rect 4228 55462 4258 55514
rect 4282 55462 4292 55514
rect 4292 55462 4338 55514
rect 4362 55462 4408 55514
rect 4408 55462 4418 55514
rect 4442 55462 4472 55514
rect 4472 55462 4498 55514
rect 4202 55460 4258 55462
rect 4282 55460 4338 55462
rect 4362 55460 4418 55462
rect 4442 55460 4498 55462
rect 4202 54426 4258 54428
rect 4282 54426 4338 54428
rect 4362 54426 4418 54428
rect 4442 54426 4498 54428
rect 4202 54374 4228 54426
rect 4228 54374 4258 54426
rect 4282 54374 4292 54426
rect 4292 54374 4338 54426
rect 4362 54374 4408 54426
rect 4408 54374 4418 54426
rect 4442 54374 4472 54426
rect 4472 54374 4498 54426
rect 4202 54372 4258 54374
rect 4282 54372 4338 54374
rect 4362 54372 4418 54374
rect 4442 54372 4498 54374
rect 4202 53338 4258 53340
rect 4282 53338 4338 53340
rect 4362 53338 4418 53340
rect 4442 53338 4498 53340
rect 4202 53286 4228 53338
rect 4228 53286 4258 53338
rect 4282 53286 4292 53338
rect 4292 53286 4338 53338
rect 4362 53286 4408 53338
rect 4408 53286 4418 53338
rect 4442 53286 4472 53338
rect 4472 53286 4498 53338
rect 4202 53284 4258 53286
rect 4282 53284 4338 53286
rect 4362 53284 4418 53286
rect 4442 53284 4498 53286
rect 4202 52250 4258 52252
rect 4282 52250 4338 52252
rect 4362 52250 4418 52252
rect 4442 52250 4498 52252
rect 4202 52198 4228 52250
rect 4228 52198 4258 52250
rect 4282 52198 4292 52250
rect 4292 52198 4338 52250
rect 4362 52198 4408 52250
rect 4408 52198 4418 52250
rect 4442 52198 4472 52250
rect 4472 52198 4498 52250
rect 4202 52196 4258 52198
rect 4282 52196 4338 52198
rect 4362 52196 4418 52198
rect 4442 52196 4498 52198
rect 4202 51162 4258 51164
rect 4282 51162 4338 51164
rect 4362 51162 4418 51164
rect 4442 51162 4498 51164
rect 4202 51110 4228 51162
rect 4228 51110 4258 51162
rect 4282 51110 4292 51162
rect 4292 51110 4338 51162
rect 4362 51110 4408 51162
rect 4408 51110 4418 51162
rect 4442 51110 4472 51162
rect 4472 51110 4498 51162
rect 4202 51108 4258 51110
rect 4282 51108 4338 51110
rect 4362 51108 4418 51110
rect 4442 51108 4498 51110
rect 4202 50074 4258 50076
rect 4282 50074 4338 50076
rect 4362 50074 4418 50076
rect 4442 50074 4498 50076
rect 4202 50022 4228 50074
rect 4228 50022 4258 50074
rect 4282 50022 4292 50074
rect 4292 50022 4338 50074
rect 4362 50022 4408 50074
rect 4408 50022 4418 50074
rect 4442 50022 4472 50074
rect 4472 50022 4498 50074
rect 4202 50020 4258 50022
rect 4282 50020 4338 50022
rect 4362 50020 4418 50022
rect 4442 50020 4498 50022
rect 4202 48986 4258 48988
rect 4282 48986 4338 48988
rect 4362 48986 4418 48988
rect 4442 48986 4498 48988
rect 4202 48934 4228 48986
rect 4228 48934 4258 48986
rect 4282 48934 4292 48986
rect 4292 48934 4338 48986
rect 4362 48934 4408 48986
rect 4408 48934 4418 48986
rect 4442 48934 4472 48986
rect 4472 48934 4498 48986
rect 4202 48932 4258 48934
rect 4282 48932 4338 48934
rect 4362 48932 4418 48934
rect 4442 48932 4498 48934
rect 4202 47898 4258 47900
rect 4282 47898 4338 47900
rect 4362 47898 4418 47900
rect 4442 47898 4498 47900
rect 4202 47846 4228 47898
rect 4228 47846 4258 47898
rect 4282 47846 4292 47898
rect 4292 47846 4338 47898
rect 4362 47846 4408 47898
rect 4408 47846 4418 47898
rect 4442 47846 4472 47898
rect 4472 47846 4498 47898
rect 4202 47844 4258 47846
rect 4282 47844 4338 47846
rect 4362 47844 4418 47846
rect 4442 47844 4498 47846
rect 4202 46810 4258 46812
rect 4282 46810 4338 46812
rect 4362 46810 4418 46812
rect 4442 46810 4498 46812
rect 4202 46758 4228 46810
rect 4228 46758 4258 46810
rect 4282 46758 4292 46810
rect 4292 46758 4338 46810
rect 4362 46758 4408 46810
rect 4408 46758 4418 46810
rect 4442 46758 4472 46810
rect 4472 46758 4498 46810
rect 4202 46756 4258 46758
rect 4282 46756 4338 46758
rect 4362 46756 4418 46758
rect 4442 46756 4498 46758
rect 4202 45722 4258 45724
rect 4282 45722 4338 45724
rect 4362 45722 4418 45724
rect 4442 45722 4498 45724
rect 4202 45670 4228 45722
rect 4228 45670 4258 45722
rect 4282 45670 4292 45722
rect 4292 45670 4338 45722
rect 4362 45670 4408 45722
rect 4408 45670 4418 45722
rect 4442 45670 4472 45722
rect 4472 45670 4498 45722
rect 4202 45668 4258 45670
rect 4282 45668 4338 45670
rect 4362 45668 4418 45670
rect 4442 45668 4498 45670
rect 4202 44634 4258 44636
rect 4282 44634 4338 44636
rect 4362 44634 4418 44636
rect 4442 44634 4498 44636
rect 4202 44582 4228 44634
rect 4228 44582 4258 44634
rect 4282 44582 4292 44634
rect 4292 44582 4338 44634
rect 4362 44582 4408 44634
rect 4408 44582 4418 44634
rect 4442 44582 4472 44634
rect 4472 44582 4498 44634
rect 4202 44580 4258 44582
rect 4282 44580 4338 44582
rect 4362 44580 4418 44582
rect 4442 44580 4498 44582
rect 4202 43546 4258 43548
rect 4282 43546 4338 43548
rect 4362 43546 4418 43548
rect 4442 43546 4498 43548
rect 4202 43494 4228 43546
rect 4228 43494 4258 43546
rect 4282 43494 4292 43546
rect 4292 43494 4338 43546
rect 4362 43494 4408 43546
rect 4408 43494 4418 43546
rect 4442 43494 4472 43546
rect 4472 43494 4498 43546
rect 4202 43492 4258 43494
rect 4282 43492 4338 43494
rect 4362 43492 4418 43494
rect 4442 43492 4498 43494
rect 4202 42458 4258 42460
rect 4282 42458 4338 42460
rect 4362 42458 4418 42460
rect 4442 42458 4498 42460
rect 4202 42406 4228 42458
rect 4228 42406 4258 42458
rect 4282 42406 4292 42458
rect 4292 42406 4338 42458
rect 4362 42406 4408 42458
rect 4408 42406 4418 42458
rect 4442 42406 4472 42458
rect 4472 42406 4498 42458
rect 4202 42404 4258 42406
rect 4282 42404 4338 42406
rect 4362 42404 4418 42406
rect 4442 42404 4498 42406
rect 4202 41370 4258 41372
rect 4282 41370 4338 41372
rect 4362 41370 4418 41372
rect 4442 41370 4498 41372
rect 4202 41318 4228 41370
rect 4228 41318 4258 41370
rect 4282 41318 4292 41370
rect 4292 41318 4338 41370
rect 4362 41318 4408 41370
rect 4408 41318 4418 41370
rect 4442 41318 4472 41370
rect 4472 41318 4498 41370
rect 4202 41316 4258 41318
rect 4282 41316 4338 41318
rect 4362 41316 4418 41318
rect 4442 41316 4498 41318
rect 4202 40282 4258 40284
rect 4282 40282 4338 40284
rect 4362 40282 4418 40284
rect 4442 40282 4498 40284
rect 4202 40230 4228 40282
rect 4228 40230 4258 40282
rect 4282 40230 4292 40282
rect 4292 40230 4338 40282
rect 4362 40230 4408 40282
rect 4408 40230 4418 40282
rect 4442 40230 4472 40282
rect 4472 40230 4498 40282
rect 4202 40228 4258 40230
rect 4282 40228 4338 40230
rect 4362 40228 4418 40230
rect 4442 40228 4498 40230
rect 4202 39194 4258 39196
rect 4282 39194 4338 39196
rect 4362 39194 4418 39196
rect 4442 39194 4498 39196
rect 4202 39142 4228 39194
rect 4228 39142 4258 39194
rect 4282 39142 4292 39194
rect 4292 39142 4338 39194
rect 4362 39142 4408 39194
rect 4408 39142 4418 39194
rect 4442 39142 4472 39194
rect 4472 39142 4498 39194
rect 4202 39140 4258 39142
rect 4282 39140 4338 39142
rect 4362 39140 4418 39142
rect 4442 39140 4498 39142
rect 4202 38106 4258 38108
rect 4282 38106 4338 38108
rect 4362 38106 4418 38108
rect 4442 38106 4498 38108
rect 4202 38054 4228 38106
rect 4228 38054 4258 38106
rect 4282 38054 4292 38106
rect 4292 38054 4338 38106
rect 4362 38054 4408 38106
rect 4408 38054 4418 38106
rect 4442 38054 4472 38106
rect 4472 38054 4498 38106
rect 4202 38052 4258 38054
rect 4282 38052 4338 38054
rect 4362 38052 4418 38054
rect 4442 38052 4498 38054
rect 4202 37018 4258 37020
rect 4282 37018 4338 37020
rect 4362 37018 4418 37020
rect 4442 37018 4498 37020
rect 4202 36966 4228 37018
rect 4228 36966 4258 37018
rect 4282 36966 4292 37018
rect 4292 36966 4338 37018
rect 4362 36966 4408 37018
rect 4408 36966 4418 37018
rect 4442 36966 4472 37018
rect 4472 36966 4498 37018
rect 4202 36964 4258 36966
rect 4282 36964 4338 36966
rect 4362 36964 4418 36966
rect 4442 36964 4498 36966
rect 4202 35930 4258 35932
rect 4282 35930 4338 35932
rect 4362 35930 4418 35932
rect 4442 35930 4498 35932
rect 4202 35878 4228 35930
rect 4228 35878 4258 35930
rect 4282 35878 4292 35930
rect 4292 35878 4338 35930
rect 4362 35878 4408 35930
rect 4408 35878 4418 35930
rect 4442 35878 4472 35930
rect 4472 35878 4498 35930
rect 4202 35876 4258 35878
rect 4282 35876 4338 35878
rect 4362 35876 4418 35878
rect 4442 35876 4498 35878
rect 4202 34842 4258 34844
rect 4282 34842 4338 34844
rect 4362 34842 4418 34844
rect 4442 34842 4498 34844
rect 4202 34790 4228 34842
rect 4228 34790 4258 34842
rect 4282 34790 4292 34842
rect 4292 34790 4338 34842
rect 4362 34790 4408 34842
rect 4408 34790 4418 34842
rect 4442 34790 4472 34842
rect 4472 34790 4498 34842
rect 4202 34788 4258 34790
rect 4282 34788 4338 34790
rect 4362 34788 4418 34790
rect 4442 34788 4498 34790
rect 4202 33754 4258 33756
rect 4282 33754 4338 33756
rect 4362 33754 4418 33756
rect 4442 33754 4498 33756
rect 4202 33702 4228 33754
rect 4228 33702 4258 33754
rect 4282 33702 4292 33754
rect 4292 33702 4338 33754
rect 4362 33702 4408 33754
rect 4408 33702 4418 33754
rect 4442 33702 4472 33754
rect 4472 33702 4498 33754
rect 4202 33700 4258 33702
rect 4282 33700 4338 33702
rect 4362 33700 4418 33702
rect 4442 33700 4498 33702
rect 4202 32666 4258 32668
rect 4282 32666 4338 32668
rect 4362 32666 4418 32668
rect 4442 32666 4498 32668
rect 4202 32614 4228 32666
rect 4228 32614 4258 32666
rect 4282 32614 4292 32666
rect 4292 32614 4338 32666
rect 4362 32614 4408 32666
rect 4408 32614 4418 32666
rect 4442 32614 4472 32666
rect 4472 32614 4498 32666
rect 4202 32612 4258 32614
rect 4282 32612 4338 32614
rect 4362 32612 4418 32614
rect 4442 32612 4498 32614
rect 4202 31578 4258 31580
rect 4282 31578 4338 31580
rect 4362 31578 4418 31580
rect 4442 31578 4498 31580
rect 4202 31526 4228 31578
rect 4228 31526 4258 31578
rect 4282 31526 4292 31578
rect 4292 31526 4338 31578
rect 4362 31526 4408 31578
rect 4408 31526 4418 31578
rect 4442 31526 4472 31578
rect 4472 31526 4498 31578
rect 4202 31524 4258 31526
rect 4282 31524 4338 31526
rect 4362 31524 4418 31526
rect 4442 31524 4498 31526
rect 4202 30490 4258 30492
rect 4282 30490 4338 30492
rect 4362 30490 4418 30492
rect 4442 30490 4498 30492
rect 4202 30438 4228 30490
rect 4228 30438 4258 30490
rect 4282 30438 4292 30490
rect 4292 30438 4338 30490
rect 4362 30438 4408 30490
rect 4408 30438 4418 30490
rect 4442 30438 4472 30490
rect 4472 30438 4498 30490
rect 4202 30436 4258 30438
rect 4282 30436 4338 30438
rect 4362 30436 4418 30438
rect 4442 30436 4498 30438
rect 4202 29402 4258 29404
rect 4282 29402 4338 29404
rect 4362 29402 4418 29404
rect 4442 29402 4498 29404
rect 4202 29350 4228 29402
rect 4228 29350 4258 29402
rect 4282 29350 4292 29402
rect 4292 29350 4338 29402
rect 4362 29350 4408 29402
rect 4408 29350 4418 29402
rect 4442 29350 4472 29402
rect 4472 29350 4498 29402
rect 4202 29348 4258 29350
rect 4282 29348 4338 29350
rect 4362 29348 4418 29350
rect 4442 29348 4498 29350
rect 4202 28314 4258 28316
rect 4282 28314 4338 28316
rect 4362 28314 4418 28316
rect 4442 28314 4498 28316
rect 4202 28262 4228 28314
rect 4228 28262 4258 28314
rect 4282 28262 4292 28314
rect 4292 28262 4338 28314
rect 4362 28262 4408 28314
rect 4408 28262 4418 28314
rect 4442 28262 4472 28314
rect 4472 28262 4498 28314
rect 4202 28260 4258 28262
rect 4282 28260 4338 28262
rect 4362 28260 4418 28262
rect 4442 28260 4498 28262
rect 4202 27226 4258 27228
rect 4282 27226 4338 27228
rect 4362 27226 4418 27228
rect 4442 27226 4498 27228
rect 4202 27174 4228 27226
rect 4228 27174 4258 27226
rect 4282 27174 4292 27226
rect 4292 27174 4338 27226
rect 4362 27174 4408 27226
rect 4408 27174 4418 27226
rect 4442 27174 4472 27226
rect 4472 27174 4498 27226
rect 4202 27172 4258 27174
rect 4282 27172 4338 27174
rect 4362 27172 4418 27174
rect 4442 27172 4498 27174
rect 4202 26138 4258 26140
rect 4282 26138 4338 26140
rect 4362 26138 4418 26140
rect 4442 26138 4498 26140
rect 4202 26086 4228 26138
rect 4228 26086 4258 26138
rect 4282 26086 4292 26138
rect 4292 26086 4338 26138
rect 4362 26086 4408 26138
rect 4408 26086 4418 26138
rect 4442 26086 4472 26138
rect 4472 26086 4498 26138
rect 4202 26084 4258 26086
rect 4282 26084 4338 26086
rect 4362 26084 4418 26086
rect 4442 26084 4498 26086
rect 4202 25050 4258 25052
rect 4282 25050 4338 25052
rect 4362 25050 4418 25052
rect 4442 25050 4498 25052
rect 4202 24998 4228 25050
rect 4228 24998 4258 25050
rect 4282 24998 4292 25050
rect 4292 24998 4338 25050
rect 4362 24998 4408 25050
rect 4408 24998 4418 25050
rect 4442 24998 4472 25050
rect 4472 24998 4498 25050
rect 4202 24996 4258 24998
rect 4282 24996 4338 24998
rect 4362 24996 4418 24998
rect 4442 24996 4498 24998
rect 4202 23962 4258 23964
rect 4282 23962 4338 23964
rect 4362 23962 4418 23964
rect 4442 23962 4498 23964
rect 4202 23910 4228 23962
rect 4228 23910 4258 23962
rect 4282 23910 4292 23962
rect 4292 23910 4338 23962
rect 4362 23910 4408 23962
rect 4408 23910 4418 23962
rect 4442 23910 4472 23962
rect 4472 23910 4498 23962
rect 4202 23908 4258 23910
rect 4282 23908 4338 23910
rect 4362 23908 4418 23910
rect 4442 23908 4498 23910
rect 4202 22874 4258 22876
rect 4282 22874 4338 22876
rect 4362 22874 4418 22876
rect 4442 22874 4498 22876
rect 4202 22822 4228 22874
rect 4228 22822 4258 22874
rect 4282 22822 4292 22874
rect 4292 22822 4338 22874
rect 4362 22822 4408 22874
rect 4408 22822 4418 22874
rect 4442 22822 4472 22874
rect 4472 22822 4498 22874
rect 4202 22820 4258 22822
rect 4282 22820 4338 22822
rect 4362 22820 4418 22822
rect 4442 22820 4498 22822
rect 4202 21786 4258 21788
rect 4282 21786 4338 21788
rect 4362 21786 4418 21788
rect 4442 21786 4498 21788
rect 4202 21734 4228 21786
rect 4228 21734 4258 21786
rect 4282 21734 4292 21786
rect 4292 21734 4338 21786
rect 4362 21734 4408 21786
rect 4408 21734 4418 21786
rect 4442 21734 4472 21786
rect 4472 21734 4498 21786
rect 4202 21732 4258 21734
rect 4282 21732 4338 21734
rect 4362 21732 4418 21734
rect 4442 21732 4498 21734
rect 4202 20698 4258 20700
rect 4282 20698 4338 20700
rect 4362 20698 4418 20700
rect 4442 20698 4498 20700
rect 4202 20646 4228 20698
rect 4228 20646 4258 20698
rect 4282 20646 4292 20698
rect 4292 20646 4338 20698
rect 4362 20646 4408 20698
rect 4408 20646 4418 20698
rect 4442 20646 4472 20698
rect 4472 20646 4498 20698
rect 4202 20644 4258 20646
rect 4282 20644 4338 20646
rect 4362 20644 4418 20646
rect 4442 20644 4498 20646
rect 4202 19610 4258 19612
rect 4282 19610 4338 19612
rect 4362 19610 4418 19612
rect 4442 19610 4498 19612
rect 4202 19558 4228 19610
rect 4228 19558 4258 19610
rect 4282 19558 4292 19610
rect 4292 19558 4338 19610
rect 4362 19558 4408 19610
rect 4408 19558 4418 19610
rect 4442 19558 4472 19610
rect 4472 19558 4498 19610
rect 4202 19556 4258 19558
rect 4282 19556 4338 19558
rect 4362 19556 4418 19558
rect 4442 19556 4498 19558
rect 4202 18522 4258 18524
rect 4282 18522 4338 18524
rect 4362 18522 4418 18524
rect 4442 18522 4498 18524
rect 4202 18470 4228 18522
rect 4228 18470 4258 18522
rect 4282 18470 4292 18522
rect 4292 18470 4338 18522
rect 4362 18470 4408 18522
rect 4408 18470 4418 18522
rect 4442 18470 4472 18522
rect 4472 18470 4498 18522
rect 4202 18468 4258 18470
rect 4282 18468 4338 18470
rect 4362 18468 4418 18470
rect 4442 18468 4498 18470
rect 4202 17434 4258 17436
rect 4282 17434 4338 17436
rect 4362 17434 4418 17436
rect 4442 17434 4498 17436
rect 4202 17382 4228 17434
rect 4228 17382 4258 17434
rect 4282 17382 4292 17434
rect 4292 17382 4338 17434
rect 4362 17382 4408 17434
rect 4408 17382 4418 17434
rect 4442 17382 4472 17434
rect 4472 17382 4498 17434
rect 4202 17380 4258 17382
rect 4282 17380 4338 17382
rect 4362 17380 4418 17382
rect 4442 17380 4498 17382
rect 4202 16346 4258 16348
rect 4282 16346 4338 16348
rect 4362 16346 4418 16348
rect 4442 16346 4498 16348
rect 4202 16294 4228 16346
rect 4228 16294 4258 16346
rect 4282 16294 4292 16346
rect 4292 16294 4338 16346
rect 4362 16294 4408 16346
rect 4408 16294 4418 16346
rect 4442 16294 4472 16346
rect 4472 16294 4498 16346
rect 4202 16292 4258 16294
rect 4282 16292 4338 16294
rect 4362 16292 4418 16294
rect 4442 16292 4498 16294
rect 4202 15258 4258 15260
rect 4282 15258 4338 15260
rect 4362 15258 4418 15260
rect 4442 15258 4498 15260
rect 4202 15206 4228 15258
rect 4228 15206 4258 15258
rect 4282 15206 4292 15258
rect 4292 15206 4338 15258
rect 4362 15206 4408 15258
rect 4408 15206 4418 15258
rect 4442 15206 4472 15258
rect 4472 15206 4498 15258
rect 4202 15204 4258 15206
rect 4282 15204 4338 15206
rect 4362 15204 4418 15206
rect 4442 15204 4498 15206
rect 4202 14170 4258 14172
rect 4282 14170 4338 14172
rect 4362 14170 4418 14172
rect 4442 14170 4498 14172
rect 4202 14118 4228 14170
rect 4228 14118 4258 14170
rect 4282 14118 4292 14170
rect 4292 14118 4338 14170
rect 4362 14118 4408 14170
rect 4408 14118 4418 14170
rect 4442 14118 4472 14170
rect 4472 14118 4498 14170
rect 4202 14116 4258 14118
rect 4282 14116 4338 14118
rect 4362 14116 4418 14118
rect 4442 14116 4498 14118
rect 4202 13082 4258 13084
rect 4282 13082 4338 13084
rect 4362 13082 4418 13084
rect 4442 13082 4498 13084
rect 4202 13030 4228 13082
rect 4228 13030 4258 13082
rect 4282 13030 4292 13082
rect 4292 13030 4338 13082
rect 4362 13030 4408 13082
rect 4408 13030 4418 13082
rect 4442 13030 4472 13082
rect 4472 13030 4498 13082
rect 4202 13028 4258 13030
rect 4282 13028 4338 13030
rect 4362 13028 4418 13030
rect 4442 13028 4498 13030
rect 4202 11994 4258 11996
rect 4282 11994 4338 11996
rect 4362 11994 4418 11996
rect 4442 11994 4498 11996
rect 4202 11942 4228 11994
rect 4228 11942 4258 11994
rect 4282 11942 4292 11994
rect 4292 11942 4338 11994
rect 4362 11942 4408 11994
rect 4408 11942 4418 11994
rect 4442 11942 4472 11994
rect 4472 11942 4498 11994
rect 4202 11940 4258 11942
rect 4282 11940 4338 11942
rect 4362 11940 4418 11942
rect 4442 11940 4498 11942
rect 4202 10906 4258 10908
rect 4282 10906 4338 10908
rect 4362 10906 4418 10908
rect 4442 10906 4498 10908
rect 4202 10854 4228 10906
rect 4228 10854 4258 10906
rect 4282 10854 4292 10906
rect 4292 10854 4338 10906
rect 4362 10854 4408 10906
rect 4408 10854 4418 10906
rect 4442 10854 4472 10906
rect 4472 10854 4498 10906
rect 4202 10852 4258 10854
rect 4282 10852 4338 10854
rect 4362 10852 4418 10854
rect 4442 10852 4498 10854
rect 4202 9818 4258 9820
rect 4282 9818 4338 9820
rect 4362 9818 4418 9820
rect 4442 9818 4498 9820
rect 4202 9766 4228 9818
rect 4228 9766 4258 9818
rect 4282 9766 4292 9818
rect 4292 9766 4338 9818
rect 4362 9766 4408 9818
rect 4408 9766 4418 9818
rect 4442 9766 4472 9818
rect 4472 9766 4498 9818
rect 4202 9764 4258 9766
rect 4282 9764 4338 9766
rect 4362 9764 4418 9766
rect 4442 9764 4498 9766
rect 4202 8730 4258 8732
rect 4282 8730 4338 8732
rect 4362 8730 4418 8732
rect 4442 8730 4498 8732
rect 4202 8678 4228 8730
rect 4228 8678 4258 8730
rect 4282 8678 4292 8730
rect 4292 8678 4338 8730
rect 4362 8678 4408 8730
rect 4408 8678 4418 8730
rect 4442 8678 4472 8730
rect 4472 8678 4498 8730
rect 4202 8676 4258 8678
rect 4282 8676 4338 8678
rect 4362 8676 4418 8678
rect 4442 8676 4498 8678
rect 4202 7642 4258 7644
rect 4282 7642 4338 7644
rect 4362 7642 4418 7644
rect 4442 7642 4498 7644
rect 4202 7590 4228 7642
rect 4228 7590 4258 7642
rect 4282 7590 4292 7642
rect 4292 7590 4338 7642
rect 4362 7590 4408 7642
rect 4408 7590 4418 7642
rect 4442 7590 4472 7642
rect 4472 7590 4498 7642
rect 4202 7588 4258 7590
rect 4282 7588 4338 7590
rect 4362 7588 4418 7590
rect 4442 7588 4498 7590
rect 4202 6554 4258 6556
rect 4282 6554 4338 6556
rect 4362 6554 4418 6556
rect 4442 6554 4498 6556
rect 4202 6502 4228 6554
rect 4228 6502 4258 6554
rect 4282 6502 4292 6554
rect 4292 6502 4338 6554
rect 4362 6502 4408 6554
rect 4408 6502 4418 6554
rect 4442 6502 4472 6554
rect 4472 6502 4498 6554
rect 4202 6500 4258 6502
rect 4282 6500 4338 6502
rect 4362 6500 4418 6502
rect 4442 6500 4498 6502
rect 4202 5466 4258 5468
rect 4282 5466 4338 5468
rect 4362 5466 4418 5468
rect 4442 5466 4498 5468
rect 4202 5414 4228 5466
rect 4228 5414 4258 5466
rect 4282 5414 4292 5466
rect 4292 5414 4338 5466
rect 4362 5414 4408 5466
rect 4408 5414 4418 5466
rect 4442 5414 4472 5466
rect 4472 5414 4498 5466
rect 4202 5412 4258 5414
rect 4282 5412 4338 5414
rect 4362 5412 4418 5414
rect 4442 5412 4498 5414
rect 4202 4378 4258 4380
rect 4282 4378 4338 4380
rect 4362 4378 4418 4380
rect 4442 4378 4498 4380
rect 4202 4326 4228 4378
rect 4228 4326 4258 4378
rect 4282 4326 4292 4378
rect 4292 4326 4338 4378
rect 4362 4326 4408 4378
rect 4408 4326 4418 4378
rect 4442 4326 4472 4378
rect 4472 4326 4498 4378
rect 4202 4324 4258 4326
rect 4282 4324 4338 4326
rect 4362 4324 4418 4326
rect 4442 4324 4498 4326
rect 4202 3290 4258 3292
rect 4282 3290 4338 3292
rect 4362 3290 4418 3292
rect 4442 3290 4498 3292
rect 4202 3238 4228 3290
rect 4228 3238 4258 3290
rect 4282 3238 4292 3290
rect 4292 3238 4338 3290
rect 4362 3238 4408 3290
rect 4408 3238 4418 3290
rect 4442 3238 4472 3290
rect 4472 3238 4498 3290
rect 4202 3236 4258 3238
rect 4282 3236 4338 3238
rect 4362 3236 4418 3238
rect 4442 3236 4498 3238
rect 4202 2202 4258 2204
rect 4282 2202 4338 2204
rect 4362 2202 4418 2204
rect 4442 2202 4498 2204
rect 4202 2150 4228 2202
rect 4228 2150 4258 2202
rect 4282 2150 4292 2202
rect 4292 2150 4338 2202
rect 4362 2150 4408 2202
rect 4408 2150 4418 2202
rect 4442 2150 4472 2202
rect 4472 2150 4498 2202
rect 4202 2148 4258 2150
rect 4282 2148 4338 2150
rect 4362 2148 4418 2150
rect 4442 2148 4498 2150
rect 5244 17992 5300 18048
rect 5428 17992 5484 18048
rect 8004 19252 8006 19272
rect 8006 19252 8058 19272
rect 8058 19252 8060 19272
rect 8004 19216 8060 19252
rect 8004 13932 8060 13968
rect 8004 13912 8006 13932
rect 8006 13912 8058 13932
rect 8058 13912 8060 13932
rect 8464 23604 8466 23624
rect 8466 23604 8518 23624
rect 8518 23604 8520 23624
rect 8464 23568 8520 23604
rect 8924 19216 8980 19272
rect 8832 18420 8888 18456
rect 8832 18400 8834 18420
rect 8834 18400 8886 18420
rect 8886 18400 8888 18420
rect 9016 18420 9072 18456
rect 9016 18400 9018 18420
rect 9018 18400 9070 18420
rect 9070 18400 9072 18420
rect 8280 14918 8336 14920
rect 8280 14866 8282 14918
rect 8282 14866 8334 14918
rect 8334 14866 8336 14918
rect 8280 14864 8336 14866
rect 8648 14864 8704 14920
rect 8832 13912 8888 13968
rect 9108 17176 9164 17232
rect 8234 7302 8290 7304
rect 8234 7250 8236 7302
rect 8236 7250 8288 7302
rect 8288 7250 8290 7302
rect 8234 7248 8290 7250
rect 9568 17212 9570 17232
rect 9570 17212 9622 17232
rect 9622 17212 9624 17232
rect 9568 17176 9624 17212
rect 11776 23568 11832 23624
rect 12696 7248 12752 7304
rect 14168 35944 14224 36000
rect 14352 35944 14408 36000
rect 19562 57146 19618 57148
rect 19642 57146 19698 57148
rect 19722 57146 19778 57148
rect 19802 57146 19858 57148
rect 19562 57094 19588 57146
rect 19588 57094 19618 57146
rect 19642 57094 19652 57146
rect 19652 57094 19698 57146
rect 19722 57094 19768 57146
rect 19768 57094 19778 57146
rect 19802 57094 19832 57146
rect 19832 57094 19858 57146
rect 19562 57092 19618 57094
rect 19642 57092 19698 57094
rect 19722 57092 19778 57094
rect 19802 57092 19858 57094
rect 19562 56058 19618 56060
rect 19642 56058 19698 56060
rect 19722 56058 19778 56060
rect 19802 56058 19858 56060
rect 19562 56006 19588 56058
rect 19588 56006 19618 56058
rect 19642 56006 19652 56058
rect 19652 56006 19698 56058
rect 19722 56006 19768 56058
rect 19768 56006 19778 56058
rect 19802 56006 19832 56058
rect 19832 56006 19858 56058
rect 19562 56004 19618 56006
rect 19642 56004 19698 56006
rect 19722 56004 19778 56006
rect 19802 56004 19858 56006
rect 19136 37168 19192 37224
rect 19562 54970 19618 54972
rect 19642 54970 19698 54972
rect 19722 54970 19778 54972
rect 19802 54970 19858 54972
rect 19562 54918 19588 54970
rect 19588 54918 19618 54970
rect 19642 54918 19652 54970
rect 19652 54918 19698 54970
rect 19722 54918 19768 54970
rect 19768 54918 19778 54970
rect 19802 54918 19832 54970
rect 19832 54918 19858 54970
rect 19562 54916 19618 54918
rect 19642 54916 19698 54918
rect 19722 54916 19778 54918
rect 19802 54916 19858 54918
rect 19562 53882 19618 53884
rect 19642 53882 19698 53884
rect 19722 53882 19778 53884
rect 19802 53882 19858 53884
rect 19562 53830 19588 53882
rect 19588 53830 19618 53882
rect 19642 53830 19652 53882
rect 19652 53830 19698 53882
rect 19722 53830 19768 53882
rect 19768 53830 19778 53882
rect 19802 53830 19832 53882
rect 19832 53830 19858 53882
rect 19562 53828 19618 53830
rect 19642 53828 19698 53830
rect 19722 53828 19778 53830
rect 19802 53828 19858 53830
rect 19562 52794 19618 52796
rect 19642 52794 19698 52796
rect 19722 52794 19778 52796
rect 19802 52794 19858 52796
rect 19562 52742 19588 52794
rect 19588 52742 19618 52794
rect 19642 52742 19652 52794
rect 19652 52742 19698 52794
rect 19722 52742 19768 52794
rect 19768 52742 19778 52794
rect 19802 52742 19832 52794
rect 19832 52742 19858 52794
rect 19562 52740 19618 52742
rect 19642 52740 19698 52742
rect 19722 52740 19778 52742
rect 19802 52740 19858 52742
rect 19562 51706 19618 51708
rect 19642 51706 19698 51708
rect 19722 51706 19778 51708
rect 19802 51706 19858 51708
rect 19562 51654 19588 51706
rect 19588 51654 19618 51706
rect 19642 51654 19652 51706
rect 19652 51654 19698 51706
rect 19722 51654 19768 51706
rect 19768 51654 19778 51706
rect 19802 51654 19832 51706
rect 19832 51654 19858 51706
rect 19562 51652 19618 51654
rect 19642 51652 19698 51654
rect 19722 51652 19778 51654
rect 19802 51652 19858 51654
rect 19562 50618 19618 50620
rect 19642 50618 19698 50620
rect 19722 50618 19778 50620
rect 19802 50618 19858 50620
rect 19562 50566 19588 50618
rect 19588 50566 19618 50618
rect 19642 50566 19652 50618
rect 19652 50566 19698 50618
rect 19722 50566 19768 50618
rect 19768 50566 19778 50618
rect 19802 50566 19832 50618
rect 19832 50566 19858 50618
rect 19562 50564 19618 50566
rect 19642 50564 19698 50566
rect 19722 50564 19778 50566
rect 19802 50564 19858 50566
rect 19562 49530 19618 49532
rect 19642 49530 19698 49532
rect 19722 49530 19778 49532
rect 19802 49530 19858 49532
rect 19562 49478 19588 49530
rect 19588 49478 19618 49530
rect 19642 49478 19652 49530
rect 19652 49478 19698 49530
rect 19722 49478 19768 49530
rect 19768 49478 19778 49530
rect 19802 49478 19832 49530
rect 19832 49478 19858 49530
rect 19562 49476 19618 49478
rect 19642 49476 19698 49478
rect 19722 49476 19778 49478
rect 19802 49476 19858 49478
rect 19562 48442 19618 48444
rect 19642 48442 19698 48444
rect 19722 48442 19778 48444
rect 19802 48442 19858 48444
rect 19562 48390 19588 48442
rect 19588 48390 19618 48442
rect 19642 48390 19652 48442
rect 19652 48390 19698 48442
rect 19722 48390 19768 48442
rect 19768 48390 19778 48442
rect 19802 48390 19832 48442
rect 19832 48390 19858 48442
rect 19562 48388 19618 48390
rect 19642 48388 19698 48390
rect 19722 48388 19778 48390
rect 19802 48388 19858 48390
rect 19562 47354 19618 47356
rect 19642 47354 19698 47356
rect 19722 47354 19778 47356
rect 19802 47354 19858 47356
rect 19562 47302 19588 47354
rect 19588 47302 19618 47354
rect 19642 47302 19652 47354
rect 19652 47302 19698 47354
rect 19722 47302 19768 47354
rect 19768 47302 19778 47354
rect 19802 47302 19832 47354
rect 19832 47302 19858 47354
rect 19562 47300 19618 47302
rect 19642 47300 19698 47302
rect 19722 47300 19778 47302
rect 19802 47300 19858 47302
rect 19562 46266 19618 46268
rect 19642 46266 19698 46268
rect 19722 46266 19778 46268
rect 19802 46266 19858 46268
rect 19562 46214 19588 46266
rect 19588 46214 19618 46266
rect 19642 46214 19652 46266
rect 19652 46214 19698 46266
rect 19722 46214 19768 46266
rect 19768 46214 19778 46266
rect 19802 46214 19832 46266
rect 19832 46214 19858 46266
rect 19562 46212 19618 46214
rect 19642 46212 19698 46214
rect 19722 46212 19778 46214
rect 19802 46212 19858 46214
rect 19562 45178 19618 45180
rect 19642 45178 19698 45180
rect 19722 45178 19778 45180
rect 19802 45178 19858 45180
rect 19562 45126 19588 45178
rect 19588 45126 19618 45178
rect 19642 45126 19652 45178
rect 19652 45126 19698 45178
rect 19722 45126 19768 45178
rect 19768 45126 19778 45178
rect 19802 45126 19832 45178
rect 19832 45126 19858 45178
rect 19562 45124 19618 45126
rect 19642 45124 19698 45126
rect 19722 45124 19778 45126
rect 19802 45124 19858 45126
rect 19562 44090 19618 44092
rect 19642 44090 19698 44092
rect 19722 44090 19778 44092
rect 19802 44090 19858 44092
rect 19562 44038 19588 44090
rect 19588 44038 19618 44090
rect 19642 44038 19652 44090
rect 19652 44038 19698 44090
rect 19722 44038 19768 44090
rect 19768 44038 19778 44090
rect 19802 44038 19832 44090
rect 19832 44038 19858 44090
rect 19562 44036 19618 44038
rect 19642 44036 19698 44038
rect 19722 44036 19778 44038
rect 19802 44036 19858 44038
rect 19562 43002 19618 43004
rect 19642 43002 19698 43004
rect 19722 43002 19778 43004
rect 19802 43002 19858 43004
rect 19562 42950 19588 43002
rect 19588 42950 19618 43002
rect 19642 42950 19652 43002
rect 19652 42950 19698 43002
rect 19722 42950 19768 43002
rect 19768 42950 19778 43002
rect 19802 42950 19832 43002
rect 19832 42950 19858 43002
rect 19562 42948 19618 42950
rect 19642 42948 19698 42950
rect 19722 42948 19778 42950
rect 19802 42948 19858 42950
rect 19562 41914 19618 41916
rect 19642 41914 19698 41916
rect 19722 41914 19778 41916
rect 19802 41914 19858 41916
rect 19562 41862 19588 41914
rect 19588 41862 19618 41914
rect 19642 41862 19652 41914
rect 19652 41862 19698 41914
rect 19722 41862 19768 41914
rect 19768 41862 19778 41914
rect 19802 41862 19832 41914
rect 19832 41862 19858 41914
rect 19562 41860 19618 41862
rect 19642 41860 19698 41862
rect 19722 41860 19778 41862
rect 19802 41860 19858 41862
rect 19562 40826 19618 40828
rect 19642 40826 19698 40828
rect 19722 40826 19778 40828
rect 19802 40826 19858 40828
rect 19562 40774 19588 40826
rect 19588 40774 19618 40826
rect 19642 40774 19652 40826
rect 19652 40774 19698 40826
rect 19722 40774 19768 40826
rect 19768 40774 19778 40826
rect 19802 40774 19832 40826
rect 19832 40774 19858 40826
rect 19562 40772 19618 40774
rect 19642 40772 19698 40774
rect 19722 40772 19778 40774
rect 19802 40772 19858 40774
rect 19562 39738 19618 39740
rect 19642 39738 19698 39740
rect 19722 39738 19778 39740
rect 19802 39738 19858 39740
rect 19562 39686 19588 39738
rect 19588 39686 19618 39738
rect 19642 39686 19652 39738
rect 19652 39686 19698 39738
rect 19722 39686 19768 39738
rect 19768 39686 19778 39738
rect 19802 39686 19832 39738
rect 19832 39686 19858 39738
rect 19562 39684 19618 39686
rect 19642 39684 19698 39686
rect 19722 39684 19778 39686
rect 19802 39684 19858 39686
rect 19562 38650 19618 38652
rect 19642 38650 19698 38652
rect 19722 38650 19778 38652
rect 19802 38650 19858 38652
rect 19562 38598 19588 38650
rect 19588 38598 19618 38650
rect 19642 38598 19652 38650
rect 19652 38598 19698 38650
rect 19722 38598 19768 38650
rect 19768 38598 19778 38650
rect 19802 38598 19832 38650
rect 19832 38598 19858 38650
rect 19562 38596 19618 38598
rect 19642 38596 19698 38598
rect 19722 38596 19778 38598
rect 19802 38596 19858 38598
rect 19562 37562 19618 37564
rect 19642 37562 19698 37564
rect 19722 37562 19778 37564
rect 19802 37562 19858 37564
rect 19562 37510 19588 37562
rect 19588 37510 19618 37562
rect 19642 37510 19652 37562
rect 19652 37510 19698 37562
rect 19722 37510 19768 37562
rect 19768 37510 19778 37562
rect 19802 37510 19832 37562
rect 19832 37510 19858 37562
rect 19562 37508 19618 37510
rect 19642 37508 19698 37510
rect 19722 37508 19778 37510
rect 19802 37508 19858 37510
rect 19562 36474 19618 36476
rect 19642 36474 19698 36476
rect 19722 36474 19778 36476
rect 19802 36474 19858 36476
rect 19562 36422 19588 36474
rect 19588 36422 19618 36474
rect 19642 36422 19652 36474
rect 19652 36422 19698 36474
rect 19722 36422 19768 36474
rect 19768 36422 19778 36474
rect 19802 36422 19832 36474
rect 19832 36422 19858 36474
rect 19562 36420 19618 36422
rect 19642 36420 19698 36422
rect 19722 36420 19778 36422
rect 19802 36420 19858 36422
rect 19562 35386 19618 35388
rect 19642 35386 19698 35388
rect 19722 35386 19778 35388
rect 19802 35386 19858 35388
rect 19562 35334 19588 35386
rect 19588 35334 19618 35386
rect 19642 35334 19652 35386
rect 19652 35334 19698 35386
rect 19722 35334 19768 35386
rect 19768 35334 19778 35386
rect 19802 35334 19832 35386
rect 19832 35334 19858 35386
rect 19562 35332 19618 35334
rect 19642 35332 19698 35334
rect 19722 35332 19778 35334
rect 19802 35332 19858 35334
rect 19562 34298 19618 34300
rect 19642 34298 19698 34300
rect 19722 34298 19778 34300
rect 19802 34298 19858 34300
rect 19562 34246 19588 34298
rect 19588 34246 19618 34298
rect 19642 34246 19652 34298
rect 19652 34246 19698 34298
rect 19722 34246 19768 34298
rect 19768 34246 19778 34298
rect 19802 34246 19832 34298
rect 19832 34246 19858 34298
rect 19562 34244 19618 34246
rect 19642 34244 19698 34246
rect 19722 34244 19778 34246
rect 19802 34244 19858 34246
rect 19562 33210 19618 33212
rect 19642 33210 19698 33212
rect 19722 33210 19778 33212
rect 19802 33210 19858 33212
rect 19562 33158 19588 33210
rect 19588 33158 19618 33210
rect 19642 33158 19652 33210
rect 19652 33158 19698 33210
rect 19722 33158 19768 33210
rect 19768 33158 19778 33210
rect 19802 33158 19832 33210
rect 19832 33158 19858 33210
rect 19562 33156 19618 33158
rect 19642 33156 19698 33158
rect 19722 33156 19778 33158
rect 19802 33156 19858 33158
rect 19562 32122 19618 32124
rect 19642 32122 19698 32124
rect 19722 32122 19778 32124
rect 19802 32122 19858 32124
rect 19562 32070 19588 32122
rect 19588 32070 19618 32122
rect 19642 32070 19652 32122
rect 19652 32070 19698 32122
rect 19722 32070 19768 32122
rect 19768 32070 19778 32122
rect 19802 32070 19832 32122
rect 19832 32070 19858 32122
rect 19562 32068 19618 32070
rect 19642 32068 19698 32070
rect 19722 32068 19778 32070
rect 19802 32068 19858 32070
rect 19562 31034 19618 31036
rect 19642 31034 19698 31036
rect 19722 31034 19778 31036
rect 19802 31034 19858 31036
rect 19562 30982 19588 31034
rect 19588 30982 19618 31034
rect 19642 30982 19652 31034
rect 19652 30982 19698 31034
rect 19722 30982 19768 31034
rect 19768 30982 19778 31034
rect 19802 30982 19832 31034
rect 19832 30982 19858 31034
rect 19562 30980 19618 30982
rect 19642 30980 19698 30982
rect 19722 30980 19778 30982
rect 19802 30980 19858 30982
rect 19562 29946 19618 29948
rect 19642 29946 19698 29948
rect 19722 29946 19778 29948
rect 19802 29946 19858 29948
rect 19562 29894 19588 29946
rect 19588 29894 19618 29946
rect 19642 29894 19652 29946
rect 19652 29894 19698 29946
rect 19722 29894 19768 29946
rect 19768 29894 19778 29946
rect 19802 29894 19832 29946
rect 19832 29894 19858 29946
rect 19562 29892 19618 29894
rect 19642 29892 19698 29894
rect 19722 29892 19778 29894
rect 19802 29892 19858 29894
rect 19562 28858 19618 28860
rect 19642 28858 19698 28860
rect 19722 28858 19778 28860
rect 19802 28858 19858 28860
rect 19562 28806 19588 28858
rect 19588 28806 19618 28858
rect 19642 28806 19652 28858
rect 19652 28806 19698 28858
rect 19722 28806 19768 28858
rect 19768 28806 19778 28858
rect 19802 28806 19832 28858
rect 19832 28806 19858 28858
rect 19562 28804 19618 28806
rect 19642 28804 19698 28806
rect 19722 28804 19778 28806
rect 19802 28804 19858 28806
rect 19562 27770 19618 27772
rect 19642 27770 19698 27772
rect 19722 27770 19778 27772
rect 19802 27770 19858 27772
rect 19562 27718 19588 27770
rect 19588 27718 19618 27770
rect 19642 27718 19652 27770
rect 19652 27718 19698 27770
rect 19722 27718 19768 27770
rect 19768 27718 19778 27770
rect 19802 27718 19832 27770
rect 19832 27718 19858 27770
rect 19562 27716 19618 27718
rect 19642 27716 19698 27718
rect 19722 27716 19778 27718
rect 19802 27716 19858 27718
rect 19562 26682 19618 26684
rect 19642 26682 19698 26684
rect 19722 26682 19778 26684
rect 19802 26682 19858 26684
rect 19562 26630 19588 26682
rect 19588 26630 19618 26682
rect 19642 26630 19652 26682
rect 19652 26630 19698 26682
rect 19722 26630 19768 26682
rect 19768 26630 19778 26682
rect 19802 26630 19832 26682
rect 19832 26630 19858 26682
rect 19562 26628 19618 26630
rect 19642 26628 19698 26630
rect 19722 26628 19778 26630
rect 19802 26628 19858 26630
rect 19562 25594 19618 25596
rect 19642 25594 19698 25596
rect 19722 25594 19778 25596
rect 19802 25594 19858 25596
rect 19562 25542 19588 25594
rect 19588 25542 19618 25594
rect 19642 25542 19652 25594
rect 19652 25542 19698 25594
rect 19722 25542 19768 25594
rect 19768 25542 19778 25594
rect 19802 25542 19832 25594
rect 19832 25542 19858 25594
rect 19562 25540 19618 25542
rect 19642 25540 19698 25542
rect 19722 25540 19778 25542
rect 19802 25540 19858 25542
rect 19562 24506 19618 24508
rect 19642 24506 19698 24508
rect 19722 24506 19778 24508
rect 19802 24506 19858 24508
rect 19562 24454 19588 24506
rect 19588 24454 19618 24506
rect 19642 24454 19652 24506
rect 19652 24454 19698 24506
rect 19722 24454 19768 24506
rect 19768 24454 19778 24506
rect 19802 24454 19832 24506
rect 19832 24454 19858 24506
rect 19562 24452 19618 24454
rect 19642 24452 19698 24454
rect 19722 24452 19778 24454
rect 19802 24452 19858 24454
rect 19562 23418 19618 23420
rect 19642 23418 19698 23420
rect 19722 23418 19778 23420
rect 19802 23418 19858 23420
rect 19562 23366 19588 23418
rect 19588 23366 19618 23418
rect 19642 23366 19652 23418
rect 19652 23366 19698 23418
rect 19722 23366 19768 23418
rect 19768 23366 19778 23418
rect 19802 23366 19832 23418
rect 19832 23366 19858 23418
rect 19562 23364 19618 23366
rect 19642 23364 19698 23366
rect 19722 23364 19778 23366
rect 19802 23364 19858 23366
rect 19562 22330 19618 22332
rect 19642 22330 19698 22332
rect 19722 22330 19778 22332
rect 19802 22330 19858 22332
rect 19562 22278 19588 22330
rect 19588 22278 19618 22330
rect 19642 22278 19652 22330
rect 19652 22278 19698 22330
rect 19722 22278 19768 22330
rect 19768 22278 19778 22330
rect 19802 22278 19832 22330
rect 19832 22278 19858 22330
rect 19562 22276 19618 22278
rect 19642 22276 19698 22278
rect 19722 22276 19778 22278
rect 19802 22276 19858 22278
rect 19562 21242 19618 21244
rect 19642 21242 19698 21244
rect 19722 21242 19778 21244
rect 19802 21242 19858 21244
rect 19562 21190 19588 21242
rect 19588 21190 19618 21242
rect 19642 21190 19652 21242
rect 19652 21190 19698 21242
rect 19722 21190 19768 21242
rect 19768 21190 19778 21242
rect 19802 21190 19832 21242
rect 19832 21190 19858 21242
rect 19562 21188 19618 21190
rect 19642 21188 19698 21190
rect 19722 21188 19778 21190
rect 19802 21188 19858 21190
rect 19562 20154 19618 20156
rect 19642 20154 19698 20156
rect 19722 20154 19778 20156
rect 19802 20154 19858 20156
rect 19562 20102 19588 20154
rect 19588 20102 19618 20154
rect 19642 20102 19652 20154
rect 19652 20102 19698 20154
rect 19722 20102 19768 20154
rect 19768 20102 19778 20154
rect 19802 20102 19832 20154
rect 19832 20102 19858 20154
rect 19562 20100 19618 20102
rect 19642 20100 19698 20102
rect 19722 20100 19778 20102
rect 19802 20100 19858 20102
rect 19562 19066 19618 19068
rect 19642 19066 19698 19068
rect 19722 19066 19778 19068
rect 19802 19066 19858 19068
rect 19562 19014 19588 19066
rect 19588 19014 19618 19066
rect 19642 19014 19652 19066
rect 19652 19014 19698 19066
rect 19722 19014 19768 19066
rect 19768 19014 19778 19066
rect 19802 19014 19832 19066
rect 19832 19014 19858 19066
rect 19562 19012 19618 19014
rect 19642 19012 19698 19014
rect 19722 19012 19778 19014
rect 19802 19012 19858 19014
rect 19562 17978 19618 17980
rect 19642 17978 19698 17980
rect 19722 17978 19778 17980
rect 19802 17978 19858 17980
rect 19562 17926 19588 17978
rect 19588 17926 19618 17978
rect 19642 17926 19652 17978
rect 19652 17926 19698 17978
rect 19722 17926 19768 17978
rect 19768 17926 19778 17978
rect 19802 17926 19832 17978
rect 19832 17926 19858 17978
rect 19562 17924 19618 17926
rect 19642 17924 19698 17926
rect 19722 17924 19778 17926
rect 19802 17924 19858 17926
rect 19562 16890 19618 16892
rect 19642 16890 19698 16892
rect 19722 16890 19778 16892
rect 19802 16890 19858 16892
rect 19562 16838 19588 16890
rect 19588 16838 19618 16890
rect 19642 16838 19652 16890
rect 19652 16838 19698 16890
rect 19722 16838 19768 16890
rect 19768 16838 19778 16890
rect 19802 16838 19832 16890
rect 19832 16838 19858 16890
rect 19562 16836 19618 16838
rect 19642 16836 19698 16838
rect 19722 16836 19778 16838
rect 19802 16836 19858 16838
rect 19562 15802 19618 15804
rect 19642 15802 19698 15804
rect 19722 15802 19778 15804
rect 19802 15802 19858 15804
rect 19562 15750 19588 15802
rect 19588 15750 19618 15802
rect 19642 15750 19652 15802
rect 19652 15750 19698 15802
rect 19722 15750 19768 15802
rect 19768 15750 19778 15802
rect 19802 15750 19832 15802
rect 19832 15750 19858 15802
rect 19562 15748 19618 15750
rect 19642 15748 19698 15750
rect 19722 15748 19778 15750
rect 19802 15748 19858 15750
rect 19562 14714 19618 14716
rect 19642 14714 19698 14716
rect 19722 14714 19778 14716
rect 19802 14714 19858 14716
rect 19562 14662 19588 14714
rect 19588 14662 19618 14714
rect 19642 14662 19652 14714
rect 19652 14662 19698 14714
rect 19722 14662 19768 14714
rect 19768 14662 19778 14714
rect 19802 14662 19832 14714
rect 19832 14662 19858 14714
rect 19562 14660 19618 14662
rect 19642 14660 19698 14662
rect 19722 14660 19778 14662
rect 19802 14660 19858 14662
rect 19562 13626 19618 13628
rect 19642 13626 19698 13628
rect 19722 13626 19778 13628
rect 19802 13626 19858 13628
rect 19562 13574 19588 13626
rect 19588 13574 19618 13626
rect 19642 13574 19652 13626
rect 19652 13574 19698 13626
rect 19722 13574 19768 13626
rect 19768 13574 19778 13626
rect 19802 13574 19832 13626
rect 19832 13574 19858 13626
rect 19562 13572 19618 13574
rect 19642 13572 19698 13574
rect 19722 13572 19778 13574
rect 19802 13572 19858 13574
rect 19562 12538 19618 12540
rect 19642 12538 19698 12540
rect 19722 12538 19778 12540
rect 19802 12538 19858 12540
rect 19562 12486 19588 12538
rect 19588 12486 19618 12538
rect 19642 12486 19652 12538
rect 19652 12486 19698 12538
rect 19722 12486 19768 12538
rect 19768 12486 19778 12538
rect 19802 12486 19832 12538
rect 19832 12486 19858 12538
rect 19562 12484 19618 12486
rect 19642 12484 19698 12486
rect 19722 12484 19778 12486
rect 19802 12484 19858 12486
rect 19562 11450 19618 11452
rect 19642 11450 19698 11452
rect 19722 11450 19778 11452
rect 19802 11450 19858 11452
rect 19562 11398 19588 11450
rect 19588 11398 19618 11450
rect 19642 11398 19652 11450
rect 19652 11398 19698 11450
rect 19722 11398 19768 11450
rect 19768 11398 19778 11450
rect 19802 11398 19832 11450
rect 19832 11398 19858 11450
rect 19562 11396 19618 11398
rect 19642 11396 19698 11398
rect 19722 11396 19778 11398
rect 19802 11396 19858 11398
rect 19562 10362 19618 10364
rect 19642 10362 19698 10364
rect 19722 10362 19778 10364
rect 19802 10362 19858 10364
rect 19562 10310 19588 10362
rect 19588 10310 19618 10362
rect 19642 10310 19652 10362
rect 19652 10310 19698 10362
rect 19722 10310 19768 10362
rect 19768 10310 19778 10362
rect 19802 10310 19832 10362
rect 19832 10310 19858 10362
rect 19562 10308 19618 10310
rect 19642 10308 19698 10310
rect 19722 10308 19778 10310
rect 19802 10308 19858 10310
rect 19562 9274 19618 9276
rect 19642 9274 19698 9276
rect 19722 9274 19778 9276
rect 19802 9274 19858 9276
rect 19562 9222 19588 9274
rect 19588 9222 19618 9274
rect 19642 9222 19652 9274
rect 19652 9222 19698 9274
rect 19722 9222 19768 9274
rect 19768 9222 19778 9274
rect 19802 9222 19832 9274
rect 19832 9222 19858 9274
rect 19562 9220 19618 9222
rect 19642 9220 19698 9222
rect 19722 9220 19778 9222
rect 19802 9220 19858 9222
rect 19562 8186 19618 8188
rect 19642 8186 19698 8188
rect 19722 8186 19778 8188
rect 19802 8186 19858 8188
rect 19562 8134 19588 8186
rect 19588 8134 19618 8186
rect 19642 8134 19652 8186
rect 19652 8134 19698 8186
rect 19722 8134 19768 8186
rect 19768 8134 19778 8186
rect 19802 8134 19832 8186
rect 19832 8134 19858 8186
rect 19562 8132 19618 8134
rect 19642 8132 19698 8134
rect 19722 8132 19778 8134
rect 19802 8132 19858 8134
rect 19562 7098 19618 7100
rect 19642 7098 19698 7100
rect 19722 7098 19778 7100
rect 19802 7098 19858 7100
rect 19562 7046 19588 7098
rect 19588 7046 19618 7098
rect 19642 7046 19652 7098
rect 19652 7046 19698 7098
rect 19722 7046 19768 7098
rect 19768 7046 19778 7098
rect 19802 7046 19832 7098
rect 19832 7046 19858 7098
rect 19562 7044 19618 7046
rect 19642 7044 19698 7046
rect 19722 7044 19778 7046
rect 19802 7044 19858 7046
rect 19562 6010 19618 6012
rect 19642 6010 19698 6012
rect 19722 6010 19778 6012
rect 19802 6010 19858 6012
rect 19562 5958 19588 6010
rect 19588 5958 19618 6010
rect 19642 5958 19652 6010
rect 19652 5958 19698 6010
rect 19722 5958 19768 6010
rect 19768 5958 19778 6010
rect 19802 5958 19832 6010
rect 19832 5958 19858 6010
rect 19562 5956 19618 5958
rect 19642 5956 19698 5958
rect 19722 5956 19778 5958
rect 19802 5956 19858 5958
rect 19562 4922 19618 4924
rect 19642 4922 19698 4924
rect 19722 4922 19778 4924
rect 19802 4922 19858 4924
rect 19562 4870 19588 4922
rect 19588 4870 19618 4922
rect 19642 4870 19652 4922
rect 19652 4870 19698 4922
rect 19722 4870 19768 4922
rect 19768 4870 19778 4922
rect 19802 4870 19832 4922
rect 19832 4870 19858 4922
rect 19562 4868 19618 4870
rect 19642 4868 19698 4870
rect 19722 4868 19778 4870
rect 19802 4868 19858 4870
rect 19562 3834 19618 3836
rect 19642 3834 19698 3836
rect 19722 3834 19778 3836
rect 19802 3834 19858 3836
rect 19562 3782 19588 3834
rect 19588 3782 19618 3834
rect 19642 3782 19652 3834
rect 19652 3782 19698 3834
rect 19722 3782 19768 3834
rect 19768 3782 19778 3834
rect 19802 3782 19832 3834
rect 19832 3782 19858 3834
rect 19562 3780 19618 3782
rect 19642 3780 19698 3782
rect 19722 3780 19778 3782
rect 19802 3780 19858 3782
rect 19562 2746 19618 2748
rect 19642 2746 19698 2748
rect 19722 2746 19778 2748
rect 19802 2746 19858 2748
rect 19562 2694 19588 2746
rect 19588 2694 19618 2746
rect 19642 2694 19652 2746
rect 19652 2694 19698 2746
rect 19722 2694 19768 2746
rect 19768 2694 19778 2746
rect 19802 2694 19832 2746
rect 19832 2694 19858 2746
rect 19562 2692 19618 2694
rect 19642 2692 19698 2694
rect 19722 2692 19778 2694
rect 19802 2692 19858 2694
rect 25484 56208 25540 56264
rect 25852 17992 25908 18048
rect 25852 17856 25908 17912
rect 27784 37204 27786 37224
rect 27786 37204 27838 37224
rect 27838 37204 27840 37224
rect 27784 37168 27840 37204
rect 31648 56208 31704 56264
rect 32568 56072 32624 56128
rect 31280 55936 31336 55992
rect 31832 55936 31888 55992
rect 32476 55936 32532 55992
rect 33856 56208 33912 56264
rect 34922 57690 34978 57692
rect 35002 57690 35058 57692
rect 35082 57690 35138 57692
rect 35162 57690 35218 57692
rect 34922 57638 34948 57690
rect 34948 57638 34978 57690
rect 35002 57638 35012 57690
rect 35012 57638 35058 57690
rect 35082 57638 35128 57690
rect 35128 57638 35138 57690
rect 35162 57638 35192 57690
rect 35192 57638 35218 57690
rect 34922 57636 34978 57638
rect 35002 57636 35058 57638
rect 35082 57636 35138 57638
rect 35162 57636 35218 57638
rect 34922 56602 34978 56604
rect 35002 56602 35058 56604
rect 35082 56602 35138 56604
rect 35162 56602 35218 56604
rect 34922 56550 34948 56602
rect 34948 56550 34978 56602
rect 35002 56550 35012 56602
rect 35012 56550 35058 56602
rect 35082 56550 35128 56602
rect 35128 56550 35138 56602
rect 35162 56550 35192 56602
rect 35192 56550 35218 56602
rect 34922 56548 34978 56550
rect 35002 56548 35058 56550
rect 35082 56548 35138 56550
rect 35162 56548 35218 56550
rect 34922 55514 34978 55516
rect 35002 55514 35058 55516
rect 35082 55514 35138 55516
rect 35162 55514 35218 55516
rect 34922 55462 34948 55514
rect 34948 55462 34978 55514
rect 35002 55462 35012 55514
rect 35012 55462 35058 55514
rect 35082 55462 35128 55514
rect 35128 55462 35138 55514
rect 35162 55462 35192 55514
rect 35192 55462 35218 55514
rect 34922 55460 34978 55462
rect 35002 55460 35058 55462
rect 35082 55460 35138 55462
rect 35162 55460 35218 55462
rect 35972 56244 35974 56264
rect 35974 56244 36026 56264
rect 36026 56244 36028 56264
rect 35972 56208 36028 56244
rect 34922 54426 34978 54428
rect 35002 54426 35058 54428
rect 35082 54426 35138 54428
rect 35162 54426 35218 54428
rect 34922 54374 34948 54426
rect 34948 54374 34978 54426
rect 35002 54374 35012 54426
rect 35012 54374 35058 54426
rect 35082 54374 35128 54426
rect 35128 54374 35138 54426
rect 35162 54374 35192 54426
rect 35192 54374 35218 54426
rect 34922 54372 34978 54374
rect 35002 54372 35058 54374
rect 35082 54372 35138 54374
rect 35162 54372 35218 54374
rect 34922 53338 34978 53340
rect 35002 53338 35058 53340
rect 35082 53338 35138 53340
rect 35162 53338 35218 53340
rect 34922 53286 34948 53338
rect 34948 53286 34978 53338
rect 35002 53286 35012 53338
rect 35012 53286 35058 53338
rect 35082 53286 35128 53338
rect 35128 53286 35138 53338
rect 35162 53286 35192 53338
rect 35192 53286 35218 53338
rect 34922 53284 34978 53286
rect 35002 53284 35058 53286
rect 35082 53284 35138 53286
rect 35162 53284 35218 53286
rect 34922 52250 34978 52252
rect 35002 52250 35058 52252
rect 35082 52250 35138 52252
rect 35162 52250 35218 52252
rect 34922 52198 34948 52250
rect 34948 52198 34978 52250
rect 35002 52198 35012 52250
rect 35012 52198 35058 52250
rect 35082 52198 35128 52250
rect 35128 52198 35138 52250
rect 35162 52198 35192 52250
rect 35192 52198 35218 52250
rect 34922 52196 34978 52198
rect 35002 52196 35058 52198
rect 35082 52196 35138 52198
rect 35162 52196 35218 52198
rect 34922 51162 34978 51164
rect 35002 51162 35058 51164
rect 35082 51162 35138 51164
rect 35162 51162 35218 51164
rect 34922 51110 34948 51162
rect 34948 51110 34978 51162
rect 35002 51110 35012 51162
rect 35012 51110 35058 51162
rect 35082 51110 35128 51162
rect 35128 51110 35138 51162
rect 35162 51110 35192 51162
rect 35192 51110 35218 51162
rect 34922 51108 34978 51110
rect 35002 51108 35058 51110
rect 35082 51108 35138 51110
rect 35162 51108 35218 51110
rect 34922 50074 34978 50076
rect 35002 50074 35058 50076
rect 35082 50074 35138 50076
rect 35162 50074 35218 50076
rect 34922 50022 34948 50074
rect 34948 50022 34978 50074
rect 35002 50022 35012 50074
rect 35012 50022 35058 50074
rect 35082 50022 35128 50074
rect 35128 50022 35138 50074
rect 35162 50022 35192 50074
rect 35192 50022 35218 50074
rect 34922 50020 34978 50022
rect 35002 50020 35058 50022
rect 35082 50020 35138 50022
rect 35162 50020 35218 50022
rect 34922 48986 34978 48988
rect 35002 48986 35058 48988
rect 35082 48986 35138 48988
rect 35162 48986 35218 48988
rect 34922 48934 34948 48986
rect 34948 48934 34978 48986
rect 35002 48934 35012 48986
rect 35012 48934 35058 48986
rect 35082 48934 35128 48986
rect 35128 48934 35138 48986
rect 35162 48934 35192 48986
rect 35192 48934 35218 48986
rect 34922 48932 34978 48934
rect 35002 48932 35058 48934
rect 35082 48932 35138 48934
rect 35162 48932 35218 48934
rect 34922 47898 34978 47900
rect 35002 47898 35058 47900
rect 35082 47898 35138 47900
rect 35162 47898 35218 47900
rect 34922 47846 34948 47898
rect 34948 47846 34978 47898
rect 35002 47846 35012 47898
rect 35012 47846 35058 47898
rect 35082 47846 35128 47898
rect 35128 47846 35138 47898
rect 35162 47846 35192 47898
rect 35192 47846 35218 47898
rect 34922 47844 34978 47846
rect 35002 47844 35058 47846
rect 35082 47844 35138 47846
rect 35162 47844 35218 47846
rect 34922 46810 34978 46812
rect 35002 46810 35058 46812
rect 35082 46810 35138 46812
rect 35162 46810 35218 46812
rect 34922 46758 34948 46810
rect 34948 46758 34978 46810
rect 35002 46758 35012 46810
rect 35012 46758 35058 46810
rect 35082 46758 35128 46810
rect 35128 46758 35138 46810
rect 35162 46758 35192 46810
rect 35192 46758 35218 46810
rect 34922 46756 34978 46758
rect 35002 46756 35058 46758
rect 35082 46756 35138 46758
rect 35162 46756 35218 46758
rect 34922 45722 34978 45724
rect 35002 45722 35058 45724
rect 35082 45722 35138 45724
rect 35162 45722 35218 45724
rect 34922 45670 34948 45722
rect 34948 45670 34978 45722
rect 35002 45670 35012 45722
rect 35012 45670 35058 45722
rect 35082 45670 35128 45722
rect 35128 45670 35138 45722
rect 35162 45670 35192 45722
rect 35192 45670 35218 45722
rect 34922 45668 34978 45670
rect 35002 45668 35058 45670
rect 35082 45668 35138 45670
rect 35162 45668 35218 45670
rect 34922 44634 34978 44636
rect 35002 44634 35058 44636
rect 35082 44634 35138 44636
rect 35162 44634 35218 44636
rect 34922 44582 34948 44634
rect 34948 44582 34978 44634
rect 35002 44582 35012 44634
rect 35012 44582 35058 44634
rect 35082 44582 35128 44634
rect 35128 44582 35138 44634
rect 35162 44582 35192 44634
rect 35192 44582 35218 44634
rect 34922 44580 34978 44582
rect 35002 44580 35058 44582
rect 35082 44580 35138 44582
rect 35162 44580 35218 44582
rect 34922 43546 34978 43548
rect 35002 43546 35058 43548
rect 35082 43546 35138 43548
rect 35162 43546 35218 43548
rect 34922 43494 34948 43546
rect 34948 43494 34978 43546
rect 35002 43494 35012 43546
rect 35012 43494 35058 43546
rect 35082 43494 35128 43546
rect 35128 43494 35138 43546
rect 35162 43494 35192 43546
rect 35192 43494 35218 43546
rect 34922 43492 34978 43494
rect 35002 43492 35058 43494
rect 35082 43492 35138 43494
rect 35162 43492 35218 43494
rect 34922 42458 34978 42460
rect 35002 42458 35058 42460
rect 35082 42458 35138 42460
rect 35162 42458 35218 42460
rect 34922 42406 34948 42458
rect 34948 42406 34978 42458
rect 35002 42406 35012 42458
rect 35012 42406 35058 42458
rect 35082 42406 35128 42458
rect 35128 42406 35138 42458
rect 35162 42406 35192 42458
rect 35192 42406 35218 42458
rect 34922 42404 34978 42406
rect 35002 42404 35058 42406
rect 35082 42404 35138 42406
rect 35162 42404 35218 42406
rect 34922 41370 34978 41372
rect 35002 41370 35058 41372
rect 35082 41370 35138 41372
rect 35162 41370 35218 41372
rect 34922 41318 34948 41370
rect 34948 41318 34978 41370
rect 35002 41318 35012 41370
rect 35012 41318 35058 41370
rect 35082 41318 35128 41370
rect 35128 41318 35138 41370
rect 35162 41318 35192 41370
rect 35192 41318 35218 41370
rect 34922 41316 34978 41318
rect 35002 41316 35058 41318
rect 35082 41316 35138 41318
rect 35162 41316 35218 41318
rect 34922 40282 34978 40284
rect 35002 40282 35058 40284
rect 35082 40282 35138 40284
rect 35162 40282 35218 40284
rect 34922 40230 34948 40282
rect 34948 40230 34978 40282
rect 35002 40230 35012 40282
rect 35012 40230 35058 40282
rect 35082 40230 35128 40282
rect 35128 40230 35138 40282
rect 35162 40230 35192 40282
rect 35192 40230 35218 40282
rect 34922 40228 34978 40230
rect 35002 40228 35058 40230
rect 35082 40228 35138 40230
rect 35162 40228 35218 40230
rect 34922 39194 34978 39196
rect 35002 39194 35058 39196
rect 35082 39194 35138 39196
rect 35162 39194 35218 39196
rect 34922 39142 34948 39194
rect 34948 39142 34978 39194
rect 35002 39142 35012 39194
rect 35012 39142 35058 39194
rect 35082 39142 35128 39194
rect 35128 39142 35138 39194
rect 35162 39142 35192 39194
rect 35192 39142 35218 39194
rect 34922 39140 34978 39142
rect 35002 39140 35058 39142
rect 35082 39140 35138 39142
rect 35162 39140 35218 39142
rect 34922 38106 34978 38108
rect 35002 38106 35058 38108
rect 35082 38106 35138 38108
rect 35162 38106 35218 38108
rect 34922 38054 34948 38106
rect 34948 38054 34978 38106
rect 35002 38054 35012 38106
rect 35012 38054 35058 38106
rect 35082 38054 35128 38106
rect 35128 38054 35138 38106
rect 35162 38054 35192 38106
rect 35192 38054 35218 38106
rect 34922 38052 34978 38054
rect 35002 38052 35058 38054
rect 35082 38052 35138 38054
rect 35162 38052 35218 38054
rect 34922 37018 34978 37020
rect 35002 37018 35058 37020
rect 35082 37018 35138 37020
rect 35162 37018 35218 37020
rect 34922 36966 34948 37018
rect 34948 36966 34978 37018
rect 35002 36966 35012 37018
rect 35012 36966 35058 37018
rect 35082 36966 35128 37018
rect 35128 36966 35138 37018
rect 35162 36966 35192 37018
rect 35192 36966 35218 37018
rect 34922 36964 34978 36966
rect 35002 36964 35058 36966
rect 35082 36964 35138 36966
rect 35162 36964 35218 36966
rect 34316 36080 34372 36136
rect 34500 35944 34556 36000
rect 34922 35930 34978 35932
rect 35002 35930 35058 35932
rect 35082 35930 35138 35932
rect 35162 35930 35218 35932
rect 34922 35878 34948 35930
rect 34948 35878 34978 35930
rect 35002 35878 35012 35930
rect 35012 35878 35058 35930
rect 35082 35878 35128 35930
rect 35128 35878 35138 35930
rect 35162 35878 35192 35930
rect 35192 35878 35218 35930
rect 34922 35876 34978 35878
rect 35002 35876 35058 35878
rect 35082 35876 35138 35878
rect 35162 35876 35218 35878
rect 34922 34842 34978 34844
rect 35002 34842 35058 34844
rect 35082 34842 35138 34844
rect 35162 34842 35218 34844
rect 34922 34790 34948 34842
rect 34948 34790 34978 34842
rect 35002 34790 35012 34842
rect 35012 34790 35058 34842
rect 35082 34790 35128 34842
rect 35128 34790 35138 34842
rect 35162 34790 35192 34842
rect 35192 34790 35218 34842
rect 34922 34788 34978 34790
rect 35002 34788 35058 34790
rect 35082 34788 35138 34790
rect 35162 34788 35218 34790
rect 34922 33754 34978 33756
rect 35002 33754 35058 33756
rect 35082 33754 35138 33756
rect 35162 33754 35218 33756
rect 34922 33702 34948 33754
rect 34948 33702 34978 33754
rect 35002 33702 35012 33754
rect 35012 33702 35058 33754
rect 35082 33702 35128 33754
rect 35128 33702 35138 33754
rect 35162 33702 35192 33754
rect 35192 33702 35218 33754
rect 34922 33700 34978 33702
rect 35002 33700 35058 33702
rect 35082 33700 35138 33702
rect 35162 33700 35218 33702
rect 34922 32666 34978 32668
rect 35002 32666 35058 32668
rect 35082 32666 35138 32668
rect 35162 32666 35218 32668
rect 34922 32614 34948 32666
rect 34948 32614 34978 32666
rect 35002 32614 35012 32666
rect 35012 32614 35058 32666
rect 35082 32614 35128 32666
rect 35128 32614 35138 32666
rect 35162 32614 35192 32666
rect 35192 32614 35218 32666
rect 34922 32612 34978 32614
rect 35002 32612 35058 32614
rect 35082 32612 35138 32614
rect 35162 32612 35218 32614
rect 34922 31578 34978 31580
rect 35002 31578 35058 31580
rect 35082 31578 35138 31580
rect 35162 31578 35218 31580
rect 34922 31526 34948 31578
rect 34948 31526 34978 31578
rect 35002 31526 35012 31578
rect 35012 31526 35058 31578
rect 35082 31526 35128 31578
rect 35128 31526 35138 31578
rect 35162 31526 35192 31578
rect 35192 31526 35218 31578
rect 34922 31524 34978 31526
rect 35002 31524 35058 31526
rect 35082 31524 35138 31526
rect 35162 31524 35218 31526
rect 34922 30490 34978 30492
rect 35002 30490 35058 30492
rect 35082 30490 35138 30492
rect 35162 30490 35218 30492
rect 34922 30438 34948 30490
rect 34948 30438 34978 30490
rect 35002 30438 35012 30490
rect 35012 30438 35058 30490
rect 35082 30438 35128 30490
rect 35128 30438 35138 30490
rect 35162 30438 35192 30490
rect 35192 30438 35218 30490
rect 34922 30436 34978 30438
rect 35002 30436 35058 30438
rect 35082 30436 35138 30438
rect 35162 30436 35218 30438
rect 34922 29402 34978 29404
rect 35002 29402 35058 29404
rect 35082 29402 35138 29404
rect 35162 29402 35218 29404
rect 34922 29350 34948 29402
rect 34948 29350 34978 29402
rect 35002 29350 35012 29402
rect 35012 29350 35058 29402
rect 35082 29350 35128 29402
rect 35128 29350 35138 29402
rect 35162 29350 35192 29402
rect 35192 29350 35218 29402
rect 34922 29348 34978 29350
rect 35002 29348 35058 29350
rect 35082 29348 35138 29350
rect 35162 29348 35218 29350
rect 34922 28314 34978 28316
rect 35002 28314 35058 28316
rect 35082 28314 35138 28316
rect 35162 28314 35218 28316
rect 34922 28262 34948 28314
rect 34948 28262 34978 28314
rect 35002 28262 35012 28314
rect 35012 28262 35058 28314
rect 35082 28262 35128 28314
rect 35128 28262 35138 28314
rect 35162 28262 35192 28314
rect 35192 28262 35218 28314
rect 34922 28260 34978 28262
rect 35002 28260 35058 28262
rect 35082 28260 35138 28262
rect 35162 28260 35218 28262
rect 34922 27226 34978 27228
rect 35002 27226 35058 27228
rect 35082 27226 35138 27228
rect 35162 27226 35218 27228
rect 34922 27174 34948 27226
rect 34948 27174 34978 27226
rect 35002 27174 35012 27226
rect 35012 27174 35058 27226
rect 35082 27174 35128 27226
rect 35128 27174 35138 27226
rect 35162 27174 35192 27226
rect 35192 27174 35218 27226
rect 34922 27172 34978 27174
rect 35002 27172 35058 27174
rect 35082 27172 35138 27174
rect 35162 27172 35218 27174
rect 34922 26138 34978 26140
rect 35002 26138 35058 26140
rect 35082 26138 35138 26140
rect 35162 26138 35218 26140
rect 34922 26086 34948 26138
rect 34948 26086 34978 26138
rect 35002 26086 35012 26138
rect 35012 26086 35058 26138
rect 35082 26086 35128 26138
rect 35128 26086 35138 26138
rect 35162 26086 35192 26138
rect 35192 26086 35218 26138
rect 34922 26084 34978 26086
rect 35002 26084 35058 26086
rect 35082 26084 35138 26086
rect 35162 26084 35218 26086
rect 34922 25050 34978 25052
rect 35002 25050 35058 25052
rect 35082 25050 35138 25052
rect 35162 25050 35218 25052
rect 34922 24998 34948 25050
rect 34948 24998 34978 25050
rect 35002 24998 35012 25050
rect 35012 24998 35058 25050
rect 35082 24998 35128 25050
rect 35128 24998 35138 25050
rect 35162 24998 35192 25050
rect 35192 24998 35218 25050
rect 34922 24996 34978 24998
rect 35002 24996 35058 24998
rect 35082 24996 35138 24998
rect 35162 24996 35218 24998
rect 34922 23962 34978 23964
rect 35002 23962 35058 23964
rect 35082 23962 35138 23964
rect 35162 23962 35218 23964
rect 34922 23910 34948 23962
rect 34948 23910 34978 23962
rect 35002 23910 35012 23962
rect 35012 23910 35058 23962
rect 35082 23910 35128 23962
rect 35128 23910 35138 23962
rect 35162 23910 35192 23962
rect 35192 23910 35218 23962
rect 34922 23908 34978 23910
rect 35002 23908 35058 23910
rect 35082 23908 35138 23910
rect 35162 23908 35218 23910
rect 34922 22874 34978 22876
rect 35002 22874 35058 22876
rect 35082 22874 35138 22876
rect 35162 22874 35218 22876
rect 34922 22822 34948 22874
rect 34948 22822 34978 22874
rect 35002 22822 35012 22874
rect 35012 22822 35058 22874
rect 35082 22822 35128 22874
rect 35128 22822 35138 22874
rect 35162 22822 35192 22874
rect 35192 22822 35218 22874
rect 34922 22820 34978 22822
rect 35002 22820 35058 22822
rect 35082 22820 35138 22822
rect 35162 22820 35218 22822
rect 34922 21786 34978 21788
rect 35002 21786 35058 21788
rect 35082 21786 35138 21788
rect 35162 21786 35218 21788
rect 34922 21734 34948 21786
rect 34948 21734 34978 21786
rect 35002 21734 35012 21786
rect 35012 21734 35058 21786
rect 35082 21734 35128 21786
rect 35128 21734 35138 21786
rect 35162 21734 35192 21786
rect 35192 21734 35218 21786
rect 34922 21732 34978 21734
rect 35002 21732 35058 21734
rect 35082 21732 35138 21734
rect 35162 21732 35218 21734
rect 34922 20698 34978 20700
rect 35002 20698 35058 20700
rect 35082 20698 35138 20700
rect 35162 20698 35218 20700
rect 34922 20646 34948 20698
rect 34948 20646 34978 20698
rect 35002 20646 35012 20698
rect 35012 20646 35058 20698
rect 35082 20646 35128 20698
rect 35128 20646 35138 20698
rect 35162 20646 35192 20698
rect 35192 20646 35218 20698
rect 34922 20644 34978 20646
rect 35002 20644 35058 20646
rect 35082 20644 35138 20646
rect 35162 20644 35218 20646
rect 34922 19610 34978 19612
rect 35002 19610 35058 19612
rect 35082 19610 35138 19612
rect 35162 19610 35218 19612
rect 34922 19558 34948 19610
rect 34948 19558 34978 19610
rect 35002 19558 35012 19610
rect 35012 19558 35058 19610
rect 35082 19558 35128 19610
rect 35128 19558 35138 19610
rect 35162 19558 35192 19610
rect 35192 19558 35218 19610
rect 34922 19556 34978 19558
rect 35002 19556 35058 19558
rect 35082 19556 35138 19558
rect 35162 19556 35218 19558
rect 34922 18522 34978 18524
rect 35002 18522 35058 18524
rect 35082 18522 35138 18524
rect 35162 18522 35218 18524
rect 34922 18470 34948 18522
rect 34948 18470 34978 18522
rect 35002 18470 35012 18522
rect 35012 18470 35058 18522
rect 35082 18470 35128 18522
rect 35128 18470 35138 18522
rect 35162 18470 35192 18522
rect 35192 18470 35218 18522
rect 34922 18468 34978 18470
rect 35002 18468 35058 18470
rect 35082 18468 35138 18470
rect 35162 18468 35218 18470
rect 34922 17434 34978 17436
rect 35002 17434 35058 17436
rect 35082 17434 35138 17436
rect 35162 17434 35218 17436
rect 34922 17382 34948 17434
rect 34948 17382 34978 17434
rect 35002 17382 35012 17434
rect 35012 17382 35058 17434
rect 35082 17382 35128 17434
rect 35128 17382 35138 17434
rect 35162 17382 35192 17434
rect 35192 17382 35218 17434
rect 34922 17380 34978 17382
rect 35002 17380 35058 17382
rect 35082 17380 35138 17382
rect 35162 17380 35218 17382
rect 34922 16346 34978 16348
rect 35002 16346 35058 16348
rect 35082 16346 35138 16348
rect 35162 16346 35218 16348
rect 34922 16294 34948 16346
rect 34948 16294 34978 16346
rect 35002 16294 35012 16346
rect 35012 16294 35058 16346
rect 35082 16294 35128 16346
rect 35128 16294 35138 16346
rect 35162 16294 35192 16346
rect 35192 16294 35218 16346
rect 34922 16292 34978 16294
rect 35002 16292 35058 16294
rect 35082 16292 35138 16294
rect 35162 16292 35218 16294
rect 34922 15258 34978 15260
rect 35002 15258 35058 15260
rect 35082 15258 35138 15260
rect 35162 15258 35218 15260
rect 34922 15206 34948 15258
rect 34948 15206 34978 15258
rect 35002 15206 35012 15258
rect 35012 15206 35058 15258
rect 35082 15206 35128 15258
rect 35128 15206 35138 15258
rect 35162 15206 35192 15258
rect 35192 15206 35218 15258
rect 34922 15204 34978 15206
rect 35002 15204 35058 15206
rect 35082 15204 35138 15206
rect 35162 15204 35218 15206
rect 34922 14170 34978 14172
rect 35002 14170 35058 14172
rect 35082 14170 35138 14172
rect 35162 14170 35218 14172
rect 34922 14118 34948 14170
rect 34948 14118 34978 14170
rect 35002 14118 35012 14170
rect 35012 14118 35058 14170
rect 35082 14118 35128 14170
rect 35128 14118 35138 14170
rect 35162 14118 35192 14170
rect 35192 14118 35218 14170
rect 34922 14116 34978 14118
rect 35002 14116 35058 14118
rect 35082 14116 35138 14118
rect 35162 14116 35218 14118
rect 34922 13082 34978 13084
rect 35002 13082 35058 13084
rect 35082 13082 35138 13084
rect 35162 13082 35218 13084
rect 34922 13030 34948 13082
rect 34948 13030 34978 13082
rect 35002 13030 35012 13082
rect 35012 13030 35058 13082
rect 35082 13030 35128 13082
rect 35128 13030 35138 13082
rect 35162 13030 35192 13082
rect 35192 13030 35218 13082
rect 34922 13028 34978 13030
rect 35002 13028 35058 13030
rect 35082 13028 35138 13030
rect 35162 13028 35218 13030
rect 34922 11994 34978 11996
rect 35002 11994 35058 11996
rect 35082 11994 35138 11996
rect 35162 11994 35218 11996
rect 34922 11942 34948 11994
rect 34948 11942 34978 11994
rect 35002 11942 35012 11994
rect 35012 11942 35058 11994
rect 35082 11942 35128 11994
rect 35128 11942 35138 11994
rect 35162 11942 35192 11994
rect 35192 11942 35218 11994
rect 34922 11940 34978 11942
rect 35002 11940 35058 11942
rect 35082 11940 35138 11942
rect 35162 11940 35218 11942
rect 34922 10906 34978 10908
rect 35002 10906 35058 10908
rect 35082 10906 35138 10908
rect 35162 10906 35218 10908
rect 34922 10854 34948 10906
rect 34948 10854 34978 10906
rect 35002 10854 35012 10906
rect 35012 10854 35058 10906
rect 35082 10854 35128 10906
rect 35128 10854 35138 10906
rect 35162 10854 35192 10906
rect 35192 10854 35218 10906
rect 34922 10852 34978 10854
rect 35002 10852 35058 10854
rect 35082 10852 35138 10854
rect 35162 10852 35218 10854
rect 34922 9818 34978 9820
rect 35002 9818 35058 9820
rect 35082 9818 35138 9820
rect 35162 9818 35218 9820
rect 34922 9766 34948 9818
rect 34948 9766 34978 9818
rect 35002 9766 35012 9818
rect 35012 9766 35058 9818
rect 35082 9766 35128 9818
rect 35128 9766 35138 9818
rect 35162 9766 35192 9818
rect 35192 9766 35218 9818
rect 34922 9764 34978 9766
rect 35002 9764 35058 9766
rect 35082 9764 35138 9766
rect 35162 9764 35218 9766
rect 34922 8730 34978 8732
rect 35002 8730 35058 8732
rect 35082 8730 35138 8732
rect 35162 8730 35218 8732
rect 34922 8678 34948 8730
rect 34948 8678 34978 8730
rect 35002 8678 35012 8730
rect 35012 8678 35058 8730
rect 35082 8678 35128 8730
rect 35128 8678 35138 8730
rect 35162 8678 35192 8730
rect 35192 8678 35218 8730
rect 34922 8676 34978 8678
rect 35002 8676 35058 8678
rect 35082 8676 35138 8678
rect 35162 8676 35218 8678
rect 34922 7642 34978 7644
rect 35002 7642 35058 7644
rect 35082 7642 35138 7644
rect 35162 7642 35218 7644
rect 34922 7590 34948 7642
rect 34948 7590 34978 7642
rect 35002 7590 35012 7642
rect 35012 7590 35058 7642
rect 35082 7590 35128 7642
rect 35128 7590 35138 7642
rect 35162 7590 35192 7642
rect 35192 7590 35218 7642
rect 34922 7588 34978 7590
rect 35002 7588 35058 7590
rect 35082 7588 35138 7590
rect 35162 7588 35218 7590
rect 34922 6554 34978 6556
rect 35002 6554 35058 6556
rect 35082 6554 35138 6556
rect 35162 6554 35218 6556
rect 34922 6502 34948 6554
rect 34948 6502 34978 6554
rect 35002 6502 35012 6554
rect 35012 6502 35058 6554
rect 35082 6502 35128 6554
rect 35128 6502 35138 6554
rect 35162 6502 35192 6554
rect 35192 6502 35218 6554
rect 34922 6500 34978 6502
rect 35002 6500 35058 6502
rect 35082 6500 35138 6502
rect 35162 6500 35218 6502
rect 34922 5466 34978 5468
rect 35002 5466 35058 5468
rect 35082 5466 35138 5468
rect 35162 5466 35218 5468
rect 34922 5414 34948 5466
rect 34948 5414 34978 5466
rect 35002 5414 35012 5466
rect 35012 5414 35058 5466
rect 35082 5414 35128 5466
rect 35128 5414 35138 5466
rect 35162 5414 35192 5466
rect 35192 5414 35218 5466
rect 34922 5412 34978 5414
rect 35002 5412 35058 5414
rect 35082 5412 35138 5414
rect 35162 5412 35218 5414
rect 34922 4378 34978 4380
rect 35002 4378 35058 4380
rect 35082 4378 35138 4380
rect 35162 4378 35218 4380
rect 34922 4326 34948 4378
rect 34948 4326 34978 4378
rect 35002 4326 35012 4378
rect 35012 4326 35058 4378
rect 35082 4326 35128 4378
rect 35128 4326 35138 4378
rect 35162 4326 35192 4378
rect 35192 4326 35218 4378
rect 34922 4324 34978 4326
rect 35002 4324 35058 4326
rect 35082 4324 35138 4326
rect 35162 4324 35218 4326
rect 34922 3290 34978 3292
rect 35002 3290 35058 3292
rect 35082 3290 35138 3292
rect 35162 3290 35218 3292
rect 34922 3238 34948 3290
rect 34948 3238 34978 3290
rect 35002 3238 35012 3290
rect 35012 3238 35058 3290
rect 35082 3238 35128 3290
rect 35128 3238 35138 3290
rect 35162 3238 35192 3290
rect 35192 3238 35218 3290
rect 34922 3236 34978 3238
rect 35002 3236 35058 3238
rect 35082 3236 35138 3238
rect 35162 3236 35218 3238
rect 34922 2202 34978 2204
rect 35002 2202 35058 2204
rect 35082 2202 35138 2204
rect 35162 2202 35218 2204
rect 34922 2150 34948 2202
rect 34948 2150 34978 2202
rect 35002 2150 35012 2202
rect 35012 2150 35058 2202
rect 35082 2150 35128 2202
rect 35128 2150 35138 2202
rect 35162 2150 35192 2202
rect 35192 2150 35218 2202
rect 34922 2148 34978 2150
rect 35002 2148 35058 2150
rect 35082 2148 35138 2150
rect 35162 2148 35218 2150
rect 38640 56364 38696 56400
rect 38640 56344 38642 56364
rect 38642 56344 38694 56364
rect 38694 56344 38696 56364
rect 36340 2796 36342 2816
rect 36342 2796 36394 2816
rect 36394 2796 36396 2816
rect 36340 2760 36396 2796
rect 36892 856 36948 912
rect 37168 856 37224 912
rect 40940 56072 40996 56128
rect 41216 56072 41272 56128
rect 41400 56108 41402 56128
rect 41402 56108 41454 56128
rect 41454 56108 41456 56128
rect 41400 56072 41456 56108
rect 41492 55936 41548 55992
rect 41400 55700 41402 55720
rect 41402 55700 41454 55720
rect 41454 55700 41456 55720
rect 41400 55664 41456 55700
rect 39836 38800 39892 38856
rect 39652 38664 39708 38720
rect 43884 55664 43940 55720
rect 42596 26288 42652 26344
rect 42872 26288 42928 26344
rect 41308 2896 41364 2952
rect 41492 2932 41494 2952
rect 41494 2932 41546 2952
rect 41546 2932 41548 2952
rect 41492 2896 41548 2932
rect 41308 2760 41364 2816
rect 46184 56380 46186 56400
rect 46186 56380 46238 56400
rect 46238 56380 46240 56400
rect 46184 56344 46240 56380
rect 47012 55800 47068 55856
rect 45908 3712 45964 3768
rect 46920 3712 46976 3768
rect 50282 57146 50338 57148
rect 50362 57146 50418 57148
rect 50442 57146 50498 57148
rect 50522 57146 50578 57148
rect 50282 57094 50308 57146
rect 50308 57094 50338 57146
rect 50362 57094 50372 57146
rect 50372 57094 50418 57146
rect 50442 57094 50488 57146
rect 50488 57094 50498 57146
rect 50522 57094 50552 57146
rect 50552 57094 50578 57146
rect 50282 57092 50338 57094
rect 50362 57092 50418 57094
rect 50442 57092 50498 57094
rect 50522 57092 50578 57094
rect 50282 56058 50338 56060
rect 50362 56058 50418 56060
rect 50442 56058 50498 56060
rect 50522 56058 50578 56060
rect 50282 56006 50308 56058
rect 50308 56006 50338 56058
rect 50362 56006 50372 56058
rect 50372 56006 50418 56058
rect 50442 56006 50488 56058
rect 50488 56006 50498 56058
rect 50522 56006 50552 56058
rect 50552 56006 50578 56058
rect 50282 56004 50338 56006
rect 50362 56004 50418 56006
rect 50442 56004 50498 56006
rect 50522 56004 50578 56006
rect 51244 56616 51300 56672
rect 50282 54970 50338 54972
rect 50362 54970 50418 54972
rect 50442 54970 50498 54972
rect 50522 54970 50578 54972
rect 50282 54918 50308 54970
rect 50308 54918 50338 54970
rect 50362 54918 50372 54970
rect 50372 54918 50418 54970
rect 50442 54918 50488 54970
rect 50488 54918 50498 54970
rect 50522 54918 50552 54970
rect 50552 54918 50578 54970
rect 50282 54916 50338 54918
rect 50362 54916 50418 54918
rect 50442 54916 50498 54918
rect 50522 54916 50578 54918
rect 50282 53882 50338 53884
rect 50362 53882 50418 53884
rect 50442 53882 50498 53884
rect 50522 53882 50578 53884
rect 50282 53830 50308 53882
rect 50308 53830 50338 53882
rect 50362 53830 50372 53882
rect 50372 53830 50418 53882
rect 50442 53830 50488 53882
rect 50488 53830 50498 53882
rect 50522 53830 50552 53882
rect 50552 53830 50578 53882
rect 50282 53828 50338 53830
rect 50362 53828 50418 53830
rect 50442 53828 50498 53830
rect 50522 53828 50578 53830
rect 50282 52794 50338 52796
rect 50362 52794 50418 52796
rect 50442 52794 50498 52796
rect 50522 52794 50578 52796
rect 50282 52742 50308 52794
rect 50308 52742 50338 52794
rect 50362 52742 50372 52794
rect 50372 52742 50418 52794
rect 50442 52742 50488 52794
rect 50488 52742 50498 52794
rect 50522 52742 50552 52794
rect 50552 52742 50578 52794
rect 50282 52740 50338 52742
rect 50362 52740 50418 52742
rect 50442 52740 50498 52742
rect 50522 52740 50578 52742
rect 50282 51706 50338 51708
rect 50362 51706 50418 51708
rect 50442 51706 50498 51708
rect 50522 51706 50578 51708
rect 50282 51654 50308 51706
rect 50308 51654 50338 51706
rect 50362 51654 50372 51706
rect 50372 51654 50418 51706
rect 50442 51654 50488 51706
rect 50488 51654 50498 51706
rect 50522 51654 50552 51706
rect 50552 51654 50578 51706
rect 50282 51652 50338 51654
rect 50362 51652 50418 51654
rect 50442 51652 50498 51654
rect 50522 51652 50578 51654
rect 49496 38664 49552 38720
rect 49588 38528 49644 38584
rect 50282 50618 50338 50620
rect 50362 50618 50418 50620
rect 50442 50618 50498 50620
rect 50522 50618 50578 50620
rect 50282 50566 50308 50618
rect 50308 50566 50338 50618
rect 50362 50566 50372 50618
rect 50372 50566 50418 50618
rect 50442 50566 50488 50618
rect 50488 50566 50498 50618
rect 50522 50566 50552 50618
rect 50552 50566 50578 50618
rect 50282 50564 50338 50566
rect 50362 50564 50418 50566
rect 50442 50564 50498 50566
rect 50522 50564 50578 50566
rect 50282 49530 50338 49532
rect 50362 49530 50418 49532
rect 50442 49530 50498 49532
rect 50522 49530 50578 49532
rect 50282 49478 50308 49530
rect 50308 49478 50338 49530
rect 50362 49478 50372 49530
rect 50372 49478 50418 49530
rect 50442 49478 50488 49530
rect 50488 49478 50498 49530
rect 50522 49478 50552 49530
rect 50552 49478 50578 49530
rect 50282 49476 50338 49478
rect 50362 49476 50418 49478
rect 50442 49476 50498 49478
rect 50522 49476 50578 49478
rect 50282 48442 50338 48444
rect 50362 48442 50418 48444
rect 50442 48442 50498 48444
rect 50522 48442 50578 48444
rect 50282 48390 50308 48442
rect 50308 48390 50338 48442
rect 50362 48390 50372 48442
rect 50372 48390 50418 48442
rect 50442 48390 50488 48442
rect 50488 48390 50498 48442
rect 50522 48390 50552 48442
rect 50552 48390 50578 48442
rect 50282 48388 50338 48390
rect 50362 48388 50418 48390
rect 50442 48388 50498 48390
rect 50522 48388 50578 48390
rect 50282 47354 50338 47356
rect 50362 47354 50418 47356
rect 50442 47354 50498 47356
rect 50522 47354 50578 47356
rect 50282 47302 50308 47354
rect 50308 47302 50338 47354
rect 50362 47302 50372 47354
rect 50372 47302 50418 47354
rect 50442 47302 50488 47354
rect 50488 47302 50498 47354
rect 50522 47302 50552 47354
rect 50552 47302 50578 47354
rect 50282 47300 50338 47302
rect 50362 47300 50418 47302
rect 50442 47300 50498 47302
rect 50522 47300 50578 47302
rect 50282 46266 50338 46268
rect 50362 46266 50418 46268
rect 50442 46266 50498 46268
rect 50522 46266 50578 46268
rect 50282 46214 50308 46266
rect 50308 46214 50338 46266
rect 50362 46214 50372 46266
rect 50372 46214 50418 46266
rect 50442 46214 50488 46266
rect 50488 46214 50498 46266
rect 50522 46214 50552 46266
rect 50552 46214 50578 46266
rect 50282 46212 50338 46214
rect 50362 46212 50418 46214
rect 50442 46212 50498 46214
rect 50522 46212 50578 46214
rect 50282 45178 50338 45180
rect 50362 45178 50418 45180
rect 50442 45178 50498 45180
rect 50522 45178 50578 45180
rect 50282 45126 50308 45178
rect 50308 45126 50338 45178
rect 50362 45126 50372 45178
rect 50372 45126 50418 45178
rect 50442 45126 50488 45178
rect 50488 45126 50498 45178
rect 50522 45126 50552 45178
rect 50552 45126 50578 45178
rect 50282 45124 50338 45126
rect 50362 45124 50418 45126
rect 50442 45124 50498 45126
rect 50522 45124 50578 45126
rect 50282 44090 50338 44092
rect 50362 44090 50418 44092
rect 50442 44090 50498 44092
rect 50522 44090 50578 44092
rect 50282 44038 50308 44090
rect 50308 44038 50338 44090
rect 50362 44038 50372 44090
rect 50372 44038 50418 44090
rect 50442 44038 50488 44090
rect 50488 44038 50498 44090
rect 50522 44038 50552 44090
rect 50552 44038 50578 44090
rect 50282 44036 50338 44038
rect 50362 44036 50418 44038
rect 50442 44036 50498 44038
rect 50522 44036 50578 44038
rect 50282 43002 50338 43004
rect 50362 43002 50418 43004
rect 50442 43002 50498 43004
rect 50522 43002 50578 43004
rect 50282 42950 50308 43002
rect 50308 42950 50338 43002
rect 50362 42950 50372 43002
rect 50372 42950 50418 43002
rect 50442 42950 50488 43002
rect 50488 42950 50498 43002
rect 50522 42950 50552 43002
rect 50552 42950 50578 43002
rect 50282 42948 50338 42950
rect 50362 42948 50418 42950
rect 50442 42948 50498 42950
rect 50522 42948 50578 42950
rect 50282 41914 50338 41916
rect 50362 41914 50418 41916
rect 50442 41914 50498 41916
rect 50522 41914 50578 41916
rect 50282 41862 50308 41914
rect 50308 41862 50338 41914
rect 50362 41862 50372 41914
rect 50372 41862 50418 41914
rect 50442 41862 50488 41914
rect 50488 41862 50498 41914
rect 50522 41862 50552 41914
rect 50552 41862 50578 41914
rect 50282 41860 50338 41862
rect 50362 41860 50418 41862
rect 50442 41860 50498 41862
rect 50522 41860 50578 41862
rect 50282 40826 50338 40828
rect 50362 40826 50418 40828
rect 50442 40826 50498 40828
rect 50522 40826 50578 40828
rect 50282 40774 50308 40826
rect 50308 40774 50338 40826
rect 50362 40774 50372 40826
rect 50372 40774 50418 40826
rect 50442 40774 50488 40826
rect 50488 40774 50498 40826
rect 50522 40774 50552 40826
rect 50552 40774 50578 40826
rect 50282 40772 50338 40774
rect 50362 40772 50418 40774
rect 50442 40772 50498 40774
rect 50522 40772 50578 40774
rect 50282 39738 50338 39740
rect 50362 39738 50418 39740
rect 50442 39738 50498 39740
rect 50522 39738 50578 39740
rect 50282 39686 50308 39738
rect 50308 39686 50338 39738
rect 50362 39686 50372 39738
rect 50372 39686 50418 39738
rect 50442 39686 50488 39738
rect 50488 39686 50498 39738
rect 50522 39686 50552 39738
rect 50552 39686 50578 39738
rect 50282 39684 50338 39686
rect 50362 39684 50418 39686
rect 50442 39684 50498 39686
rect 50522 39684 50578 39686
rect 50282 38650 50338 38652
rect 50362 38650 50418 38652
rect 50442 38650 50498 38652
rect 50522 38650 50578 38652
rect 50282 38598 50308 38650
rect 50308 38598 50338 38650
rect 50362 38598 50372 38650
rect 50372 38598 50418 38650
rect 50442 38598 50488 38650
rect 50488 38598 50498 38650
rect 50522 38598 50552 38650
rect 50552 38598 50578 38650
rect 50282 38596 50338 38598
rect 50362 38596 50418 38598
rect 50442 38596 50498 38598
rect 50522 38596 50578 38598
rect 50282 37562 50338 37564
rect 50362 37562 50418 37564
rect 50442 37562 50498 37564
rect 50522 37562 50578 37564
rect 50282 37510 50308 37562
rect 50308 37510 50338 37562
rect 50362 37510 50372 37562
rect 50372 37510 50418 37562
rect 50442 37510 50488 37562
rect 50488 37510 50498 37562
rect 50522 37510 50552 37562
rect 50552 37510 50578 37562
rect 50282 37508 50338 37510
rect 50362 37508 50418 37510
rect 50442 37508 50498 37510
rect 50522 37508 50578 37510
rect 50282 36474 50338 36476
rect 50362 36474 50418 36476
rect 50442 36474 50498 36476
rect 50522 36474 50578 36476
rect 50282 36422 50308 36474
rect 50308 36422 50338 36474
rect 50362 36422 50372 36474
rect 50372 36422 50418 36474
rect 50442 36422 50488 36474
rect 50488 36422 50498 36474
rect 50522 36422 50552 36474
rect 50552 36422 50578 36474
rect 50282 36420 50338 36422
rect 50362 36420 50418 36422
rect 50442 36420 50498 36422
rect 50522 36420 50578 36422
rect 50282 35386 50338 35388
rect 50362 35386 50418 35388
rect 50442 35386 50498 35388
rect 50522 35386 50578 35388
rect 50282 35334 50308 35386
rect 50308 35334 50338 35386
rect 50362 35334 50372 35386
rect 50372 35334 50418 35386
rect 50442 35334 50488 35386
rect 50488 35334 50498 35386
rect 50522 35334 50552 35386
rect 50552 35334 50578 35386
rect 50282 35332 50338 35334
rect 50362 35332 50418 35334
rect 50442 35332 50498 35334
rect 50522 35332 50578 35334
rect 50282 34298 50338 34300
rect 50362 34298 50418 34300
rect 50442 34298 50498 34300
rect 50522 34298 50578 34300
rect 50282 34246 50308 34298
rect 50308 34246 50338 34298
rect 50362 34246 50372 34298
rect 50372 34246 50418 34298
rect 50442 34246 50488 34298
rect 50488 34246 50498 34298
rect 50522 34246 50552 34298
rect 50552 34246 50578 34298
rect 50282 34244 50338 34246
rect 50362 34244 50418 34246
rect 50442 34244 50498 34246
rect 50522 34244 50578 34246
rect 50282 33210 50338 33212
rect 50362 33210 50418 33212
rect 50442 33210 50498 33212
rect 50522 33210 50578 33212
rect 50282 33158 50308 33210
rect 50308 33158 50338 33210
rect 50362 33158 50372 33210
rect 50372 33158 50418 33210
rect 50442 33158 50488 33210
rect 50488 33158 50498 33210
rect 50522 33158 50552 33210
rect 50552 33158 50578 33210
rect 50282 33156 50338 33158
rect 50362 33156 50418 33158
rect 50442 33156 50498 33158
rect 50522 33156 50578 33158
rect 50282 32122 50338 32124
rect 50362 32122 50418 32124
rect 50442 32122 50498 32124
rect 50522 32122 50578 32124
rect 50282 32070 50308 32122
rect 50308 32070 50338 32122
rect 50362 32070 50372 32122
rect 50372 32070 50418 32122
rect 50442 32070 50488 32122
rect 50488 32070 50498 32122
rect 50522 32070 50552 32122
rect 50552 32070 50578 32122
rect 50282 32068 50338 32070
rect 50362 32068 50418 32070
rect 50442 32068 50498 32070
rect 50522 32068 50578 32070
rect 50282 31034 50338 31036
rect 50362 31034 50418 31036
rect 50442 31034 50498 31036
rect 50522 31034 50578 31036
rect 50282 30982 50308 31034
rect 50308 30982 50338 31034
rect 50362 30982 50372 31034
rect 50372 30982 50418 31034
rect 50442 30982 50488 31034
rect 50488 30982 50498 31034
rect 50522 30982 50552 31034
rect 50552 30982 50578 31034
rect 50282 30980 50338 30982
rect 50362 30980 50418 30982
rect 50442 30980 50498 30982
rect 50522 30980 50578 30982
rect 50282 29946 50338 29948
rect 50362 29946 50418 29948
rect 50442 29946 50498 29948
rect 50522 29946 50578 29948
rect 50282 29894 50308 29946
rect 50308 29894 50338 29946
rect 50362 29894 50372 29946
rect 50372 29894 50418 29946
rect 50442 29894 50488 29946
rect 50488 29894 50498 29946
rect 50522 29894 50552 29946
rect 50552 29894 50578 29946
rect 50282 29892 50338 29894
rect 50362 29892 50418 29894
rect 50442 29892 50498 29894
rect 50522 29892 50578 29894
rect 50282 28858 50338 28860
rect 50362 28858 50418 28860
rect 50442 28858 50498 28860
rect 50522 28858 50578 28860
rect 50282 28806 50308 28858
rect 50308 28806 50338 28858
rect 50362 28806 50372 28858
rect 50372 28806 50418 28858
rect 50442 28806 50488 28858
rect 50488 28806 50498 28858
rect 50522 28806 50552 28858
rect 50552 28806 50578 28858
rect 50282 28804 50338 28806
rect 50362 28804 50418 28806
rect 50442 28804 50498 28806
rect 50522 28804 50578 28806
rect 50282 27770 50338 27772
rect 50362 27770 50418 27772
rect 50442 27770 50498 27772
rect 50522 27770 50578 27772
rect 50282 27718 50308 27770
rect 50308 27718 50338 27770
rect 50362 27718 50372 27770
rect 50372 27718 50418 27770
rect 50442 27718 50488 27770
rect 50488 27718 50498 27770
rect 50522 27718 50552 27770
rect 50552 27718 50578 27770
rect 50282 27716 50338 27718
rect 50362 27716 50418 27718
rect 50442 27716 50498 27718
rect 50522 27716 50578 27718
rect 50282 26682 50338 26684
rect 50362 26682 50418 26684
rect 50442 26682 50498 26684
rect 50522 26682 50578 26684
rect 50282 26630 50308 26682
rect 50308 26630 50338 26682
rect 50362 26630 50372 26682
rect 50372 26630 50418 26682
rect 50442 26630 50488 26682
rect 50488 26630 50498 26682
rect 50522 26630 50552 26682
rect 50552 26630 50578 26682
rect 50282 26628 50338 26630
rect 50362 26628 50418 26630
rect 50442 26628 50498 26630
rect 50522 26628 50578 26630
rect 50282 25594 50338 25596
rect 50362 25594 50418 25596
rect 50442 25594 50498 25596
rect 50522 25594 50578 25596
rect 50282 25542 50308 25594
rect 50308 25542 50338 25594
rect 50362 25542 50372 25594
rect 50372 25542 50418 25594
rect 50442 25542 50488 25594
rect 50488 25542 50498 25594
rect 50522 25542 50552 25594
rect 50552 25542 50578 25594
rect 50282 25540 50338 25542
rect 50362 25540 50418 25542
rect 50442 25540 50498 25542
rect 50522 25540 50578 25542
rect 50282 24506 50338 24508
rect 50362 24506 50418 24508
rect 50442 24506 50498 24508
rect 50522 24506 50578 24508
rect 50282 24454 50308 24506
rect 50308 24454 50338 24506
rect 50362 24454 50372 24506
rect 50372 24454 50418 24506
rect 50442 24454 50488 24506
rect 50488 24454 50498 24506
rect 50522 24454 50552 24506
rect 50552 24454 50578 24506
rect 50282 24452 50338 24454
rect 50362 24452 50418 24454
rect 50442 24452 50498 24454
rect 50522 24452 50578 24454
rect 50282 23418 50338 23420
rect 50362 23418 50418 23420
rect 50442 23418 50498 23420
rect 50522 23418 50578 23420
rect 50282 23366 50308 23418
rect 50308 23366 50338 23418
rect 50362 23366 50372 23418
rect 50372 23366 50418 23418
rect 50442 23366 50488 23418
rect 50488 23366 50498 23418
rect 50522 23366 50552 23418
rect 50552 23366 50578 23418
rect 50282 23364 50338 23366
rect 50362 23364 50418 23366
rect 50442 23364 50498 23366
rect 50522 23364 50578 23366
rect 50282 22330 50338 22332
rect 50362 22330 50418 22332
rect 50442 22330 50498 22332
rect 50522 22330 50578 22332
rect 50282 22278 50308 22330
rect 50308 22278 50338 22330
rect 50362 22278 50372 22330
rect 50372 22278 50418 22330
rect 50442 22278 50488 22330
rect 50488 22278 50498 22330
rect 50522 22278 50552 22330
rect 50552 22278 50578 22330
rect 50282 22276 50338 22278
rect 50362 22276 50418 22278
rect 50442 22276 50498 22278
rect 50522 22276 50578 22278
rect 50282 21242 50338 21244
rect 50362 21242 50418 21244
rect 50442 21242 50498 21244
rect 50522 21242 50578 21244
rect 50282 21190 50308 21242
rect 50308 21190 50338 21242
rect 50362 21190 50372 21242
rect 50372 21190 50418 21242
rect 50442 21190 50488 21242
rect 50488 21190 50498 21242
rect 50522 21190 50552 21242
rect 50552 21190 50578 21242
rect 50282 21188 50338 21190
rect 50362 21188 50418 21190
rect 50442 21188 50498 21190
rect 50522 21188 50578 21190
rect 50282 20154 50338 20156
rect 50362 20154 50418 20156
rect 50442 20154 50498 20156
rect 50522 20154 50578 20156
rect 50282 20102 50308 20154
rect 50308 20102 50338 20154
rect 50362 20102 50372 20154
rect 50372 20102 50418 20154
rect 50442 20102 50488 20154
rect 50488 20102 50498 20154
rect 50522 20102 50552 20154
rect 50552 20102 50578 20154
rect 50282 20100 50338 20102
rect 50362 20100 50418 20102
rect 50442 20100 50498 20102
rect 50522 20100 50578 20102
rect 50282 19066 50338 19068
rect 50362 19066 50418 19068
rect 50442 19066 50498 19068
rect 50522 19066 50578 19068
rect 50282 19014 50308 19066
rect 50308 19014 50338 19066
rect 50362 19014 50372 19066
rect 50372 19014 50418 19066
rect 50442 19014 50488 19066
rect 50488 19014 50498 19066
rect 50522 19014 50552 19066
rect 50552 19014 50578 19066
rect 50282 19012 50338 19014
rect 50362 19012 50418 19014
rect 50442 19012 50498 19014
rect 50522 19012 50578 19014
rect 50282 17978 50338 17980
rect 50362 17978 50418 17980
rect 50442 17978 50498 17980
rect 50522 17978 50578 17980
rect 50282 17926 50308 17978
rect 50308 17926 50338 17978
rect 50362 17926 50372 17978
rect 50372 17926 50418 17978
rect 50442 17926 50488 17978
rect 50488 17926 50498 17978
rect 50522 17926 50552 17978
rect 50552 17926 50578 17978
rect 50282 17924 50338 17926
rect 50362 17924 50418 17926
rect 50442 17924 50498 17926
rect 50522 17924 50578 17926
rect 50282 16890 50338 16892
rect 50362 16890 50418 16892
rect 50442 16890 50498 16892
rect 50522 16890 50578 16892
rect 50282 16838 50308 16890
rect 50308 16838 50338 16890
rect 50362 16838 50372 16890
rect 50372 16838 50418 16890
rect 50442 16838 50488 16890
rect 50488 16838 50498 16890
rect 50522 16838 50552 16890
rect 50552 16838 50578 16890
rect 50282 16836 50338 16838
rect 50362 16836 50418 16838
rect 50442 16836 50498 16838
rect 50522 16836 50578 16838
rect 50282 15802 50338 15804
rect 50362 15802 50418 15804
rect 50442 15802 50498 15804
rect 50522 15802 50578 15804
rect 50282 15750 50308 15802
rect 50308 15750 50338 15802
rect 50362 15750 50372 15802
rect 50372 15750 50418 15802
rect 50442 15750 50488 15802
rect 50488 15750 50498 15802
rect 50522 15750 50552 15802
rect 50552 15750 50578 15802
rect 50282 15748 50338 15750
rect 50362 15748 50418 15750
rect 50442 15748 50498 15750
rect 50522 15748 50578 15750
rect 50282 14714 50338 14716
rect 50362 14714 50418 14716
rect 50442 14714 50498 14716
rect 50522 14714 50578 14716
rect 50282 14662 50308 14714
rect 50308 14662 50338 14714
rect 50362 14662 50372 14714
rect 50372 14662 50418 14714
rect 50442 14662 50488 14714
rect 50488 14662 50498 14714
rect 50522 14662 50552 14714
rect 50552 14662 50578 14714
rect 50282 14660 50338 14662
rect 50362 14660 50418 14662
rect 50442 14660 50498 14662
rect 50522 14660 50578 14662
rect 50282 13626 50338 13628
rect 50362 13626 50418 13628
rect 50442 13626 50498 13628
rect 50522 13626 50578 13628
rect 50282 13574 50308 13626
rect 50308 13574 50338 13626
rect 50362 13574 50372 13626
rect 50372 13574 50418 13626
rect 50442 13574 50488 13626
rect 50488 13574 50498 13626
rect 50522 13574 50552 13626
rect 50552 13574 50578 13626
rect 50282 13572 50338 13574
rect 50362 13572 50418 13574
rect 50442 13572 50498 13574
rect 50522 13572 50578 13574
rect 50282 12538 50338 12540
rect 50362 12538 50418 12540
rect 50442 12538 50498 12540
rect 50522 12538 50578 12540
rect 50282 12486 50308 12538
rect 50308 12486 50338 12538
rect 50362 12486 50372 12538
rect 50372 12486 50418 12538
rect 50442 12486 50488 12538
rect 50488 12486 50498 12538
rect 50522 12486 50552 12538
rect 50552 12486 50578 12538
rect 50282 12484 50338 12486
rect 50362 12484 50418 12486
rect 50442 12484 50498 12486
rect 50522 12484 50578 12486
rect 50282 11450 50338 11452
rect 50362 11450 50418 11452
rect 50442 11450 50498 11452
rect 50522 11450 50578 11452
rect 50282 11398 50308 11450
rect 50308 11398 50338 11450
rect 50362 11398 50372 11450
rect 50372 11398 50418 11450
rect 50442 11398 50488 11450
rect 50488 11398 50498 11450
rect 50522 11398 50552 11450
rect 50552 11398 50578 11450
rect 50282 11396 50338 11398
rect 50362 11396 50418 11398
rect 50442 11396 50498 11398
rect 50522 11396 50578 11398
rect 50282 10362 50338 10364
rect 50362 10362 50418 10364
rect 50442 10362 50498 10364
rect 50522 10362 50578 10364
rect 50282 10310 50308 10362
rect 50308 10310 50338 10362
rect 50362 10310 50372 10362
rect 50372 10310 50418 10362
rect 50442 10310 50488 10362
rect 50488 10310 50498 10362
rect 50522 10310 50552 10362
rect 50552 10310 50578 10362
rect 50282 10308 50338 10310
rect 50362 10308 50418 10310
rect 50442 10308 50498 10310
rect 50522 10308 50578 10310
rect 50282 9274 50338 9276
rect 50362 9274 50418 9276
rect 50442 9274 50498 9276
rect 50522 9274 50578 9276
rect 50282 9222 50308 9274
rect 50308 9222 50338 9274
rect 50362 9222 50372 9274
rect 50372 9222 50418 9274
rect 50442 9222 50488 9274
rect 50488 9222 50498 9274
rect 50522 9222 50552 9274
rect 50552 9222 50578 9274
rect 50282 9220 50338 9222
rect 50362 9220 50418 9222
rect 50442 9220 50498 9222
rect 50522 9220 50578 9222
rect 50282 8186 50338 8188
rect 50362 8186 50418 8188
rect 50442 8186 50498 8188
rect 50522 8186 50578 8188
rect 50282 8134 50308 8186
rect 50308 8134 50338 8186
rect 50362 8134 50372 8186
rect 50372 8134 50418 8186
rect 50442 8134 50488 8186
rect 50488 8134 50498 8186
rect 50522 8134 50552 8186
rect 50552 8134 50578 8186
rect 50282 8132 50338 8134
rect 50362 8132 50418 8134
rect 50442 8132 50498 8134
rect 50522 8132 50578 8134
rect 50282 7098 50338 7100
rect 50362 7098 50418 7100
rect 50442 7098 50498 7100
rect 50522 7098 50578 7100
rect 50282 7046 50308 7098
rect 50308 7046 50338 7098
rect 50362 7046 50372 7098
rect 50372 7046 50418 7098
rect 50442 7046 50488 7098
rect 50488 7046 50498 7098
rect 50522 7046 50552 7098
rect 50552 7046 50578 7098
rect 50282 7044 50338 7046
rect 50362 7044 50418 7046
rect 50442 7044 50498 7046
rect 50522 7044 50578 7046
rect 50282 6010 50338 6012
rect 50362 6010 50418 6012
rect 50442 6010 50498 6012
rect 50522 6010 50578 6012
rect 50282 5958 50308 6010
rect 50308 5958 50338 6010
rect 50362 5958 50372 6010
rect 50372 5958 50418 6010
rect 50442 5958 50488 6010
rect 50488 5958 50498 6010
rect 50522 5958 50552 6010
rect 50552 5958 50578 6010
rect 50282 5956 50338 5958
rect 50362 5956 50418 5958
rect 50442 5956 50498 5958
rect 50522 5956 50578 5958
rect 50282 4922 50338 4924
rect 50362 4922 50418 4924
rect 50442 4922 50498 4924
rect 50522 4922 50578 4924
rect 50282 4870 50308 4922
rect 50308 4870 50338 4922
rect 50362 4870 50372 4922
rect 50372 4870 50418 4922
rect 50442 4870 50488 4922
rect 50488 4870 50498 4922
rect 50522 4870 50552 4922
rect 50552 4870 50578 4922
rect 50282 4868 50338 4870
rect 50362 4868 50418 4870
rect 50442 4868 50498 4870
rect 50522 4868 50578 4870
rect 52256 56752 52312 56808
rect 50282 3834 50338 3836
rect 50362 3834 50418 3836
rect 50442 3834 50498 3836
rect 50522 3834 50578 3836
rect 50282 3782 50308 3834
rect 50308 3782 50338 3834
rect 50362 3782 50372 3834
rect 50372 3782 50418 3834
rect 50442 3782 50488 3834
rect 50488 3782 50498 3834
rect 50522 3782 50552 3834
rect 50552 3782 50578 3834
rect 50282 3780 50338 3782
rect 50362 3780 50418 3782
rect 50442 3780 50498 3782
rect 50522 3780 50578 3782
rect 50282 2746 50338 2748
rect 50362 2746 50418 2748
rect 50442 2746 50498 2748
rect 50522 2746 50578 2748
rect 50282 2694 50308 2746
rect 50308 2694 50338 2746
rect 50362 2694 50372 2746
rect 50372 2694 50418 2746
rect 50442 2694 50488 2746
rect 50488 2694 50498 2746
rect 50522 2694 50552 2746
rect 50552 2694 50578 2746
rect 50282 2692 50338 2694
rect 50362 2692 50418 2694
rect 50442 2692 50498 2694
rect 50522 2692 50578 2694
<< metal3 >>
rect 4190 57696 4510 57697
rect 4190 57632 4198 57696
rect 4262 57632 4278 57696
rect 4342 57632 4358 57696
rect 4422 57632 4438 57696
rect 4502 57632 4510 57696
rect 4190 57631 4510 57632
rect 34910 57696 35230 57697
rect 34910 57632 34918 57696
rect 34982 57632 34998 57696
rect 35062 57632 35078 57696
rect 35142 57632 35158 57696
rect 35222 57632 35230 57696
rect 34910 57631 35230 57632
rect 19550 57152 19870 57153
rect 19550 57088 19558 57152
rect 19622 57088 19638 57152
rect 19702 57088 19718 57152
rect 19782 57088 19798 57152
rect 19862 57088 19870 57152
rect 19550 57087 19870 57088
rect 50270 57152 50590 57153
rect 50270 57088 50278 57152
rect 50342 57088 50358 57152
rect 50422 57088 50438 57152
rect 50502 57088 50518 57152
rect 50582 57088 50590 57152
rect 50270 57087 50590 57088
rect 52251 56810 52317 56813
rect 51196 56808 52317 56810
rect 51196 56752 52256 56808
rect 52312 56752 52317 56808
rect 51196 56750 52317 56752
rect 51196 56677 51256 56750
rect 52251 56747 52317 56750
rect 51196 56672 51305 56677
rect 51196 56616 51244 56672
rect 51300 56616 51305 56672
rect 51196 56614 51305 56616
rect 51239 56611 51305 56614
rect 4190 56608 4510 56609
rect 4190 56544 4198 56608
rect 4262 56544 4278 56608
rect 4342 56544 4358 56608
rect 4422 56544 4438 56608
rect 4502 56544 4510 56608
rect 4190 56543 4510 56544
rect 34910 56608 35230 56609
rect 34910 56544 34918 56608
rect 34982 56544 34998 56608
rect 35062 56544 35078 56608
rect 35142 56544 35158 56608
rect 35222 56544 35230 56608
rect 34910 56543 35230 56544
rect 38635 56402 38701 56405
rect 46179 56402 46245 56405
rect 38635 56400 46245 56402
rect 38635 56344 38640 56400
rect 38696 56344 46184 56400
rect 46240 56344 46245 56400
rect 38635 56342 46245 56344
rect 38635 56339 38701 56342
rect 46179 56339 46245 56342
rect 25479 56266 25545 56269
rect 31643 56266 31709 56269
rect 25479 56264 31709 56266
rect 25479 56208 25484 56264
rect 25540 56208 31648 56264
rect 31704 56208 31709 56264
rect 25479 56206 31709 56208
rect 25479 56203 25545 56206
rect 31643 56203 31709 56206
rect 33851 56266 33917 56269
rect 35967 56266 36033 56269
rect 33851 56264 36033 56266
rect 33851 56208 33856 56264
rect 33912 56208 35972 56264
rect 36028 56208 36033 56264
rect 33851 56206 36033 56208
rect 33851 56203 33917 56206
rect 35967 56203 36033 56206
rect 32563 56130 32629 56133
rect 40935 56130 41001 56133
rect 32563 56128 41001 56130
rect 32563 56072 32568 56128
rect 32624 56072 40940 56128
rect 40996 56072 41001 56128
rect 32563 56070 41001 56072
rect 32563 56067 32629 56070
rect 40935 56067 41001 56070
rect 41211 56130 41277 56133
rect 41395 56130 41461 56133
rect 41211 56128 41461 56130
rect 41211 56072 41216 56128
rect 41272 56072 41400 56128
rect 41456 56072 41461 56128
rect 41211 56070 41461 56072
rect 41211 56067 41277 56070
rect 41395 56067 41461 56070
rect 19550 56064 19870 56065
rect 19550 56000 19558 56064
rect 19622 56000 19638 56064
rect 19702 56000 19718 56064
rect 19782 56000 19798 56064
rect 19862 56000 19870 56064
rect 19550 55999 19870 56000
rect 50270 56064 50590 56065
rect 50270 56000 50278 56064
rect 50342 56000 50358 56064
rect 50422 56000 50438 56064
rect 50502 56000 50518 56064
rect 50582 56000 50590 56064
rect 50270 55999 50590 56000
rect 31275 55994 31341 55997
rect 31827 55994 31893 55997
rect 31275 55992 31893 55994
rect 31275 55936 31280 55992
rect 31336 55936 31832 55992
rect 31888 55936 31893 55992
rect 31275 55934 31893 55936
rect 31275 55931 31341 55934
rect 31827 55931 31893 55934
rect 32471 55994 32537 55997
rect 41487 55994 41553 55997
rect 32471 55992 41553 55994
rect 32471 55936 32476 55992
rect 32532 55936 41492 55992
rect 41548 55936 41553 55992
rect 32471 55934 41553 55936
rect 32471 55931 32537 55934
rect 41487 55931 41553 55934
rect 2111 55858 2177 55861
rect 47007 55858 47073 55861
rect 2111 55856 47073 55858
rect 2111 55800 2116 55856
rect 2172 55800 47012 55856
rect 47068 55800 47073 55856
rect 2111 55798 47073 55800
rect 2111 55795 2177 55798
rect 47007 55795 47073 55798
rect 41395 55722 41461 55725
rect 43879 55722 43945 55725
rect 41395 55720 43945 55722
rect 41395 55664 41400 55720
rect 41456 55664 43884 55720
rect 43940 55664 43945 55720
rect 41395 55662 43945 55664
rect 41395 55659 41461 55662
rect 43879 55659 43945 55662
rect 4190 55520 4510 55521
rect 4190 55456 4198 55520
rect 4262 55456 4278 55520
rect 4342 55456 4358 55520
rect 4422 55456 4438 55520
rect 4502 55456 4510 55520
rect 4190 55455 4510 55456
rect 34910 55520 35230 55521
rect 34910 55456 34918 55520
rect 34982 55456 34998 55520
rect 35062 55456 35078 55520
rect 35142 55456 35158 55520
rect 35222 55456 35230 55520
rect 34910 55455 35230 55456
rect 19550 54976 19870 54977
rect 19550 54912 19558 54976
rect 19622 54912 19638 54976
rect 19702 54912 19718 54976
rect 19782 54912 19798 54976
rect 19862 54912 19870 54976
rect 19550 54911 19870 54912
rect 50270 54976 50590 54977
rect 50270 54912 50278 54976
rect 50342 54912 50358 54976
rect 50422 54912 50438 54976
rect 50502 54912 50518 54976
rect 50582 54912 50590 54976
rect 50270 54911 50590 54912
rect 4190 54432 4510 54433
rect 4190 54368 4198 54432
rect 4262 54368 4278 54432
rect 4342 54368 4358 54432
rect 4422 54368 4438 54432
rect 4502 54368 4510 54432
rect 4190 54367 4510 54368
rect 34910 54432 35230 54433
rect 34910 54368 34918 54432
rect 34982 54368 34998 54432
rect 35062 54368 35078 54432
rect 35142 54368 35158 54432
rect 35222 54368 35230 54432
rect 34910 54367 35230 54368
rect 19550 53888 19870 53889
rect 19550 53824 19558 53888
rect 19622 53824 19638 53888
rect 19702 53824 19718 53888
rect 19782 53824 19798 53888
rect 19862 53824 19870 53888
rect 19550 53823 19870 53824
rect 50270 53888 50590 53889
rect 50270 53824 50278 53888
rect 50342 53824 50358 53888
rect 50422 53824 50438 53888
rect 50502 53824 50518 53888
rect 50582 53824 50590 53888
rect 50270 53823 50590 53824
rect 4190 53344 4510 53345
rect 4190 53280 4198 53344
rect 4262 53280 4278 53344
rect 4342 53280 4358 53344
rect 4422 53280 4438 53344
rect 4502 53280 4510 53344
rect 4190 53279 4510 53280
rect 34910 53344 35230 53345
rect 34910 53280 34918 53344
rect 34982 53280 34998 53344
rect 35062 53280 35078 53344
rect 35142 53280 35158 53344
rect 35222 53280 35230 53344
rect 34910 53279 35230 53280
rect 19550 52800 19870 52801
rect 19550 52736 19558 52800
rect 19622 52736 19638 52800
rect 19702 52736 19718 52800
rect 19782 52736 19798 52800
rect 19862 52736 19870 52800
rect 19550 52735 19870 52736
rect 50270 52800 50590 52801
rect 50270 52736 50278 52800
rect 50342 52736 50358 52800
rect 50422 52736 50438 52800
rect 50502 52736 50518 52800
rect 50582 52736 50590 52800
rect 50270 52735 50590 52736
rect 4190 52256 4510 52257
rect 4190 52192 4198 52256
rect 4262 52192 4278 52256
rect 4342 52192 4358 52256
rect 4422 52192 4438 52256
rect 4502 52192 4510 52256
rect 4190 52191 4510 52192
rect 34910 52256 35230 52257
rect 34910 52192 34918 52256
rect 34982 52192 34998 52256
rect 35062 52192 35078 52256
rect 35142 52192 35158 52256
rect 35222 52192 35230 52256
rect 34910 52191 35230 52192
rect 19550 51712 19870 51713
rect 19550 51648 19558 51712
rect 19622 51648 19638 51712
rect 19702 51648 19718 51712
rect 19782 51648 19798 51712
rect 19862 51648 19870 51712
rect 19550 51647 19870 51648
rect 50270 51712 50590 51713
rect 50270 51648 50278 51712
rect 50342 51648 50358 51712
rect 50422 51648 50438 51712
rect 50502 51648 50518 51712
rect 50582 51648 50590 51712
rect 50270 51647 50590 51648
rect 4190 51168 4510 51169
rect 4190 51104 4198 51168
rect 4262 51104 4278 51168
rect 4342 51104 4358 51168
rect 4422 51104 4438 51168
rect 4502 51104 4510 51168
rect 4190 51103 4510 51104
rect 34910 51168 35230 51169
rect 34910 51104 34918 51168
rect 34982 51104 34998 51168
rect 35062 51104 35078 51168
rect 35142 51104 35158 51168
rect 35222 51104 35230 51168
rect 34910 51103 35230 51104
rect 19550 50624 19870 50625
rect 19550 50560 19558 50624
rect 19622 50560 19638 50624
rect 19702 50560 19718 50624
rect 19782 50560 19798 50624
rect 19862 50560 19870 50624
rect 19550 50559 19870 50560
rect 50270 50624 50590 50625
rect 50270 50560 50278 50624
rect 50342 50560 50358 50624
rect 50422 50560 50438 50624
rect 50502 50560 50518 50624
rect 50582 50560 50590 50624
rect 50270 50559 50590 50560
rect 4190 50080 4510 50081
rect 4190 50016 4198 50080
rect 4262 50016 4278 50080
rect 4342 50016 4358 50080
rect 4422 50016 4438 50080
rect 4502 50016 4510 50080
rect 4190 50015 4510 50016
rect 34910 50080 35230 50081
rect 34910 50016 34918 50080
rect 34982 50016 34998 50080
rect 35062 50016 35078 50080
rect 35142 50016 35158 50080
rect 35222 50016 35230 50080
rect 34910 50015 35230 50016
rect 19550 49536 19870 49537
rect 19550 49472 19558 49536
rect 19622 49472 19638 49536
rect 19702 49472 19718 49536
rect 19782 49472 19798 49536
rect 19862 49472 19870 49536
rect 19550 49471 19870 49472
rect 50270 49536 50590 49537
rect 50270 49472 50278 49536
rect 50342 49472 50358 49536
rect 50422 49472 50438 49536
rect 50502 49472 50518 49536
rect 50582 49472 50590 49536
rect 50270 49471 50590 49472
rect 4190 48992 4510 48993
rect 4190 48928 4198 48992
rect 4262 48928 4278 48992
rect 4342 48928 4358 48992
rect 4422 48928 4438 48992
rect 4502 48928 4510 48992
rect 4190 48927 4510 48928
rect 34910 48992 35230 48993
rect 34910 48928 34918 48992
rect 34982 48928 34998 48992
rect 35062 48928 35078 48992
rect 35142 48928 35158 48992
rect 35222 48928 35230 48992
rect 34910 48927 35230 48928
rect 19550 48448 19870 48449
rect 19550 48384 19558 48448
rect 19622 48384 19638 48448
rect 19702 48384 19718 48448
rect 19782 48384 19798 48448
rect 19862 48384 19870 48448
rect 19550 48383 19870 48384
rect 50270 48448 50590 48449
rect 50270 48384 50278 48448
rect 50342 48384 50358 48448
rect 50422 48384 50438 48448
rect 50502 48384 50518 48448
rect 50582 48384 50590 48448
rect 50270 48383 50590 48384
rect 4190 47904 4510 47905
rect 4190 47840 4198 47904
rect 4262 47840 4278 47904
rect 4342 47840 4358 47904
rect 4422 47840 4438 47904
rect 4502 47840 4510 47904
rect 4190 47839 4510 47840
rect 34910 47904 35230 47905
rect 34910 47840 34918 47904
rect 34982 47840 34998 47904
rect 35062 47840 35078 47904
rect 35142 47840 35158 47904
rect 35222 47840 35230 47904
rect 34910 47839 35230 47840
rect 19550 47360 19870 47361
rect 19550 47296 19558 47360
rect 19622 47296 19638 47360
rect 19702 47296 19718 47360
rect 19782 47296 19798 47360
rect 19862 47296 19870 47360
rect 19550 47295 19870 47296
rect 50270 47360 50590 47361
rect 50270 47296 50278 47360
rect 50342 47296 50358 47360
rect 50422 47296 50438 47360
rect 50502 47296 50518 47360
rect 50582 47296 50590 47360
rect 50270 47295 50590 47296
rect 4190 46816 4510 46817
rect 4190 46752 4198 46816
rect 4262 46752 4278 46816
rect 4342 46752 4358 46816
rect 4422 46752 4438 46816
rect 4502 46752 4510 46816
rect 4190 46751 4510 46752
rect 34910 46816 35230 46817
rect 34910 46752 34918 46816
rect 34982 46752 34998 46816
rect 35062 46752 35078 46816
rect 35142 46752 35158 46816
rect 35222 46752 35230 46816
rect 34910 46751 35230 46752
rect 19550 46272 19870 46273
rect 19550 46208 19558 46272
rect 19622 46208 19638 46272
rect 19702 46208 19718 46272
rect 19782 46208 19798 46272
rect 19862 46208 19870 46272
rect 19550 46207 19870 46208
rect 50270 46272 50590 46273
rect 50270 46208 50278 46272
rect 50342 46208 50358 46272
rect 50422 46208 50438 46272
rect 50502 46208 50518 46272
rect 50582 46208 50590 46272
rect 50270 46207 50590 46208
rect 4190 45728 4510 45729
rect 4190 45664 4198 45728
rect 4262 45664 4278 45728
rect 4342 45664 4358 45728
rect 4422 45664 4438 45728
rect 4502 45664 4510 45728
rect 4190 45663 4510 45664
rect 34910 45728 35230 45729
rect 34910 45664 34918 45728
rect 34982 45664 34998 45728
rect 35062 45664 35078 45728
rect 35142 45664 35158 45728
rect 35222 45664 35230 45728
rect 34910 45663 35230 45664
rect 19550 45184 19870 45185
rect 19550 45120 19558 45184
rect 19622 45120 19638 45184
rect 19702 45120 19718 45184
rect 19782 45120 19798 45184
rect 19862 45120 19870 45184
rect 19550 45119 19870 45120
rect 50270 45184 50590 45185
rect 50270 45120 50278 45184
rect 50342 45120 50358 45184
rect 50422 45120 50438 45184
rect 50502 45120 50518 45184
rect 50582 45120 50590 45184
rect 50270 45119 50590 45120
rect 4190 44640 4510 44641
rect 4190 44576 4198 44640
rect 4262 44576 4278 44640
rect 4342 44576 4358 44640
rect 4422 44576 4438 44640
rect 4502 44576 4510 44640
rect 4190 44575 4510 44576
rect 34910 44640 35230 44641
rect 34910 44576 34918 44640
rect 34982 44576 34998 44640
rect 35062 44576 35078 44640
rect 35142 44576 35158 44640
rect 35222 44576 35230 44640
rect 34910 44575 35230 44576
rect 19550 44096 19870 44097
rect 19550 44032 19558 44096
rect 19622 44032 19638 44096
rect 19702 44032 19718 44096
rect 19782 44032 19798 44096
rect 19862 44032 19870 44096
rect 19550 44031 19870 44032
rect 50270 44096 50590 44097
rect 50270 44032 50278 44096
rect 50342 44032 50358 44096
rect 50422 44032 50438 44096
rect 50502 44032 50518 44096
rect 50582 44032 50590 44096
rect 50270 44031 50590 44032
rect 4190 43552 4510 43553
rect 4190 43488 4198 43552
rect 4262 43488 4278 43552
rect 4342 43488 4358 43552
rect 4422 43488 4438 43552
rect 4502 43488 4510 43552
rect 4190 43487 4510 43488
rect 34910 43552 35230 43553
rect 34910 43488 34918 43552
rect 34982 43488 34998 43552
rect 35062 43488 35078 43552
rect 35142 43488 35158 43552
rect 35222 43488 35230 43552
rect 34910 43487 35230 43488
rect 19550 43008 19870 43009
rect 19550 42944 19558 43008
rect 19622 42944 19638 43008
rect 19702 42944 19718 43008
rect 19782 42944 19798 43008
rect 19862 42944 19870 43008
rect 19550 42943 19870 42944
rect 50270 43008 50590 43009
rect 50270 42944 50278 43008
rect 50342 42944 50358 43008
rect 50422 42944 50438 43008
rect 50502 42944 50518 43008
rect 50582 42944 50590 43008
rect 50270 42943 50590 42944
rect 4190 42464 4510 42465
rect 4190 42400 4198 42464
rect 4262 42400 4278 42464
rect 4342 42400 4358 42464
rect 4422 42400 4438 42464
rect 4502 42400 4510 42464
rect 4190 42399 4510 42400
rect 34910 42464 35230 42465
rect 34910 42400 34918 42464
rect 34982 42400 34998 42464
rect 35062 42400 35078 42464
rect 35142 42400 35158 42464
rect 35222 42400 35230 42464
rect 34910 42399 35230 42400
rect 19550 41920 19870 41921
rect 19550 41856 19558 41920
rect 19622 41856 19638 41920
rect 19702 41856 19718 41920
rect 19782 41856 19798 41920
rect 19862 41856 19870 41920
rect 19550 41855 19870 41856
rect 50270 41920 50590 41921
rect 50270 41856 50278 41920
rect 50342 41856 50358 41920
rect 50422 41856 50438 41920
rect 50502 41856 50518 41920
rect 50582 41856 50590 41920
rect 50270 41855 50590 41856
rect 4190 41376 4510 41377
rect 4190 41312 4198 41376
rect 4262 41312 4278 41376
rect 4342 41312 4358 41376
rect 4422 41312 4438 41376
rect 4502 41312 4510 41376
rect 4190 41311 4510 41312
rect 34910 41376 35230 41377
rect 34910 41312 34918 41376
rect 34982 41312 34998 41376
rect 35062 41312 35078 41376
rect 35142 41312 35158 41376
rect 35222 41312 35230 41376
rect 34910 41311 35230 41312
rect 19550 40832 19870 40833
rect 19550 40768 19558 40832
rect 19622 40768 19638 40832
rect 19702 40768 19718 40832
rect 19782 40768 19798 40832
rect 19862 40768 19870 40832
rect 19550 40767 19870 40768
rect 50270 40832 50590 40833
rect 50270 40768 50278 40832
rect 50342 40768 50358 40832
rect 50422 40768 50438 40832
rect 50502 40768 50518 40832
rect 50582 40768 50590 40832
rect 50270 40767 50590 40768
rect 4190 40288 4510 40289
rect 4190 40224 4198 40288
rect 4262 40224 4278 40288
rect 4342 40224 4358 40288
rect 4422 40224 4438 40288
rect 4502 40224 4510 40288
rect 4190 40223 4510 40224
rect 34910 40288 35230 40289
rect 34910 40224 34918 40288
rect 34982 40224 34998 40288
rect 35062 40224 35078 40288
rect 35142 40224 35158 40288
rect 35222 40224 35230 40288
rect 34910 40223 35230 40224
rect 19550 39744 19870 39745
rect 19550 39680 19558 39744
rect 19622 39680 19638 39744
rect 19702 39680 19718 39744
rect 19782 39680 19798 39744
rect 19862 39680 19870 39744
rect 19550 39679 19870 39680
rect 50270 39744 50590 39745
rect 50270 39680 50278 39744
rect 50342 39680 50358 39744
rect 50422 39680 50438 39744
rect 50502 39680 50518 39744
rect 50582 39680 50590 39744
rect 50270 39679 50590 39680
rect 4190 39200 4510 39201
rect 4190 39136 4198 39200
rect 4262 39136 4278 39200
rect 4342 39136 4358 39200
rect 4422 39136 4438 39200
rect 4502 39136 4510 39200
rect 4190 39135 4510 39136
rect 34910 39200 35230 39201
rect 34910 39136 34918 39200
rect 34982 39136 34998 39200
rect 35062 39136 35078 39200
rect 35142 39136 35158 39200
rect 35222 39136 35230 39200
rect 34910 39135 35230 39136
rect 39831 38858 39897 38861
rect 39604 38856 39897 38858
rect 39604 38800 39836 38856
rect 39892 38800 39897 38856
rect 39604 38798 39897 38800
rect 39604 38725 39664 38798
rect 39831 38795 39897 38798
rect 39604 38720 39713 38725
rect 39604 38664 39652 38720
rect 39708 38664 39713 38720
rect 39604 38662 39713 38664
rect 39647 38659 39713 38662
rect 49491 38722 49557 38725
rect 49491 38720 49600 38722
rect 49491 38664 49496 38720
rect 49552 38664 49600 38720
rect 49491 38659 49600 38664
rect 19550 38656 19870 38657
rect 19550 38592 19558 38656
rect 19622 38592 19638 38656
rect 19702 38592 19718 38656
rect 19782 38592 19798 38656
rect 19862 38592 19870 38656
rect 19550 38591 19870 38592
rect 49540 38589 49600 38659
rect 50270 38656 50590 38657
rect 50270 38592 50278 38656
rect 50342 38592 50358 38656
rect 50422 38592 50438 38656
rect 50502 38592 50518 38656
rect 50582 38592 50590 38656
rect 50270 38591 50590 38592
rect 49540 38584 49649 38589
rect 49540 38528 49588 38584
rect 49644 38528 49649 38584
rect 49540 38526 49649 38528
rect 49583 38523 49649 38526
rect 4190 38112 4510 38113
rect 4190 38048 4198 38112
rect 4262 38048 4278 38112
rect 4342 38048 4358 38112
rect 4422 38048 4438 38112
rect 4502 38048 4510 38112
rect 4190 38047 4510 38048
rect 34910 38112 35230 38113
rect 34910 38048 34918 38112
rect 34982 38048 34998 38112
rect 35062 38048 35078 38112
rect 35142 38048 35158 38112
rect 35222 38048 35230 38112
rect 34910 38047 35230 38048
rect 19550 37568 19870 37569
rect 19550 37504 19558 37568
rect 19622 37504 19638 37568
rect 19702 37504 19718 37568
rect 19782 37504 19798 37568
rect 19862 37504 19870 37568
rect 19550 37503 19870 37504
rect 50270 37568 50590 37569
rect 50270 37504 50278 37568
rect 50342 37504 50358 37568
rect 50422 37504 50438 37568
rect 50502 37504 50518 37568
rect 50582 37504 50590 37568
rect 50270 37503 50590 37504
rect 19131 37226 19197 37229
rect 27779 37226 27845 37229
rect 19131 37224 27845 37226
rect 19131 37168 19136 37224
rect 19192 37168 27784 37224
rect 27840 37168 27845 37224
rect 19131 37166 27845 37168
rect 19131 37163 19197 37166
rect 27779 37163 27845 37166
rect 4190 37024 4510 37025
rect 4190 36960 4198 37024
rect 4262 36960 4278 37024
rect 4342 36960 4358 37024
rect 4422 36960 4438 37024
rect 4502 36960 4510 37024
rect 4190 36959 4510 36960
rect 34910 37024 35230 37025
rect 34910 36960 34918 37024
rect 34982 36960 34998 37024
rect 35062 36960 35078 37024
rect 35142 36960 35158 37024
rect 35222 36960 35230 37024
rect 34910 36959 35230 36960
rect 19550 36480 19870 36481
rect 19550 36416 19558 36480
rect 19622 36416 19638 36480
rect 19702 36416 19718 36480
rect 19782 36416 19798 36480
rect 19862 36416 19870 36480
rect 19550 36415 19870 36416
rect 50270 36480 50590 36481
rect 50270 36416 50278 36480
rect 50342 36416 50358 36480
rect 50422 36416 50438 36480
rect 50502 36416 50518 36480
rect 50582 36416 50590 36480
rect 50270 36415 50590 36416
rect 34311 36138 34377 36141
rect 34311 36136 34558 36138
rect 34311 36080 34316 36136
rect 34372 36080 34558 36136
rect 34311 36078 34558 36080
rect 34311 36075 34377 36078
rect 34498 36005 34558 36078
rect 14163 36002 14229 36005
rect 14347 36002 14413 36005
rect 14163 36000 14413 36002
rect 14163 35944 14168 36000
rect 14224 35944 14352 36000
rect 14408 35944 14413 36000
rect 14163 35942 14413 35944
rect 14163 35939 14229 35942
rect 14347 35939 14413 35942
rect 34495 36000 34561 36005
rect 34495 35944 34500 36000
rect 34556 35944 34561 36000
rect 34495 35939 34561 35944
rect 4190 35936 4510 35937
rect 4190 35872 4198 35936
rect 4262 35872 4278 35936
rect 4342 35872 4358 35936
rect 4422 35872 4438 35936
rect 4502 35872 4510 35936
rect 4190 35871 4510 35872
rect 34910 35936 35230 35937
rect 34910 35872 34918 35936
rect 34982 35872 34998 35936
rect 35062 35872 35078 35936
rect 35142 35872 35158 35936
rect 35222 35872 35230 35936
rect 34910 35871 35230 35872
rect 19550 35392 19870 35393
rect 19550 35328 19558 35392
rect 19622 35328 19638 35392
rect 19702 35328 19718 35392
rect 19782 35328 19798 35392
rect 19862 35328 19870 35392
rect 19550 35327 19870 35328
rect 50270 35392 50590 35393
rect 50270 35328 50278 35392
rect 50342 35328 50358 35392
rect 50422 35328 50438 35392
rect 50502 35328 50518 35392
rect 50582 35328 50590 35392
rect 50270 35327 50590 35328
rect 4190 34848 4510 34849
rect 4190 34784 4198 34848
rect 4262 34784 4278 34848
rect 4342 34784 4358 34848
rect 4422 34784 4438 34848
rect 4502 34784 4510 34848
rect 4190 34783 4510 34784
rect 34910 34848 35230 34849
rect 34910 34784 34918 34848
rect 34982 34784 34998 34848
rect 35062 34784 35078 34848
rect 35142 34784 35158 34848
rect 35222 34784 35230 34848
rect 34910 34783 35230 34784
rect 19550 34304 19870 34305
rect 19550 34240 19558 34304
rect 19622 34240 19638 34304
rect 19702 34240 19718 34304
rect 19782 34240 19798 34304
rect 19862 34240 19870 34304
rect 19550 34239 19870 34240
rect 50270 34304 50590 34305
rect 50270 34240 50278 34304
rect 50342 34240 50358 34304
rect 50422 34240 50438 34304
rect 50502 34240 50518 34304
rect 50582 34240 50590 34304
rect 50270 34239 50590 34240
rect 4190 33760 4510 33761
rect 4190 33696 4198 33760
rect 4262 33696 4278 33760
rect 4342 33696 4358 33760
rect 4422 33696 4438 33760
rect 4502 33696 4510 33760
rect 4190 33695 4510 33696
rect 34910 33760 35230 33761
rect 34910 33696 34918 33760
rect 34982 33696 34998 33760
rect 35062 33696 35078 33760
rect 35142 33696 35158 33760
rect 35222 33696 35230 33760
rect 34910 33695 35230 33696
rect 19550 33216 19870 33217
rect 19550 33152 19558 33216
rect 19622 33152 19638 33216
rect 19702 33152 19718 33216
rect 19782 33152 19798 33216
rect 19862 33152 19870 33216
rect 19550 33151 19870 33152
rect 50270 33216 50590 33217
rect 50270 33152 50278 33216
rect 50342 33152 50358 33216
rect 50422 33152 50438 33216
rect 50502 33152 50518 33216
rect 50582 33152 50590 33216
rect 50270 33151 50590 33152
rect 4190 32672 4510 32673
rect 4190 32608 4198 32672
rect 4262 32608 4278 32672
rect 4342 32608 4358 32672
rect 4422 32608 4438 32672
rect 4502 32608 4510 32672
rect 4190 32607 4510 32608
rect 34910 32672 35230 32673
rect 34910 32608 34918 32672
rect 34982 32608 34998 32672
rect 35062 32608 35078 32672
rect 35142 32608 35158 32672
rect 35222 32608 35230 32672
rect 34910 32607 35230 32608
rect 19550 32128 19870 32129
rect 19550 32064 19558 32128
rect 19622 32064 19638 32128
rect 19702 32064 19718 32128
rect 19782 32064 19798 32128
rect 19862 32064 19870 32128
rect 19550 32063 19870 32064
rect 50270 32128 50590 32129
rect 50270 32064 50278 32128
rect 50342 32064 50358 32128
rect 50422 32064 50438 32128
rect 50502 32064 50518 32128
rect 50582 32064 50590 32128
rect 50270 32063 50590 32064
rect 4190 31584 4510 31585
rect 4190 31520 4198 31584
rect 4262 31520 4278 31584
rect 4342 31520 4358 31584
rect 4422 31520 4438 31584
rect 4502 31520 4510 31584
rect 4190 31519 4510 31520
rect 34910 31584 35230 31585
rect 34910 31520 34918 31584
rect 34982 31520 34998 31584
rect 35062 31520 35078 31584
rect 35142 31520 35158 31584
rect 35222 31520 35230 31584
rect 34910 31519 35230 31520
rect 19550 31040 19870 31041
rect 19550 30976 19558 31040
rect 19622 30976 19638 31040
rect 19702 30976 19718 31040
rect 19782 30976 19798 31040
rect 19862 30976 19870 31040
rect 19550 30975 19870 30976
rect 50270 31040 50590 31041
rect 50270 30976 50278 31040
rect 50342 30976 50358 31040
rect 50422 30976 50438 31040
rect 50502 30976 50518 31040
rect 50582 30976 50590 31040
rect 50270 30975 50590 30976
rect 4190 30496 4510 30497
rect 4190 30432 4198 30496
rect 4262 30432 4278 30496
rect 4342 30432 4358 30496
rect 4422 30432 4438 30496
rect 4502 30432 4510 30496
rect 4190 30431 4510 30432
rect 34910 30496 35230 30497
rect 34910 30432 34918 30496
rect 34982 30432 34998 30496
rect 35062 30432 35078 30496
rect 35142 30432 35158 30496
rect 35222 30432 35230 30496
rect 34910 30431 35230 30432
rect 19550 29952 19870 29953
rect 19550 29888 19558 29952
rect 19622 29888 19638 29952
rect 19702 29888 19718 29952
rect 19782 29888 19798 29952
rect 19862 29888 19870 29952
rect 19550 29887 19870 29888
rect 50270 29952 50590 29953
rect 50270 29888 50278 29952
rect 50342 29888 50358 29952
rect 50422 29888 50438 29952
rect 50502 29888 50518 29952
rect 50582 29888 50590 29952
rect 50270 29887 50590 29888
rect 4190 29408 4510 29409
rect 4190 29344 4198 29408
rect 4262 29344 4278 29408
rect 4342 29344 4358 29408
rect 4422 29344 4438 29408
rect 4502 29344 4510 29408
rect 4190 29343 4510 29344
rect 34910 29408 35230 29409
rect 34910 29344 34918 29408
rect 34982 29344 34998 29408
rect 35062 29344 35078 29408
rect 35142 29344 35158 29408
rect 35222 29344 35230 29408
rect 34910 29343 35230 29344
rect 19550 28864 19870 28865
rect 19550 28800 19558 28864
rect 19622 28800 19638 28864
rect 19702 28800 19718 28864
rect 19782 28800 19798 28864
rect 19862 28800 19870 28864
rect 19550 28799 19870 28800
rect 50270 28864 50590 28865
rect 50270 28800 50278 28864
rect 50342 28800 50358 28864
rect 50422 28800 50438 28864
rect 50502 28800 50518 28864
rect 50582 28800 50590 28864
rect 50270 28799 50590 28800
rect 4190 28320 4510 28321
rect 4190 28256 4198 28320
rect 4262 28256 4278 28320
rect 4342 28256 4358 28320
rect 4422 28256 4438 28320
rect 4502 28256 4510 28320
rect 4190 28255 4510 28256
rect 34910 28320 35230 28321
rect 34910 28256 34918 28320
rect 34982 28256 34998 28320
rect 35062 28256 35078 28320
rect 35142 28256 35158 28320
rect 35222 28256 35230 28320
rect 34910 28255 35230 28256
rect 19550 27776 19870 27777
rect 19550 27712 19558 27776
rect 19622 27712 19638 27776
rect 19702 27712 19718 27776
rect 19782 27712 19798 27776
rect 19862 27712 19870 27776
rect 19550 27711 19870 27712
rect 50270 27776 50590 27777
rect 50270 27712 50278 27776
rect 50342 27712 50358 27776
rect 50422 27712 50438 27776
rect 50502 27712 50518 27776
rect 50582 27712 50590 27776
rect 50270 27711 50590 27712
rect 4190 27232 4510 27233
rect 4190 27168 4198 27232
rect 4262 27168 4278 27232
rect 4342 27168 4358 27232
rect 4422 27168 4438 27232
rect 4502 27168 4510 27232
rect 4190 27167 4510 27168
rect 34910 27232 35230 27233
rect 34910 27168 34918 27232
rect 34982 27168 34998 27232
rect 35062 27168 35078 27232
rect 35142 27168 35158 27232
rect 35222 27168 35230 27232
rect 34910 27167 35230 27168
rect 19550 26688 19870 26689
rect 19550 26624 19558 26688
rect 19622 26624 19638 26688
rect 19702 26624 19718 26688
rect 19782 26624 19798 26688
rect 19862 26624 19870 26688
rect 19550 26623 19870 26624
rect 50270 26688 50590 26689
rect 50270 26624 50278 26688
rect 50342 26624 50358 26688
rect 50422 26624 50438 26688
rect 50502 26624 50518 26688
rect 50582 26624 50590 26688
rect 50270 26623 50590 26624
rect 42591 26346 42657 26349
rect 42867 26346 42933 26349
rect 42591 26344 42933 26346
rect 42591 26288 42596 26344
rect 42652 26288 42872 26344
rect 42928 26288 42933 26344
rect 42591 26286 42933 26288
rect 42591 26283 42657 26286
rect 42867 26283 42933 26286
rect 4190 26144 4510 26145
rect 4190 26080 4198 26144
rect 4262 26080 4278 26144
rect 4342 26080 4358 26144
rect 4422 26080 4438 26144
rect 4502 26080 4510 26144
rect 4190 26079 4510 26080
rect 34910 26144 35230 26145
rect 34910 26080 34918 26144
rect 34982 26080 34998 26144
rect 35062 26080 35078 26144
rect 35142 26080 35158 26144
rect 35222 26080 35230 26144
rect 34910 26079 35230 26080
rect 19550 25600 19870 25601
rect 19550 25536 19558 25600
rect 19622 25536 19638 25600
rect 19702 25536 19718 25600
rect 19782 25536 19798 25600
rect 19862 25536 19870 25600
rect 19550 25535 19870 25536
rect 50270 25600 50590 25601
rect 50270 25536 50278 25600
rect 50342 25536 50358 25600
rect 50422 25536 50438 25600
rect 50502 25536 50518 25600
rect 50582 25536 50590 25600
rect 50270 25535 50590 25536
rect 4190 25056 4510 25057
rect 4190 24992 4198 25056
rect 4262 24992 4278 25056
rect 4342 24992 4358 25056
rect 4422 24992 4438 25056
rect 4502 24992 4510 25056
rect 4190 24991 4510 24992
rect 34910 25056 35230 25057
rect 34910 24992 34918 25056
rect 34982 24992 34998 25056
rect 35062 24992 35078 25056
rect 35142 24992 35158 25056
rect 35222 24992 35230 25056
rect 34910 24991 35230 24992
rect 19550 24512 19870 24513
rect 19550 24448 19558 24512
rect 19622 24448 19638 24512
rect 19702 24448 19718 24512
rect 19782 24448 19798 24512
rect 19862 24448 19870 24512
rect 19550 24447 19870 24448
rect 50270 24512 50590 24513
rect 50270 24448 50278 24512
rect 50342 24448 50358 24512
rect 50422 24448 50438 24512
rect 50502 24448 50518 24512
rect 50582 24448 50590 24512
rect 50270 24447 50590 24448
rect 4190 23968 4510 23969
rect 4190 23904 4198 23968
rect 4262 23904 4278 23968
rect 4342 23904 4358 23968
rect 4422 23904 4438 23968
rect 4502 23904 4510 23968
rect 4190 23903 4510 23904
rect 34910 23968 35230 23969
rect 34910 23904 34918 23968
rect 34982 23904 34998 23968
rect 35062 23904 35078 23968
rect 35142 23904 35158 23968
rect 35222 23904 35230 23968
rect 34910 23903 35230 23904
rect 8459 23626 8525 23629
rect 11771 23626 11837 23629
rect 8459 23624 11837 23626
rect 8459 23568 8464 23624
rect 8520 23568 11776 23624
rect 11832 23568 11837 23624
rect 8459 23566 11837 23568
rect 8459 23563 8525 23566
rect 11771 23563 11837 23566
rect 19550 23424 19870 23425
rect 19550 23360 19558 23424
rect 19622 23360 19638 23424
rect 19702 23360 19718 23424
rect 19782 23360 19798 23424
rect 19862 23360 19870 23424
rect 19550 23359 19870 23360
rect 50270 23424 50590 23425
rect 50270 23360 50278 23424
rect 50342 23360 50358 23424
rect 50422 23360 50438 23424
rect 50502 23360 50518 23424
rect 50582 23360 50590 23424
rect 50270 23359 50590 23360
rect 4190 22880 4510 22881
rect 4190 22816 4198 22880
rect 4262 22816 4278 22880
rect 4342 22816 4358 22880
rect 4422 22816 4438 22880
rect 4502 22816 4510 22880
rect 4190 22815 4510 22816
rect 34910 22880 35230 22881
rect 34910 22816 34918 22880
rect 34982 22816 34998 22880
rect 35062 22816 35078 22880
rect 35142 22816 35158 22880
rect 35222 22816 35230 22880
rect 34910 22815 35230 22816
rect 19550 22336 19870 22337
rect 19550 22272 19558 22336
rect 19622 22272 19638 22336
rect 19702 22272 19718 22336
rect 19782 22272 19798 22336
rect 19862 22272 19870 22336
rect 19550 22271 19870 22272
rect 50270 22336 50590 22337
rect 50270 22272 50278 22336
rect 50342 22272 50358 22336
rect 50422 22272 50438 22336
rect 50502 22272 50518 22336
rect 50582 22272 50590 22336
rect 50270 22271 50590 22272
rect 4190 21792 4510 21793
rect 4190 21728 4198 21792
rect 4262 21728 4278 21792
rect 4342 21728 4358 21792
rect 4422 21728 4438 21792
rect 4502 21728 4510 21792
rect 4190 21727 4510 21728
rect 34910 21792 35230 21793
rect 34910 21728 34918 21792
rect 34982 21728 34998 21792
rect 35062 21728 35078 21792
rect 35142 21728 35158 21792
rect 35222 21728 35230 21792
rect 34910 21727 35230 21728
rect 19550 21248 19870 21249
rect 19550 21184 19558 21248
rect 19622 21184 19638 21248
rect 19702 21184 19718 21248
rect 19782 21184 19798 21248
rect 19862 21184 19870 21248
rect 19550 21183 19870 21184
rect 50270 21248 50590 21249
rect 50270 21184 50278 21248
rect 50342 21184 50358 21248
rect 50422 21184 50438 21248
rect 50502 21184 50518 21248
rect 50582 21184 50590 21248
rect 50270 21183 50590 21184
rect 4190 20704 4510 20705
rect 4190 20640 4198 20704
rect 4262 20640 4278 20704
rect 4342 20640 4358 20704
rect 4422 20640 4438 20704
rect 4502 20640 4510 20704
rect 4190 20639 4510 20640
rect 34910 20704 35230 20705
rect 34910 20640 34918 20704
rect 34982 20640 34998 20704
rect 35062 20640 35078 20704
rect 35142 20640 35158 20704
rect 35222 20640 35230 20704
rect 34910 20639 35230 20640
rect 19550 20160 19870 20161
rect 19550 20096 19558 20160
rect 19622 20096 19638 20160
rect 19702 20096 19718 20160
rect 19782 20096 19798 20160
rect 19862 20096 19870 20160
rect 19550 20095 19870 20096
rect 50270 20160 50590 20161
rect 50270 20096 50278 20160
rect 50342 20096 50358 20160
rect 50422 20096 50438 20160
rect 50502 20096 50518 20160
rect 50582 20096 50590 20160
rect 50270 20095 50590 20096
rect 4190 19616 4510 19617
rect 4190 19552 4198 19616
rect 4262 19552 4278 19616
rect 4342 19552 4358 19616
rect 4422 19552 4438 19616
rect 4502 19552 4510 19616
rect 4190 19551 4510 19552
rect 34910 19616 35230 19617
rect 34910 19552 34918 19616
rect 34982 19552 34998 19616
rect 35062 19552 35078 19616
rect 35142 19552 35158 19616
rect 35222 19552 35230 19616
rect 34910 19551 35230 19552
rect 7999 19274 8065 19277
rect 8919 19274 8985 19277
rect 7999 19272 8985 19274
rect 7999 19216 8004 19272
rect 8060 19216 8924 19272
rect 8980 19216 8985 19272
rect 7999 19214 8985 19216
rect 7999 19211 8065 19214
rect 8919 19211 8985 19214
rect 19550 19072 19870 19073
rect 19550 19008 19558 19072
rect 19622 19008 19638 19072
rect 19702 19008 19718 19072
rect 19782 19008 19798 19072
rect 19862 19008 19870 19072
rect 19550 19007 19870 19008
rect 50270 19072 50590 19073
rect 50270 19008 50278 19072
rect 50342 19008 50358 19072
rect 50422 19008 50438 19072
rect 50502 19008 50518 19072
rect 50582 19008 50590 19072
rect 50270 19007 50590 19008
rect 4190 18528 4510 18529
rect 4190 18464 4198 18528
rect 4262 18464 4278 18528
rect 4342 18464 4358 18528
rect 4422 18464 4438 18528
rect 4502 18464 4510 18528
rect 4190 18463 4510 18464
rect 34910 18528 35230 18529
rect 34910 18464 34918 18528
rect 34982 18464 34998 18528
rect 35062 18464 35078 18528
rect 35142 18464 35158 18528
rect 35222 18464 35230 18528
rect 34910 18463 35230 18464
rect 8827 18458 8893 18461
rect 9011 18458 9077 18461
rect 8827 18456 9077 18458
rect 8827 18400 8832 18456
rect 8888 18400 9016 18456
rect 9072 18400 9077 18456
rect 8827 18398 9077 18400
rect 8827 18395 8893 18398
rect 9011 18395 9077 18398
rect 3399 18186 3465 18189
rect 3399 18184 3784 18186
rect 3399 18128 3404 18184
rect 3460 18128 3784 18184
rect 3399 18126 3784 18128
rect 3399 18123 3465 18126
rect 3583 18050 3649 18053
rect 3724 18050 3784 18126
rect 3583 18048 3784 18050
rect 3583 17992 3588 18048
rect 3644 17992 3784 18048
rect 3583 17990 3784 17992
rect 5239 18050 5305 18053
rect 5423 18050 5489 18053
rect 25847 18050 25913 18053
rect 5239 18048 5489 18050
rect 5239 17992 5244 18048
rect 5300 17992 5428 18048
rect 5484 17992 5489 18048
rect 5239 17990 5489 17992
rect 3583 17987 3649 17990
rect 5239 17987 5305 17990
rect 5423 17987 5489 17990
rect 25804 18048 25913 18050
rect 25804 17992 25852 18048
rect 25908 17992 25913 18048
rect 25804 17987 25913 17992
rect 19550 17984 19870 17985
rect 19550 17920 19558 17984
rect 19622 17920 19638 17984
rect 19702 17920 19718 17984
rect 19782 17920 19798 17984
rect 19862 17920 19870 17984
rect 19550 17919 19870 17920
rect 25804 17917 25864 17987
rect 50270 17984 50590 17985
rect 50270 17920 50278 17984
rect 50342 17920 50358 17984
rect 50422 17920 50438 17984
rect 50502 17920 50518 17984
rect 50582 17920 50590 17984
rect 50270 17919 50590 17920
rect 25804 17912 25913 17917
rect 25804 17856 25852 17912
rect 25908 17856 25913 17912
rect 25804 17854 25913 17856
rect 25847 17851 25913 17854
rect 4190 17440 4510 17441
rect 4190 17376 4198 17440
rect 4262 17376 4278 17440
rect 4342 17376 4358 17440
rect 4422 17376 4438 17440
rect 4502 17376 4510 17440
rect 4190 17375 4510 17376
rect 34910 17440 35230 17441
rect 34910 17376 34918 17440
rect 34982 17376 34998 17440
rect 35062 17376 35078 17440
rect 35142 17376 35158 17440
rect 35222 17376 35230 17440
rect 34910 17375 35230 17376
rect 9103 17234 9169 17237
rect 9563 17234 9629 17237
rect 9103 17232 9629 17234
rect 9103 17176 9108 17232
rect 9164 17176 9568 17232
rect 9624 17176 9629 17232
rect 9103 17174 9629 17176
rect 9103 17171 9169 17174
rect 9563 17171 9629 17174
rect 19550 16896 19870 16897
rect 19550 16832 19558 16896
rect 19622 16832 19638 16896
rect 19702 16832 19718 16896
rect 19782 16832 19798 16896
rect 19862 16832 19870 16896
rect 19550 16831 19870 16832
rect 50270 16896 50590 16897
rect 50270 16832 50278 16896
rect 50342 16832 50358 16896
rect 50422 16832 50438 16896
rect 50502 16832 50518 16896
rect 50582 16832 50590 16896
rect 50270 16831 50590 16832
rect 4190 16352 4510 16353
rect 4190 16288 4198 16352
rect 4262 16288 4278 16352
rect 4342 16288 4358 16352
rect 4422 16288 4438 16352
rect 4502 16288 4510 16352
rect 4190 16287 4510 16288
rect 34910 16352 35230 16353
rect 34910 16288 34918 16352
rect 34982 16288 34998 16352
rect 35062 16288 35078 16352
rect 35142 16288 35158 16352
rect 35222 16288 35230 16352
rect 34910 16287 35230 16288
rect 19550 15808 19870 15809
rect 19550 15744 19558 15808
rect 19622 15744 19638 15808
rect 19702 15744 19718 15808
rect 19782 15744 19798 15808
rect 19862 15744 19870 15808
rect 19550 15743 19870 15744
rect 50270 15808 50590 15809
rect 50270 15744 50278 15808
rect 50342 15744 50358 15808
rect 50422 15744 50438 15808
rect 50502 15744 50518 15808
rect 50582 15744 50590 15808
rect 50270 15743 50590 15744
rect 4190 15264 4510 15265
rect 4190 15200 4198 15264
rect 4262 15200 4278 15264
rect 4342 15200 4358 15264
rect 4422 15200 4438 15264
rect 4502 15200 4510 15264
rect 4190 15199 4510 15200
rect 34910 15264 35230 15265
rect 34910 15200 34918 15264
rect 34982 15200 34998 15264
rect 35062 15200 35078 15264
rect 35142 15200 35158 15264
rect 35222 15200 35230 15264
rect 34910 15199 35230 15200
rect 8275 14922 8341 14925
rect 8643 14922 8709 14925
rect 8275 14920 8709 14922
rect 8275 14864 8280 14920
rect 8336 14864 8648 14920
rect 8704 14864 8709 14920
rect 8275 14862 8709 14864
rect 8275 14859 8341 14862
rect 8643 14859 8709 14862
rect 19550 14720 19870 14721
rect 19550 14656 19558 14720
rect 19622 14656 19638 14720
rect 19702 14656 19718 14720
rect 19782 14656 19798 14720
rect 19862 14656 19870 14720
rect 19550 14655 19870 14656
rect 50270 14720 50590 14721
rect 50270 14656 50278 14720
rect 50342 14656 50358 14720
rect 50422 14656 50438 14720
rect 50502 14656 50518 14720
rect 50582 14656 50590 14720
rect 50270 14655 50590 14656
rect 4190 14176 4510 14177
rect 4190 14112 4198 14176
rect 4262 14112 4278 14176
rect 4342 14112 4358 14176
rect 4422 14112 4438 14176
rect 4502 14112 4510 14176
rect 4190 14111 4510 14112
rect 34910 14176 35230 14177
rect 34910 14112 34918 14176
rect 34982 14112 34998 14176
rect 35062 14112 35078 14176
rect 35142 14112 35158 14176
rect 35222 14112 35230 14176
rect 34910 14111 35230 14112
rect 7999 13970 8065 13973
rect 8827 13970 8893 13973
rect 7999 13968 8893 13970
rect 7999 13912 8004 13968
rect 8060 13912 8832 13968
rect 8888 13912 8893 13968
rect 7999 13910 8893 13912
rect 7999 13907 8065 13910
rect 8827 13907 8893 13910
rect 19550 13632 19870 13633
rect 19550 13568 19558 13632
rect 19622 13568 19638 13632
rect 19702 13568 19718 13632
rect 19782 13568 19798 13632
rect 19862 13568 19870 13632
rect 19550 13567 19870 13568
rect 50270 13632 50590 13633
rect 50270 13568 50278 13632
rect 50342 13568 50358 13632
rect 50422 13568 50438 13632
rect 50502 13568 50518 13632
rect 50582 13568 50590 13632
rect 50270 13567 50590 13568
rect 4190 13088 4510 13089
rect 4190 13024 4198 13088
rect 4262 13024 4278 13088
rect 4342 13024 4358 13088
rect 4422 13024 4438 13088
rect 4502 13024 4510 13088
rect 4190 13023 4510 13024
rect 34910 13088 35230 13089
rect 34910 13024 34918 13088
rect 34982 13024 34998 13088
rect 35062 13024 35078 13088
rect 35142 13024 35158 13088
rect 35222 13024 35230 13088
rect 34910 13023 35230 13024
rect 19550 12544 19870 12545
rect 19550 12480 19558 12544
rect 19622 12480 19638 12544
rect 19702 12480 19718 12544
rect 19782 12480 19798 12544
rect 19862 12480 19870 12544
rect 19550 12479 19870 12480
rect 50270 12544 50590 12545
rect 50270 12480 50278 12544
rect 50342 12480 50358 12544
rect 50422 12480 50438 12544
rect 50502 12480 50518 12544
rect 50582 12480 50590 12544
rect 50270 12479 50590 12480
rect 4190 12000 4510 12001
rect 4190 11936 4198 12000
rect 4262 11936 4278 12000
rect 4342 11936 4358 12000
rect 4422 11936 4438 12000
rect 4502 11936 4510 12000
rect 4190 11935 4510 11936
rect 34910 12000 35230 12001
rect 34910 11936 34918 12000
rect 34982 11936 34998 12000
rect 35062 11936 35078 12000
rect 35142 11936 35158 12000
rect 35222 11936 35230 12000
rect 34910 11935 35230 11936
rect 19550 11456 19870 11457
rect 19550 11392 19558 11456
rect 19622 11392 19638 11456
rect 19702 11392 19718 11456
rect 19782 11392 19798 11456
rect 19862 11392 19870 11456
rect 19550 11391 19870 11392
rect 50270 11456 50590 11457
rect 50270 11392 50278 11456
rect 50342 11392 50358 11456
rect 50422 11392 50438 11456
rect 50502 11392 50518 11456
rect 50582 11392 50590 11456
rect 50270 11391 50590 11392
rect 4190 10912 4510 10913
rect 4190 10848 4198 10912
rect 4262 10848 4278 10912
rect 4342 10848 4358 10912
rect 4422 10848 4438 10912
rect 4502 10848 4510 10912
rect 4190 10847 4510 10848
rect 34910 10912 35230 10913
rect 34910 10848 34918 10912
rect 34982 10848 34998 10912
rect 35062 10848 35078 10912
rect 35142 10848 35158 10912
rect 35222 10848 35230 10912
rect 34910 10847 35230 10848
rect 19550 10368 19870 10369
rect 19550 10304 19558 10368
rect 19622 10304 19638 10368
rect 19702 10304 19718 10368
rect 19782 10304 19798 10368
rect 19862 10304 19870 10368
rect 19550 10303 19870 10304
rect 50270 10368 50590 10369
rect 50270 10304 50278 10368
rect 50342 10304 50358 10368
rect 50422 10304 50438 10368
rect 50502 10304 50518 10368
rect 50582 10304 50590 10368
rect 50270 10303 50590 10304
rect 4190 9824 4510 9825
rect 4190 9760 4198 9824
rect 4262 9760 4278 9824
rect 4342 9760 4358 9824
rect 4422 9760 4438 9824
rect 4502 9760 4510 9824
rect 4190 9759 4510 9760
rect 34910 9824 35230 9825
rect 34910 9760 34918 9824
rect 34982 9760 34998 9824
rect 35062 9760 35078 9824
rect 35142 9760 35158 9824
rect 35222 9760 35230 9824
rect 34910 9759 35230 9760
rect 19550 9280 19870 9281
rect 19550 9216 19558 9280
rect 19622 9216 19638 9280
rect 19702 9216 19718 9280
rect 19782 9216 19798 9280
rect 19862 9216 19870 9280
rect 19550 9215 19870 9216
rect 50270 9280 50590 9281
rect 50270 9216 50278 9280
rect 50342 9216 50358 9280
rect 50422 9216 50438 9280
rect 50502 9216 50518 9280
rect 50582 9216 50590 9280
rect 50270 9215 50590 9216
rect 4190 8736 4510 8737
rect 4190 8672 4198 8736
rect 4262 8672 4278 8736
rect 4342 8672 4358 8736
rect 4422 8672 4438 8736
rect 4502 8672 4510 8736
rect 4190 8671 4510 8672
rect 34910 8736 35230 8737
rect 34910 8672 34918 8736
rect 34982 8672 34998 8736
rect 35062 8672 35078 8736
rect 35142 8672 35158 8736
rect 35222 8672 35230 8736
rect 34910 8671 35230 8672
rect 19550 8192 19870 8193
rect 19550 8128 19558 8192
rect 19622 8128 19638 8192
rect 19702 8128 19718 8192
rect 19782 8128 19798 8192
rect 19862 8128 19870 8192
rect 19550 8127 19870 8128
rect 50270 8192 50590 8193
rect 50270 8128 50278 8192
rect 50342 8128 50358 8192
rect 50422 8128 50438 8192
rect 50502 8128 50518 8192
rect 50582 8128 50590 8192
rect 50270 8127 50590 8128
rect 4190 7648 4510 7649
rect 4190 7584 4198 7648
rect 4262 7584 4278 7648
rect 4342 7584 4358 7648
rect 4422 7584 4438 7648
rect 4502 7584 4510 7648
rect 4190 7583 4510 7584
rect 34910 7648 35230 7649
rect 34910 7584 34918 7648
rect 34982 7584 34998 7648
rect 35062 7584 35078 7648
rect 35142 7584 35158 7648
rect 35222 7584 35230 7648
rect 34910 7583 35230 7584
rect 8229 7306 8295 7309
rect 12691 7306 12757 7309
rect 8229 7304 12757 7306
rect 8229 7248 8234 7304
rect 8290 7248 12696 7304
rect 12752 7248 12757 7304
rect 8229 7246 12757 7248
rect 8229 7243 8295 7246
rect 12691 7243 12757 7246
rect 19550 7104 19870 7105
rect 19550 7040 19558 7104
rect 19622 7040 19638 7104
rect 19702 7040 19718 7104
rect 19782 7040 19798 7104
rect 19862 7040 19870 7104
rect 19550 7039 19870 7040
rect 50270 7104 50590 7105
rect 50270 7040 50278 7104
rect 50342 7040 50358 7104
rect 50422 7040 50438 7104
rect 50502 7040 50518 7104
rect 50582 7040 50590 7104
rect 50270 7039 50590 7040
rect 4190 6560 4510 6561
rect 4190 6496 4198 6560
rect 4262 6496 4278 6560
rect 4342 6496 4358 6560
rect 4422 6496 4438 6560
rect 4502 6496 4510 6560
rect 4190 6495 4510 6496
rect 34910 6560 35230 6561
rect 34910 6496 34918 6560
rect 34982 6496 34998 6560
rect 35062 6496 35078 6560
rect 35142 6496 35158 6560
rect 35222 6496 35230 6560
rect 34910 6495 35230 6496
rect 19550 6016 19870 6017
rect 19550 5952 19558 6016
rect 19622 5952 19638 6016
rect 19702 5952 19718 6016
rect 19782 5952 19798 6016
rect 19862 5952 19870 6016
rect 19550 5951 19870 5952
rect 50270 6016 50590 6017
rect 50270 5952 50278 6016
rect 50342 5952 50358 6016
rect 50422 5952 50438 6016
rect 50502 5952 50518 6016
rect 50582 5952 50590 6016
rect 50270 5951 50590 5952
rect 4190 5472 4510 5473
rect 4190 5408 4198 5472
rect 4262 5408 4278 5472
rect 4342 5408 4358 5472
rect 4422 5408 4438 5472
rect 4502 5408 4510 5472
rect 4190 5407 4510 5408
rect 34910 5472 35230 5473
rect 34910 5408 34918 5472
rect 34982 5408 34998 5472
rect 35062 5408 35078 5472
rect 35142 5408 35158 5472
rect 35222 5408 35230 5472
rect 34910 5407 35230 5408
rect 19550 4928 19870 4929
rect 19550 4864 19558 4928
rect 19622 4864 19638 4928
rect 19702 4864 19718 4928
rect 19782 4864 19798 4928
rect 19862 4864 19870 4928
rect 19550 4863 19870 4864
rect 50270 4928 50590 4929
rect 50270 4864 50278 4928
rect 50342 4864 50358 4928
rect 50422 4864 50438 4928
rect 50502 4864 50518 4928
rect 50582 4864 50590 4928
rect 50270 4863 50590 4864
rect 4190 4384 4510 4385
rect 4190 4320 4198 4384
rect 4262 4320 4278 4384
rect 4342 4320 4358 4384
rect 4422 4320 4438 4384
rect 4502 4320 4510 4384
rect 4190 4319 4510 4320
rect 34910 4384 35230 4385
rect 34910 4320 34918 4384
rect 34982 4320 34998 4384
rect 35062 4320 35078 4384
rect 35142 4320 35158 4384
rect 35222 4320 35230 4384
rect 34910 4319 35230 4320
rect 19550 3840 19870 3841
rect 19550 3776 19558 3840
rect 19622 3776 19638 3840
rect 19702 3776 19718 3840
rect 19782 3776 19798 3840
rect 19862 3776 19870 3840
rect 19550 3775 19870 3776
rect 50270 3840 50590 3841
rect 50270 3776 50278 3840
rect 50342 3776 50358 3840
rect 50422 3776 50438 3840
rect 50502 3776 50518 3840
rect 50582 3776 50590 3840
rect 50270 3775 50590 3776
rect 45903 3770 45969 3773
rect 46915 3770 46981 3773
rect 45903 3768 46981 3770
rect 45903 3712 45908 3768
rect 45964 3712 46920 3768
rect 46976 3712 46981 3768
rect 45903 3710 46981 3712
rect 45903 3707 45969 3710
rect 46915 3707 46981 3710
rect 4190 3296 4510 3297
rect 4190 3232 4198 3296
rect 4262 3232 4278 3296
rect 4342 3232 4358 3296
rect 4422 3232 4438 3296
rect 4502 3232 4510 3296
rect 4190 3231 4510 3232
rect 34910 3296 35230 3297
rect 34910 3232 34918 3296
rect 34982 3232 34998 3296
rect 35062 3232 35078 3296
rect 35142 3232 35158 3296
rect 35222 3232 35230 3296
rect 34910 3231 35230 3232
rect 41303 2954 41369 2957
rect 41487 2954 41553 2957
rect 41303 2952 41553 2954
rect 41303 2896 41308 2952
rect 41364 2896 41492 2952
rect 41548 2896 41553 2952
rect 41303 2894 41553 2896
rect 41303 2891 41369 2894
rect 41487 2891 41553 2894
rect 36335 2818 36401 2821
rect 41303 2818 41369 2821
rect 36335 2816 41369 2818
rect 36335 2760 36340 2816
rect 36396 2760 41308 2816
rect 41364 2760 41369 2816
rect 36335 2758 41369 2760
rect 36335 2755 36401 2758
rect 41303 2755 41369 2758
rect 19550 2752 19870 2753
rect 19550 2688 19558 2752
rect 19622 2688 19638 2752
rect 19702 2688 19718 2752
rect 19782 2688 19798 2752
rect 19862 2688 19870 2752
rect 19550 2687 19870 2688
rect 50270 2752 50590 2753
rect 50270 2688 50278 2752
rect 50342 2688 50358 2752
rect 50422 2688 50438 2752
rect 50502 2688 50518 2752
rect 50582 2688 50590 2752
rect 50270 2687 50590 2688
rect 4190 2208 4510 2209
rect 4190 2144 4198 2208
rect 4262 2144 4278 2208
rect 4342 2144 4358 2208
rect 4422 2144 4438 2208
rect 4502 2144 4510 2208
rect 4190 2143 4510 2144
rect 34910 2208 35230 2209
rect 34910 2144 34918 2208
rect 34982 2144 34998 2208
rect 35062 2144 35078 2208
rect 35142 2144 35158 2208
rect 35222 2144 35230 2208
rect 34910 2143 35230 2144
rect 36887 914 36953 917
rect 37163 914 37229 917
rect 36887 912 37229 914
rect 36887 856 36892 912
rect 36948 856 37168 912
rect 37224 856 37229 912
rect 36887 854 37229 856
rect 36887 851 36953 854
rect 37163 851 37229 854
<< via3 >>
rect 4198 57692 4262 57696
rect 4198 57636 4202 57692
rect 4202 57636 4258 57692
rect 4258 57636 4262 57692
rect 4198 57632 4262 57636
rect 4278 57692 4342 57696
rect 4278 57636 4282 57692
rect 4282 57636 4338 57692
rect 4338 57636 4342 57692
rect 4278 57632 4342 57636
rect 4358 57692 4422 57696
rect 4358 57636 4362 57692
rect 4362 57636 4418 57692
rect 4418 57636 4422 57692
rect 4358 57632 4422 57636
rect 4438 57692 4502 57696
rect 4438 57636 4442 57692
rect 4442 57636 4498 57692
rect 4498 57636 4502 57692
rect 4438 57632 4502 57636
rect 34918 57692 34982 57696
rect 34918 57636 34922 57692
rect 34922 57636 34978 57692
rect 34978 57636 34982 57692
rect 34918 57632 34982 57636
rect 34998 57692 35062 57696
rect 34998 57636 35002 57692
rect 35002 57636 35058 57692
rect 35058 57636 35062 57692
rect 34998 57632 35062 57636
rect 35078 57692 35142 57696
rect 35078 57636 35082 57692
rect 35082 57636 35138 57692
rect 35138 57636 35142 57692
rect 35078 57632 35142 57636
rect 35158 57692 35222 57696
rect 35158 57636 35162 57692
rect 35162 57636 35218 57692
rect 35218 57636 35222 57692
rect 35158 57632 35222 57636
rect 19558 57148 19622 57152
rect 19558 57092 19562 57148
rect 19562 57092 19618 57148
rect 19618 57092 19622 57148
rect 19558 57088 19622 57092
rect 19638 57148 19702 57152
rect 19638 57092 19642 57148
rect 19642 57092 19698 57148
rect 19698 57092 19702 57148
rect 19638 57088 19702 57092
rect 19718 57148 19782 57152
rect 19718 57092 19722 57148
rect 19722 57092 19778 57148
rect 19778 57092 19782 57148
rect 19718 57088 19782 57092
rect 19798 57148 19862 57152
rect 19798 57092 19802 57148
rect 19802 57092 19858 57148
rect 19858 57092 19862 57148
rect 19798 57088 19862 57092
rect 50278 57148 50342 57152
rect 50278 57092 50282 57148
rect 50282 57092 50338 57148
rect 50338 57092 50342 57148
rect 50278 57088 50342 57092
rect 50358 57148 50422 57152
rect 50358 57092 50362 57148
rect 50362 57092 50418 57148
rect 50418 57092 50422 57148
rect 50358 57088 50422 57092
rect 50438 57148 50502 57152
rect 50438 57092 50442 57148
rect 50442 57092 50498 57148
rect 50498 57092 50502 57148
rect 50438 57088 50502 57092
rect 50518 57148 50582 57152
rect 50518 57092 50522 57148
rect 50522 57092 50578 57148
rect 50578 57092 50582 57148
rect 50518 57088 50582 57092
rect 4198 56604 4262 56608
rect 4198 56548 4202 56604
rect 4202 56548 4258 56604
rect 4258 56548 4262 56604
rect 4198 56544 4262 56548
rect 4278 56604 4342 56608
rect 4278 56548 4282 56604
rect 4282 56548 4338 56604
rect 4338 56548 4342 56604
rect 4278 56544 4342 56548
rect 4358 56604 4422 56608
rect 4358 56548 4362 56604
rect 4362 56548 4418 56604
rect 4418 56548 4422 56604
rect 4358 56544 4422 56548
rect 4438 56604 4502 56608
rect 4438 56548 4442 56604
rect 4442 56548 4498 56604
rect 4498 56548 4502 56604
rect 4438 56544 4502 56548
rect 34918 56604 34982 56608
rect 34918 56548 34922 56604
rect 34922 56548 34978 56604
rect 34978 56548 34982 56604
rect 34918 56544 34982 56548
rect 34998 56604 35062 56608
rect 34998 56548 35002 56604
rect 35002 56548 35058 56604
rect 35058 56548 35062 56604
rect 34998 56544 35062 56548
rect 35078 56604 35142 56608
rect 35078 56548 35082 56604
rect 35082 56548 35138 56604
rect 35138 56548 35142 56604
rect 35078 56544 35142 56548
rect 35158 56604 35222 56608
rect 35158 56548 35162 56604
rect 35162 56548 35218 56604
rect 35218 56548 35222 56604
rect 35158 56544 35222 56548
rect 19558 56060 19622 56064
rect 19558 56004 19562 56060
rect 19562 56004 19618 56060
rect 19618 56004 19622 56060
rect 19558 56000 19622 56004
rect 19638 56060 19702 56064
rect 19638 56004 19642 56060
rect 19642 56004 19698 56060
rect 19698 56004 19702 56060
rect 19638 56000 19702 56004
rect 19718 56060 19782 56064
rect 19718 56004 19722 56060
rect 19722 56004 19778 56060
rect 19778 56004 19782 56060
rect 19718 56000 19782 56004
rect 19798 56060 19862 56064
rect 19798 56004 19802 56060
rect 19802 56004 19858 56060
rect 19858 56004 19862 56060
rect 19798 56000 19862 56004
rect 50278 56060 50342 56064
rect 50278 56004 50282 56060
rect 50282 56004 50338 56060
rect 50338 56004 50342 56060
rect 50278 56000 50342 56004
rect 50358 56060 50422 56064
rect 50358 56004 50362 56060
rect 50362 56004 50418 56060
rect 50418 56004 50422 56060
rect 50358 56000 50422 56004
rect 50438 56060 50502 56064
rect 50438 56004 50442 56060
rect 50442 56004 50498 56060
rect 50498 56004 50502 56060
rect 50438 56000 50502 56004
rect 50518 56060 50582 56064
rect 50518 56004 50522 56060
rect 50522 56004 50578 56060
rect 50578 56004 50582 56060
rect 50518 56000 50582 56004
rect 4198 55516 4262 55520
rect 4198 55460 4202 55516
rect 4202 55460 4258 55516
rect 4258 55460 4262 55516
rect 4198 55456 4262 55460
rect 4278 55516 4342 55520
rect 4278 55460 4282 55516
rect 4282 55460 4338 55516
rect 4338 55460 4342 55516
rect 4278 55456 4342 55460
rect 4358 55516 4422 55520
rect 4358 55460 4362 55516
rect 4362 55460 4418 55516
rect 4418 55460 4422 55516
rect 4358 55456 4422 55460
rect 4438 55516 4502 55520
rect 4438 55460 4442 55516
rect 4442 55460 4498 55516
rect 4498 55460 4502 55516
rect 4438 55456 4502 55460
rect 34918 55516 34982 55520
rect 34918 55460 34922 55516
rect 34922 55460 34978 55516
rect 34978 55460 34982 55516
rect 34918 55456 34982 55460
rect 34998 55516 35062 55520
rect 34998 55460 35002 55516
rect 35002 55460 35058 55516
rect 35058 55460 35062 55516
rect 34998 55456 35062 55460
rect 35078 55516 35142 55520
rect 35078 55460 35082 55516
rect 35082 55460 35138 55516
rect 35138 55460 35142 55516
rect 35078 55456 35142 55460
rect 35158 55516 35222 55520
rect 35158 55460 35162 55516
rect 35162 55460 35218 55516
rect 35218 55460 35222 55516
rect 35158 55456 35222 55460
rect 19558 54972 19622 54976
rect 19558 54916 19562 54972
rect 19562 54916 19618 54972
rect 19618 54916 19622 54972
rect 19558 54912 19622 54916
rect 19638 54972 19702 54976
rect 19638 54916 19642 54972
rect 19642 54916 19698 54972
rect 19698 54916 19702 54972
rect 19638 54912 19702 54916
rect 19718 54972 19782 54976
rect 19718 54916 19722 54972
rect 19722 54916 19778 54972
rect 19778 54916 19782 54972
rect 19718 54912 19782 54916
rect 19798 54972 19862 54976
rect 19798 54916 19802 54972
rect 19802 54916 19858 54972
rect 19858 54916 19862 54972
rect 19798 54912 19862 54916
rect 50278 54972 50342 54976
rect 50278 54916 50282 54972
rect 50282 54916 50338 54972
rect 50338 54916 50342 54972
rect 50278 54912 50342 54916
rect 50358 54972 50422 54976
rect 50358 54916 50362 54972
rect 50362 54916 50418 54972
rect 50418 54916 50422 54972
rect 50358 54912 50422 54916
rect 50438 54972 50502 54976
rect 50438 54916 50442 54972
rect 50442 54916 50498 54972
rect 50498 54916 50502 54972
rect 50438 54912 50502 54916
rect 50518 54972 50582 54976
rect 50518 54916 50522 54972
rect 50522 54916 50578 54972
rect 50578 54916 50582 54972
rect 50518 54912 50582 54916
rect 4198 54428 4262 54432
rect 4198 54372 4202 54428
rect 4202 54372 4258 54428
rect 4258 54372 4262 54428
rect 4198 54368 4262 54372
rect 4278 54428 4342 54432
rect 4278 54372 4282 54428
rect 4282 54372 4338 54428
rect 4338 54372 4342 54428
rect 4278 54368 4342 54372
rect 4358 54428 4422 54432
rect 4358 54372 4362 54428
rect 4362 54372 4418 54428
rect 4418 54372 4422 54428
rect 4358 54368 4422 54372
rect 4438 54428 4502 54432
rect 4438 54372 4442 54428
rect 4442 54372 4498 54428
rect 4498 54372 4502 54428
rect 4438 54368 4502 54372
rect 34918 54428 34982 54432
rect 34918 54372 34922 54428
rect 34922 54372 34978 54428
rect 34978 54372 34982 54428
rect 34918 54368 34982 54372
rect 34998 54428 35062 54432
rect 34998 54372 35002 54428
rect 35002 54372 35058 54428
rect 35058 54372 35062 54428
rect 34998 54368 35062 54372
rect 35078 54428 35142 54432
rect 35078 54372 35082 54428
rect 35082 54372 35138 54428
rect 35138 54372 35142 54428
rect 35078 54368 35142 54372
rect 35158 54428 35222 54432
rect 35158 54372 35162 54428
rect 35162 54372 35218 54428
rect 35218 54372 35222 54428
rect 35158 54368 35222 54372
rect 19558 53884 19622 53888
rect 19558 53828 19562 53884
rect 19562 53828 19618 53884
rect 19618 53828 19622 53884
rect 19558 53824 19622 53828
rect 19638 53884 19702 53888
rect 19638 53828 19642 53884
rect 19642 53828 19698 53884
rect 19698 53828 19702 53884
rect 19638 53824 19702 53828
rect 19718 53884 19782 53888
rect 19718 53828 19722 53884
rect 19722 53828 19778 53884
rect 19778 53828 19782 53884
rect 19718 53824 19782 53828
rect 19798 53884 19862 53888
rect 19798 53828 19802 53884
rect 19802 53828 19858 53884
rect 19858 53828 19862 53884
rect 19798 53824 19862 53828
rect 50278 53884 50342 53888
rect 50278 53828 50282 53884
rect 50282 53828 50338 53884
rect 50338 53828 50342 53884
rect 50278 53824 50342 53828
rect 50358 53884 50422 53888
rect 50358 53828 50362 53884
rect 50362 53828 50418 53884
rect 50418 53828 50422 53884
rect 50358 53824 50422 53828
rect 50438 53884 50502 53888
rect 50438 53828 50442 53884
rect 50442 53828 50498 53884
rect 50498 53828 50502 53884
rect 50438 53824 50502 53828
rect 50518 53884 50582 53888
rect 50518 53828 50522 53884
rect 50522 53828 50578 53884
rect 50578 53828 50582 53884
rect 50518 53824 50582 53828
rect 4198 53340 4262 53344
rect 4198 53284 4202 53340
rect 4202 53284 4258 53340
rect 4258 53284 4262 53340
rect 4198 53280 4262 53284
rect 4278 53340 4342 53344
rect 4278 53284 4282 53340
rect 4282 53284 4338 53340
rect 4338 53284 4342 53340
rect 4278 53280 4342 53284
rect 4358 53340 4422 53344
rect 4358 53284 4362 53340
rect 4362 53284 4418 53340
rect 4418 53284 4422 53340
rect 4358 53280 4422 53284
rect 4438 53340 4502 53344
rect 4438 53284 4442 53340
rect 4442 53284 4498 53340
rect 4498 53284 4502 53340
rect 4438 53280 4502 53284
rect 34918 53340 34982 53344
rect 34918 53284 34922 53340
rect 34922 53284 34978 53340
rect 34978 53284 34982 53340
rect 34918 53280 34982 53284
rect 34998 53340 35062 53344
rect 34998 53284 35002 53340
rect 35002 53284 35058 53340
rect 35058 53284 35062 53340
rect 34998 53280 35062 53284
rect 35078 53340 35142 53344
rect 35078 53284 35082 53340
rect 35082 53284 35138 53340
rect 35138 53284 35142 53340
rect 35078 53280 35142 53284
rect 35158 53340 35222 53344
rect 35158 53284 35162 53340
rect 35162 53284 35218 53340
rect 35218 53284 35222 53340
rect 35158 53280 35222 53284
rect 19558 52796 19622 52800
rect 19558 52740 19562 52796
rect 19562 52740 19618 52796
rect 19618 52740 19622 52796
rect 19558 52736 19622 52740
rect 19638 52796 19702 52800
rect 19638 52740 19642 52796
rect 19642 52740 19698 52796
rect 19698 52740 19702 52796
rect 19638 52736 19702 52740
rect 19718 52796 19782 52800
rect 19718 52740 19722 52796
rect 19722 52740 19778 52796
rect 19778 52740 19782 52796
rect 19718 52736 19782 52740
rect 19798 52796 19862 52800
rect 19798 52740 19802 52796
rect 19802 52740 19858 52796
rect 19858 52740 19862 52796
rect 19798 52736 19862 52740
rect 50278 52796 50342 52800
rect 50278 52740 50282 52796
rect 50282 52740 50338 52796
rect 50338 52740 50342 52796
rect 50278 52736 50342 52740
rect 50358 52796 50422 52800
rect 50358 52740 50362 52796
rect 50362 52740 50418 52796
rect 50418 52740 50422 52796
rect 50358 52736 50422 52740
rect 50438 52796 50502 52800
rect 50438 52740 50442 52796
rect 50442 52740 50498 52796
rect 50498 52740 50502 52796
rect 50438 52736 50502 52740
rect 50518 52796 50582 52800
rect 50518 52740 50522 52796
rect 50522 52740 50578 52796
rect 50578 52740 50582 52796
rect 50518 52736 50582 52740
rect 4198 52252 4262 52256
rect 4198 52196 4202 52252
rect 4202 52196 4258 52252
rect 4258 52196 4262 52252
rect 4198 52192 4262 52196
rect 4278 52252 4342 52256
rect 4278 52196 4282 52252
rect 4282 52196 4338 52252
rect 4338 52196 4342 52252
rect 4278 52192 4342 52196
rect 4358 52252 4422 52256
rect 4358 52196 4362 52252
rect 4362 52196 4418 52252
rect 4418 52196 4422 52252
rect 4358 52192 4422 52196
rect 4438 52252 4502 52256
rect 4438 52196 4442 52252
rect 4442 52196 4498 52252
rect 4498 52196 4502 52252
rect 4438 52192 4502 52196
rect 34918 52252 34982 52256
rect 34918 52196 34922 52252
rect 34922 52196 34978 52252
rect 34978 52196 34982 52252
rect 34918 52192 34982 52196
rect 34998 52252 35062 52256
rect 34998 52196 35002 52252
rect 35002 52196 35058 52252
rect 35058 52196 35062 52252
rect 34998 52192 35062 52196
rect 35078 52252 35142 52256
rect 35078 52196 35082 52252
rect 35082 52196 35138 52252
rect 35138 52196 35142 52252
rect 35078 52192 35142 52196
rect 35158 52252 35222 52256
rect 35158 52196 35162 52252
rect 35162 52196 35218 52252
rect 35218 52196 35222 52252
rect 35158 52192 35222 52196
rect 19558 51708 19622 51712
rect 19558 51652 19562 51708
rect 19562 51652 19618 51708
rect 19618 51652 19622 51708
rect 19558 51648 19622 51652
rect 19638 51708 19702 51712
rect 19638 51652 19642 51708
rect 19642 51652 19698 51708
rect 19698 51652 19702 51708
rect 19638 51648 19702 51652
rect 19718 51708 19782 51712
rect 19718 51652 19722 51708
rect 19722 51652 19778 51708
rect 19778 51652 19782 51708
rect 19718 51648 19782 51652
rect 19798 51708 19862 51712
rect 19798 51652 19802 51708
rect 19802 51652 19858 51708
rect 19858 51652 19862 51708
rect 19798 51648 19862 51652
rect 50278 51708 50342 51712
rect 50278 51652 50282 51708
rect 50282 51652 50338 51708
rect 50338 51652 50342 51708
rect 50278 51648 50342 51652
rect 50358 51708 50422 51712
rect 50358 51652 50362 51708
rect 50362 51652 50418 51708
rect 50418 51652 50422 51708
rect 50358 51648 50422 51652
rect 50438 51708 50502 51712
rect 50438 51652 50442 51708
rect 50442 51652 50498 51708
rect 50498 51652 50502 51708
rect 50438 51648 50502 51652
rect 50518 51708 50582 51712
rect 50518 51652 50522 51708
rect 50522 51652 50578 51708
rect 50578 51652 50582 51708
rect 50518 51648 50582 51652
rect 4198 51164 4262 51168
rect 4198 51108 4202 51164
rect 4202 51108 4258 51164
rect 4258 51108 4262 51164
rect 4198 51104 4262 51108
rect 4278 51164 4342 51168
rect 4278 51108 4282 51164
rect 4282 51108 4338 51164
rect 4338 51108 4342 51164
rect 4278 51104 4342 51108
rect 4358 51164 4422 51168
rect 4358 51108 4362 51164
rect 4362 51108 4418 51164
rect 4418 51108 4422 51164
rect 4358 51104 4422 51108
rect 4438 51164 4502 51168
rect 4438 51108 4442 51164
rect 4442 51108 4498 51164
rect 4498 51108 4502 51164
rect 4438 51104 4502 51108
rect 34918 51164 34982 51168
rect 34918 51108 34922 51164
rect 34922 51108 34978 51164
rect 34978 51108 34982 51164
rect 34918 51104 34982 51108
rect 34998 51164 35062 51168
rect 34998 51108 35002 51164
rect 35002 51108 35058 51164
rect 35058 51108 35062 51164
rect 34998 51104 35062 51108
rect 35078 51164 35142 51168
rect 35078 51108 35082 51164
rect 35082 51108 35138 51164
rect 35138 51108 35142 51164
rect 35078 51104 35142 51108
rect 35158 51164 35222 51168
rect 35158 51108 35162 51164
rect 35162 51108 35218 51164
rect 35218 51108 35222 51164
rect 35158 51104 35222 51108
rect 19558 50620 19622 50624
rect 19558 50564 19562 50620
rect 19562 50564 19618 50620
rect 19618 50564 19622 50620
rect 19558 50560 19622 50564
rect 19638 50620 19702 50624
rect 19638 50564 19642 50620
rect 19642 50564 19698 50620
rect 19698 50564 19702 50620
rect 19638 50560 19702 50564
rect 19718 50620 19782 50624
rect 19718 50564 19722 50620
rect 19722 50564 19778 50620
rect 19778 50564 19782 50620
rect 19718 50560 19782 50564
rect 19798 50620 19862 50624
rect 19798 50564 19802 50620
rect 19802 50564 19858 50620
rect 19858 50564 19862 50620
rect 19798 50560 19862 50564
rect 50278 50620 50342 50624
rect 50278 50564 50282 50620
rect 50282 50564 50338 50620
rect 50338 50564 50342 50620
rect 50278 50560 50342 50564
rect 50358 50620 50422 50624
rect 50358 50564 50362 50620
rect 50362 50564 50418 50620
rect 50418 50564 50422 50620
rect 50358 50560 50422 50564
rect 50438 50620 50502 50624
rect 50438 50564 50442 50620
rect 50442 50564 50498 50620
rect 50498 50564 50502 50620
rect 50438 50560 50502 50564
rect 50518 50620 50582 50624
rect 50518 50564 50522 50620
rect 50522 50564 50578 50620
rect 50578 50564 50582 50620
rect 50518 50560 50582 50564
rect 4198 50076 4262 50080
rect 4198 50020 4202 50076
rect 4202 50020 4258 50076
rect 4258 50020 4262 50076
rect 4198 50016 4262 50020
rect 4278 50076 4342 50080
rect 4278 50020 4282 50076
rect 4282 50020 4338 50076
rect 4338 50020 4342 50076
rect 4278 50016 4342 50020
rect 4358 50076 4422 50080
rect 4358 50020 4362 50076
rect 4362 50020 4418 50076
rect 4418 50020 4422 50076
rect 4358 50016 4422 50020
rect 4438 50076 4502 50080
rect 4438 50020 4442 50076
rect 4442 50020 4498 50076
rect 4498 50020 4502 50076
rect 4438 50016 4502 50020
rect 34918 50076 34982 50080
rect 34918 50020 34922 50076
rect 34922 50020 34978 50076
rect 34978 50020 34982 50076
rect 34918 50016 34982 50020
rect 34998 50076 35062 50080
rect 34998 50020 35002 50076
rect 35002 50020 35058 50076
rect 35058 50020 35062 50076
rect 34998 50016 35062 50020
rect 35078 50076 35142 50080
rect 35078 50020 35082 50076
rect 35082 50020 35138 50076
rect 35138 50020 35142 50076
rect 35078 50016 35142 50020
rect 35158 50076 35222 50080
rect 35158 50020 35162 50076
rect 35162 50020 35218 50076
rect 35218 50020 35222 50076
rect 35158 50016 35222 50020
rect 19558 49532 19622 49536
rect 19558 49476 19562 49532
rect 19562 49476 19618 49532
rect 19618 49476 19622 49532
rect 19558 49472 19622 49476
rect 19638 49532 19702 49536
rect 19638 49476 19642 49532
rect 19642 49476 19698 49532
rect 19698 49476 19702 49532
rect 19638 49472 19702 49476
rect 19718 49532 19782 49536
rect 19718 49476 19722 49532
rect 19722 49476 19778 49532
rect 19778 49476 19782 49532
rect 19718 49472 19782 49476
rect 19798 49532 19862 49536
rect 19798 49476 19802 49532
rect 19802 49476 19858 49532
rect 19858 49476 19862 49532
rect 19798 49472 19862 49476
rect 50278 49532 50342 49536
rect 50278 49476 50282 49532
rect 50282 49476 50338 49532
rect 50338 49476 50342 49532
rect 50278 49472 50342 49476
rect 50358 49532 50422 49536
rect 50358 49476 50362 49532
rect 50362 49476 50418 49532
rect 50418 49476 50422 49532
rect 50358 49472 50422 49476
rect 50438 49532 50502 49536
rect 50438 49476 50442 49532
rect 50442 49476 50498 49532
rect 50498 49476 50502 49532
rect 50438 49472 50502 49476
rect 50518 49532 50582 49536
rect 50518 49476 50522 49532
rect 50522 49476 50578 49532
rect 50578 49476 50582 49532
rect 50518 49472 50582 49476
rect 4198 48988 4262 48992
rect 4198 48932 4202 48988
rect 4202 48932 4258 48988
rect 4258 48932 4262 48988
rect 4198 48928 4262 48932
rect 4278 48988 4342 48992
rect 4278 48932 4282 48988
rect 4282 48932 4338 48988
rect 4338 48932 4342 48988
rect 4278 48928 4342 48932
rect 4358 48988 4422 48992
rect 4358 48932 4362 48988
rect 4362 48932 4418 48988
rect 4418 48932 4422 48988
rect 4358 48928 4422 48932
rect 4438 48988 4502 48992
rect 4438 48932 4442 48988
rect 4442 48932 4498 48988
rect 4498 48932 4502 48988
rect 4438 48928 4502 48932
rect 34918 48988 34982 48992
rect 34918 48932 34922 48988
rect 34922 48932 34978 48988
rect 34978 48932 34982 48988
rect 34918 48928 34982 48932
rect 34998 48988 35062 48992
rect 34998 48932 35002 48988
rect 35002 48932 35058 48988
rect 35058 48932 35062 48988
rect 34998 48928 35062 48932
rect 35078 48988 35142 48992
rect 35078 48932 35082 48988
rect 35082 48932 35138 48988
rect 35138 48932 35142 48988
rect 35078 48928 35142 48932
rect 35158 48988 35222 48992
rect 35158 48932 35162 48988
rect 35162 48932 35218 48988
rect 35218 48932 35222 48988
rect 35158 48928 35222 48932
rect 19558 48444 19622 48448
rect 19558 48388 19562 48444
rect 19562 48388 19618 48444
rect 19618 48388 19622 48444
rect 19558 48384 19622 48388
rect 19638 48444 19702 48448
rect 19638 48388 19642 48444
rect 19642 48388 19698 48444
rect 19698 48388 19702 48444
rect 19638 48384 19702 48388
rect 19718 48444 19782 48448
rect 19718 48388 19722 48444
rect 19722 48388 19778 48444
rect 19778 48388 19782 48444
rect 19718 48384 19782 48388
rect 19798 48444 19862 48448
rect 19798 48388 19802 48444
rect 19802 48388 19858 48444
rect 19858 48388 19862 48444
rect 19798 48384 19862 48388
rect 50278 48444 50342 48448
rect 50278 48388 50282 48444
rect 50282 48388 50338 48444
rect 50338 48388 50342 48444
rect 50278 48384 50342 48388
rect 50358 48444 50422 48448
rect 50358 48388 50362 48444
rect 50362 48388 50418 48444
rect 50418 48388 50422 48444
rect 50358 48384 50422 48388
rect 50438 48444 50502 48448
rect 50438 48388 50442 48444
rect 50442 48388 50498 48444
rect 50498 48388 50502 48444
rect 50438 48384 50502 48388
rect 50518 48444 50582 48448
rect 50518 48388 50522 48444
rect 50522 48388 50578 48444
rect 50578 48388 50582 48444
rect 50518 48384 50582 48388
rect 4198 47900 4262 47904
rect 4198 47844 4202 47900
rect 4202 47844 4258 47900
rect 4258 47844 4262 47900
rect 4198 47840 4262 47844
rect 4278 47900 4342 47904
rect 4278 47844 4282 47900
rect 4282 47844 4338 47900
rect 4338 47844 4342 47900
rect 4278 47840 4342 47844
rect 4358 47900 4422 47904
rect 4358 47844 4362 47900
rect 4362 47844 4418 47900
rect 4418 47844 4422 47900
rect 4358 47840 4422 47844
rect 4438 47900 4502 47904
rect 4438 47844 4442 47900
rect 4442 47844 4498 47900
rect 4498 47844 4502 47900
rect 4438 47840 4502 47844
rect 34918 47900 34982 47904
rect 34918 47844 34922 47900
rect 34922 47844 34978 47900
rect 34978 47844 34982 47900
rect 34918 47840 34982 47844
rect 34998 47900 35062 47904
rect 34998 47844 35002 47900
rect 35002 47844 35058 47900
rect 35058 47844 35062 47900
rect 34998 47840 35062 47844
rect 35078 47900 35142 47904
rect 35078 47844 35082 47900
rect 35082 47844 35138 47900
rect 35138 47844 35142 47900
rect 35078 47840 35142 47844
rect 35158 47900 35222 47904
rect 35158 47844 35162 47900
rect 35162 47844 35218 47900
rect 35218 47844 35222 47900
rect 35158 47840 35222 47844
rect 19558 47356 19622 47360
rect 19558 47300 19562 47356
rect 19562 47300 19618 47356
rect 19618 47300 19622 47356
rect 19558 47296 19622 47300
rect 19638 47356 19702 47360
rect 19638 47300 19642 47356
rect 19642 47300 19698 47356
rect 19698 47300 19702 47356
rect 19638 47296 19702 47300
rect 19718 47356 19782 47360
rect 19718 47300 19722 47356
rect 19722 47300 19778 47356
rect 19778 47300 19782 47356
rect 19718 47296 19782 47300
rect 19798 47356 19862 47360
rect 19798 47300 19802 47356
rect 19802 47300 19858 47356
rect 19858 47300 19862 47356
rect 19798 47296 19862 47300
rect 50278 47356 50342 47360
rect 50278 47300 50282 47356
rect 50282 47300 50338 47356
rect 50338 47300 50342 47356
rect 50278 47296 50342 47300
rect 50358 47356 50422 47360
rect 50358 47300 50362 47356
rect 50362 47300 50418 47356
rect 50418 47300 50422 47356
rect 50358 47296 50422 47300
rect 50438 47356 50502 47360
rect 50438 47300 50442 47356
rect 50442 47300 50498 47356
rect 50498 47300 50502 47356
rect 50438 47296 50502 47300
rect 50518 47356 50582 47360
rect 50518 47300 50522 47356
rect 50522 47300 50578 47356
rect 50578 47300 50582 47356
rect 50518 47296 50582 47300
rect 4198 46812 4262 46816
rect 4198 46756 4202 46812
rect 4202 46756 4258 46812
rect 4258 46756 4262 46812
rect 4198 46752 4262 46756
rect 4278 46812 4342 46816
rect 4278 46756 4282 46812
rect 4282 46756 4338 46812
rect 4338 46756 4342 46812
rect 4278 46752 4342 46756
rect 4358 46812 4422 46816
rect 4358 46756 4362 46812
rect 4362 46756 4418 46812
rect 4418 46756 4422 46812
rect 4358 46752 4422 46756
rect 4438 46812 4502 46816
rect 4438 46756 4442 46812
rect 4442 46756 4498 46812
rect 4498 46756 4502 46812
rect 4438 46752 4502 46756
rect 34918 46812 34982 46816
rect 34918 46756 34922 46812
rect 34922 46756 34978 46812
rect 34978 46756 34982 46812
rect 34918 46752 34982 46756
rect 34998 46812 35062 46816
rect 34998 46756 35002 46812
rect 35002 46756 35058 46812
rect 35058 46756 35062 46812
rect 34998 46752 35062 46756
rect 35078 46812 35142 46816
rect 35078 46756 35082 46812
rect 35082 46756 35138 46812
rect 35138 46756 35142 46812
rect 35078 46752 35142 46756
rect 35158 46812 35222 46816
rect 35158 46756 35162 46812
rect 35162 46756 35218 46812
rect 35218 46756 35222 46812
rect 35158 46752 35222 46756
rect 19558 46268 19622 46272
rect 19558 46212 19562 46268
rect 19562 46212 19618 46268
rect 19618 46212 19622 46268
rect 19558 46208 19622 46212
rect 19638 46268 19702 46272
rect 19638 46212 19642 46268
rect 19642 46212 19698 46268
rect 19698 46212 19702 46268
rect 19638 46208 19702 46212
rect 19718 46268 19782 46272
rect 19718 46212 19722 46268
rect 19722 46212 19778 46268
rect 19778 46212 19782 46268
rect 19718 46208 19782 46212
rect 19798 46268 19862 46272
rect 19798 46212 19802 46268
rect 19802 46212 19858 46268
rect 19858 46212 19862 46268
rect 19798 46208 19862 46212
rect 50278 46268 50342 46272
rect 50278 46212 50282 46268
rect 50282 46212 50338 46268
rect 50338 46212 50342 46268
rect 50278 46208 50342 46212
rect 50358 46268 50422 46272
rect 50358 46212 50362 46268
rect 50362 46212 50418 46268
rect 50418 46212 50422 46268
rect 50358 46208 50422 46212
rect 50438 46268 50502 46272
rect 50438 46212 50442 46268
rect 50442 46212 50498 46268
rect 50498 46212 50502 46268
rect 50438 46208 50502 46212
rect 50518 46268 50582 46272
rect 50518 46212 50522 46268
rect 50522 46212 50578 46268
rect 50578 46212 50582 46268
rect 50518 46208 50582 46212
rect 4198 45724 4262 45728
rect 4198 45668 4202 45724
rect 4202 45668 4258 45724
rect 4258 45668 4262 45724
rect 4198 45664 4262 45668
rect 4278 45724 4342 45728
rect 4278 45668 4282 45724
rect 4282 45668 4338 45724
rect 4338 45668 4342 45724
rect 4278 45664 4342 45668
rect 4358 45724 4422 45728
rect 4358 45668 4362 45724
rect 4362 45668 4418 45724
rect 4418 45668 4422 45724
rect 4358 45664 4422 45668
rect 4438 45724 4502 45728
rect 4438 45668 4442 45724
rect 4442 45668 4498 45724
rect 4498 45668 4502 45724
rect 4438 45664 4502 45668
rect 34918 45724 34982 45728
rect 34918 45668 34922 45724
rect 34922 45668 34978 45724
rect 34978 45668 34982 45724
rect 34918 45664 34982 45668
rect 34998 45724 35062 45728
rect 34998 45668 35002 45724
rect 35002 45668 35058 45724
rect 35058 45668 35062 45724
rect 34998 45664 35062 45668
rect 35078 45724 35142 45728
rect 35078 45668 35082 45724
rect 35082 45668 35138 45724
rect 35138 45668 35142 45724
rect 35078 45664 35142 45668
rect 35158 45724 35222 45728
rect 35158 45668 35162 45724
rect 35162 45668 35218 45724
rect 35218 45668 35222 45724
rect 35158 45664 35222 45668
rect 19558 45180 19622 45184
rect 19558 45124 19562 45180
rect 19562 45124 19618 45180
rect 19618 45124 19622 45180
rect 19558 45120 19622 45124
rect 19638 45180 19702 45184
rect 19638 45124 19642 45180
rect 19642 45124 19698 45180
rect 19698 45124 19702 45180
rect 19638 45120 19702 45124
rect 19718 45180 19782 45184
rect 19718 45124 19722 45180
rect 19722 45124 19778 45180
rect 19778 45124 19782 45180
rect 19718 45120 19782 45124
rect 19798 45180 19862 45184
rect 19798 45124 19802 45180
rect 19802 45124 19858 45180
rect 19858 45124 19862 45180
rect 19798 45120 19862 45124
rect 50278 45180 50342 45184
rect 50278 45124 50282 45180
rect 50282 45124 50338 45180
rect 50338 45124 50342 45180
rect 50278 45120 50342 45124
rect 50358 45180 50422 45184
rect 50358 45124 50362 45180
rect 50362 45124 50418 45180
rect 50418 45124 50422 45180
rect 50358 45120 50422 45124
rect 50438 45180 50502 45184
rect 50438 45124 50442 45180
rect 50442 45124 50498 45180
rect 50498 45124 50502 45180
rect 50438 45120 50502 45124
rect 50518 45180 50582 45184
rect 50518 45124 50522 45180
rect 50522 45124 50578 45180
rect 50578 45124 50582 45180
rect 50518 45120 50582 45124
rect 4198 44636 4262 44640
rect 4198 44580 4202 44636
rect 4202 44580 4258 44636
rect 4258 44580 4262 44636
rect 4198 44576 4262 44580
rect 4278 44636 4342 44640
rect 4278 44580 4282 44636
rect 4282 44580 4338 44636
rect 4338 44580 4342 44636
rect 4278 44576 4342 44580
rect 4358 44636 4422 44640
rect 4358 44580 4362 44636
rect 4362 44580 4418 44636
rect 4418 44580 4422 44636
rect 4358 44576 4422 44580
rect 4438 44636 4502 44640
rect 4438 44580 4442 44636
rect 4442 44580 4498 44636
rect 4498 44580 4502 44636
rect 4438 44576 4502 44580
rect 34918 44636 34982 44640
rect 34918 44580 34922 44636
rect 34922 44580 34978 44636
rect 34978 44580 34982 44636
rect 34918 44576 34982 44580
rect 34998 44636 35062 44640
rect 34998 44580 35002 44636
rect 35002 44580 35058 44636
rect 35058 44580 35062 44636
rect 34998 44576 35062 44580
rect 35078 44636 35142 44640
rect 35078 44580 35082 44636
rect 35082 44580 35138 44636
rect 35138 44580 35142 44636
rect 35078 44576 35142 44580
rect 35158 44636 35222 44640
rect 35158 44580 35162 44636
rect 35162 44580 35218 44636
rect 35218 44580 35222 44636
rect 35158 44576 35222 44580
rect 19558 44092 19622 44096
rect 19558 44036 19562 44092
rect 19562 44036 19618 44092
rect 19618 44036 19622 44092
rect 19558 44032 19622 44036
rect 19638 44092 19702 44096
rect 19638 44036 19642 44092
rect 19642 44036 19698 44092
rect 19698 44036 19702 44092
rect 19638 44032 19702 44036
rect 19718 44092 19782 44096
rect 19718 44036 19722 44092
rect 19722 44036 19778 44092
rect 19778 44036 19782 44092
rect 19718 44032 19782 44036
rect 19798 44092 19862 44096
rect 19798 44036 19802 44092
rect 19802 44036 19858 44092
rect 19858 44036 19862 44092
rect 19798 44032 19862 44036
rect 50278 44092 50342 44096
rect 50278 44036 50282 44092
rect 50282 44036 50338 44092
rect 50338 44036 50342 44092
rect 50278 44032 50342 44036
rect 50358 44092 50422 44096
rect 50358 44036 50362 44092
rect 50362 44036 50418 44092
rect 50418 44036 50422 44092
rect 50358 44032 50422 44036
rect 50438 44092 50502 44096
rect 50438 44036 50442 44092
rect 50442 44036 50498 44092
rect 50498 44036 50502 44092
rect 50438 44032 50502 44036
rect 50518 44092 50582 44096
rect 50518 44036 50522 44092
rect 50522 44036 50578 44092
rect 50578 44036 50582 44092
rect 50518 44032 50582 44036
rect 4198 43548 4262 43552
rect 4198 43492 4202 43548
rect 4202 43492 4258 43548
rect 4258 43492 4262 43548
rect 4198 43488 4262 43492
rect 4278 43548 4342 43552
rect 4278 43492 4282 43548
rect 4282 43492 4338 43548
rect 4338 43492 4342 43548
rect 4278 43488 4342 43492
rect 4358 43548 4422 43552
rect 4358 43492 4362 43548
rect 4362 43492 4418 43548
rect 4418 43492 4422 43548
rect 4358 43488 4422 43492
rect 4438 43548 4502 43552
rect 4438 43492 4442 43548
rect 4442 43492 4498 43548
rect 4498 43492 4502 43548
rect 4438 43488 4502 43492
rect 34918 43548 34982 43552
rect 34918 43492 34922 43548
rect 34922 43492 34978 43548
rect 34978 43492 34982 43548
rect 34918 43488 34982 43492
rect 34998 43548 35062 43552
rect 34998 43492 35002 43548
rect 35002 43492 35058 43548
rect 35058 43492 35062 43548
rect 34998 43488 35062 43492
rect 35078 43548 35142 43552
rect 35078 43492 35082 43548
rect 35082 43492 35138 43548
rect 35138 43492 35142 43548
rect 35078 43488 35142 43492
rect 35158 43548 35222 43552
rect 35158 43492 35162 43548
rect 35162 43492 35218 43548
rect 35218 43492 35222 43548
rect 35158 43488 35222 43492
rect 19558 43004 19622 43008
rect 19558 42948 19562 43004
rect 19562 42948 19618 43004
rect 19618 42948 19622 43004
rect 19558 42944 19622 42948
rect 19638 43004 19702 43008
rect 19638 42948 19642 43004
rect 19642 42948 19698 43004
rect 19698 42948 19702 43004
rect 19638 42944 19702 42948
rect 19718 43004 19782 43008
rect 19718 42948 19722 43004
rect 19722 42948 19778 43004
rect 19778 42948 19782 43004
rect 19718 42944 19782 42948
rect 19798 43004 19862 43008
rect 19798 42948 19802 43004
rect 19802 42948 19858 43004
rect 19858 42948 19862 43004
rect 19798 42944 19862 42948
rect 50278 43004 50342 43008
rect 50278 42948 50282 43004
rect 50282 42948 50338 43004
rect 50338 42948 50342 43004
rect 50278 42944 50342 42948
rect 50358 43004 50422 43008
rect 50358 42948 50362 43004
rect 50362 42948 50418 43004
rect 50418 42948 50422 43004
rect 50358 42944 50422 42948
rect 50438 43004 50502 43008
rect 50438 42948 50442 43004
rect 50442 42948 50498 43004
rect 50498 42948 50502 43004
rect 50438 42944 50502 42948
rect 50518 43004 50582 43008
rect 50518 42948 50522 43004
rect 50522 42948 50578 43004
rect 50578 42948 50582 43004
rect 50518 42944 50582 42948
rect 4198 42460 4262 42464
rect 4198 42404 4202 42460
rect 4202 42404 4258 42460
rect 4258 42404 4262 42460
rect 4198 42400 4262 42404
rect 4278 42460 4342 42464
rect 4278 42404 4282 42460
rect 4282 42404 4338 42460
rect 4338 42404 4342 42460
rect 4278 42400 4342 42404
rect 4358 42460 4422 42464
rect 4358 42404 4362 42460
rect 4362 42404 4418 42460
rect 4418 42404 4422 42460
rect 4358 42400 4422 42404
rect 4438 42460 4502 42464
rect 4438 42404 4442 42460
rect 4442 42404 4498 42460
rect 4498 42404 4502 42460
rect 4438 42400 4502 42404
rect 34918 42460 34982 42464
rect 34918 42404 34922 42460
rect 34922 42404 34978 42460
rect 34978 42404 34982 42460
rect 34918 42400 34982 42404
rect 34998 42460 35062 42464
rect 34998 42404 35002 42460
rect 35002 42404 35058 42460
rect 35058 42404 35062 42460
rect 34998 42400 35062 42404
rect 35078 42460 35142 42464
rect 35078 42404 35082 42460
rect 35082 42404 35138 42460
rect 35138 42404 35142 42460
rect 35078 42400 35142 42404
rect 35158 42460 35222 42464
rect 35158 42404 35162 42460
rect 35162 42404 35218 42460
rect 35218 42404 35222 42460
rect 35158 42400 35222 42404
rect 19558 41916 19622 41920
rect 19558 41860 19562 41916
rect 19562 41860 19618 41916
rect 19618 41860 19622 41916
rect 19558 41856 19622 41860
rect 19638 41916 19702 41920
rect 19638 41860 19642 41916
rect 19642 41860 19698 41916
rect 19698 41860 19702 41916
rect 19638 41856 19702 41860
rect 19718 41916 19782 41920
rect 19718 41860 19722 41916
rect 19722 41860 19778 41916
rect 19778 41860 19782 41916
rect 19718 41856 19782 41860
rect 19798 41916 19862 41920
rect 19798 41860 19802 41916
rect 19802 41860 19858 41916
rect 19858 41860 19862 41916
rect 19798 41856 19862 41860
rect 50278 41916 50342 41920
rect 50278 41860 50282 41916
rect 50282 41860 50338 41916
rect 50338 41860 50342 41916
rect 50278 41856 50342 41860
rect 50358 41916 50422 41920
rect 50358 41860 50362 41916
rect 50362 41860 50418 41916
rect 50418 41860 50422 41916
rect 50358 41856 50422 41860
rect 50438 41916 50502 41920
rect 50438 41860 50442 41916
rect 50442 41860 50498 41916
rect 50498 41860 50502 41916
rect 50438 41856 50502 41860
rect 50518 41916 50582 41920
rect 50518 41860 50522 41916
rect 50522 41860 50578 41916
rect 50578 41860 50582 41916
rect 50518 41856 50582 41860
rect 4198 41372 4262 41376
rect 4198 41316 4202 41372
rect 4202 41316 4258 41372
rect 4258 41316 4262 41372
rect 4198 41312 4262 41316
rect 4278 41372 4342 41376
rect 4278 41316 4282 41372
rect 4282 41316 4338 41372
rect 4338 41316 4342 41372
rect 4278 41312 4342 41316
rect 4358 41372 4422 41376
rect 4358 41316 4362 41372
rect 4362 41316 4418 41372
rect 4418 41316 4422 41372
rect 4358 41312 4422 41316
rect 4438 41372 4502 41376
rect 4438 41316 4442 41372
rect 4442 41316 4498 41372
rect 4498 41316 4502 41372
rect 4438 41312 4502 41316
rect 34918 41372 34982 41376
rect 34918 41316 34922 41372
rect 34922 41316 34978 41372
rect 34978 41316 34982 41372
rect 34918 41312 34982 41316
rect 34998 41372 35062 41376
rect 34998 41316 35002 41372
rect 35002 41316 35058 41372
rect 35058 41316 35062 41372
rect 34998 41312 35062 41316
rect 35078 41372 35142 41376
rect 35078 41316 35082 41372
rect 35082 41316 35138 41372
rect 35138 41316 35142 41372
rect 35078 41312 35142 41316
rect 35158 41372 35222 41376
rect 35158 41316 35162 41372
rect 35162 41316 35218 41372
rect 35218 41316 35222 41372
rect 35158 41312 35222 41316
rect 19558 40828 19622 40832
rect 19558 40772 19562 40828
rect 19562 40772 19618 40828
rect 19618 40772 19622 40828
rect 19558 40768 19622 40772
rect 19638 40828 19702 40832
rect 19638 40772 19642 40828
rect 19642 40772 19698 40828
rect 19698 40772 19702 40828
rect 19638 40768 19702 40772
rect 19718 40828 19782 40832
rect 19718 40772 19722 40828
rect 19722 40772 19778 40828
rect 19778 40772 19782 40828
rect 19718 40768 19782 40772
rect 19798 40828 19862 40832
rect 19798 40772 19802 40828
rect 19802 40772 19858 40828
rect 19858 40772 19862 40828
rect 19798 40768 19862 40772
rect 50278 40828 50342 40832
rect 50278 40772 50282 40828
rect 50282 40772 50338 40828
rect 50338 40772 50342 40828
rect 50278 40768 50342 40772
rect 50358 40828 50422 40832
rect 50358 40772 50362 40828
rect 50362 40772 50418 40828
rect 50418 40772 50422 40828
rect 50358 40768 50422 40772
rect 50438 40828 50502 40832
rect 50438 40772 50442 40828
rect 50442 40772 50498 40828
rect 50498 40772 50502 40828
rect 50438 40768 50502 40772
rect 50518 40828 50582 40832
rect 50518 40772 50522 40828
rect 50522 40772 50578 40828
rect 50578 40772 50582 40828
rect 50518 40768 50582 40772
rect 4198 40284 4262 40288
rect 4198 40228 4202 40284
rect 4202 40228 4258 40284
rect 4258 40228 4262 40284
rect 4198 40224 4262 40228
rect 4278 40284 4342 40288
rect 4278 40228 4282 40284
rect 4282 40228 4338 40284
rect 4338 40228 4342 40284
rect 4278 40224 4342 40228
rect 4358 40284 4422 40288
rect 4358 40228 4362 40284
rect 4362 40228 4418 40284
rect 4418 40228 4422 40284
rect 4358 40224 4422 40228
rect 4438 40284 4502 40288
rect 4438 40228 4442 40284
rect 4442 40228 4498 40284
rect 4498 40228 4502 40284
rect 4438 40224 4502 40228
rect 34918 40284 34982 40288
rect 34918 40228 34922 40284
rect 34922 40228 34978 40284
rect 34978 40228 34982 40284
rect 34918 40224 34982 40228
rect 34998 40284 35062 40288
rect 34998 40228 35002 40284
rect 35002 40228 35058 40284
rect 35058 40228 35062 40284
rect 34998 40224 35062 40228
rect 35078 40284 35142 40288
rect 35078 40228 35082 40284
rect 35082 40228 35138 40284
rect 35138 40228 35142 40284
rect 35078 40224 35142 40228
rect 35158 40284 35222 40288
rect 35158 40228 35162 40284
rect 35162 40228 35218 40284
rect 35218 40228 35222 40284
rect 35158 40224 35222 40228
rect 19558 39740 19622 39744
rect 19558 39684 19562 39740
rect 19562 39684 19618 39740
rect 19618 39684 19622 39740
rect 19558 39680 19622 39684
rect 19638 39740 19702 39744
rect 19638 39684 19642 39740
rect 19642 39684 19698 39740
rect 19698 39684 19702 39740
rect 19638 39680 19702 39684
rect 19718 39740 19782 39744
rect 19718 39684 19722 39740
rect 19722 39684 19778 39740
rect 19778 39684 19782 39740
rect 19718 39680 19782 39684
rect 19798 39740 19862 39744
rect 19798 39684 19802 39740
rect 19802 39684 19858 39740
rect 19858 39684 19862 39740
rect 19798 39680 19862 39684
rect 50278 39740 50342 39744
rect 50278 39684 50282 39740
rect 50282 39684 50338 39740
rect 50338 39684 50342 39740
rect 50278 39680 50342 39684
rect 50358 39740 50422 39744
rect 50358 39684 50362 39740
rect 50362 39684 50418 39740
rect 50418 39684 50422 39740
rect 50358 39680 50422 39684
rect 50438 39740 50502 39744
rect 50438 39684 50442 39740
rect 50442 39684 50498 39740
rect 50498 39684 50502 39740
rect 50438 39680 50502 39684
rect 50518 39740 50582 39744
rect 50518 39684 50522 39740
rect 50522 39684 50578 39740
rect 50578 39684 50582 39740
rect 50518 39680 50582 39684
rect 4198 39196 4262 39200
rect 4198 39140 4202 39196
rect 4202 39140 4258 39196
rect 4258 39140 4262 39196
rect 4198 39136 4262 39140
rect 4278 39196 4342 39200
rect 4278 39140 4282 39196
rect 4282 39140 4338 39196
rect 4338 39140 4342 39196
rect 4278 39136 4342 39140
rect 4358 39196 4422 39200
rect 4358 39140 4362 39196
rect 4362 39140 4418 39196
rect 4418 39140 4422 39196
rect 4358 39136 4422 39140
rect 4438 39196 4502 39200
rect 4438 39140 4442 39196
rect 4442 39140 4498 39196
rect 4498 39140 4502 39196
rect 4438 39136 4502 39140
rect 34918 39196 34982 39200
rect 34918 39140 34922 39196
rect 34922 39140 34978 39196
rect 34978 39140 34982 39196
rect 34918 39136 34982 39140
rect 34998 39196 35062 39200
rect 34998 39140 35002 39196
rect 35002 39140 35058 39196
rect 35058 39140 35062 39196
rect 34998 39136 35062 39140
rect 35078 39196 35142 39200
rect 35078 39140 35082 39196
rect 35082 39140 35138 39196
rect 35138 39140 35142 39196
rect 35078 39136 35142 39140
rect 35158 39196 35222 39200
rect 35158 39140 35162 39196
rect 35162 39140 35218 39196
rect 35218 39140 35222 39196
rect 35158 39136 35222 39140
rect 19558 38652 19622 38656
rect 19558 38596 19562 38652
rect 19562 38596 19618 38652
rect 19618 38596 19622 38652
rect 19558 38592 19622 38596
rect 19638 38652 19702 38656
rect 19638 38596 19642 38652
rect 19642 38596 19698 38652
rect 19698 38596 19702 38652
rect 19638 38592 19702 38596
rect 19718 38652 19782 38656
rect 19718 38596 19722 38652
rect 19722 38596 19778 38652
rect 19778 38596 19782 38652
rect 19718 38592 19782 38596
rect 19798 38652 19862 38656
rect 19798 38596 19802 38652
rect 19802 38596 19858 38652
rect 19858 38596 19862 38652
rect 19798 38592 19862 38596
rect 50278 38652 50342 38656
rect 50278 38596 50282 38652
rect 50282 38596 50338 38652
rect 50338 38596 50342 38652
rect 50278 38592 50342 38596
rect 50358 38652 50422 38656
rect 50358 38596 50362 38652
rect 50362 38596 50418 38652
rect 50418 38596 50422 38652
rect 50358 38592 50422 38596
rect 50438 38652 50502 38656
rect 50438 38596 50442 38652
rect 50442 38596 50498 38652
rect 50498 38596 50502 38652
rect 50438 38592 50502 38596
rect 50518 38652 50582 38656
rect 50518 38596 50522 38652
rect 50522 38596 50578 38652
rect 50578 38596 50582 38652
rect 50518 38592 50582 38596
rect 4198 38108 4262 38112
rect 4198 38052 4202 38108
rect 4202 38052 4258 38108
rect 4258 38052 4262 38108
rect 4198 38048 4262 38052
rect 4278 38108 4342 38112
rect 4278 38052 4282 38108
rect 4282 38052 4338 38108
rect 4338 38052 4342 38108
rect 4278 38048 4342 38052
rect 4358 38108 4422 38112
rect 4358 38052 4362 38108
rect 4362 38052 4418 38108
rect 4418 38052 4422 38108
rect 4358 38048 4422 38052
rect 4438 38108 4502 38112
rect 4438 38052 4442 38108
rect 4442 38052 4498 38108
rect 4498 38052 4502 38108
rect 4438 38048 4502 38052
rect 34918 38108 34982 38112
rect 34918 38052 34922 38108
rect 34922 38052 34978 38108
rect 34978 38052 34982 38108
rect 34918 38048 34982 38052
rect 34998 38108 35062 38112
rect 34998 38052 35002 38108
rect 35002 38052 35058 38108
rect 35058 38052 35062 38108
rect 34998 38048 35062 38052
rect 35078 38108 35142 38112
rect 35078 38052 35082 38108
rect 35082 38052 35138 38108
rect 35138 38052 35142 38108
rect 35078 38048 35142 38052
rect 35158 38108 35222 38112
rect 35158 38052 35162 38108
rect 35162 38052 35218 38108
rect 35218 38052 35222 38108
rect 35158 38048 35222 38052
rect 19558 37564 19622 37568
rect 19558 37508 19562 37564
rect 19562 37508 19618 37564
rect 19618 37508 19622 37564
rect 19558 37504 19622 37508
rect 19638 37564 19702 37568
rect 19638 37508 19642 37564
rect 19642 37508 19698 37564
rect 19698 37508 19702 37564
rect 19638 37504 19702 37508
rect 19718 37564 19782 37568
rect 19718 37508 19722 37564
rect 19722 37508 19778 37564
rect 19778 37508 19782 37564
rect 19718 37504 19782 37508
rect 19798 37564 19862 37568
rect 19798 37508 19802 37564
rect 19802 37508 19858 37564
rect 19858 37508 19862 37564
rect 19798 37504 19862 37508
rect 50278 37564 50342 37568
rect 50278 37508 50282 37564
rect 50282 37508 50338 37564
rect 50338 37508 50342 37564
rect 50278 37504 50342 37508
rect 50358 37564 50422 37568
rect 50358 37508 50362 37564
rect 50362 37508 50418 37564
rect 50418 37508 50422 37564
rect 50358 37504 50422 37508
rect 50438 37564 50502 37568
rect 50438 37508 50442 37564
rect 50442 37508 50498 37564
rect 50498 37508 50502 37564
rect 50438 37504 50502 37508
rect 50518 37564 50582 37568
rect 50518 37508 50522 37564
rect 50522 37508 50578 37564
rect 50578 37508 50582 37564
rect 50518 37504 50582 37508
rect 4198 37020 4262 37024
rect 4198 36964 4202 37020
rect 4202 36964 4258 37020
rect 4258 36964 4262 37020
rect 4198 36960 4262 36964
rect 4278 37020 4342 37024
rect 4278 36964 4282 37020
rect 4282 36964 4338 37020
rect 4338 36964 4342 37020
rect 4278 36960 4342 36964
rect 4358 37020 4422 37024
rect 4358 36964 4362 37020
rect 4362 36964 4418 37020
rect 4418 36964 4422 37020
rect 4358 36960 4422 36964
rect 4438 37020 4502 37024
rect 4438 36964 4442 37020
rect 4442 36964 4498 37020
rect 4498 36964 4502 37020
rect 4438 36960 4502 36964
rect 34918 37020 34982 37024
rect 34918 36964 34922 37020
rect 34922 36964 34978 37020
rect 34978 36964 34982 37020
rect 34918 36960 34982 36964
rect 34998 37020 35062 37024
rect 34998 36964 35002 37020
rect 35002 36964 35058 37020
rect 35058 36964 35062 37020
rect 34998 36960 35062 36964
rect 35078 37020 35142 37024
rect 35078 36964 35082 37020
rect 35082 36964 35138 37020
rect 35138 36964 35142 37020
rect 35078 36960 35142 36964
rect 35158 37020 35222 37024
rect 35158 36964 35162 37020
rect 35162 36964 35218 37020
rect 35218 36964 35222 37020
rect 35158 36960 35222 36964
rect 19558 36476 19622 36480
rect 19558 36420 19562 36476
rect 19562 36420 19618 36476
rect 19618 36420 19622 36476
rect 19558 36416 19622 36420
rect 19638 36476 19702 36480
rect 19638 36420 19642 36476
rect 19642 36420 19698 36476
rect 19698 36420 19702 36476
rect 19638 36416 19702 36420
rect 19718 36476 19782 36480
rect 19718 36420 19722 36476
rect 19722 36420 19778 36476
rect 19778 36420 19782 36476
rect 19718 36416 19782 36420
rect 19798 36476 19862 36480
rect 19798 36420 19802 36476
rect 19802 36420 19858 36476
rect 19858 36420 19862 36476
rect 19798 36416 19862 36420
rect 50278 36476 50342 36480
rect 50278 36420 50282 36476
rect 50282 36420 50338 36476
rect 50338 36420 50342 36476
rect 50278 36416 50342 36420
rect 50358 36476 50422 36480
rect 50358 36420 50362 36476
rect 50362 36420 50418 36476
rect 50418 36420 50422 36476
rect 50358 36416 50422 36420
rect 50438 36476 50502 36480
rect 50438 36420 50442 36476
rect 50442 36420 50498 36476
rect 50498 36420 50502 36476
rect 50438 36416 50502 36420
rect 50518 36476 50582 36480
rect 50518 36420 50522 36476
rect 50522 36420 50578 36476
rect 50578 36420 50582 36476
rect 50518 36416 50582 36420
rect 4198 35932 4262 35936
rect 4198 35876 4202 35932
rect 4202 35876 4258 35932
rect 4258 35876 4262 35932
rect 4198 35872 4262 35876
rect 4278 35932 4342 35936
rect 4278 35876 4282 35932
rect 4282 35876 4338 35932
rect 4338 35876 4342 35932
rect 4278 35872 4342 35876
rect 4358 35932 4422 35936
rect 4358 35876 4362 35932
rect 4362 35876 4418 35932
rect 4418 35876 4422 35932
rect 4358 35872 4422 35876
rect 4438 35932 4502 35936
rect 4438 35876 4442 35932
rect 4442 35876 4498 35932
rect 4498 35876 4502 35932
rect 4438 35872 4502 35876
rect 34918 35932 34982 35936
rect 34918 35876 34922 35932
rect 34922 35876 34978 35932
rect 34978 35876 34982 35932
rect 34918 35872 34982 35876
rect 34998 35932 35062 35936
rect 34998 35876 35002 35932
rect 35002 35876 35058 35932
rect 35058 35876 35062 35932
rect 34998 35872 35062 35876
rect 35078 35932 35142 35936
rect 35078 35876 35082 35932
rect 35082 35876 35138 35932
rect 35138 35876 35142 35932
rect 35078 35872 35142 35876
rect 35158 35932 35222 35936
rect 35158 35876 35162 35932
rect 35162 35876 35218 35932
rect 35218 35876 35222 35932
rect 35158 35872 35222 35876
rect 19558 35388 19622 35392
rect 19558 35332 19562 35388
rect 19562 35332 19618 35388
rect 19618 35332 19622 35388
rect 19558 35328 19622 35332
rect 19638 35388 19702 35392
rect 19638 35332 19642 35388
rect 19642 35332 19698 35388
rect 19698 35332 19702 35388
rect 19638 35328 19702 35332
rect 19718 35388 19782 35392
rect 19718 35332 19722 35388
rect 19722 35332 19778 35388
rect 19778 35332 19782 35388
rect 19718 35328 19782 35332
rect 19798 35388 19862 35392
rect 19798 35332 19802 35388
rect 19802 35332 19858 35388
rect 19858 35332 19862 35388
rect 19798 35328 19862 35332
rect 50278 35388 50342 35392
rect 50278 35332 50282 35388
rect 50282 35332 50338 35388
rect 50338 35332 50342 35388
rect 50278 35328 50342 35332
rect 50358 35388 50422 35392
rect 50358 35332 50362 35388
rect 50362 35332 50418 35388
rect 50418 35332 50422 35388
rect 50358 35328 50422 35332
rect 50438 35388 50502 35392
rect 50438 35332 50442 35388
rect 50442 35332 50498 35388
rect 50498 35332 50502 35388
rect 50438 35328 50502 35332
rect 50518 35388 50582 35392
rect 50518 35332 50522 35388
rect 50522 35332 50578 35388
rect 50578 35332 50582 35388
rect 50518 35328 50582 35332
rect 4198 34844 4262 34848
rect 4198 34788 4202 34844
rect 4202 34788 4258 34844
rect 4258 34788 4262 34844
rect 4198 34784 4262 34788
rect 4278 34844 4342 34848
rect 4278 34788 4282 34844
rect 4282 34788 4338 34844
rect 4338 34788 4342 34844
rect 4278 34784 4342 34788
rect 4358 34844 4422 34848
rect 4358 34788 4362 34844
rect 4362 34788 4418 34844
rect 4418 34788 4422 34844
rect 4358 34784 4422 34788
rect 4438 34844 4502 34848
rect 4438 34788 4442 34844
rect 4442 34788 4498 34844
rect 4498 34788 4502 34844
rect 4438 34784 4502 34788
rect 34918 34844 34982 34848
rect 34918 34788 34922 34844
rect 34922 34788 34978 34844
rect 34978 34788 34982 34844
rect 34918 34784 34982 34788
rect 34998 34844 35062 34848
rect 34998 34788 35002 34844
rect 35002 34788 35058 34844
rect 35058 34788 35062 34844
rect 34998 34784 35062 34788
rect 35078 34844 35142 34848
rect 35078 34788 35082 34844
rect 35082 34788 35138 34844
rect 35138 34788 35142 34844
rect 35078 34784 35142 34788
rect 35158 34844 35222 34848
rect 35158 34788 35162 34844
rect 35162 34788 35218 34844
rect 35218 34788 35222 34844
rect 35158 34784 35222 34788
rect 19558 34300 19622 34304
rect 19558 34244 19562 34300
rect 19562 34244 19618 34300
rect 19618 34244 19622 34300
rect 19558 34240 19622 34244
rect 19638 34300 19702 34304
rect 19638 34244 19642 34300
rect 19642 34244 19698 34300
rect 19698 34244 19702 34300
rect 19638 34240 19702 34244
rect 19718 34300 19782 34304
rect 19718 34244 19722 34300
rect 19722 34244 19778 34300
rect 19778 34244 19782 34300
rect 19718 34240 19782 34244
rect 19798 34300 19862 34304
rect 19798 34244 19802 34300
rect 19802 34244 19858 34300
rect 19858 34244 19862 34300
rect 19798 34240 19862 34244
rect 50278 34300 50342 34304
rect 50278 34244 50282 34300
rect 50282 34244 50338 34300
rect 50338 34244 50342 34300
rect 50278 34240 50342 34244
rect 50358 34300 50422 34304
rect 50358 34244 50362 34300
rect 50362 34244 50418 34300
rect 50418 34244 50422 34300
rect 50358 34240 50422 34244
rect 50438 34300 50502 34304
rect 50438 34244 50442 34300
rect 50442 34244 50498 34300
rect 50498 34244 50502 34300
rect 50438 34240 50502 34244
rect 50518 34300 50582 34304
rect 50518 34244 50522 34300
rect 50522 34244 50578 34300
rect 50578 34244 50582 34300
rect 50518 34240 50582 34244
rect 4198 33756 4262 33760
rect 4198 33700 4202 33756
rect 4202 33700 4258 33756
rect 4258 33700 4262 33756
rect 4198 33696 4262 33700
rect 4278 33756 4342 33760
rect 4278 33700 4282 33756
rect 4282 33700 4338 33756
rect 4338 33700 4342 33756
rect 4278 33696 4342 33700
rect 4358 33756 4422 33760
rect 4358 33700 4362 33756
rect 4362 33700 4418 33756
rect 4418 33700 4422 33756
rect 4358 33696 4422 33700
rect 4438 33756 4502 33760
rect 4438 33700 4442 33756
rect 4442 33700 4498 33756
rect 4498 33700 4502 33756
rect 4438 33696 4502 33700
rect 34918 33756 34982 33760
rect 34918 33700 34922 33756
rect 34922 33700 34978 33756
rect 34978 33700 34982 33756
rect 34918 33696 34982 33700
rect 34998 33756 35062 33760
rect 34998 33700 35002 33756
rect 35002 33700 35058 33756
rect 35058 33700 35062 33756
rect 34998 33696 35062 33700
rect 35078 33756 35142 33760
rect 35078 33700 35082 33756
rect 35082 33700 35138 33756
rect 35138 33700 35142 33756
rect 35078 33696 35142 33700
rect 35158 33756 35222 33760
rect 35158 33700 35162 33756
rect 35162 33700 35218 33756
rect 35218 33700 35222 33756
rect 35158 33696 35222 33700
rect 19558 33212 19622 33216
rect 19558 33156 19562 33212
rect 19562 33156 19618 33212
rect 19618 33156 19622 33212
rect 19558 33152 19622 33156
rect 19638 33212 19702 33216
rect 19638 33156 19642 33212
rect 19642 33156 19698 33212
rect 19698 33156 19702 33212
rect 19638 33152 19702 33156
rect 19718 33212 19782 33216
rect 19718 33156 19722 33212
rect 19722 33156 19778 33212
rect 19778 33156 19782 33212
rect 19718 33152 19782 33156
rect 19798 33212 19862 33216
rect 19798 33156 19802 33212
rect 19802 33156 19858 33212
rect 19858 33156 19862 33212
rect 19798 33152 19862 33156
rect 50278 33212 50342 33216
rect 50278 33156 50282 33212
rect 50282 33156 50338 33212
rect 50338 33156 50342 33212
rect 50278 33152 50342 33156
rect 50358 33212 50422 33216
rect 50358 33156 50362 33212
rect 50362 33156 50418 33212
rect 50418 33156 50422 33212
rect 50358 33152 50422 33156
rect 50438 33212 50502 33216
rect 50438 33156 50442 33212
rect 50442 33156 50498 33212
rect 50498 33156 50502 33212
rect 50438 33152 50502 33156
rect 50518 33212 50582 33216
rect 50518 33156 50522 33212
rect 50522 33156 50578 33212
rect 50578 33156 50582 33212
rect 50518 33152 50582 33156
rect 4198 32668 4262 32672
rect 4198 32612 4202 32668
rect 4202 32612 4258 32668
rect 4258 32612 4262 32668
rect 4198 32608 4262 32612
rect 4278 32668 4342 32672
rect 4278 32612 4282 32668
rect 4282 32612 4338 32668
rect 4338 32612 4342 32668
rect 4278 32608 4342 32612
rect 4358 32668 4422 32672
rect 4358 32612 4362 32668
rect 4362 32612 4418 32668
rect 4418 32612 4422 32668
rect 4358 32608 4422 32612
rect 4438 32668 4502 32672
rect 4438 32612 4442 32668
rect 4442 32612 4498 32668
rect 4498 32612 4502 32668
rect 4438 32608 4502 32612
rect 34918 32668 34982 32672
rect 34918 32612 34922 32668
rect 34922 32612 34978 32668
rect 34978 32612 34982 32668
rect 34918 32608 34982 32612
rect 34998 32668 35062 32672
rect 34998 32612 35002 32668
rect 35002 32612 35058 32668
rect 35058 32612 35062 32668
rect 34998 32608 35062 32612
rect 35078 32668 35142 32672
rect 35078 32612 35082 32668
rect 35082 32612 35138 32668
rect 35138 32612 35142 32668
rect 35078 32608 35142 32612
rect 35158 32668 35222 32672
rect 35158 32612 35162 32668
rect 35162 32612 35218 32668
rect 35218 32612 35222 32668
rect 35158 32608 35222 32612
rect 19558 32124 19622 32128
rect 19558 32068 19562 32124
rect 19562 32068 19618 32124
rect 19618 32068 19622 32124
rect 19558 32064 19622 32068
rect 19638 32124 19702 32128
rect 19638 32068 19642 32124
rect 19642 32068 19698 32124
rect 19698 32068 19702 32124
rect 19638 32064 19702 32068
rect 19718 32124 19782 32128
rect 19718 32068 19722 32124
rect 19722 32068 19778 32124
rect 19778 32068 19782 32124
rect 19718 32064 19782 32068
rect 19798 32124 19862 32128
rect 19798 32068 19802 32124
rect 19802 32068 19858 32124
rect 19858 32068 19862 32124
rect 19798 32064 19862 32068
rect 50278 32124 50342 32128
rect 50278 32068 50282 32124
rect 50282 32068 50338 32124
rect 50338 32068 50342 32124
rect 50278 32064 50342 32068
rect 50358 32124 50422 32128
rect 50358 32068 50362 32124
rect 50362 32068 50418 32124
rect 50418 32068 50422 32124
rect 50358 32064 50422 32068
rect 50438 32124 50502 32128
rect 50438 32068 50442 32124
rect 50442 32068 50498 32124
rect 50498 32068 50502 32124
rect 50438 32064 50502 32068
rect 50518 32124 50582 32128
rect 50518 32068 50522 32124
rect 50522 32068 50578 32124
rect 50578 32068 50582 32124
rect 50518 32064 50582 32068
rect 4198 31580 4262 31584
rect 4198 31524 4202 31580
rect 4202 31524 4258 31580
rect 4258 31524 4262 31580
rect 4198 31520 4262 31524
rect 4278 31580 4342 31584
rect 4278 31524 4282 31580
rect 4282 31524 4338 31580
rect 4338 31524 4342 31580
rect 4278 31520 4342 31524
rect 4358 31580 4422 31584
rect 4358 31524 4362 31580
rect 4362 31524 4418 31580
rect 4418 31524 4422 31580
rect 4358 31520 4422 31524
rect 4438 31580 4502 31584
rect 4438 31524 4442 31580
rect 4442 31524 4498 31580
rect 4498 31524 4502 31580
rect 4438 31520 4502 31524
rect 34918 31580 34982 31584
rect 34918 31524 34922 31580
rect 34922 31524 34978 31580
rect 34978 31524 34982 31580
rect 34918 31520 34982 31524
rect 34998 31580 35062 31584
rect 34998 31524 35002 31580
rect 35002 31524 35058 31580
rect 35058 31524 35062 31580
rect 34998 31520 35062 31524
rect 35078 31580 35142 31584
rect 35078 31524 35082 31580
rect 35082 31524 35138 31580
rect 35138 31524 35142 31580
rect 35078 31520 35142 31524
rect 35158 31580 35222 31584
rect 35158 31524 35162 31580
rect 35162 31524 35218 31580
rect 35218 31524 35222 31580
rect 35158 31520 35222 31524
rect 19558 31036 19622 31040
rect 19558 30980 19562 31036
rect 19562 30980 19618 31036
rect 19618 30980 19622 31036
rect 19558 30976 19622 30980
rect 19638 31036 19702 31040
rect 19638 30980 19642 31036
rect 19642 30980 19698 31036
rect 19698 30980 19702 31036
rect 19638 30976 19702 30980
rect 19718 31036 19782 31040
rect 19718 30980 19722 31036
rect 19722 30980 19778 31036
rect 19778 30980 19782 31036
rect 19718 30976 19782 30980
rect 19798 31036 19862 31040
rect 19798 30980 19802 31036
rect 19802 30980 19858 31036
rect 19858 30980 19862 31036
rect 19798 30976 19862 30980
rect 50278 31036 50342 31040
rect 50278 30980 50282 31036
rect 50282 30980 50338 31036
rect 50338 30980 50342 31036
rect 50278 30976 50342 30980
rect 50358 31036 50422 31040
rect 50358 30980 50362 31036
rect 50362 30980 50418 31036
rect 50418 30980 50422 31036
rect 50358 30976 50422 30980
rect 50438 31036 50502 31040
rect 50438 30980 50442 31036
rect 50442 30980 50498 31036
rect 50498 30980 50502 31036
rect 50438 30976 50502 30980
rect 50518 31036 50582 31040
rect 50518 30980 50522 31036
rect 50522 30980 50578 31036
rect 50578 30980 50582 31036
rect 50518 30976 50582 30980
rect 4198 30492 4262 30496
rect 4198 30436 4202 30492
rect 4202 30436 4258 30492
rect 4258 30436 4262 30492
rect 4198 30432 4262 30436
rect 4278 30492 4342 30496
rect 4278 30436 4282 30492
rect 4282 30436 4338 30492
rect 4338 30436 4342 30492
rect 4278 30432 4342 30436
rect 4358 30492 4422 30496
rect 4358 30436 4362 30492
rect 4362 30436 4418 30492
rect 4418 30436 4422 30492
rect 4358 30432 4422 30436
rect 4438 30492 4502 30496
rect 4438 30436 4442 30492
rect 4442 30436 4498 30492
rect 4498 30436 4502 30492
rect 4438 30432 4502 30436
rect 34918 30492 34982 30496
rect 34918 30436 34922 30492
rect 34922 30436 34978 30492
rect 34978 30436 34982 30492
rect 34918 30432 34982 30436
rect 34998 30492 35062 30496
rect 34998 30436 35002 30492
rect 35002 30436 35058 30492
rect 35058 30436 35062 30492
rect 34998 30432 35062 30436
rect 35078 30492 35142 30496
rect 35078 30436 35082 30492
rect 35082 30436 35138 30492
rect 35138 30436 35142 30492
rect 35078 30432 35142 30436
rect 35158 30492 35222 30496
rect 35158 30436 35162 30492
rect 35162 30436 35218 30492
rect 35218 30436 35222 30492
rect 35158 30432 35222 30436
rect 19558 29948 19622 29952
rect 19558 29892 19562 29948
rect 19562 29892 19618 29948
rect 19618 29892 19622 29948
rect 19558 29888 19622 29892
rect 19638 29948 19702 29952
rect 19638 29892 19642 29948
rect 19642 29892 19698 29948
rect 19698 29892 19702 29948
rect 19638 29888 19702 29892
rect 19718 29948 19782 29952
rect 19718 29892 19722 29948
rect 19722 29892 19778 29948
rect 19778 29892 19782 29948
rect 19718 29888 19782 29892
rect 19798 29948 19862 29952
rect 19798 29892 19802 29948
rect 19802 29892 19858 29948
rect 19858 29892 19862 29948
rect 19798 29888 19862 29892
rect 50278 29948 50342 29952
rect 50278 29892 50282 29948
rect 50282 29892 50338 29948
rect 50338 29892 50342 29948
rect 50278 29888 50342 29892
rect 50358 29948 50422 29952
rect 50358 29892 50362 29948
rect 50362 29892 50418 29948
rect 50418 29892 50422 29948
rect 50358 29888 50422 29892
rect 50438 29948 50502 29952
rect 50438 29892 50442 29948
rect 50442 29892 50498 29948
rect 50498 29892 50502 29948
rect 50438 29888 50502 29892
rect 50518 29948 50582 29952
rect 50518 29892 50522 29948
rect 50522 29892 50578 29948
rect 50578 29892 50582 29948
rect 50518 29888 50582 29892
rect 4198 29404 4262 29408
rect 4198 29348 4202 29404
rect 4202 29348 4258 29404
rect 4258 29348 4262 29404
rect 4198 29344 4262 29348
rect 4278 29404 4342 29408
rect 4278 29348 4282 29404
rect 4282 29348 4338 29404
rect 4338 29348 4342 29404
rect 4278 29344 4342 29348
rect 4358 29404 4422 29408
rect 4358 29348 4362 29404
rect 4362 29348 4418 29404
rect 4418 29348 4422 29404
rect 4358 29344 4422 29348
rect 4438 29404 4502 29408
rect 4438 29348 4442 29404
rect 4442 29348 4498 29404
rect 4498 29348 4502 29404
rect 4438 29344 4502 29348
rect 34918 29404 34982 29408
rect 34918 29348 34922 29404
rect 34922 29348 34978 29404
rect 34978 29348 34982 29404
rect 34918 29344 34982 29348
rect 34998 29404 35062 29408
rect 34998 29348 35002 29404
rect 35002 29348 35058 29404
rect 35058 29348 35062 29404
rect 34998 29344 35062 29348
rect 35078 29404 35142 29408
rect 35078 29348 35082 29404
rect 35082 29348 35138 29404
rect 35138 29348 35142 29404
rect 35078 29344 35142 29348
rect 35158 29404 35222 29408
rect 35158 29348 35162 29404
rect 35162 29348 35218 29404
rect 35218 29348 35222 29404
rect 35158 29344 35222 29348
rect 19558 28860 19622 28864
rect 19558 28804 19562 28860
rect 19562 28804 19618 28860
rect 19618 28804 19622 28860
rect 19558 28800 19622 28804
rect 19638 28860 19702 28864
rect 19638 28804 19642 28860
rect 19642 28804 19698 28860
rect 19698 28804 19702 28860
rect 19638 28800 19702 28804
rect 19718 28860 19782 28864
rect 19718 28804 19722 28860
rect 19722 28804 19778 28860
rect 19778 28804 19782 28860
rect 19718 28800 19782 28804
rect 19798 28860 19862 28864
rect 19798 28804 19802 28860
rect 19802 28804 19858 28860
rect 19858 28804 19862 28860
rect 19798 28800 19862 28804
rect 50278 28860 50342 28864
rect 50278 28804 50282 28860
rect 50282 28804 50338 28860
rect 50338 28804 50342 28860
rect 50278 28800 50342 28804
rect 50358 28860 50422 28864
rect 50358 28804 50362 28860
rect 50362 28804 50418 28860
rect 50418 28804 50422 28860
rect 50358 28800 50422 28804
rect 50438 28860 50502 28864
rect 50438 28804 50442 28860
rect 50442 28804 50498 28860
rect 50498 28804 50502 28860
rect 50438 28800 50502 28804
rect 50518 28860 50582 28864
rect 50518 28804 50522 28860
rect 50522 28804 50578 28860
rect 50578 28804 50582 28860
rect 50518 28800 50582 28804
rect 4198 28316 4262 28320
rect 4198 28260 4202 28316
rect 4202 28260 4258 28316
rect 4258 28260 4262 28316
rect 4198 28256 4262 28260
rect 4278 28316 4342 28320
rect 4278 28260 4282 28316
rect 4282 28260 4338 28316
rect 4338 28260 4342 28316
rect 4278 28256 4342 28260
rect 4358 28316 4422 28320
rect 4358 28260 4362 28316
rect 4362 28260 4418 28316
rect 4418 28260 4422 28316
rect 4358 28256 4422 28260
rect 4438 28316 4502 28320
rect 4438 28260 4442 28316
rect 4442 28260 4498 28316
rect 4498 28260 4502 28316
rect 4438 28256 4502 28260
rect 34918 28316 34982 28320
rect 34918 28260 34922 28316
rect 34922 28260 34978 28316
rect 34978 28260 34982 28316
rect 34918 28256 34982 28260
rect 34998 28316 35062 28320
rect 34998 28260 35002 28316
rect 35002 28260 35058 28316
rect 35058 28260 35062 28316
rect 34998 28256 35062 28260
rect 35078 28316 35142 28320
rect 35078 28260 35082 28316
rect 35082 28260 35138 28316
rect 35138 28260 35142 28316
rect 35078 28256 35142 28260
rect 35158 28316 35222 28320
rect 35158 28260 35162 28316
rect 35162 28260 35218 28316
rect 35218 28260 35222 28316
rect 35158 28256 35222 28260
rect 19558 27772 19622 27776
rect 19558 27716 19562 27772
rect 19562 27716 19618 27772
rect 19618 27716 19622 27772
rect 19558 27712 19622 27716
rect 19638 27772 19702 27776
rect 19638 27716 19642 27772
rect 19642 27716 19698 27772
rect 19698 27716 19702 27772
rect 19638 27712 19702 27716
rect 19718 27772 19782 27776
rect 19718 27716 19722 27772
rect 19722 27716 19778 27772
rect 19778 27716 19782 27772
rect 19718 27712 19782 27716
rect 19798 27772 19862 27776
rect 19798 27716 19802 27772
rect 19802 27716 19858 27772
rect 19858 27716 19862 27772
rect 19798 27712 19862 27716
rect 50278 27772 50342 27776
rect 50278 27716 50282 27772
rect 50282 27716 50338 27772
rect 50338 27716 50342 27772
rect 50278 27712 50342 27716
rect 50358 27772 50422 27776
rect 50358 27716 50362 27772
rect 50362 27716 50418 27772
rect 50418 27716 50422 27772
rect 50358 27712 50422 27716
rect 50438 27772 50502 27776
rect 50438 27716 50442 27772
rect 50442 27716 50498 27772
rect 50498 27716 50502 27772
rect 50438 27712 50502 27716
rect 50518 27772 50582 27776
rect 50518 27716 50522 27772
rect 50522 27716 50578 27772
rect 50578 27716 50582 27772
rect 50518 27712 50582 27716
rect 4198 27228 4262 27232
rect 4198 27172 4202 27228
rect 4202 27172 4258 27228
rect 4258 27172 4262 27228
rect 4198 27168 4262 27172
rect 4278 27228 4342 27232
rect 4278 27172 4282 27228
rect 4282 27172 4338 27228
rect 4338 27172 4342 27228
rect 4278 27168 4342 27172
rect 4358 27228 4422 27232
rect 4358 27172 4362 27228
rect 4362 27172 4418 27228
rect 4418 27172 4422 27228
rect 4358 27168 4422 27172
rect 4438 27228 4502 27232
rect 4438 27172 4442 27228
rect 4442 27172 4498 27228
rect 4498 27172 4502 27228
rect 4438 27168 4502 27172
rect 34918 27228 34982 27232
rect 34918 27172 34922 27228
rect 34922 27172 34978 27228
rect 34978 27172 34982 27228
rect 34918 27168 34982 27172
rect 34998 27228 35062 27232
rect 34998 27172 35002 27228
rect 35002 27172 35058 27228
rect 35058 27172 35062 27228
rect 34998 27168 35062 27172
rect 35078 27228 35142 27232
rect 35078 27172 35082 27228
rect 35082 27172 35138 27228
rect 35138 27172 35142 27228
rect 35078 27168 35142 27172
rect 35158 27228 35222 27232
rect 35158 27172 35162 27228
rect 35162 27172 35218 27228
rect 35218 27172 35222 27228
rect 35158 27168 35222 27172
rect 19558 26684 19622 26688
rect 19558 26628 19562 26684
rect 19562 26628 19618 26684
rect 19618 26628 19622 26684
rect 19558 26624 19622 26628
rect 19638 26684 19702 26688
rect 19638 26628 19642 26684
rect 19642 26628 19698 26684
rect 19698 26628 19702 26684
rect 19638 26624 19702 26628
rect 19718 26684 19782 26688
rect 19718 26628 19722 26684
rect 19722 26628 19778 26684
rect 19778 26628 19782 26684
rect 19718 26624 19782 26628
rect 19798 26684 19862 26688
rect 19798 26628 19802 26684
rect 19802 26628 19858 26684
rect 19858 26628 19862 26684
rect 19798 26624 19862 26628
rect 50278 26684 50342 26688
rect 50278 26628 50282 26684
rect 50282 26628 50338 26684
rect 50338 26628 50342 26684
rect 50278 26624 50342 26628
rect 50358 26684 50422 26688
rect 50358 26628 50362 26684
rect 50362 26628 50418 26684
rect 50418 26628 50422 26684
rect 50358 26624 50422 26628
rect 50438 26684 50502 26688
rect 50438 26628 50442 26684
rect 50442 26628 50498 26684
rect 50498 26628 50502 26684
rect 50438 26624 50502 26628
rect 50518 26684 50582 26688
rect 50518 26628 50522 26684
rect 50522 26628 50578 26684
rect 50578 26628 50582 26684
rect 50518 26624 50582 26628
rect 4198 26140 4262 26144
rect 4198 26084 4202 26140
rect 4202 26084 4258 26140
rect 4258 26084 4262 26140
rect 4198 26080 4262 26084
rect 4278 26140 4342 26144
rect 4278 26084 4282 26140
rect 4282 26084 4338 26140
rect 4338 26084 4342 26140
rect 4278 26080 4342 26084
rect 4358 26140 4422 26144
rect 4358 26084 4362 26140
rect 4362 26084 4418 26140
rect 4418 26084 4422 26140
rect 4358 26080 4422 26084
rect 4438 26140 4502 26144
rect 4438 26084 4442 26140
rect 4442 26084 4498 26140
rect 4498 26084 4502 26140
rect 4438 26080 4502 26084
rect 34918 26140 34982 26144
rect 34918 26084 34922 26140
rect 34922 26084 34978 26140
rect 34978 26084 34982 26140
rect 34918 26080 34982 26084
rect 34998 26140 35062 26144
rect 34998 26084 35002 26140
rect 35002 26084 35058 26140
rect 35058 26084 35062 26140
rect 34998 26080 35062 26084
rect 35078 26140 35142 26144
rect 35078 26084 35082 26140
rect 35082 26084 35138 26140
rect 35138 26084 35142 26140
rect 35078 26080 35142 26084
rect 35158 26140 35222 26144
rect 35158 26084 35162 26140
rect 35162 26084 35218 26140
rect 35218 26084 35222 26140
rect 35158 26080 35222 26084
rect 19558 25596 19622 25600
rect 19558 25540 19562 25596
rect 19562 25540 19618 25596
rect 19618 25540 19622 25596
rect 19558 25536 19622 25540
rect 19638 25596 19702 25600
rect 19638 25540 19642 25596
rect 19642 25540 19698 25596
rect 19698 25540 19702 25596
rect 19638 25536 19702 25540
rect 19718 25596 19782 25600
rect 19718 25540 19722 25596
rect 19722 25540 19778 25596
rect 19778 25540 19782 25596
rect 19718 25536 19782 25540
rect 19798 25596 19862 25600
rect 19798 25540 19802 25596
rect 19802 25540 19858 25596
rect 19858 25540 19862 25596
rect 19798 25536 19862 25540
rect 50278 25596 50342 25600
rect 50278 25540 50282 25596
rect 50282 25540 50338 25596
rect 50338 25540 50342 25596
rect 50278 25536 50342 25540
rect 50358 25596 50422 25600
rect 50358 25540 50362 25596
rect 50362 25540 50418 25596
rect 50418 25540 50422 25596
rect 50358 25536 50422 25540
rect 50438 25596 50502 25600
rect 50438 25540 50442 25596
rect 50442 25540 50498 25596
rect 50498 25540 50502 25596
rect 50438 25536 50502 25540
rect 50518 25596 50582 25600
rect 50518 25540 50522 25596
rect 50522 25540 50578 25596
rect 50578 25540 50582 25596
rect 50518 25536 50582 25540
rect 4198 25052 4262 25056
rect 4198 24996 4202 25052
rect 4202 24996 4258 25052
rect 4258 24996 4262 25052
rect 4198 24992 4262 24996
rect 4278 25052 4342 25056
rect 4278 24996 4282 25052
rect 4282 24996 4338 25052
rect 4338 24996 4342 25052
rect 4278 24992 4342 24996
rect 4358 25052 4422 25056
rect 4358 24996 4362 25052
rect 4362 24996 4418 25052
rect 4418 24996 4422 25052
rect 4358 24992 4422 24996
rect 4438 25052 4502 25056
rect 4438 24996 4442 25052
rect 4442 24996 4498 25052
rect 4498 24996 4502 25052
rect 4438 24992 4502 24996
rect 34918 25052 34982 25056
rect 34918 24996 34922 25052
rect 34922 24996 34978 25052
rect 34978 24996 34982 25052
rect 34918 24992 34982 24996
rect 34998 25052 35062 25056
rect 34998 24996 35002 25052
rect 35002 24996 35058 25052
rect 35058 24996 35062 25052
rect 34998 24992 35062 24996
rect 35078 25052 35142 25056
rect 35078 24996 35082 25052
rect 35082 24996 35138 25052
rect 35138 24996 35142 25052
rect 35078 24992 35142 24996
rect 35158 25052 35222 25056
rect 35158 24996 35162 25052
rect 35162 24996 35218 25052
rect 35218 24996 35222 25052
rect 35158 24992 35222 24996
rect 19558 24508 19622 24512
rect 19558 24452 19562 24508
rect 19562 24452 19618 24508
rect 19618 24452 19622 24508
rect 19558 24448 19622 24452
rect 19638 24508 19702 24512
rect 19638 24452 19642 24508
rect 19642 24452 19698 24508
rect 19698 24452 19702 24508
rect 19638 24448 19702 24452
rect 19718 24508 19782 24512
rect 19718 24452 19722 24508
rect 19722 24452 19778 24508
rect 19778 24452 19782 24508
rect 19718 24448 19782 24452
rect 19798 24508 19862 24512
rect 19798 24452 19802 24508
rect 19802 24452 19858 24508
rect 19858 24452 19862 24508
rect 19798 24448 19862 24452
rect 50278 24508 50342 24512
rect 50278 24452 50282 24508
rect 50282 24452 50338 24508
rect 50338 24452 50342 24508
rect 50278 24448 50342 24452
rect 50358 24508 50422 24512
rect 50358 24452 50362 24508
rect 50362 24452 50418 24508
rect 50418 24452 50422 24508
rect 50358 24448 50422 24452
rect 50438 24508 50502 24512
rect 50438 24452 50442 24508
rect 50442 24452 50498 24508
rect 50498 24452 50502 24508
rect 50438 24448 50502 24452
rect 50518 24508 50582 24512
rect 50518 24452 50522 24508
rect 50522 24452 50578 24508
rect 50578 24452 50582 24508
rect 50518 24448 50582 24452
rect 4198 23964 4262 23968
rect 4198 23908 4202 23964
rect 4202 23908 4258 23964
rect 4258 23908 4262 23964
rect 4198 23904 4262 23908
rect 4278 23964 4342 23968
rect 4278 23908 4282 23964
rect 4282 23908 4338 23964
rect 4338 23908 4342 23964
rect 4278 23904 4342 23908
rect 4358 23964 4422 23968
rect 4358 23908 4362 23964
rect 4362 23908 4418 23964
rect 4418 23908 4422 23964
rect 4358 23904 4422 23908
rect 4438 23964 4502 23968
rect 4438 23908 4442 23964
rect 4442 23908 4498 23964
rect 4498 23908 4502 23964
rect 4438 23904 4502 23908
rect 34918 23964 34982 23968
rect 34918 23908 34922 23964
rect 34922 23908 34978 23964
rect 34978 23908 34982 23964
rect 34918 23904 34982 23908
rect 34998 23964 35062 23968
rect 34998 23908 35002 23964
rect 35002 23908 35058 23964
rect 35058 23908 35062 23964
rect 34998 23904 35062 23908
rect 35078 23964 35142 23968
rect 35078 23908 35082 23964
rect 35082 23908 35138 23964
rect 35138 23908 35142 23964
rect 35078 23904 35142 23908
rect 35158 23964 35222 23968
rect 35158 23908 35162 23964
rect 35162 23908 35218 23964
rect 35218 23908 35222 23964
rect 35158 23904 35222 23908
rect 19558 23420 19622 23424
rect 19558 23364 19562 23420
rect 19562 23364 19618 23420
rect 19618 23364 19622 23420
rect 19558 23360 19622 23364
rect 19638 23420 19702 23424
rect 19638 23364 19642 23420
rect 19642 23364 19698 23420
rect 19698 23364 19702 23420
rect 19638 23360 19702 23364
rect 19718 23420 19782 23424
rect 19718 23364 19722 23420
rect 19722 23364 19778 23420
rect 19778 23364 19782 23420
rect 19718 23360 19782 23364
rect 19798 23420 19862 23424
rect 19798 23364 19802 23420
rect 19802 23364 19858 23420
rect 19858 23364 19862 23420
rect 19798 23360 19862 23364
rect 50278 23420 50342 23424
rect 50278 23364 50282 23420
rect 50282 23364 50338 23420
rect 50338 23364 50342 23420
rect 50278 23360 50342 23364
rect 50358 23420 50422 23424
rect 50358 23364 50362 23420
rect 50362 23364 50418 23420
rect 50418 23364 50422 23420
rect 50358 23360 50422 23364
rect 50438 23420 50502 23424
rect 50438 23364 50442 23420
rect 50442 23364 50498 23420
rect 50498 23364 50502 23420
rect 50438 23360 50502 23364
rect 50518 23420 50582 23424
rect 50518 23364 50522 23420
rect 50522 23364 50578 23420
rect 50578 23364 50582 23420
rect 50518 23360 50582 23364
rect 4198 22876 4262 22880
rect 4198 22820 4202 22876
rect 4202 22820 4258 22876
rect 4258 22820 4262 22876
rect 4198 22816 4262 22820
rect 4278 22876 4342 22880
rect 4278 22820 4282 22876
rect 4282 22820 4338 22876
rect 4338 22820 4342 22876
rect 4278 22816 4342 22820
rect 4358 22876 4422 22880
rect 4358 22820 4362 22876
rect 4362 22820 4418 22876
rect 4418 22820 4422 22876
rect 4358 22816 4422 22820
rect 4438 22876 4502 22880
rect 4438 22820 4442 22876
rect 4442 22820 4498 22876
rect 4498 22820 4502 22876
rect 4438 22816 4502 22820
rect 34918 22876 34982 22880
rect 34918 22820 34922 22876
rect 34922 22820 34978 22876
rect 34978 22820 34982 22876
rect 34918 22816 34982 22820
rect 34998 22876 35062 22880
rect 34998 22820 35002 22876
rect 35002 22820 35058 22876
rect 35058 22820 35062 22876
rect 34998 22816 35062 22820
rect 35078 22876 35142 22880
rect 35078 22820 35082 22876
rect 35082 22820 35138 22876
rect 35138 22820 35142 22876
rect 35078 22816 35142 22820
rect 35158 22876 35222 22880
rect 35158 22820 35162 22876
rect 35162 22820 35218 22876
rect 35218 22820 35222 22876
rect 35158 22816 35222 22820
rect 19558 22332 19622 22336
rect 19558 22276 19562 22332
rect 19562 22276 19618 22332
rect 19618 22276 19622 22332
rect 19558 22272 19622 22276
rect 19638 22332 19702 22336
rect 19638 22276 19642 22332
rect 19642 22276 19698 22332
rect 19698 22276 19702 22332
rect 19638 22272 19702 22276
rect 19718 22332 19782 22336
rect 19718 22276 19722 22332
rect 19722 22276 19778 22332
rect 19778 22276 19782 22332
rect 19718 22272 19782 22276
rect 19798 22332 19862 22336
rect 19798 22276 19802 22332
rect 19802 22276 19858 22332
rect 19858 22276 19862 22332
rect 19798 22272 19862 22276
rect 50278 22332 50342 22336
rect 50278 22276 50282 22332
rect 50282 22276 50338 22332
rect 50338 22276 50342 22332
rect 50278 22272 50342 22276
rect 50358 22332 50422 22336
rect 50358 22276 50362 22332
rect 50362 22276 50418 22332
rect 50418 22276 50422 22332
rect 50358 22272 50422 22276
rect 50438 22332 50502 22336
rect 50438 22276 50442 22332
rect 50442 22276 50498 22332
rect 50498 22276 50502 22332
rect 50438 22272 50502 22276
rect 50518 22332 50582 22336
rect 50518 22276 50522 22332
rect 50522 22276 50578 22332
rect 50578 22276 50582 22332
rect 50518 22272 50582 22276
rect 4198 21788 4262 21792
rect 4198 21732 4202 21788
rect 4202 21732 4258 21788
rect 4258 21732 4262 21788
rect 4198 21728 4262 21732
rect 4278 21788 4342 21792
rect 4278 21732 4282 21788
rect 4282 21732 4338 21788
rect 4338 21732 4342 21788
rect 4278 21728 4342 21732
rect 4358 21788 4422 21792
rect 4358 21732 4362 21788
rect 4362 21732 4418 21788
rect 4418 21732 4422 21788
rect 4358 21728 4422 21732
rect 4438 21788 4502 21792
rect 4438 21732 4442 21788
rect 4442 21732 4498 21788
rect 4498 21732 4502 21788
rect 4438 21728 4502 21732
rect 34918 21788 34982 21792
rect 34918 21732 34922 21788
rect 34922 21732 34978 21788
rect 34978 21732 34982 21788
rect 34918 21728 34982 21732
rect 34998 21788 35062 21792
rect 34998 21732 35002 21788
rect 35002 21732 35058 21788
rect 35058 21732 35062 21788
rect 34998 21728 35062 21732
rect 35078 21788 35142 21792
rect 35078 21732 35082 21788
rect 35082 21732 35138 21788
rect 35138 21732 35142 21788
rect 35078 21728 35142 21732
rect 35158 21788 35222 21792
rect 35158 21732 35162 21788
rect 35162 21732 35218 21788
rect 35218 21732 35222 21788
rect 35158 21728 35222 21732
rect 19558 21244 19622 21248
rect 19558 21188 19562 21244
rect 19562 21188 19618 21244
rect 19618 21188 19622 21244
rect 19558 21184 19622 21188
rect 19638 21244 19702 21248
rect 19638 21188 19642 21244
rect 19642 21188 19698 21244
rect 19698 21188 19702 21244
rect 19638 21184 19702 21188
rect 19718 21244 19782 21248
rect 19718 21188 19722 21244
rect 19722 21188 19778 21244
rect 19778 21188 19782 21244
rect 19718 21184 19782 21188
rect 19798 21244 19862 21248
rect 19798 21188 19802 21244
rect 19802 21188 19858 21244
rect 19858 21188 19862 21244
rect 19798 21184 19862 21188
rect 50278 21244 50342 21248
rect 50278 21188 50282 21244
rect 50282 21188 50338 21244
rect 50338 21188 50342 21244
rect 50278 21184 50342 21188
rect 50358 21244 50422 21248
rect 50358 21188 50362 21244
rect 50362 21188 50418 21244
rect 50418 21188 50422 21244
rect 50358 21184 50422 21188
rect 50438 21244 50502 21248
rect 50438 21188 50442 21244
rect 50442 21188 50498 21244
rect 50498 21188 50502 21244
rect 50438 21184 50502 21188
rect 50518 21244 50582 21248
rect 50518 21188 50522 21244
rect 50522 21188 50578 21244
rect 50578 21188 50582 21244
rect 50518 21184 50582 21188
rect 4198 20700 4262 20704
rect 4198 20644 4202 20700
rect 4202 20644 4258 20700
rect 4258 20644 4262 20700
rect 4198 20640 4262 20644
rect 4278 20700 4342 20704
rect 4278 20644 4282 20700
rect 4282 20644 4338 20700
rect 4338 20644 4342 20700
rect 4278 20640 4342 20644
rect 4358 20700 4422 20704
rect 4358 20644 4362 20700
rect 4362 20644 4418 20700
rect 4418 20644 4422 20700
rect 4358 20640 4422 20644
rect 4438 20700 4502 20704
rect 4438 20644 4442 20700
rect 4442 20644 4498 20700
rect 4498 20644 4502 20700
rect 4438 20640 4502 20644
rect 34918 20700 34982 20704
rect 34918 20644 34922 20700
rect 34922 20644 34978 20700
rect 34978 20644 34982 20700
rect 34918 20640 34982 20644
rect 34998 20700 35062 20704
rect 34998 20644 35002 20700
rect 35002 20644 35058 20700
rect 35058 20644 35062 20700
rect 34998 20640 35062 20644
rect 35078 20700 35142 20704
rect 35078 20644 35082 20700
rect 35082 20644 35138 20700
rect 35138 20644 35142 20700
rect 35078 20640 35142 20644
rect 35158 20700 35222 20704
rect 35158 20644 35162 20700
rect 35162 20644 35218 20700
rect 35218 20644 35222 20700
rect 35158 20640 35222 20644
rect 19558 20156 19622 20160
rect 19558 20100 19562 20156
rect 19562 20100 19618 20156
rect 19618 20100 19622 20156
rect 19558 20096 19622 20100
rect 19638 20156 19702 20160
rect 19638 20100 19642 20156
rect 19642 20100 19698 20156
rect 19698 20100 19702 20156
rect 19638 20096 19702 20100
rect 19718 20156 19782 20160
rect 19718 20100 19722 20156
rect 19722 20100 19778 20156
rect 19778 20100 19782 20156
rect 19718 20096 19782 20100
rect 19798 20156 19862 20160
rect 19798 20100 19802 20156
rect 19802 20100 19858 20156
rect 19858 20100 19862 20156
rect 19798 20096 19862 20100
rect 50278 20156 50342 20160
rect 50278 20100 50282 20156
rect 50282 20100 50338 20156
rect 50338 20100 50342 20156
rect 50278 20096 50342 20100
rect 50358 20156 50422 20160
rect 50358 20100 50362 20156
rect 50362 20100 50418 20156
rect 50418 20100 50422 20156
rect 50358 20096 50422 20100
rect 50438 20156 50502 20160
rect 50438 20100 50442 20156
rect 50442 20100 50498 20156
rect 50498 20100 50502 20156
rect 50438 20096 50502 20100
rect 50518 20156 50582 20160
rect 50518 20100 50522 20156
rect 50522 20100 50578 20156
rect 50578 20100 50582 20156
rect 50518 20096 50582 20100
rect 4198 19612 4262 19616
rect 4198 19556 4202 19612
rect 4202 19556 4258 19612
rect 4258 19556 4262 19612
rect 4198 19552 4262 19556
rect 4278 19612 4342 19616
rect 4278 19556 4282 19612
rect 4282 19556 4338 19612
rect 4338 19556 4342 19612
rect 4278 19552 4342 19556
rect 4358 19612 4422 19616
rect 4358 19556 4362 19612
rect 4362 19556 4418 19612
rect 4418 19556 4422 19612
rect 4358 19552 4422 19556
rect 4438 19612 4502 19616
rect 4438 19556 4442 19612
rect 4442 19556 4498 19612
rect 4498 19556 4502 19612
rect 4438 19552 4502 19556
rect 34918 19612 34982 19616
rect 34918 19556 34922 19612
rect 34922 19556 34978 19612
rect 34978 19556 34982 19612
rect 34918 19552 34982 19556
rect 34998 19612 35062 19616
rect 34998 19556 35002 19612
rect 35002 19556 35058 19612
rect 35058 19556 35062 19612
rect 34998 19552 35062 19556
rect 35078 19612 35142 19616
rect 35078 19556 35082 19612
rect 35082 19556 35138 19612
rect 35138 19556 35142 19612
rect 35078 19552 35142 19556
rect 35158 19612 35222 19616
rect 35158 19556 35162 19612
rect 35162 19556 35218 19612
rect 35218 19556 35222 19612
rect 35158 19552 35222 19556
rect 19558 19068 19622 19072
rect 19558 19012 19562 19068
rect 19562 19012 19618 19068
rect 19618 19012 19622 19068
rect 19558 19008 19622 19012
rect 19638 19068 19702 19072
rect 19638 19012 19642 19068
rect 19642 19012 19698 19068
rect 19698 19012 19702 19068
rect 19638 19008 19702 19012
rect 19718 19068 19782 19072
rect 19718 19012 19722 19068
rect 19722 19012 19778 19068
rect 19778 19012 19782 19068
rect 19718 19008 19782 19012
rect 19798 19068 19862 19072
rect 19798 19012 19802 19068
rect 19802 19012 19858 19068
rect 19858 19012 19862 19068
rect 19798 19008 19862 19012
rect 50278 19068 50342 19072
rect 50278 19012 50282 19068
rect 50282 19012 50338 19068
rect 50338 19012 50342 19068
rect 50278 19008 50342 19012
rect 50358 19068 50422 19072
rect 50358 19012 50362 19068
rect 50362 19012 50418 19068
rect 50418 19012 50422 19068
rect 50358 19008 50422 19012
rect 50438 19068 50502 19072
rect 50438 19012 50442 19068
rect 50442 19012 50498 19068
rect 50498 19012 50502 19068
rect 50438 19008 50502 19012
rect 50518 19068 50582 19072
rect 50518 19012 50522 19068
rect 50522 19012 50578 19068
rect 50578 19012 50582 19068
rect 50518 19008 50582 19012
rect 4198 18524 4262 18528
rect 4198 18468 4202 18524
rect 4202 18468 4258 18524
rect 4258 18468 4262 18524
rect 4198 18464 4262 18468
rect 4278 18524 4342 18528
rect 4278 18468 4282 18524
rect 4282 18468 4338 18524
rect 4338 18468 4342 18524
rect 4278 18464 4342 18468
rect 4358 18524 4422 18528
rect 4358 18468 4362 18524
rect 4362 18468 4418 18524
rect 4418 18468 4422 18524
rect 4358 18464 4422 18468
rect 4438 18524 4502 18528
rect 4438 18468 4442 18524
rect 4442 18468 4498 18524
rect 4498 18468 4502 18524
rect 4438 18464 4502 18468
rect 34918 18524 34982 18528
rect 34918 18468 34922 18524
rect 34922 18468 34978 18524
rect 34978 18468 34982 18524
rect 34918 18464 34982 18468
rect 34998 18524 35062 18528
rect 34998 18468 35002 18524
rect 35002 18468 35058 18524
rect 35058 18468 35062 18524
rect 34998 18464 35062 18468
rect 35078 18524 35142 18528
rect 35078 18468 35082 18524
rect 35082 18468 35138 18524
rect 35138 18468 35142 18524
rect 35078 18464 35142 18468
rect 35158 18524 35222 18528
rect 35158 18468 35162 18524
rect 35162 18468 35218 18524
rect 35218 18468 35222 18524
rect 35158 18464 35222 18468
rect 19558 17980 19622 17984
rect 19558 17924 19562 17980
rect 19562 17924 19618 17980
rect 19618 17924 19622 17980
rect 19558 17920 19622 17924
rect 19638 17980 19702 17984
rect 19638 17924 19642 17980
rect 19642 17924 19698 17980
rect 19698 17924 19702 17980
rect 19638 17920 19702 17924
rect 19718 17980 19782 17984
rect 19718 17924 19722 17980
rect 19722 17924 19778 17980
rect 19778 17924 19782 17980
rect 19718 17920 19782 17924
rect 19798 17980 19862 17984
rect 19798 17924 19802 17980
rect 19802 17924 19858 17980
rect 19858 17924 19862 17980
rect 19798 17920 19862 17924
rect 50278 17980 50342 17984
rect 50278 17924 50282 17980
rect 50282 17924 50338 17980
rect 50338 17924 50342 17980
rect 50278 17920 50342 17924
rect 50358 17980 50422 17984
rect 50358 17924 50362 17980
rect 50362 17924 50418 17980
rect 50418 17924 50422 17980
rect 50358 17920 50422 17924
rect 50438 17980 50502 17984
rect 50438 17924 50442 17980
rect 50442 17924 50498 17980
rect 50498 17924 50502 17980
rect 50438 17920 50502 17924
rect 50518 17980 50582 17984
rect 50518 17924 50522 17980
rect 50522 17924 50578 17980
rect 50578 17924 50582 17980
rect 50518 17920 50582 17924
rect 4198 17436 4262 17440
rect 4198 17380 4202 17436
rect 4202 17380 4258 17436
rect 4258 17380 4262 17436
rect 4198 17376 4262 17380
rect 4278 17436 4342 17440
rect 4278 17380 4282 17436
rect 4282 17380 4338 17436
rect 4338 17380 4342 17436
rect 4278 17376 4342 17380
rect 4358 17436 4422 17440
rect 4358 17380 4362 17436
rect 4362 17380 4418 17436
rect 4418 17380 4422 17436
rect 4358 17376 4422 17380
rect 4438 17436 4502 17440
rect 4438 17380 4442 17436
rect 4442 17380 4498 17436
rect 4498 17380 4502 17436
rect 4438 17376 4502 17380
rect 34918 17436 34982 17440
rect 34918 17380 34922 17436
rect 34922 17380 34978 17436
rect 34978 17380 34982 17436
rect 34918 17376 34982 17380
rect 34998 17436 35062 17440
rect 34998 17380 35002 17436
rect 35002 17380 35058 17436
rect 35058 17380 35062 17436
rect 34998 17376 35062 17380
rect 35078 17436 35142 17440
rect 35078 17380 35082 17436
rect 35082 17380 35138 17436
rect 35138 17380 35142 17436
rect 35078 17376 35142 17380
rect 35158 17436 35222 17440
rect 35158 17380 35162 17436
rect 35162 17380 35218 17436
rect 35218 17380 35222 17436
rect 35158 17376 35222 17380
rect 19558 16892 19622 16896
rect 19558 16836 19562 16892
rect 19562 16836 19618 16892
rect 19618 16836 19622 16892
rect 19558 16832 19622 16836
rect 19638 16892 19702 16896
rect 19638 16836 19642 16892
rect 19642 16836 19698 16892
rect 19698 16836 19702 16892
rect 19638 16832 19702 16836
rect 19718 16892 19782 16896
rect 19718 16836 19722 16892
rect 19722 16836 19778 16892
rect 19778 16836 19782 16892
rect 19718 16832 19782 16836
rect 19798 16892 19862 16896
rect 19798 16836 19802 16892
rect 19802 16836 19858 16892
rect 19858 16836 19862 16892
rect 19798 16832 19862 16836
rect 50278 16892 50342 16896
rect 50278 16836 50282 16892
rect 50282 16836 50338 16892
rect 50338 16836 50342 16892
rect 50278 16832 50342 16836
rect 50358 16892 50422 16896
rect 50358 16836 50362 16892
rect 50362 16836 50418 16892
rect 50418 16836 50422 16892
rect 50358 16832 50422 16836
rect 50438 16892 50502 16896
rect 50438 16836 50442 16892
rect 50442 16836 50498 16892
rect 50498 16836 50502 16892
rect 50438 16832 50502 16836
rect 50518 16892 50582 16896
rect 50518 16836 50522 16892
rect 50522 16836 50578 16892
rect 50578 16836 50582 16892
rect 50518 16832 50582 16836
rect 4198 16348 4262 16352
rect 4198 16292 4202 16348
rect 4202 16292 4258 16348
rect 4258 16292 4262 16348
rect 4198 16288 4262 16292
rect 4278 16348 4342 16352
rect 4278 16292 4282 16348
rect 4282 16292 4338 16348
rect 4338 16292 4342 16348
rect 4278 16288 4342 16292
rect 4358 16348 4422 16352
rect 4358 16292 4362 16348
rect 4362 16292 4418 16348
rect 4418 16292 4422 16348
rect 4358 16288 4422 16292
rect 4438 16348 4502 16352
rect 4438 16292 4442 16348
rect 4442 16292 4498 16348
rect 4498 16292 4502 16348
rect 4438 16288 4502 16292
rect 34918 16348 34982 16352
rect 34918 16292 34922 16348
rect 34922 16292 34978 16348
rect 34978 16292 34982 16348
rect 34918 16288 34982 16292
rect 34998 16348 35062 16352
rect 34998 16292 35002 16348
rect 35002 16292 35058 16348
rect 35058 16292 35062 16348
rect 34998 16288 35062 16292
rect 35078 16348 35142 16352
rect 35078 16292 35082 16348
rect 35082 16292 35138 16348
rect 35138 16292 35142 16348
rect 35078 16288 35142 16292
rect 35158 16348 35222 16352
rect 35158 16292 35162 16348
rect 35162 16292 35218 16348
rect 35218 16292 35222 16348
rect 35158 16288 35222 16292
rect 19558 15804 19622 15808
rect 19558 15748 19562 15804
rect 19562 15748 19618 15804
rect 19618 15748 19622 15804
rect 19558 15744 19622 15748
rect 19638 15804 19702 15808
rect 19638 15748 19642 15804
rect 19642 15748 19698 15804
rect 19698 15748 19702 15804
rect 19638 15744 19702 15748
rect 19718 15804 19782 15808
rect 19718 15748 19722 15804
rect 19722 15748 19778 15804
rect 19778 15748 19782 15804
rect 19718 15744 19782 15748
rect 19798 15804 19862 15808
rect 19798 15748 19802 15804
rect 19802 15748 19858 15804
rect 19858 15748 19862 15804
rect 19798 15744 19862 15748
rect 50278 15804 50342 15808
rect 50278 15748 50282 15804
rect 50282 15748 50338 15804
rect 50338 15748 50342 15804
rect 50278 15744 50342 15748
rect 50358 15804 50422 15808
rect 50358 15748 50362 15804
rect 50362 15748 50418 15804
rect 50418 15748 50422 15804
rect 50358 15744 50422 15748
rect 50438 15804 50502 15808
rect 50438 15748 50442 15804
rect 50442 15748 50498 15804
rect 50498 15748 50502 15804
rect 50438 15744 50502 15748
rect 50518 15804 50582 15808
rect 50518 15748 50522 15804
rect 50522 15748 50578 15804
rect 50578 15748 50582 15804
rect 50518 15744 50582 15748
rect 4198 15260 4262 15264
rect 4198 15204 4202 15260
rect 4202 15204 4258 15260
rect 4258 15204 4262 15260
rect 4198 15200 4262 15204
rect 4278 15260 4342 15264
rect 4278 15204 4282 15260
rect 4282 15204 4338 15260
rect 4338 15204 4342 15260
rect 4278 15200 4342 15204
rect 4358 15260 4422 15264
rect 4358 15204 4362 15260
rect 4362 15204 4418 15260
rect 4418 15204 4422 15260
rect 4358 15200 4422 15204
rect 4438 15260 4502 15264
rect 4438 15204 4442 15260
rect 4442 15204 4498 15260
rect 4498 15204 4502 15260
rect 4438 15200 4502 15204
rect 34918 15260 34982 15264
rect 34918 15204 34922 15260
rect 34922 15204 34978 15260
rect 34978 15204 34982 15260
rect 34918 15200 34982 15204
rect 34998 15260 35062 15264
rect 34998 15204 35002 15260
rect 35002 15204 35058 15260
rect 35058 15204 35062 15260
rect 34998 15200 35062 15204
rect 35078 15260 35142 15264
rect 35078 15204 35082 15260
rect 35082 15204 35138 15260
rect 35138 15204 35142 15260
rect 35078 15200 35142 15204
rect 35158 15260 35222 15264
rect 35158 15204 35162 15260
rect 35162 15204 35218 15260
rect 35218 15204 35222 15260
rect 35158 15200 35222 15204
rect 19558 14716 19622 14720
rect 19558 14660 19562 14716
rect 19562 14660 19618 14716
rect 19618 14660 19622 14716
rect 19558 14656 19622 14660
rect 19638 14716 19702 14720
rect 19638 14660 19642 14716
rect 19642 14660 19698 14716
rect 19698 14660 19702 14716
rect 19638 14656 19702 14660
rect 19718 14716 19782 14720
rect 19718 14660 19722 14716
rect 19722 14660 19778 14716
rect 19778 14660 19782 14716
rect 19718 14656 19782 14660
rect 19798 14716 19862 14720
rect 19798 14660 19802 14716
rect 19802 14660 19858 14716
rect 19858 14660 19862 14716
rect 19798 14656 19862 14660
rect 50278 14716 50342 14720
rect 50278 14660 50282 14716
rect 50282 14660 50338 14716
rect 50338 14660 50342 14716
rect 50278 14656 50342 14660
rect 50358 14716 50422 14720
rect 50358 14660 50362 14716
rect 50362 14660 50418 14716
rect 50418 14660 50422 14716
rect 50358 14656 50422 14660
rect 50438 14716 50502 14720
rect 50438 14660 50442 14716
rect 50442 14660 50498 14716
rect 50498 14660 50502 14716
rect 50438 14656 50502 14660
rect 50518 14716 50582 14720
rect 50518 14660 50522 14716
rect 50522 14660 50578 14716
rect 50578 14660 50582 14716
rect 50518 14656 50582 14660
rect 4198 14172 4262 14176
rect 4198 14116 4202 14172
rect 4202 14116 4258 14172
rect 4258 14116 4262 14172
rect 4198 14112 4262 14116
rect 4278 14172 4342 14176
rect 4278 14116 4282 14172
rect 4282 14116 4338 14172
rect 4338 14116 4342 14172
rect 4278 14112 4342 14116
rect 4358 14172 4422 14176
rect 4358 14116 4362 14172
rect 4362 14116 4418 14172
rect 4418 14116 4422 14172
rect 4358 14112 4422 14116
rect 4438 14172 4502 14176
rect 4438 14116 4442 14172
rect 4442 14116 4498 14172
rect 4498 14116 4502 14172
rect 4438 14112 4502 14116
rect 34918 14172 34982 14176
rect 34918 14116 34922 14172
rect 34922 14116 34978 14172
rect 34978 14116 34982 14172
rect 34918 14112 34982 14116
rect 34998 14172 35062 14176
rect 34998 14116 35002 14172
rect 35002 14116 35058 14172
rect 35058 14116 35062 14172
rect 34998 14112 35062 14116
rect 35078 14172 35142 14176
rect 35078 14116 35082 14172
rect 35082 14116 35138 14172
rect 35138 14116 35142 14172
rect 35078 14112 35142 14116
rect 35158 14172 35222 14176
rect 35158 14116 35162 14172
rect 35162 14116 35218 14172
rect 35218 14116 35222 14172
rect 35158 14112 35222 14116
rect 19558 13628 19622 13632
rect 19558 13572 19562 13628
rect 19562 13572 19618 13628
rect 19618 13572 19622 13628
rect 19558 13568 19622 13572
rect 19638 13628 19702 13632
rect 19638 13572 19642 13628
rect 19642 13572 19698 13628
rect 19698 13572 19702 13628
rect 19638 13568 19702 13572
rect 19718 13628 19782 13632
rect 19718 13572 19722 13628
rect 19722 13572 19778 13628
rect 19778 13572 19782 13628
rect 19718 13568 19782 13572
rect 19798 13628 19862 13632
rect 19798 13572 19802 13628
rect 19802 13572 19858 13628
rect 19858 13572 19862 13628
rect 19798 13568 19862 13572
rect 50278 13628 50342 13632
rect 50278 13572 50282 13628
rect 50282 13572 50338 13628
rect 50338 13572 50342 13628
rect 50278 13568 50342 13572
rect 50358 13628 50422 13632
rect 50358 13572 50362 13628
rect 50362 13572 50418 13628
rect 50418 13572 50422 13628
rect 50358 13568 50422 13572
rect 50438 13628 50502 13632
rect 50438 13572 50442 13628
rect 50442 13572 50498 13628
rect 50498 13572 50502 13628
rect 50438 13568 50502 13572
rect 50518 13628 50582 13632
rect 50518 13572 50522 13628
rect 50522 13572 50578 13628
rect 50578 13572 50582 13628
rect 50518 13568 50582 13572
rect 4198 13084 4262 13088
rect 4198 13028 4202 13084
rect 4202 13028 4258 13084
rect 4258 13028 4262 13084
rect 4198 13024 4262 13028
rect 4278 13084 4342 13088
rect 4278 13028 4282 13084
rect 4282 13028 4338 13084
rect 4338 13028 4342 13084
rect 4278 13024 4342 13028
rect 4358 13084 4422 13088
rect 4358 13028 4362 13084
rect 4362 13028 4418 13084
rect 4418 13028 4422 13084
rect 4358 13024 4422 13028
rect 4438 13084 4502 13088
rect 4438 13028 4442 13084
rect 4442 13028 4498 13084
rect 4498 13028 4502 13084
rect 4438 13024 4502 13028
rect 34918 13084 34982 13088
rect 34918 13028 34922 13084
rect 34922 13028 34978 13084
rect 34978 13028 34982 13084
rect 34918 13024 34982 13028
rect 34998 13084 35062 13088
rect 34998 13028 35002 13084
rect 35002 13028 35058 13084
rect 35058 13028 35062 13084
rect 34998 13024 35062 13028
rect 35078 13084 35142 13088
rect 35078 13028 35082 13084
rect 35082 13028 35138 13084
rect 35138 13028 35142 13084
rect 35078 13024 35142 13028
rect 35158 13084 35222 13088
rect 35158 13028 35162 13084
rect 35162 13028 35218 13084
rect 35218 13028 35222 13084
rect 35158 13024 35222 13028
rect 19558 12540 19622 12544
rect 19558 12484 19562 12540
rect 19562 12484 19618 12540
rect 19618 12484 19622 12540
rect 19558 12480 19622 12484
rect 19638 12540 19702 12544
rect 19638 12484 19642 12540
rect 19642 12484 19698 12540
rect 19698 12484 19702 12540
rect 19638 12480 19702 12484
rect 19718 12540 19782 12544
rect 19718 12484 19722 12540
rect 19722 12484 19778 12540
rect 19778 12484 19782 12540
rect 19718 12480 19782 12484
rect 19798 12540 19862 12544
rect 19798 12484 19802 12540
rect 19802 12484 19858 12540
rect 19858 12484 19862 12540
rect 19798 12480 19862 12484
rect 50278 12540 50342 12544
rect 50278 12484 50282 12540
rect 50282 12484 50338 12540
rect 50338 12484 50342 12540
rect 50278 12480 50342 12484
rect 50358 12540 50422 12544
rect 50358 12484 50362 12540
rect 50362 12484 50418 12540
rect 50418 12484 50422 12540
rect 50358 12480 50422 12484
rect 50438 12540 50502 12544
rect 50438 12484 50442 12540
rect 50442 12484 50498 12540
rect 50498 12484 50502 12540
rect 50438 12480 50502 12484
rect 50518 12540 50582 12544
rect 50518 12484 50522 12540
rect 50522 12484 50578 12540
rect 50578 12484 50582 12540
rect 50518 12480 50582 12484
rect 4198 11996 4262 12000
rect 4198 11940 4202 11996
rect 4202 11940 4258 11996
rect 4258 11940 4262 11996
rect 4198 11936 4262 11940
rect 4278 11996 4342 12000
rect 4278 11940 4282 11996
rect 4282 11940 4338 11996
rect 4338 11940 4342 11996
rect 4278 11936 4342 11940
rect 4358 11996 4422 12000
rect 4358 11940 4362 11996
rect 4362 11940 4418 11996
rect 4418 11940 4422 11996
rect 4358 11936 4422 11940
rect 4438 11996 4502 12000
rect 4438 11940 4442 11996
rect 4442 11940 4498 11996
rect 4498 11940 4502 11996
rect 4438 11936 4502 11940
rect 34918 11996 34982 12000
rect 34918 11940 34922 11996
rect 34922 11940 34978 11996
rect 34978 11940 34982 11996
rect 34918 11936 34982 11940
rect 34998 11996 35062 12000
rect 34998 11940 35002 11996
rect 35002 11940 35058 11996
rect 35058 11940 35062 11996
rect 34998 11936 35062 11940
rect 35078 11996 35142 12000
rect 35078 11940 35082 11996
rect 35082 11940 35138 11996
rect 35138 11940 35142 11996
rect 35078 11936 35142 11940
rect 35158 11996 35222 12000
rect 35158 11940 35162 11996
rect 35162 11940 35218 11996
rect 35218 11940 35222 11996
rect 35158 11936 35222 11940
rect 19558 11452 19622 11456
rect 19558 11396 19562 11452
rect 19562 11396 19618 11452
rect 19618 11396 19622 11452
rect 19558 11392 19622 11396
rect 19638 11452 19702 11456
rect 19638 11396 19642 11452
rect 19642 11396 19698 11452
rect 19698 11396 19702 11452
rect 19638 11392 19702 11396
rect 19718 11452 19782 11456
rect 19718 11396 19722 11452
rect 19722 11396 19778 11452
rect 19778 11396 19782 11452
rect 19718 11392 19782 11396
rect 19798 11452 19862 11456
rect 19798 11396 19802 11452
rect 19802 11396 19858 11452
rect 19858 11396 19862 11452
rect 19798 11392 19862 11396
rect 50278 11452 50342 11456
rect 50278 11396 50282 11452
rect 50282 11396 50338 11452
rect 50338 11396 50342 11452
rect 50278 11392 50342 11396
rect 50358 11452 50422 11456
rect 50358 11396 50362 11452
rect 50362 11396 50418 11452
rect 50418 11396 50422 11452
rect 50358 11392 50422 11396
rect 50438 11452 50502 11456
rect 50438 11396 50442 11452
rect 50442 11396 50498 11452
rect 50498 11396 50502 11452
rect 50438 11392 50502 11396
rect 50518 11452 50582 11456
rect 50518 11396 50522 11452
rect 50522 11396 50578 11452
rect 50578 11396 50582 11452
rect 50518 11392 50582 11396
rect 4198 10908 4262 10912
rect 4198 10852 4202 10908
rect 4202 10852 4258 10908
rect 4258 10852 4262 10908
rect 4198 10848 4262 10852
rect 4278 10908 4342 10912
rect 4278 10852 4282 10908
rect 4282 10852 4338 10908
rect 4338 10852 4342 10908
rect 4278 10848 4342 10852
rect 4358 10908 4422 10912
rect 4358 10852 4362 10908
rect 4362 10852 4418 10908
rect 4418 10852 4422 10908
rect 4358 10848 4422 10852
rect 4438 10908 4502 10912
rect 4438 10852 4442 10908
rect 4442 10852 4498 10908
rect 4498 10852 4502 10908
rect 4438 10848 4502 10852
rect 34918 10908 34982 10912
rect 34918 10852 34922 10908
rect 34922 10852 34978 10908
rect 34978 10852 34982 10908
rect 34918 10848 34982 10852
rect 34998 10908 35062 10912
rect 34998 10852 35002 10908
rect 35002 10852 35058 10908
rect 35058 10852 35062 10908
rect 34998 10848 35062 10852
rect 35078 10908 35142 10912
rect 35078 10852 35082 10908
rect 35082 10852 35138 10908
rect 35138 10852 35142 10908
rect 35078 10848 35142 10852
rect 35158 10908 35222 10912
rect 35158 10852 35162 10908
rect 35162 10852 35218 10908
rect 35218 10852 35222 10908
rect 35158 10848 35222 10852
rect 19558 10364 19622 10368
rect 19558 10308 19562 10364
rect 19562 10308 19618 10364
rect 19618 10308 19622 10364
rect 19558 10304 19622 10308
rect 19638 10364 19702 10368
rect 19638 10308 19642 10364
rect 19642 10308 19698 10364
rect 19698 10308 19702 10364
rect 19638 10304 19702 10308
rect 19718 10364 19782 10368
rect 19718 10308 19722 10364
rect 19722 10308 19778 10364
rect 19778 10308 19782 10364
rect 19718 10304 19782 10308
rect 19798 10364 19862 10368
rect 19798 10308 19802 10364
rect 19802 10308 19858 10364
rect 19858 10308 19862 10364
rect 19798 10304 19862 10308
rect 50278 10364 50342 10368
rect 50278 10308 50282 10364
rect 50282 10308 50338 10364
rect 50338 10308 50342 10364
rect 50278 10304 50342 10308
rect 50358 10364 50422 10368
rect 50358 10308 50362 10364
rect 50362 10308 50418 10364
rect 50418 10308 50422 10364
rect 50358 10304 50422 10308
rect 50438 10364 50502 10368
rect 50438 10308 50442 10364
rect 50442 10308 50498 10364
rect 50498 10308 50502 10364
rect 50438 10304 50502 10308
rect 50518 10364 50582 10368
rect 50518 10308 50522 10364
rect 50522 10308 50578 10364
rect 50578 10308 50582 10364
rect 50518 10304 50582 10308
rect 4198 9820 4262 9824
rect 4198 9764 4202 9820
rect 4202 9764 4258 9820
rect 4258 9764 4262 9820
rect 4198 9760 4262 9764
rect 4278 9820 4342 9824
rect 4278 9764 4282 9820
rect 4282 9764 4338 9820
rect 4338 9764 4342 9820
rect 4278 9760 4342 9764
rect 4358 9820 4422 9824
rect 4358 9764 4362 9820
rect 4362 9764 4418 9820
rect 4418 9764 4422 9820
rect 4358 9760 4422 9764
rect 4438 9820 4502 9824
rect 4438 9764 4442 9820
rect 4442 9764 4498 9820
rect 4498 9764 4502 9820
rect 4438 9760 4502 9764
rect 34918 9820 34982 9824
rect 34918 9764 34922 9820
rect 34922 9764 34978 9820
rect 34978 9764 34982 9820
rect 34918 9760 34982 9764
rect 34998 9820 35062 9824
rect 34998 9764 35002 9820
rect 35002 9764 35058 9820
rect 35058 9764 35062 9820
rect 34998 9760 35062 9764
rect 35078 9820 35142 9824
rect 35078 9764 35082 9820
rect 35082 9764 35138 9820
rect 35138 9764 35142 9820
rect 35078 9760 35142 9764
rect 35158 9820 35222 9824
rect 35158 9764 35162 9820
rect 35162 9764 35218 9820
rect 35218 9764 35222 9820
rect 35158 9760 35222 9764
rect 19558 9276 19622 9280
rect 19558 9220 19562 9276
rect 19562 9220 19618 9276
rect 19618 9220 19622 9276
rect 19558 9216 19622 9220
rect 19638 9276 19702 9280
rect 19638 9220 19642 9276
rect 19642 9220 19698 9276
rect 19698 9220 19702 9276
rect 19638 9216 19702 9220
rect 19718 9276 19782 9280
rect 19718 9220 19722 9276
rect 19722 9220 19778 9276
rect 19778 9220 19782 9276
rect 19718 9216 19782 9220
rect 19798 9276 19862 9280
rect 19798 9220 19802 9276
rect 19802 9220 19858 9276
rect 19858 9220 19862 9276
rect 19798 9216 19862 9220
rect 50278 9276 50342 9280
rect 50278 9220 50282 9276
rect 50282 9220 50338 9276
rect 50338 9220 50342 9276
rect 50278 9216 50342 9220
rect 50358 9276 50422 9280
rect 50358 9220 50362 9276
rect 50362 9220 50418 9276
rect 50418 9220 50422 9276
rect 50358 9216 50422 9220
rect 50438 9276 50502 9280
rect 50438 9220 50442 9276
rect 50442 9220 50498 9276
rect 50498 9220 50502 9276
rect 50438 9216 50502 9220
rect 50518 9276 50582 9280
rect 50518 9220 50522 9276
rect 50522 9220 50578 9276
rect 50578 9220 50582 9276
rect 50518 9216 50582 9220
rect 4198 8732 4262 8736
rect 4198 8676 4202 8732
rect 4202 8676 4258 8732
rect 4258 8676 4262 8732
rect 4198 8672 4262 8676
rect 4278 8732 4342 8736
rect 4278 8676 4282 8732
rect 4282 8676 4338 8732
rect 4338 8676 4342 8732
rect 4278 8672 4342 8676
rect 4358 8732 4422 8736
rect 4358 8676 4362 8732
rect 4362 8676 4418 8732
rect 4418 8676 4422 8732
rect 4358 8672 4422 8676
rect 4438 8732 4502 8736
rect 4438 8676 4442 8732
rect 4442 8676 4498 8732
rect 4498 8676 4502 8732
rect 4438 8672 4502 8676
rect 34918 8732 34982 8736
rect 34918 8676 34922 8732
rect 34922 8676 34978 8732
rect 34978 8676 34982 8732
rect 34918 8672 34982 8676
rect 34998 8732 35062 8736
rect 34998 8676 35002 8732
rect 35002 8676 35058 8732
rect 35058 8676 35062 8732
rect 34998 8672 35062 8676
rect 35078 8732 35142 8736
rect 35078 8676 35082 8732
rect 35082 8676 35138 8732
rect 35138 8676 35142 8732
rect 35078 8672 35142 8676
rect 35158 8732 35222 8736
rect 35158 8676 35162 8732
rect 35162 8676 35218 8732
rect 35218 8676 35222 8732
rect 35158 8672 35222 8676
rect 19558 8188 19622 8192
rect 19558 8132 19562 8188
rect 19562 8132 19618 8188
rect 19618 8132 19622 8188
rect 19558 8128 19622 8132
rect 19638 8188 19702 8192
rect 19638 8132 19642 8188
rect 19642 8132 19698 8188
rect 19698 8132 19702 8188
rect 19638 8128 19702 8132
rect 19718 8188 19782 8192
rect 19718 8132 19722 8188
rect 19722 8132 19778 8188
rect 19778 8132 19782 8188
rect 19718 8128 19782 8132
rect 19798 8188 19862 8192
rect 19798 8132 19802 8188
rect 19802 8132 19858 8188
rect 19858 8132 19862 8188
rect 19798 8128 19862 8132
rect 50278 8188 50342 8192
rect 50278 8132 50282 8188
rect 50282 8132 50338 8188
rect 50338 8132 50342 8188
rect 50278 8128 50342 8132
rect 50358 8188 50422 8192
rect 50358 8132 50362 8188
rect 50362 8132 50418 8188
rect 50418 8132 50422 8188
rect 50358 8128 50422 8132
rect 50438 8188 50502 8192
rect 50438 8132 50442 8188
rect 50442 8132 50498 8188
rect 50498 8132 50502 8188
rect 50438 8128 50502 8132
rect 50518 8188 50582 8192
rect 50518 8132 50522 8188
rect 50522 8132 50578 8188
rect 50578 8132 50582 8188
rect 50518 8128 50582 8132
rect 4198 7644 4262 7648
rect 4198 7588 4202 7644
rect 4202 7588 4258 7644
rect 4258 7588 4262 7644
rect 4198 7584 4262 7588
rect 4278 7644 4342 7648
rect 4278 7588 4282 7644
rect 4282 7588 4338 7644
rect 4338 7588 4342 7644
rect 4278 7584 4342 7588
rect 4358 7644 4422 7648
rect 4358 7588 4362 7644
rect 4362 7588 4418 7644
rect 4418 7588 4422 7644
rect 4358 7584 4422 7588
rect 4438 7644 4502 7648
rect 4438 7588 4442 7644
rect 4442 7588 4498 7644
rect 4498 7588 4502 7644
rect 4438 7584 4502 7588
rect 34918 7644 34982 7648
rect 34918 7588 34922 7644
rect 34922 7588 34978 7644
rect 34978 7588 34982 7644
rect 34918 7584 34982 7588
rect 34998 7644 35062 7648
rect 34998 7588 35002 7644
rect 35002 7588 35058 7644
rect 35058 7588 35062 7644
rect 34998 7584 35062 7588
rect 35078 7644 35142 7648
rect 35078 7588 35082 7644
rect 35082 7588 35138 7644
rect 35138 7588 35142 7644
rect 35078 7584 35142 7588
rect 35158 7644 35222 7648
rect 35158 7588 35162 7644
rect 35162 7588 35218 7644
rect 35218 7588 35222 7644
rect 35158 7584 35222 7588
rect 19558 7100 19622 7104
rect 19558 7044 19562 7100
rect 19562 7044 19618 7100
rect 19618 7044 19622 7100
rect 19558 7040 19622 7044
rect 19638 7100 19702 7104
rect 19638 7044 19642 7100
rect 19642 7044 19698 7100
rect 19698 7044 19702 7100
rect 19638 7040 19702 7044
rect 19718 7100 19782 7104
rect 19718 7044 19722 7100
rect 19722 7044 19778 7100
rect 19778 7044 19782 7100
rect 19718 7040 19782 7044
rect 19798 7100 19862 7104
rect 19798 7044 19802 7100
rect 19802 7044 19858 7100
rect 19858 7044 19862 7100
rect 19798 7040 19862 7044
rect 50278 7100 50342 7104
rect 50278 7044 50282 7100
rect 50282 7044 50338 7100
rect 50338 7044 50342 7100
rect 50278 7040 50342 7044
rect 50358 7100 50422 7104
rect 50358 7044 50362 7100
rect 50362 7044 50418 7100
rect 50418 7044 50422 7100
rect 50358 7040 50422 7044
rect 50438 7100 50502 7104
rect 50438 7044 50442 7100
rect 50442 7044 50498 7100
rect 50498 7044 50502 7100
rect 50438 7040 50502 7044
rect 50518 7100 50582 7104
rect 50518 7044 50522 7100
rect 50522 7044 50578 7100
rect 50578 7044 50582 7100
rect 50518 7040 50582 7044
rect 4198 6556 4262 6560
rect 4198 6500 4202 6556
rect 4202 6500 4258 6556
rect 4258 6500 4262 6556
rect 4198 6496 4262 6500
rect 4278 6556 4342 6560
rect 4278 6500 4282 6556
rect 4282 6500 4338 6556
rect 4338 6500 4342 6556
rect 4278 6496 4342 6500
rect 4358 6556 4422 6560
rect 4358 6500 4362 6556
rect 4362 6500 4418 6556
rect 4418 6500 4422 6556
rect 4358 6496 4422 6500
rect 4438 6556 4502 6560
rect 4438 6500 4442 6556
rect 4442 6500 4498 6556
rect 4498 6500 4502 6556
rect 4438 6496 4502 6500
rect 34918 6556 34982 6560
rect 34918 6500 34922 6556
rect 34922 6500 34978 6556
rect 34978 6500 34982 6556
rect 34918 6496 34982 6500
rect 34998 6556 35062 6560
rect 34998 6500 35002 6556
rect 35002 6500 35058 6556
rect 35058 6500 35062 6556
rect 34998 6496 35062 6500
rect 35078 6556 35142 6560
rect 35078 6500 35082 6556
rect 35082 6500 35138 6556
rect 35138 6500 35142 6556
rect 35078 6496 35142 6500
rect 35158 6556 35222 6560
rect 35158 6500 35162 6556
rect 35162 6500 35218 6556
rect 35218 6500 35222 6556
rect 35158 6496 35222 6500
rect 19558 6012 19622 6016
rect 19558 5956 19562 6012
rect 19562 5956 19618 6012
rect 19618 5956 19622 6012
rect 19558 5952 19622 5956
rect 19638 6012 19702 6016
rect 19638 5956 19642 6012
rect 19642 5956 19698 6012
rect 19698 5956 19702 6012
rect 19638 5952 19702 5956
rect 19718 6012 19782 6016
rect 19718 5956 19722 6012
rect 19722 5956 19778 6012
rect 19778 5956 19782 6012
rect 19718 5952 19782 5956
rect 19798 6012 19862 6016
rect 19798 5956 19802 6012
rect 19802 5956 19858 6012
rect 19858 5956 19862 6012
rect 19798 5952 19862 5956
rect 50278 6012 50342 6016
rect 50278 5956 50282 6012
rect 50282 5956 50338 6012
rect 50338 5956 50342 6012
rect 50278 5952 50342 5956
rect 50358 6012 50422 6016
rect 50358 5956 50362 6012
rect 50362 5956 50418 6012
rect 50418 5956 50422 6012
rect 50358 5952 50422 5956
rect 50438 6012 50502 6016
rect 50438 5956 50442 6012
rect 50442 5956 50498 6012
rect 50498 5956 50502 6012
rect 50438 5952 50502 5956
rect 50518 6012 50582 6016
rect 50518 5956 50522 6012
rect 50522 5956 50578 6012
rect 50578 5956 50582 6012
rect 50518 5952 50582 5956
rect 4198 5468 4262 5472
rect 4198 5412 4202 5468
rect 4202 5412 4258 5468
rect 4258 5412 4262 5468
rect 4198 5408 4262 5412
rect 4278 5468 4342 5472
rect 4278 5412 4282 5468
rect 4282 5412 4338 5468
rect 4338 5412 4342 5468
rect 4278 5408 4342 5412
rect 4358 5468 4422 5472
rect 4358 5412 4362 5468
rect 4362 5412 4418 5468
rect 4418 5412 4422 5468
rect 4358 5408 4422 5412
rect 4438 5468 4502 5472
rect 4438 5412 4442 5468
rect 4442 5412 4498 5468
rect 4498 5412 4502 5468
rect 4438 5408 4502 5412
rect 34918 5468 34982 5472
rect 34918 5412 34922 5468
rect 34922 5412 34978 5468
rect 34978 5412 34982 5468
rect 34918 5408 34982 5412
rect 34998 5468 35062 5472
rect 34998 5412 35002 5468
rect 35002 5412 35058 5468
rect 35058 5412 35062 5468
rect 34998 5408 35062 5412
rect 35078 5468 35142 5472
rect 35078 5412 35082 5468
rect 35082 5412 35138 5468
rect 35138 5412 35142 5468
rect 35078 5408 35142 5412
rect 35158 5468 35222 5472
rect 35158 5412 35162 5468
rect 35162 5412 35218 5468
rect 35218 5412 35222 5468
rect 35158 5408 35222 5412
rect 19558 4924 19622 4928
rect 19558 4868 19562 4924
rect 19562 4868 19618 4924
rect 19618 4868 19622 4924
rect 19558 4864 19622 4868
rect 19638 4924 19702 4928
rect 19638 4868 19642 4924
rect 19642 4868 19698 4924
rect 19698 4868 19702 4924
rect 19638 4864 19702 4868
rect 19718 4924 19782 4928
rect 19718 4868 19722 4924
rect 19722 4868 19778 4924
rect 19778 4868 19782 4924
rect 19718 4864 19782 4868
rect 19798 4924 19862 4928
rect 19798 4868 19802 4924
rect 19802 4868 19858 4924
rect 19858 4868 19862 4924
rect 19798 4864 19862 4868
rect 50278 4924 50342 4928
rect 50278 4868 50282 4924
rect 50282 4868 50338 4924
rect 50338 4868 50342 4924
rect 50278 4864 50342 4868
rect 50358 4924 50422 4928
rect 50358 4868 50362 4924
rect 50362 4868 50418 4924
rect 50418 4868 50422 4924
rect 50358 4864 50422 4868
rect 50438 4924 50502 4928
rect 50438 4868 50442 4924
rect 50442 4868 50498 4924
rect 50498 4868 50502 4924
rect 50438 4864 50502 4868
rect 50518 4924 50582 4928
rect 50518 4868 50522 4924
rect 50522 4868 50578 4924
rect 50578 4868 50582 4924
rect 50518 4864 50582 4868
rect 4198 4380 4262 4384
rect 4198 4324 4202 4380
rect 4202 4324 4258 4380
rect 4258 4324 4262 4380
rect 4198 4320 4262 4324
rect 4278 4380 4342 4384
rect 4278 4324 4282 4380
rect 4282 4324 4338 4380
rect 4338 4324 4342 4380
rect 4278 4320 4342 4324
rect 4358 4380 4422 4384
rect 4358 4324 4362 4380
rect 4362 4324 4418 4380
rect 4418 4324 4422 4380
rect 4358 4320 4422 4324
rect 4438 4380 4502 4384
rect 4438 4324 4442 4380
rect 4442 4324 4498 4380
rect 4498 4324 4502 4380
rect 4438 4320 4502 4324
rect 34918 4380 34982 4384
rect 34918 4324 34922 4380
rect 34922 4324 34978 4380
rect 34978 4324 34982 4380
rect 34918 4320 34982 4324
rect 34998 4380 35062 4384
rect 34998 4324 35002 4380
rect 35002 4324 35058 4380
rect 35058 4324 35062 4380
rect 34998 4320 35062 4324
rect 35078 4380 35142 4384
rect 35078 4324 35082 4380
rect 35082 4324 35138 4380
rect 35138 4324 35142 4380
rect 35078 4320 35142 4324
rect 35158 4380 35222 4384
rect 35158 4324 35162 4380
rect 35162 4324 35218 4380
rect 35218 4324 35222 4380
rect 35158 4320 35222 4324
rect 19558 3836 19622 3840
rect 19558 3780 19562 3836
rect 19562 3780 19618 3836
rect 19618 3780 19622 3836
rect 19558 3776 19622 3780
rect 19638 3836 19702 3840
rect 19638 3780 19642 3836
rect 19642 3780 19698 3836
rect 19698 3780 19702 3836
rect 19638 3776 19702 3780
rect 19718 3836 19782 3840
rect 19718 3780 19722 3836
rect 19722 3780 19778 3836
rect 19778 3780 19782 3836
rect 19718 3776 19782 3780
rect 19798 3836 19862 3840
rect 19798 3780 19802 3836
rect 19802 3780 19858 3836
rect 19858 3780 19862 3836
rect 19798 3776 19862 3780
rect 50278 3836 50342 3840
rect 50278 3780 50282 3836
rect 50282 3780 50338 3836
rect 50338 3780 50342 3836
rect 50278 3776 50342 3780
rect 50358 3836 50422 3840
rect 50358 3780 50362 3836
rect 50362 3780 50418 3836
rect 50418 3780 50422 3836
rect 50358 3776 50422 3780
rect 50438 3836 50502 3840
rect 50438 3780 50442 3836
rect 50442 3780 50498 3836
rect 50498 3780 50502 3836
rect 50438 3776 50502 3780
rect 50518 3836 50582 3840
rect 50518 3780 50522 3836
rect 50522 3780 50578 3836
rect 50578 3780 50582 3836
rect 50518 3776 50582 3780
rect 4198 3292 4262 3296
rect 4198 3236 4202 3292
rect 4202 3236 4258 3292
rect 4258 3236 4262 3292
rect 4198 3232 4262 3236
rect 4278 3292 4342 3296
rect 4278 3236 4282 3292
rect 4282 3236 4338 3292
rect 4338 3236 4342 3292
rect 4278 3232 4342 3236
rect 4358 3292 4422 3296
rect 4358 3236 4362 3292
rect 4362 3236 4418 3292
rect 4418 3236 4422 3292
rect 4358 3232 4422 3236
rect 4438 3292 4502 3296
rect 4438 3236 4442 3292
rect 4442 3236 4498 3292
rect 4498 3236 4502 3292
rect 4438 3232 4502 3236
rect 34918 3292 34982 3296
rect 34918 3236 34922 3292
rect 34922 3236 34978 3292
rect 34978 3236 34982 3292
rect 34918 3232 34982 3236
rect 34998 3292 35062 3296
rect 34998 3236 35002 3292
rect 35002 3236 35058 3292
rect 35058 3236 35062 3292
rect 34998 3232 35062 3236
rect 35078 3292 35142 3296
rect 35078 3236 35082 3292
rect 35082 3236 35138 3292
rect 35138 3236 35142 3292
rect 35078 3232 35142 3236
rect 35158 3292 35222 3296
rect 35158 3236 35162 3292
rect 35162 3236 35218 3292
rect 35218 3236 35222 3292
rect 35158 3232 35222 3236
rect 19558 2748 19622 2752
rect 19558 2692 19562 2748
rect 19562 2692 19618 2748
rect 19618 2692 19622 2748
rect 19558 2688 19622 2692
rect 19638 2748 19702 2752
rect 19638 2692 19642 2748
rect 19642 2692 19698 2748
rect 19698 2692 19702 2748
rect 19638 2688 19702 2692
rect 19718 2748 19782 2752
rect 19718 2692 19722 2748
rect 19722 2692 19778 2748
rect 19778 2692 19782 2748
rect 19718 2688 19782 2692
rect 19798 2748 19862 2752
rect 19798 2692 19802 2748
rect 19802 2692 19858 2748
rect 19858 2692 19862 2748
rect 19798 2688 19862 2692
rect 50278 2748 50342 2752
rect 50278 2692 50282 2748
rect 50282 2692 50338 2748
rect 50338 2692 50342 2748
rect 50278 2688 50342 2692
rect 50358 2748 50422 2752
rect 50358 2692 50362 2748
rect 50362 2692 50418 2748
rect 50418 2692 50422 2748
rect 50358 2688 50422 2692
rect 50438 2748 50502 2752
rect 50438 2692 50442 2748
rect 50442 2692 50498 2748
rect 50498 2692 50502 2748
rect 50438 2688 50502 2692
rect 50518 2748 50582 2752
rect 50518 2692 50522 2748
rect 50522 2692 50578 2748
rect 50578 2692 50582 2748
rect 50518 2688 50582 2692
rect 4198 2204 4262 2208
rect 4198 2148 4202 2204
rect 4202 2148 4258 2204
rect 4258 2148 4262 2204
rect 4198 2144 4262 2148
rect 4278 2204 4342 2208
rect 4278 2148 4282 2204
rect 4282 2148 4338 2204
rect 4338 2148 4342 2204
rect 4278 2144 4342 2148
rect 4358 2204 4422 2208
rect 4358 2148 4362 2204
rect 4362 2148 4418 2204
rect 4418 2148 4422 2204
rect 4358 2144 4422 2148
rect 4438 2204 4502 2208
rect 4438 2148 4442 2204
rect 4442 2148 4498 2204
rect 4498 2148 4502 2204
rect 4438 2144 4502 2148
rect 34918 2204 34982 2208
rect 34918 2148 34922 2204
rect 34922 2148 34978 2204
rect 34978 2148 34982 2204
rect 34918 2144 34982 2148
rect 34998 2204 35062 2208
rect 34998 2148 35002 2204
rect 35002 2148 35058 2204
rect 35058 2148 35062 2204
rect 34998 2144 35062 2148
rect 35078 2204 35142 2208
rect 35078 2148 35082 2204
rect 35082 2148 35138 2204
rect 35138 2148 35142 2204
rect 35078 2144 35142 2148
rect 35158 2204 35222 2208
rect 35158 2148 35162 2204
rect 35162 2148 35218 2204
rect 35218 2148 35222 2204
rect 35158 2144 35222 2148
<< metal4 >>
rect 4190 57696 4510 57712
rect 4190 57632 4198 57696
rect 4262 57632 4278 57696
rect 4342 57632 4358 57696
rect 4422 57632 4438 57696
rect 4502 57632 4510 57696
rect 4190 56608 4510 57632
rect 4190 56544 4198 56608
rect 4262 56544 4278 56608
rect 4342 56544 4358 56608
rect 4422 56544 4438 56608
rect 4502 56544 4510 56608
rect 4190 55520 4510 56544
rect 4190 55456 4198 55520
rect 4262 55456 4278 55520
rect 4342 55456 4358 55520
rect 4422 55456 4438 55520
rect 4502 55456 4510 55520
rect 4190 54432 4510 55456
rect 4190 54368 4198 54432
rect 4262 54368 4278 54432
rect 4342 54368 4358 54432
rect 4422 54368 4438 54432
rect 4502 54368 4510 54432
rect 4190 53344 4510 54368
rect 4190 53280 4198 53344
rect 4262 53280 4278 53344
rect 4342 53280 4358 53344
rect 4422 53280 4438 53344
rect 4502 53280 4510 53344
rect 4190 52256 4510 53280
rect 4190 52192 4198 52256
rect 4262 52192 4278 52256
rect 4342 52192 4358 52256
rect 4422 52192 4438 52256
rect 4502 52192 4510 52256
rect 4190 51168 4510 52192
rect 4190 51104 4198 51168
rect 4262 51104 4278 51168
rect 4342 51104 4358 51168
rect 4422 51104 4438 51168
rect 4502 51104 4510 51168
rect 4190 50080 4510 51104
rect 4190 50016 4198 50080
rect 4262 50016 4278 50080
rect 4342 50016 4358 50080
rect 4422 50016 4438 50080
rect 4502 50016 4510 50080
rect 4190 48992 4510 50016
rect 4190 48928 4198 48992
rect 4262 48928 4278 48992
rect 4342 48928 4358 48992
rect 4422 48928 4438 48992
rect 4502 48928 4510 48992
rect 4190 47904 4510 48928
rect 4190 47840 4198 47904
rect 4262 47840 4278 47904
rect 4342 47840 4358 47904
rect 4422 47840 4438 47904
rect 4502 47840 4510 47904
rect 4190 46816 4510 47840
rect 4190 46752 4198 46816
rect 4262 46752 4278 46816
rect 4342 46752 4358 46816
rect 4422 46752 4438 46816
rect 4502 46752 4510 46816
rect 4190 45728 4510 46752
rect 4190 45664 4198 45728
rect 4262 45664 4278 45728
rect 4342 45664 4358 45728
rect 4422 45664 4438 45728
rect 4502 45664 4510 45728
rect 4190 44640 4510 45664
rect 4190 44576 4198 44640
rect 4262 44576 4278 44640
rect 4342 44576 4358 44640
rect 4422 44576 4438 44640
rect 4502 44576 4510 44640
rect 4190 43552 4510 44576
rect 4190 43488 4198 43552
rect 4262 43488 4278 43552
rect 4342 43488 4358 43552
rect 4422 43488 4438 43552
rect 4502 43488 4510 43552
rect 4190 42464 4510 43488
rect 4190 42400 4198 42464
rect 4262 42400 4278 42464
rect 4342 42400 4358 42464
rect 4422 42400 4438 42464
rect 4502 42400 4510 42464
rect 4190 41376 4510 42400
rect 4190 41312 4198 41376
rect 4262 41312 4278 41376
rect 4342 41312 4358 41376
rect 4422 41312 4438 41376
rect 4502 41312 4510 41376
rect 4190 40288 4510 41312
rect 4190 40224 4198 40288
rect 4262 40224 4278 40288
rect 4342 40224 4358 40288
rect 4422 40224 4438 40288
rect 4502 40224 4510 40288
rect 4190 39200 4510 40224
rect 4190 39136 4198 39200
rect 4262 39136 4278 39200
rect 4342 39136 4358 39200
rect 4422 39136 4438 39200
rect 4502 39136 4510 39200
rect 4190 38112 4510 39136
rect 4190 38048 4198 38112
rect 4262 38048 4278 38112
rect 4342 38048 4358 38112
rect 4422 38048 4438 38112
rect 4502 38048 4510 38112
rect 4190 37024 4510 38048
rect 4190 36960 4198 37024
rect 4262 36960 4278 37024
rect 4342 36960 4358 37024
rect 4422 36960 4438 37024
rect 4502 36960 4510 37024
rect 4190 35936 4510 36960
rect 4190 35872 4198 35936
rect 4262 35872 4278 35936
rect 4342 35872 4358 35936
rect 4422 35872 4438 35936
rect 4502 35872 4510 35936
rect 4190 34848 4510 35872
rect 4190 34784 4198 34848
rect 4262 34784 4278 34848
rect 4342 34784 4358 34848
rect 4422 34784 4438 34848
rect 4502 34784 4510 34848
rect 4190 33760 4510 34784
rect 4190 33696 4198 33760
rect 4262 33696 4278 33760
rect 4342 33696 4358 33760
rect 4422 33696 4438 33760
rect 4502 33696 4510 33760
rect 4190 32672 4510 33696
rect 4190 32608 4198 32672
rect 4262 32608 4278 32672
rect 4342 32608 4358 32672
rect 4422 32608 4438 32672
rect 4502 32608 4510 32672
rect 4190 31584 4510 32608
rect 4190 31520 4198 31584
rect 4262 31520 4278 31584
rect 4342 31520 4358 31584
rect 4422 31520 4438 31584
rect 4502 31520 4510 31584
rect 4190 30496 4510 31520
rect 4190 30432 4198 30496
rect 4262 30432 4278 30496
rect 4342 30432 4358 30496
rect 4422 30432 4438 30496
rect 4502 30432 4510 30496
rect 4190 29408 4510 30432
rect 4190 29344 4198 29408
rect 4262 29344 4278 29408
rect 4342 29344 4358 29408
rect 4422 29344 4438 29408
rect 4502 29344 4510 29408
rect 4190 28320 4510 29344
rect 4190 28256 4198 28320
rect 4262 28256 4278 28320
rect 4342 28256 4358 28320
rect 4422 28256 4438 28320
rect 4502 28256 4510 28320
rect 4190 27232 4510 28256
rect 4190 27168 4198 27232
rect 4262 27168 4278 27232
rect 4342 27168 4358 27232
rect 4422 27168 4438 27232
rect 4502 27168 4510 27232
rect 4190 26144 4510 27168
rect 4190 26080 4198 26144
rect 4262 26080 4278 26144
rect 4342 26080 4358 26144
rect 4422 26080 4438 26144
rect 4502 26080 4510 26144
rect 4190 25056 4510 26080
rect 4190 24992 4198 25056
rect 4262 24992 4278 25056
rect 4342 24992 4358 25056
rect 4422 24992 4438 25056
rect 4502 24992 4510 25056
rect 4190 23968 4510 24992
rect 4190 23904 4198 23968
rect 4262 23904 4278 23968
rect 4342 23904 4358 23968
rect 4422 23904 4438 23968
rect 4502 23904 4510 23968
rect 4190 22880 4510 23904
rect 4190 22816 4198 22880
rect 4262 22816 4278 22880
rect 4342 22816 4358 22880
rect 4422 22816 4438 22880
rect 4502 22816 4510 22880
rect 4190 21792 4510 22816
rect 4190 21728 4198 21792
rect 4262 21728 4278 21792
rect 4342 21728 4358 21792
rect 4422 21728 4438 21792
rect 4502 21728 4510 21792
rect 4190 20704 4510 21728
rect 4190 20640 4198 20704
rect 4262 20640 4278 20704
rect 4342 20640 4358 20704
rect 4422 20640 4438 20704
rect 4502 20640 4510 20704
rect 4190 19616 4510 20640
rect 4190 19552 4198 19616
rect 4262 19552 4278 19616
rect 4342 19552 4358 19616
rect 4422 19552 4438 19616
rect 4502 19552 4510 19616
rect 4190 18528 4510 19552
rect 4190 18464 4198 18528
rect 4262 18464 4278 18528
rect 4342 18464 4358 18528
rect 4422 18464 4438 18528
rect 4502 18464 4510 18528
rect 4190 17440 4510 18464
rect 4190 17376 4198 17440
rect 4262 17376 4278 17440
rect 4342 17376 4358 17440
rect 4422 17376 4438 17440
rect 4502 17376 4510 17440
rect 4190 16352 4510 17376
rect 4190 16288 4198 16352
rect 4262 16288 4278 16352
rect 4342 16288 4358 16352
rect 4422 16288 4438 16352
rect 4502 16288 4510 16352
rect 4190 15264 4510 16288
rect 4190 15200 4198 15264
rect 4262 15200 4278 15264
rect 4342 15200 4358 15264
rect 4422 15200 4438 15264
rect 4502 15200 4510 15264
rect 4190 14176 4510 15200
rect 4190 14112 4198 14176
rect 4262 14112 4278 14176
rect 4342 14112 4358 14176
rect 4422 14112 4438 14176
rect 4502 14112 4510 14176
rect 4190 13088 4510 14112
rect 4190 13024 4198 13088
rect 4262 13024 4278 13088
rect 4342 13024 4358 13088
rect 4422 13024 4438 13088
rect 4502 13024 4510 13088
rect 4190 12000 4510 13024
rect 4190 11936 4198 12000
rect 4262 11936 4278 12000
rect 4342 11936 4358 12000
rect 4422 11936 4438 12000
rect 4502 11936 4510 12000
rect 4190 10912 4510 11936
rect 4190 10848 4198 10912
rect 4262 10848 4278 10912
rect 4342 10848 4358 10912
rect 4422 10848 4438 10912
rect 4502 10848 4510 10912
rect 4190 9824 4510 10848
rect 4190 9760 4198 9824
rect 4262 9760 4278 9824
rect 4342 9760 4358 9824
rect 4422 9760 4438 9824
rect 4502 9760 4510 9824
rect 4190 8736 4510 9760
rect 4190 8672 4198 8736
rect 4262 8672 4278 8736
rect 4342 8672 4358 8736
rect 4422 8672 4438 8736
rect 4502 8672 4510 8736
rect 4190 7648 4510 8672
rect 4190 7584 4198 7648
rect 4262 7584 4278 7648
rect 4342 7584 4358 7648
rect 4422 7584 4438 7648
rect 4502 7584 4510 7648
rect 4190 6560 4510 7584
rect 4190 6496 4198 6560
rect 4262 6496 4278 6560
rect 4342 6496 4358 6560
rect 4422 6496 4438 6560
rect 4502 6496 4510 6560
rect 4190 5472 4510 6496
rect 4190 5408 4198 5472
rect 4262 5408 4278 5472
rect 4342 5408 4358 5472
rect 4422 5408 4438 5472
rect 4502 5408 4510 5472
rect 4190 4384 4510 5408
rect 4190 4320 4198 4384
rect 4262 4320 4278 4384
rect 4342 4320 4358 4384
rect 4422 4320 4438 4384
rect 4502 4320 4510 4384
rect 4190 3296 4510 4320
rect 4190 3232 4198 3296
rect 4262 3232 4278 3296
rect 4342 3232 4358 3296
rect 4422 3232 4438 3296
rect 4502 3232 4510 3296
rect 4190 2208 4510 3232
rect 4190 2144 4198 2208
rect 4262 2144 4278 2208
rect 4342 2144 4358 2208
rect 4422 2144 4438 2208
rect 4502 2144 4510 2208
rect 4190 2128 4510 2144
rect 19550 57152 19870 57712
rect 19550 57088 19558 57152
rect 19622 57088 19638 57152
rect 19702 57088 19718 57152
rect 19782 57088 19798 57152
rect 19862 57088 19870 57152
rect 19550 56064 19870 57088
rect 19550 56000 19558 56064
rect 19622 56000 19638 56064
rect 19702 56000 19718 56064
rect 19782 56000 19798 56064
rect 19862 56000 19870 56064
rect 19550 54976 19870 56000
rect 19550 54912 19558 54976
rect 19622 54912 19638 54976
rect 19702 54912 19718 54976
rect 19782 54912 19798 54976
rect 19862 54912 19870 54976
rect 19550 53888 19870 54912
rect 19550 53824 19558 53888
rect 19622 53824 19638 53888
rect 19702 53824 19718 53888
rect 19782 53824 19798 53888
rect 19862 53824 19870 53888
rect 19550 52800 19870 53824
rect 19550 52736 19558 52800
rect 19622 52736 19638 52800
rect 19702 52736 19718 52800
rect 19782 52736 19798 52800
rect 19862 52736 19870 52800
rect 19550 51712 19870 52736
rect 19550 51648 19558 51712
rect 19622 51648 19638 51712
rect 19702 51648 19718 51712
rect 19782 51648 19798 51712
rect 19862 51648 19870 51712
rect 19550 50624 19870 51648
rect 19550 50560 19558 50624
rect 19622 50560 19638 50624
rect 19702 50560 19718 50624
rect 19782 50560 19798 50624
rect 19862 50560 19870 50624
rect 19550 49536 19870 50560
rect 19550 49472 19558 49536
rect 19622 49472 19638 49536
rect 19702 49472 19718 49536
rect 19782 49472 19798 49536
rect 19862 49472 19870 49536
rect 19550 48448 19870 49472
rect 19550 48384 19558 48448
rect 19622 48384 19638 48448
rect 19702 48384 19718 48448
rect 19782 48384 19798 48448
rect 19862 48384 19870 48448
rect 19550 47360 19870 48384
rect 19550 47296 19558 47360
rect 19622 47296 19638 47360
rect 19702 47296 19718 47360
rect 19782 47296 19798 47360
rect 19862 47296 19870 47360
rect 19550 46272 19870 47296
rect 19550 46208 19558 46272
rect 19622 46208 19638 46272
rect 19702 46208 19718 46272
rect 19782 46208 19798 46272
rect 19862 46208 19870 46272
rect 19550 45184 19870 46208
rect 19550 45120 19558 45184
rect 19622 45120 19638 45184
rect 19702 45120 19718 45184
rect 19782 45120 19798 45184
rect 19862 45120 19870 45184
rect 19550 44096 19870 45120
rect 19550 44032 19558 44096
rect 19622 44032 19638 44096
rect 19702 44032 19718 44096
rect 19782 44032 19798 44096
rect 19862 44032 19870 44096
rect 19550 43008 19870 44032
rect 19550 42944 19558 43008
rect 19622 42944 19638 43008
rect 19702 42944 19718 43008
rect 19782 42944 19798 43008
rect 19862 42944 19870 43008
rect 19550 41920 19870 42944
rect 19550 41856 19558 41920
rect 19622 41856 19638 41920
rect 19702 41856 19718 41920
rect 19782 41856 19798 41920
rect 19862 41856 19870 41920
rect 19550 40832 19870 41856
rect 19550 40768 19558 40832
rect 19622 40768 19638 40832
rect 19702 40768 19718 40832
rect 19782 40768 19798 40832
rect 19862 40768 19870 40832
rect 19550 39744 19870 40768
rect 19550 39680 19558 39744
rect 19622 39680 19638 39744
rect 19702 39680 19718 39744
rect 19782 39680 19798 39744
rect 19862 39680 19870 39744
rect 19550 38656 19870 39680
rect 19550 38592 19558 38656
rect 19622 38592 19638 38656
rect 19702 38592 19718 38656
rect 19782 38592 19798 38656
rect 19862 38592 19870 38656
rect 19550 37568 19870 38592
rect 19550 37504 19558 37568
rect 19622 37504 19638 37568
rect 19702 37504 19718 37568
rect 19782 37504 19798 37568
rect 19862 37504 19870 37568
rect 19550 36480 19870 37504
rect 19550 36416 19558 36480
rect 19622 36416 19638 36480
rect 19702 36416 19718 36480
rect 19782 36416 19798 36480
rect 19862 36416 19870 36480
rect 19550 35392 19870 36416
rect 19550 35328 19558 35392
rect 19622 35328 19638 35392
rect 19702 35328 19718 35392
rect 19782 35328 19798 35392
rect 19862 35328 19870 35392
rect 19550 34304 19870 35328
rect 19550 34240 19558 34304
rect 19622 34240 19638 34304
rect 19702 34240 19718 34304
rect 19782 34240 19798 34304
rect 19862 34240 19870 34304
rect 19550 33216 19870 34240
rect 19550 33152 19558 33216
rect 19622 33152 19638 33216
rect 19702 33152 19718 33216
rect 19782 33152 19798 33216
rect 19862 33152 19870 33216
rect 19550 32128 19870 33152
rect 19550 32064 19558 32128
rect 19622 32064 19638 32128
rect 19702 32064 19718 32128
rect 19782 32064 19798 32128
rect 19862 32064 19870 32128
rect 19550 31040 19870 32064
rect 19550 30976 19558 31040
rect 19622 30976 19638 31040
rect 19702 30976 19718 31040
rect 19782 30976 19798 31040
rect 19862 30976 19870 31040
rect 19550 29952 19870 30976
rect 19550 29888 19558 29952
rect 19622 29888 19638 29952
rect 19702 29888 19718 29952
rect 19782 29888 19798 29952
rect 19862 29888 19870 29952
rect 19550 28864 19870 29888
rect 19550 28800 19558 28864
rect 19622 28800 19638 28864
rect 19702 28800 19718 28864
rect 19782 28800 19798 28864
rect 19862 28800 19870 28864
rect 19550 27776 19870 28800
rect 19550 27712 19558 27776
rect 19622 27712 19638 27776
rect 19702 27712 19718 27776
rect 19782 27712 19798 27776
rect 19862 27712 19870 27776
rect 19550 26688 19870 27712
rect 19550 26624 19558 26688
rect 19622 26624 19638 26688
rect 19702 26624 19718 26688
rect 19782 26624 19798 26688
rect 19862 26624 19870 26688
rect 19550 25600 19870 26624
rect 19550 25536 19558 25600
rect 19622 25536 19638 25600
rect 19702 25536 19718 25600
rect 19782 25536 19798 25600
rect 19862 25536 19870 25600
rect 19550 24512 19870 25536
rect 19550 24448 19558 24512
rect 19622 24448 19638 24512
rect 19702 24448 19718 24512
rect 19782 24448 19798 24512
rect 19862 24448 19870 24512
rect 19550 23424 19870 24448
rect 19550 23360 19558 23424
rect 19622 23360 19638 23424
rect 19702 23360 19718 23424
rect 19782 23360 19798 23424
rect 19862 23360 19870 23424
rect 19550 22336 19870 23360
rect 19550 22272 19558 22336
rect 19622 22272 19638 22336
rect 19702 22272 19718 22336
rect 19782 22272 19798 22336
rect 19862 22272 19870 22336
rect 19550 21248 19870 22272
rect 19550 21184 19558 21248
rect 19622 21184 19638 21248
rect 19702 21184 19718 21248
rect 19782 21184 19798 21248
rect 19862 21184 19870 21248
rect 19550 20160 19870 21184
rect 19550 20096 19558 20160
rect 19622 20096 19638 20160
rect 19702 20096 19718 20160
rect 19782 20096 19798 20160
rect 19862 20096 19870 20160
rect 19550 19072 19870 20096
rect 19550 19008 19558 19072
rect 19622 19008 19638 19072
rect 19702 19008 19718 19072
rect 19782 19008 19798 19072
rect 19862 19008 19870 19072
rect 19550 17984 19870 19008
rect 19550 17920 19558 17984
rect 19622 17920 19638 17984
rect 19702 17920 19718 17984
rect 19782 17920 19798 17984
rect 19862 17920 19870 17984
rect 19550 16896 19870 17920
rect 19550 16832 19558 16896
rect 19622 16832 19638 16896
rect 19702 16832 19718 16896
rect 19782 16832 19798 16896
rect 19862 16832 19870 16896
rect 19550 15808 19870 16832
rect 19550 15744 19558 15808
rect 19622 15744 19638 15808
rect 19702 15744 19718 15808
rect 19782 15744 19798 15808
rect 19862 15744 19870 15808
rect 19550 14720 19870 15744
rect 19550 14656 19558 14720
rect 19622 14656 19638 14720
rect 19702 14656 19718 14720
rect 19782 14656 19798 14720
rect 19862 14656 19870 14720
rect 19550 13632 19870 14656
rect 19550 13568 19558 13632
rect 19622 13568 19638 13632
rect 19702 13568 19718 13632
rect 19782 13568 19798 13632
rect 19862 13568 19870 13632
rect 19550 12544 19870 13568
rect 19550 12480 19558 12544
rect 19622 12480 19638 12544
rect 19702 12480 19718 12544
rect 19782 12480 19798 12544
rect 19862 12480 19870 12544
rect 19550 11456 19870 12480
rect 19550 11392 19558 11456
rect 19622 11392 19638 11456
rect 19702 11392 19718 11456
rect 19782 11392 19798 11456
rect 19862 11392 19870 11456
rect 19550 10368 19870 11392
rect 19550 10304 19558 10368
rect 19622 10304 19638 10368
rect 19702 10304 19718 10368
rect 19782 10304 19798 10368
rect 19862 10304 19870 10368
rect 19550 9280 19870 10304
rect 19550 9216 19558 9280
rect 19622 9216 19638 9280
rect 19702 9216 19718 9280
rect 19782 9216 19798 9280
rect 19862 9216 19870 9280
rect 19550 8192 19870 9216
rect 19550 8128 19558 8192
rect 19622 8128 19638 8192
rect 19702 8128 19718 8192
rect 19782 8128 19798 8192
rect 19862 8128 19870 8192
rect 19550 7104 19870 8128
rect 19550 7040 19558 7104
rect 19622 7040 19638 7104
rect 19702 7040 19718 7104
rect 19782 7040 19798 7104
rect 19862 7040 19870 7104
rect 19550 6016 19870 7040
rect 19550 5952 19558 6016
rect 19622 5952 19638 6016
rect 19702 5952 19718 6016
rect 19782 5952 19798 6016
rect 19862 5952 19870 6016
rect 19550 4928 19870 5952
rect 19550 4864 19558 4928
rect 19622 4864 19638 4928
rect 19702 4864 19718 4928
rect 19782 4864 19798 4928
rect 19862 4864 19870 4928
rect 19550 3840 19870 4864
rect 19550 3776 19558 3840
rect 19622 3776 19638 3840
rect 19702 3776 19718 3840
rect 19782 3776 19798 3840
rect 19862 3776 19870 3840
rect 19550 2752 19870 3776
rect 19550 2688 19558 2752
rect 19622 2688 19638 2752
rect 19702 2688 19718 2752
rect 19782 2688 19798 2752
rect 19862 2688 19870 2752
rect 19550 2128 19870 2688
rect 34910 57696 35230 57712
rect 34910 57632 34918 57696
rect 34982 57632 34998 57696
rect 35062 57632 35078 57696
rect 35142 57632 35158 57696
rect 35222 57632 35230 57696
rect 34910 56608 35230 57632
rect 34910 56544 34918 56608
rect 34982 56544 34998 56608
rect 35062 56544 35078 56608
rect 35142 56544 35158 56608
rect 35222 56544 35230 56608
rect 34910 55520 35230 56544
rect 34910 55456 34918 55520
rect 34982 55456 34998 55520
rect 35062 55456 35078 55520
rect 35142 55456 35158 55520
rect 35222 55456 35230 55520
rect 34910 54432 35230 55456
rect 34910 54368 34918 54432
rect 34982 54368 34998 54432
rect 35062 54368 35078 54432
rect 35142 54368 35158 54432
rect 35222 54368 35230 54432
rect 34910 53344 35230 54368
rect 34910 53280 34918 53344
rect 34982 53280 34998 53344
rect 35062 53280 35078 53344
rect 35142 53280 35158 53344
rect 35222 53280 35230 53344
rect 34910 52256 35230 53280
rect 34910 52192 34918 52256
rect 34982 52192 34998 52256
rect 35062 52192 35078 52256
rect 35142 52192 35158 52256
rect 35222 52192 35230 52256
rect 34910 51168 35230 52192
rect 34910 51104 34918 51168
rect 34982 51104 34998 51168
rect 35062 51104 35078 51168
rect 35142 51104 35158 51168
rect 35222 51104 35230 51168
rect 34910 50080 35230 51104
rect 34910 50016 34918 50080
rect 34982 50016 34998 50080
rect 35062 50016 35078 50080
rect 35142 50016 35158 50080
rect 35222 50016 35230 50080
rect 34910 48992 35230 50016
rect 34910 48928 34918 48992
rect 34982 48928 34998 48992
rect 35062 48928 35078 48992
rect 35142 48928 35158 48992
rect 35222 48928 35230 48992
rect 34910 47904 35230 48928
rect 34910 47840 34918 47904
rect 34982 47840 34998 47904
rect 35062 47840 35078 47904
rect 35142 47840 35158 47904
rect 35222 47840 35230 47904
rect 34910 46816 35230 47840
rect 34910 46752 34918 46816
rect 34982 46752 34998 46816
rect 35062 46752 35078 46816
rect 35142 46752 35158 46816
rect 35222 46752 35230 46816
rect 34910 45728 35230 46752
rect 34910 45664 34918 45728
rect 34982 45664 34998 45728
rect 35062 45664 35078 45728
rect 35142 45664 35158 45728
rect 35222 45664 35230 45728
rect 34910 44640 35230 45664
rect 34910 44576 34918 44640
rect 34982 44576 34998 44640
rect 35062 44576 35078 44640
rect 35142 44576 35158 44640
rect 35222 44576 35230 44640
rect 34910 43552 35230 44576
rect 34910 43488 34918 43552
rect 34982 43488 34998 43552
rect 35062 43488 35078 43552
rect 35142 43488 35158 43552
rect 35222 43488 35230 43552
rect 34910 42464 35230 43488
rect 34910 42400 34918 42464
rect 34982 42400 34998 42464
rect 35062 42400 35078 42464
rect 35142 42400 35158 42464
rect 35222 42400 35230 42464
rect 34910 41376 35230 42400
rect 34910 41312 34918 41376
rect 34982 41312 34998 41376
rect 35062 41312 35078 41376
rect 35142 41312 35158 41376
rect 35222 41312 35230 41376
rect 34910 40288 35230 41312
rect 34910 40224 34918 40288
rect 34982 40224 34998 40288
rect 35062 40224 35078 40288
rect 35142 40224 35158 40288
rect 35222 40224 35230 40288
rect 34910 39200 35230 40224
rect 34910 39136 34918 39200
rect 34982 39136 34998 39200
rect 35062 39136 35078 39200
rect 35142 39136 35158 39200
rect 35222 39136 35230 39200
rect 34910 38112 35230 39136
rect 34910 38048 34918 38112
rect 34982 38048 34998 38112
rect 35062 38048 35078 38112
rect 35142 38048 35158 38112
rect 35222 38048 35230 38112
rect 34910 37024 35230 38048
rect 34910 36960 34918 37024
rect 34982 36960 34998 37024
rect 35062 36960 35078 37024
rect 35142 36960 35158 37024
rect 35222 36960 35230 37024
rect 34910 35936 35230 36960
rect 34910 35872 34918 35936
rect 34982 35872 34998 35936
rect 35062 35872 35078 35936
rect 35142 35872 35158 35936
rect 35222 35872 35230 35936
rect 34910 34848 35230 35872
rect 34910 34784 34918 34848
rect 34982 34784 34998 34848
rect 35062 34784 35078 34848
rect 35142 34784 35158 34848
rect 35222 34784 35230 34848
rect 34910 33760 35230 34784
rect 34910 33696 34918 33760
rect 34982 33696 34998 33760
rect 35062 33696 35078 33760
rect 35142 33696 35158 33760
rect 35222 33696 35230 33760
rect 34910 32672 35230 33696
rect 34910 32608 34918 32672
rect 34982 32608 34998 32672
rect 35062 32608 35078 32672
rect 35142 32608 35158 32672
rect 35222 32608 35230 32672
rect 34910 31584 35230 32608
rect 34910 31520 34918 31584
rect 34982 31520 34998 31584
rect 35062 31520 35078 31584
rect 35142 31520 35158 31584
rect 35222 31520 35230 31584
rect 34910 30496 35230 31520
rect 34910 30432 34918 30496
rect 34982 30432 34998 30496
rect 35062 30432 35078 30496
rect 35142 30432 35158 30496
rect 35222 30432 35230 30496
rect 34910 29408 35230 30432
rect 34910 29344 34918 29408
rect 34982 29344 34998 29408
rect 35062 29344 35078 29408
rect 35142 29344 35158 29408
rect 35222 29344 35230 29408
rect 34910 28320 35230 29344
rect 34910 28256 34918 28320
rect 34982 28256 34998 28320
rect 35062 28256 35078 28320
rect 35142 28256 35158 28320
rect 35222 28256 35230 28320
rect 34910 27232 35230 28256
rect 34910 27168 34918 27232
rect 34982 27168 34998 27232
rect 35062 27168 35078 27232
rect 35142 27168 35158 27232
rect 35222 27168 35230 27232
rect 34910 26144 35230 27168
rect 34910 26080 34918 26144
rect 34982 26080 34998 26144
rect 35062 26080 35078 26144
rect 35142 26080 35158 26144
rect 35222 26080 35230 26144
rect 34910 25056 35230 26080
rect 34910 24992 34918 25056
rect 34982 24992 34998 25056
rect 35062 24992 35078 25056
rect 35142 24992 35158 25056
rect 35222 24992 35230 25056
rect 34910 23968 35230 24992
rect 34910 23904 34918 23968
rect 34982 23904 34998 23968
rect 35062 23904 35078 23968
rect 35142 23904 35158 23968
rect 35222 23904 35230 23968
rect 34910 22880 35230 23904
rect 34910 22816 34918 22880
rect 34982 22816 34998 22880
rect 35062 22816 35078 22880
rect 35142 22816 35158 22880
rect 35222 22816 35230 22880
rect 34910 21792 35230 22816
rect 34910 21728 34918 21792
rect 34982 21728 34998 21792
rect 35062 21728 35078 21792
rect 35142 21728 35158 21792
rect 35222 21728 35230 21792
rect 34910 20704 35230 21728
rect 34910 20640 34918 20704
rect 34982 20640 34998 20704
rect 35062 20640 35078 20704
rect 35142 20640 35158 20704
rect 35222 20640 35230 20704
rect 34910 19616 35230 20640
rect 34910 19552 34918 19616
rect 34982 19552 34998 19616
rect 35062 19552 35078 19616
rect 35142 19552 35158 19616
rect 35222 19552 35230 19616
rect 34910 18528 35230 19552
rect 34910 18464 34918 18528
rect 34982 18464 34998 18528
rect 35062 18464 35078 18528
rect 35142 18464 35158 18528
rect 35222 18464 35230 18528
rect 34910 17440 35230 18464
rect 34910 17376 34918 17440
rect 34982 17376 34998 17440
rect 35062 17376 35078 17440
rect 35142 17376 35158 17440
rect 35222 17376 35230 17440
rect 34910 16352 35230 17376
rect 34910 16288 34918 16352
rect 34982 16288 34998 16352
rect 35062 16288 35078 16352
rect 35142 16288 35158 16352
rect 35222 16288 35230 16352
rect 34910 15264 35230 16288
rect 34910 15200 34918 15264
rect 34982 15200 34998 15264
rect 35062 15200 35078 15264
rect 35142 15200 35158 15264
rect 35222 15200 35230 15264
rect 34910 14176 35230 15200
rect 34910 14112 34918 14176
rect 34982 14112 34998 14176
rect 35062 14112 35078 14176
rect 35142 14112 35158 14176
rect 35222 14112 35230 14176
rect 34910 13088 35230 14112
rect 34910 13024 34918 13088
rect 34982 13024 34998 13088
rect 35062 13024 35078 13088
rect 35142 13024 35158 13088
rect 35222 13024 35230 13088
rect 34910 12000 35230 13024
rect 34910 11936 34918 12000
rect 34982 11936 34998 12000
rect 35062 11936 35078 12000
rect 35142 11936 35158 12000
rect 35222 11936 35230 12000
rect 34910 10912 35230 11936
rect 34910 10848 34918 10912
rect 34982 10848 34998 10912
rect 35062 10848 35078 10912
rect 35142 10848 35158 10912
rect 35222 10848 35230 10912
rect 34910 9824 35230 10848
rect 34910 9760 34918 9824
rect 34982 9760 34998 9824
rect 35062 9760 35078 9824
rect 35142 9760 35158 9824
rect 35222 9760 35230 9824
rect 34910 8736 35230 9760
rect 34910 8672 34918 8736
rect 34982 8672 34998 8736
rect 35062 8672 35078 8736
rect 35142 8672 35158 8736
rect 35222 8672 35230 8736
rect 34910 7648 35230 8672
rect 34910 7584 34918 7648
rect 34982 7584 34998 7648
rect 35062 7584 35078 7648
rect 35142 7584 35158 7648
rect 35222 7584 35230 7648
rect 34910 6560 35230 7584
rect 34910 6496 34918 6560
rect 34982 6496 34998 6560
rect 35062 6496 35078 6560
rect 35142 6496 35158 6560
rect 35222 6496 35230 6560
rect 34910 5472 35230 6496
rect 34910 5408 34918 5472
rect 34982 5408 34998 5472
rect 35062 5408 35078 5472
rect 35142 5408 35158 5472
rect 35222 5408 35230 5472
rect 34910 4384 35230 5408
rect 34910 4320 34918 4384
rect 34982 4320 34998 4384
rect 35062 4320 35078 4384
rect 35142 4320 35158 4384
rect 35222 4320 35230 4384
rect 34910 3296 35230 4320
rect 34910 3232 34918 3296
rect 34982 3232 34998 3296
rect 35062 3232 35078 3296
rect 35142 3232 35158 3296
rect 35222 3232 35230 3296
rect 34910 2208 35230 3232
rect 34910 2144 34918 2208
rect 34982 2144 34998 2208
rect 35062 2144 35078 2208
rect 35142 2144 35158 2208
rect 35222 2144 35230 2208
rect 34910 2128 35230 2144
rect 50270 57152 50590 57712
rect 50270 57088 50278 57152
rect 50342 57088 50358 57152
rect 50422 57088 50438 57152
rect 50502 57088 50518 57152
rect 50582 57088 50590 57152
rect 50270 56064 50590 57088
rect 50270 56000 50278 56064
rect 50342 56000 50358 56064
rect 50422 56000 50438 56064
rect 50502 56000 50518 56064
rect 50582 56000 50590 56064
rect 50270 54976 50590 56000
rect 50270 54912 50278 54976
rect 50342 54912 50358 54976
rect 50422 54912 50438 54976
rect 50502 54912 50518 54976
rect 50582 54912 50590 54976
rect 50270 53888 50590 54912
rect 50270 53824 50278 53888
rect 50342 53824 50358 53888
rect 50422 53824 50438 53888
rect 50502 53824 50518 53888
rect 50582 53824 50590 53888
rect 50270 52800 50590 53824
rect 50270 52736 50278 52800
rect 50342 52736 50358 52800
rect 50422 52736 50438 52800
rect 50502 52736 50518 52800
rect 50582 52736 50590 52800
rect 50270 51712 50590 52736
rect 50270 51648 50278 51712
rect 50342 51648 50358 51712
rect 50422 51648 50438 51712
rect 50502 51648 50518 51712
rect 50582 51648 50590 51712
rect 50270 50624 50590 51648
rect 50270 50560 50278 50624
rect 50342 50560 50358 50624
rect 50422 50560 50438 50624
rect 50502 50560 50518 50624
rect 50582 50560 50590 50624
rect 50270 49536 50590 50560
rect 50270 49472 50278 49536
rect 50342 49472 50358 49536
rect 50422 49472 50438 49536
rect 50502 49472 50518 49536
rect 50582 49472 50590 49536
rect 50270 48448 50590 49472
rect 50270 48384 50278 48448
rect 50342 48384 50358 48448
rect 50422 48384 50438 48448
rect 50502 48384 50518 48448
rect 50582 48384 50590 48448
rect 50270 47360 50590 48384
rect 50270 47296 50278 47360
rect 50342 47296 50358 47360
rect 50422 47296 50438 47360
rect 50502 47296 50518 47360
rect 50582 47296 50590 47360
rect 50270 46272 50590 47296
rect 50270 46208 50278 46272
rect 50342 46208 50358 46272
rect 50422 46208 50438 46272
rect 50502 46208 50518 46272
rect 50582 46208 50590 46272
rect 50270 45184 50590 46208
rect 50270 45120 50278 45184
rect 50342 45120 50358 45184
rect 50422 45120 50438 45184
rect 50502 45120 50518 45184
rect 50582 45120 50590 45184
rect 50270 44096 50590 45120
rect 50270 44032 50278 44096
rect 50342 44032 50358 44096
rect 50422 44032 50438 44096
rect 50502 44032 50518 44096
rect 50582 44032 50590 44096
rect 50270 43008 50590 44032
rect 50270 42944 50278 43008
rect 50342 42944 50358 43008
rect 50422 42944 50438 43008
rect 50502 42944 50518 43008
rect 50582 42944 50590 43008
rect 50270 41920 50590 42944
rect 50270 41856 50278 41920
rect 50342 41856 50358 41920
rect 50422 41856 50438 41920
rect 50502 41856 50518 41920
rect 50582 41856 50590 41920
rect 50270 40832 50590 41856
rect 50270 40768 50278 40832
rect 50342 40768 50358 40832
rect 50422 40768 50438 40832
rect 50502 40768 50518 40832
rect 50582 40768 50590 40832
rect 50270 39744 50590 40768
rect 50270 39680 50278 39744
rect 50342 39680 50358 39744
rect 50422 39680 50438 39744
rect 50502 39680 50518 39744
rect 50582 39680 50590 39744
rect 50270 38656 50590 39680
rect 50270 38592 50278 38656
rect 50342 38592 50358 38656
rect 50422 38592 50438 38656
rect 50502 38592 50518 38656
rect 50582 38592 50590 38656
rect 50270 37568 50590 38592
rect 50270 37504 50278 37568
rect 50342 37504 50358 37568
rect 50422 37504 50438 37568
rect 50502 37504 50518 37568
rect 50582 37504 50590 37568
rect 50270 36480 50590 37504
rect 50270 36416 50278 36480
rect 50342 36416 50358 36480
rect 50422 36416 50438 36480
rect 50502 36416 50518 36480
rect 50582 36416 50590 36480
rect 50270 35392 50590 36416
rect 50270 35328 50278 35392
rect 50342 35328 50358 35392
rect 50422 35328 50438 35392
rect 50502 35328 50518 35392
rect 50582 35328 50590 35392
rect 50270 34304 50590 35328
rect 50270 34240 50278 34304
rect 50342 34240 50358 34304
rect 50422 34240 50438 34304
rect 50502 34240 50518 34304
rect 50582 34240 50590 34304
rect 50270 33216 50590 34240
rect 50270 33152 50278 33216
rect 50342 33152 50358 33216
rect 50422 33152 50438 33216
rect 50502 33152 50518 33216
rect 50582 33152 50590 33216
rect 50270 32128 50590 33152
rect 50270 32064 50278 32128
rect 50342 32064 50358 32128
rect 50422 32064 50438 32128
rect 50502 32064 50518 32128
rect 50582 32064 50590 32128
rect 50270 31040 50590 32064
rect 50270 30976 50278 31040
rect 50342 30976 50358 31040
rect 50422 30976 50438 31040
rect 50502 30976 50518 31040
rect 50582 30976 50590 31040
rect 50270 29952 50590 30976
rect 50270 29888 50278 29952
rect 50342 29888 50358 29952
rect 50422 29888 50438 29952
rect 50502 29888 50518 29952
rect 50582 29888 50590 29952
rect 50270 28864 50590 29888
rect 50270 28800 50278 28864
rect 50342 28800 50358 28864
rect 50422 28800 50438 28864
rect 50502 28800 50518 28864
rect 50582 28800 50590 28864
rect 50270 27776 50590 28800
rect 50270 27712 50278 27776
rect 50342 27712 50358 27776
rect 50422 27712 50438 27776
rect 50502 27712 50518 27776
rect 50582 27712 50590 27776
rect 50270 26688 50590 27712
rect 50270 26624 50278 26688
rect 50342 26624 50358 26688
rect 50422 26624 50438 26688
rect 50502 26624 50518 26688
rect 50582 26624 50590 26688
rect 50270 25600 50590 26624
rect 50270 25536 50278 25600
rect 50342 25536 50358 25600
rect 50422 25536 50438 25600
rect 50502 25536 50518 25600
rect 50582 25536 50590 25600
rect 50270 24512 50590 25536
rect 50270 24448 50278 24512
rect 50342 24448 50358 24512
rect 50422 24448 50438 24512
rect 50502 24448 50518 24512
rect 50582 24448 50590 24512
rect 50270 23424 50590 24448
rect 50270 23360 50278 23424
rect 50342 23360 50358 23424
rect 50422 23360 50438 23424
rect 50502 23360 50518 23424
rect 50582 23360 50590 23424
rect 50270 22336 50590 23360
rect 50270 22272 50278 22336
rect 50342 22272 50358 22336
rect 50422 22272 50438 22336
rect 50502 22272 50518 22336
rect 50582 22272 50590 22336
rect 50270 21248 50590 22272
rect 50270 21184 50278 21248
rect 50342 21184 50358 21248
rect 50422 21184 50438 21248
rect 50502 21184 50518 21248
rect 50582 21184 50590 21248
rect 50270 20160 50590 21184
rect 50270 20096 50278 20160
rect 50342 20096 50358 20160
rect 50422 20096 50438 20160
rect 50502 20096 50518 20160
rect 50582 20096 50590 20160
rect 50270 19072 50590 20096
rect 50270 19008 50278 19072
rect 50342 19008 50358 19072
rect 50422 19008 50438 19072
rect 50502 19008 50518 19072
rect 50582 19008 50590 19072
rect 50270 17984 50590 19008
rect 50270 17920 50278 17984
rect 50342 17920 50358 17984
rect 50422 17920 50438 17984
rect 50502 17920 50518 17984
rect 50582 17920 50590 17984
rect 50270 16896 50590 17920
rect 50270 16832 50278 16896
rect 50342 16832 50358 16896
rect 50422 16832 50438 16896
rect 50502 16832 50518 16896
rect 50582 16832 50590 16896
rect 50270 15808 50590 16832
rect 50270 15744 50278 15808
rect 50342 15744 50358 15808
rect 50422 15744 50438 15808
rect 50502 15744 50518 15808
rect 50582 15744 50590 15808
rect 50270 14720 50590 15744
rect 50270 14656 50278 14720
rect 50342 14656 50358 14720
rect 50422 14656 50438 14720
rect 50502 14656 50518 14720
rect 50582 14656 50590 14720
rect 50270 13632 50590 14656
rect 50270 13568 50278 13632
rect 50342 13568 50358 13632
rect 50422 13568 50438 13632
rect 50502 13568 50518 13632
rect 50582 13568 50590 13632
rect 50270 12544 50590 13568
rect 50270 12480 50278 12544
rect 50342 12480 50358 12544
rect 50422 12480 50438 12544
rect 50502 12480 50518 12544
rect 50582 12480 50590 12544
rect 50270 11456 50590 12480
rect 50270 11392 50278 11456
rect 50342 11392 50358 11456
rect 50422 11392 50438 11456
rect 50502 11392 50518 11456
rect 50582 11392 50590 11456
rect 50270 10368 50590 11392
rect 50270 10304 50278 10368
rect 50342 10304 50358 10368
rect 50422 10304 50438 10368
rect 50502 10304 50518 10368
rect 50582 10304 50590 10368
rect 50270 9280 50590 10304
rect 50270 9216 50278 9280
rect 50342 9216 50358 9280
rect 50422 9216 50438 9280
rect 50502 9216 50518 9280
rect 50582 9216 50590 9280
rect 50270 8192 50590 9216
rect 50270 8128 50278 8192
rect 50342 8128 50358 8192
rect 50422 8128 50438 8192
rect 50502 8128 50518 8192
rect 50582 8128 50590 8192
rect 50270 7104 50590 8128
rect 50270 7040 50278 7104
rect 50342 7040 50358 7104
rect 50422 7040 50438 7104
rect 50502 7040 50518 7104
rect 50582 7040 50590 7104
rect 50270 6016 50590 7040
rect 50270 5952 50278 6016
rect 50342 5952 50358 6016
rect 50422 5952 50438 6016
rect 50502 5952 50518 6016
rect 50582 5952 50590 6016
rect 50270 4928 50590 5952
rect 50270 4864 50278 4928
rect 50342 4864 50358 4928
rect 50422 4864 50438 4928
rect 50502 4864 50518 4928
rect 50582 4864 50590 4928
rect 50270 3840 50590 4864
rect 50270 3776 50278 3840
rect 50342 3776 50358 3840
rect 50422 3776 50438 3840
rect 50502 3776 50518 3840
rect 50582 3776 50590 3840
rect 50270 2752 50590 3776
rect 50270 2688 50278 2752
rect 50342 2688 50358 2752
rect 50422 2688 50438 2752
rect 50502 2688 50518 2752
rect 50582 2688 50590 2752
rect 50270 2128 50590 2688
use sky130_fd_sc_hd__decap_12  FILLER_1_15 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607639953
transform 1 0 2466 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_3
timestamp 1607639953
transform 1 0 1362 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1607639953
transform 1 0 2466 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3
timestamp 1607639953
transform 1 0 1362 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_2 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607639953
transform 1 0 1086 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1607639953
transform 1 0 1086 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_39
timestamp 1607639953
transform 1 0 4674 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_27
timestamp 1607639953
transform 1 0 3570 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_44
timestamp 1607639953
transform 1 0 5134 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_32
timestamp 1607639953
transform 1 0 4030 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607639953
transform 1 0 3570 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_204 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607639953
transform 1 0 3938 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_62
timestamp 1607639953
transform 1 0 6790 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_59 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607639953
transform 1 0 6514 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_51 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607639953
transform 1 0 5778 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_0_63
timestamp 1607639953
transform 1 0 6882 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607639953
transform 1 0 6238 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_224
timestamp 1607639953
transform 1 0 6698 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_205
timestamp 1607639953
transform 1 0 6790 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_84
timestamp 1607639953
transform 1 0 8814 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_74
timestamp 1607639953
transform 1 0 7894 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_87
timestamp 1607639953
transform 1 0 9090 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_75
timestamp 1607639953
transform 1 0 7986 0 -1 2720
box -38 -48 1142 592
use AND2X1  AND2X1
timestamp 1608117647
transform 1 0 8078 0 1 2720
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILLER_1_108
timestamp 1607639953
transform 1 0 11022 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_96
timestamp 1607639953
transform 1 0 9918 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_106
timestamp 1607639953
transform 1 0 10838 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_94
timestamp 1607639953
transform 1 0 9734 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_206
timestamp 1607639953
transform 1 0 9642 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_123
timestamp 1607639953
transform 1 0 12402 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_120
timestamp 1607639953
transform 1 0 12126 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1607639953
transform 1 0 12586 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_118
timestamp 1607639953
transform 1 0 11942 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_225
timestamp 1607639953
transform 1 0 12310 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_207
timestamp 1607639953
transform 1 0 12494 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_147
timestamp 1607639953
transform 1 0 14610 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_135
timestamp 1607639953
transform 1 0 13506 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_151
timestamp 1607639953
transform 1 0 14978 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_145
timestamp 1607639953
transform 1 0 14426 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_137
timestamp 1607639953
transform 1 0 13690 0 -1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _091_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607639953
transform 1 0 14702 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_171
timestamp 1607639953
transform 1 0 16818 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_159
timestamp 1607639953
transform 1 0 15714 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_168
timestamp 1607639953
transform 1 0 16542 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_156
timestamp 1607639953
transform 1 0 15438 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_208
timestamp 1607639953
transform 1 0 15346 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_196
timestamp 1607639953
transform 1 0 19118 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_184
timestamp 1607639953
transform 1 0 18014 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_187
timestamp 1607639953
transform 1 0 18290 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_180
timestamp 1607639953
transform 1 0 17646 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_226
timestamp 1607639953
transform 1 0 17922 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_209
timestamp 1607639953
transform 1 0 18198 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_220
timestamp 1607639953
transform 1 0 21326 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_208
timestamp 1607639953
transform 1 0 20222 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_218
timestamp 1607639953
transform 1 0 21142 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_211
timestamp 1607639953
transform 1 0 20498 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_199
timestamp 1607639953
transform 1 0 19394 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_210
timestamp 1607639953
transform 1 0 21050 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_232
timestamp 1607639953
transform 1 0 22430 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_242
timestamp 1607639953
transform 1 0 23350 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_230
timestamp 1607639953
transform 1 0 22246 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_257
timestamp 1607639953
transform 1 0 24730 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_245
timestamp 1607639953
transform 1 0 23626 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_261
timestamp 1607639953
transform 1 0 25098 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_249
timestamp 1607639953
transform 1 0 23994 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_227
timestamp 1607639953
transform 1 0 23534 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_211
timestamp 1607639953
transform 1 0 23902 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_281
timestamp 1607639953
transform 1 0 26938 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_269
timestamp 1607639953
transform 1 0 25834 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_280
timestamp 1607639953
transform 1 0 26846 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_273
timestamp 1607639953
transform 1 0 26202 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_212
timestamp 1607639953
transform 1 0 26754 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_306
timestamp 1607639953
transform 1 0 29238 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_293
timestamp 1607639953
transform 1 0 28042 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_304
timestamp 1607639953
transform 1 0 29054 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_292
timestamp 1607639953
transform 1 0 27950 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_228
timestamp 1607639953
transform 1 0 29146 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_330
timestamp 1607639953
transform 1 0 31446 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_318
timestamp 1607639953
transform 1 0 30342 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_323
timestamp 1607639953
transform 1 0 30802 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_311
timestamp 1607639953
transform 1 0 29698 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_213
timestamp 1607639953
transform 1 0 29606 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_342
timestamp 1607639953
transform 1 0 32550 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_342
timestamp 1607639953
transform 1 0 32550 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_335
timestamp 1607639953
transform 1 0 31906 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_214
timestamp 1607639953
transform 1 0 32458 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_367
timestamp 1607639953
transform 1 0 34850 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_354
timestamp 1607639953
transform 1 0 33654 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_373
timestamp 1607639953
transform 1 0 35402 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_366
timestamp 1607639953
transform 1 0 34758 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_354
timestamp 1607639953
transform 1 0 33654 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_229
timestamp 1607639953
transform 1 0 34758 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_215
timestamp 1607639953
transform 1 0 35310 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_391
timestamp 1607639953
transform 1 0 37058 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_379
timestamp 1607639953
transform 1 0 35954 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_385
timestamp 1607639953
transform 1 0 36506 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_415
timestamp 1607639953
transform 1 0 39266 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_403
timestamp 1607639953
transform 1 0 38162 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_416
timestamp 1607639953
transform 1 0 39358 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_404
timestamp 1607639953
transform 1 0 38254 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_397
timestamp 1607639953
transform 1 0 37610 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_216
timestamp 1607639953
transform 1 0 38162 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_440
timestamp 1607639953
transform 1 0 41566 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_428
timestamp 1607639953
transform 1 0 40462 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_435
timestamp 1607639953
transform 1 0 41106 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_428
timestamp 1607639953
transform 1 0 40462 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_230
timestamp 1607639953
transform 1 0 40370 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_217
timestamp 1607639953
transform 1 0 41014 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_452
timestamp 1607639953
transform 1 0 42670 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_459
timestamp 1607639953
transform 1 0 43314 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_447
timestamp 1607639953
transform 1 0 42210 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_476
timestamp 1607639953
transform 1 0 44878 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_464
timestamp 1607639953
transform 1 0 43774 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_478
timestamp 1607639953
transform 1 0 45062 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_466
timestamp 1607639953
transform 1 0 43958 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_218
timestamp 1607639953
transform 1 0 43866 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_501
timestamp 1607639953
transform 1 0 47178 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_489
timestamp 1607639953
transform 1 0 46074 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_497
timestamp 1607639953
transform 1 0 46810 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_490
timestamp 1607639953
transform 1 0 46166 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_231
timestamp 1607639953
transform 1 0 45982 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_219
timestamp 1607639953
transform 1 0 46718 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_525
timestamp 1607639953
transform 1 0 49386 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_513
timestamp 1607639953
transform 1 0 48282 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_528
timestamp 1607639953
transform 1 0 49662 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_521
timestamp 1607639953
transform 1 0 49018 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_509
timestamp 1607639953
transform 1 0 47914 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_220
timestamp 1607639953
transform 1 0 49570 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_550
timestamp 1607639953
transform 1 0 51686 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_537
timestamp 1607639953
transform 1 0 50490 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_540
timestamp 1607639953
transform 1 0 50766 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_232
timestamp 1607639953
transform 1 0 51594 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_562
timestamp 1607639953
transform 1 0 52790 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_571
timestamp 1607639953
transform 1 0 53618 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_559
timestamp 1607639953
transform 1 0 52514 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_552
timestamp 1607639953
transform 1 0 51870 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_221
timestamp 1607639953
transform 1 0 52422 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_586
timestamp 1607639953
transform 1 0 54998 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_574
timestamp 1607639953
transform 1 0 53894 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_590
timestamp 1607639953
transform 1 0 55366 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_583
timestamp 1607639953
transform 1 0 54722 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_222
timestamp 1607639953
transform 1 0 55274 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_611
timestamp 1607639953
transform 1 0 57298 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_598
timestamp 1607639953
transform 1 0 56102 0 1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_614
timestamp 1607639953
transform 1 0 57574 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_602
timestamp 1607639953
transform 1 0 56470 0 -1 2720
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_233
timestamp 1607639953
transform 1 0 57206 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_623
timestamp 1607639953
transform 1 0 58402 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_621
timestamp 1607639953
transform 1 0 58218 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_223
timestamp 1607639953
transform 1 0 58126 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1607639953
transform -1 0 58862 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1607639953
transform -1 0 58862 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_12
timestamp 1607639953
transform 1 0 2190 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_3
timestamp 1607639953
transform 1 0 1362 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1607639953
transform 1 0 1086 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _053_
timestamp 1607639953
transform 1 0 1914 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_44
timestamp 1607639953
transform 1 0 5134 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_32
timestamp 1607639953
transform 1 0 4030 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_30 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1607639953
transform 1 0 3846 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_24
timestamp 1607639953
transform 1 0 3294 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_234
timestamp 1607639953
transform 1 0 3938 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_56
timestamp 1607639953
transform 1 0 6238 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_80
timestamp 1607639953
transform 1 0 8446 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_68
timestamp 1607639953
transform 1 0 7342 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_105
timestamp 1607639953
transform 1 0 10746 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_93
timestamp 1607639953
transform 1 0 9642 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_235
timestamp 1607639953
transform 1 0 9550 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_125
timestamp 1607639953
transform 1 0 12586 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_121
timestamp 1607639953
transform 1 0 12218 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_117
timestamp 1607639953
transform 1 0 11850 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _150_
timestamp 1607639953
transform 1 0 12310 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_154
timestamp 1607639953
transform 1 0 15254 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_149
timestamp 1607639953
transform 1 0 14794 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_137
timestamp 1607639953
transform 1 0 13690 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_236
timestamp 1607639953
transform 1 0 15162 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_166
timestamp 1607639953
transform 1 0 16358 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_190
timestamp 1607639953
transform 1 0 18566 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_178
timestamp 1607639953
transform 1 0 17462 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_215
timestamp 1607639953
transform 1 0 20866 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_202
timestamp 1607639953
transform 1 0 19670 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_237
timestamp 1607639953
transform 1 0 20774 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_239
timestamp 1607639953
transform 1 0 23074 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_227
timestamp 1607639953
transform 1 0 21970 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_263
timestamp 1607639953
transform 1 0 25282 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_251
timestamp 1607639953
transform 1 0 24178 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_276
timestamp 1607639953
transform 1 0 26478 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_238
timestamp 1607639953
transform 1 0 26386 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_300
timestamp 1607639953
transform 1 0 28686 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_288
timestamp 1607639953
transform 1 0 27582 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_324
timestamp 1607639953
transform 1 0 30894 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_312
timestamp 1607639953
transform 1 0 29790 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_349
timestamp 1607639953
transform 1 0 33194 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_337
timestamp 1607639953
transform 1 0 32090 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_239
timestamp 1607639953
transform 1 0 31998 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_373
timestamp 1607639953
transform 1 0 35402 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_361
timestamp 1607639953
transform 1 0 34298 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_385
timestamp 1607639953
transform 1 0 36506 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_410
timestamp 1607639953
transform 1 0 38806 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_398
timestamp 1607639953
transform 1 0 37702 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_240
timestamp 1607639953
transform 1 0 37610 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_434
timestamp 1607639953
transform 1 0 41014 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_422
timestamp 1607639953
transform 1 0 39910 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_459
timestamp 1607639953
transform 1 0 43314 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_457
timestamp 1607639953
transform 1 0 43130 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_449
timestamp 1607639953
transform 1 0 42394 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_241
timestamp 1607639953
transform 1 0 43222 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _028_
timestamp 1607639953
transform 1 0 42118 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_483
timestamp 1607639953
transform 1 0 45522 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_471
timestamp 1607639953
transform 1 0 44418 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_495
timestamp 1607639953
transform 1 0 46626 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_520
timestamp 1607639953
transform 1 0 48926 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_507
timestamp 1607639953
transform 1 0 47730 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_242
timestamp 1607639953
transform 1 0 48834 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_544
timestamp 1607639953
transform 1 0 51134 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_532
timestamp 1607639953
transform 1 0 50030 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_568
timestamp 1607639953
transform 1 0 53342 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_556
timestamp 1607639953
transform 1 0 52238 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_590
timestamp 1607639953
transform 1 0 55366 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_581
timestamp 1607639953
transform 1 0 54538 0 -1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_243
timestamp 1607639953
transform 1 0 54446 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _174_
timestamp 1607639953
transform 1 0 55090 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_614
timestamp 1607639953
transform 1 0 57574 0 -1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_602
timestamp 1607639953
transform 1 0 56470 0 -1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_622
timestamp 1607639953
transform 1 0 58310 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1607639953
transform -1 0 58862 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1607639953
transform 1 0 2466 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1607639953
transform 1 0 1362 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1607639953
transform 1 0 1086 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1607639953
transform 1 0 4674 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1607639953
transform 1 0 3570 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_62
timestamp 1607639953
transform 1 0 6790 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_59
timestamp 1607639953
transform 1 0 6514 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_51
timestamp 1607639953
transform 1 0 5778 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_244
timestamp 1607639953
transform 1 0 6698 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_84
timestamp 1607639953
transform 1 0 8814 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_74
timestamp 1607639953
transform 1 0 7894 0 1 3808
box -38 -48 222 592
use AND2X2  AND2X2
timestamp 1608117647
transform 1 0 8078 0 1 3808
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILLER_3_108
timestamp 1607639953
transform 1 0 11022 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_96
timestamp 1607639953
transform 1 0 9918 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_123
timestamp 1607639953
transform 1 0 12402 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_120
timestamp 1607639953
transform 1 0 12126 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_245
timestamp 1607639953
transform 1 0 12310 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_147
timestamp 1607639953
transform 1 0 14610 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_135
timestamp 1607639953
transform 1 0 13506 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_171
timestamp 1607639953
transform 1 0 16818 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_159
timestamp 1607639953
transform 1 0 15714 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_196
timestamp 1607639953
transform 1 0 19118 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_184
timestamp 1607639953
transform 1 0 18014 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_246
timestamp 1607639953
transform 1 0 17922 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_220
timestamp 1607639953
transform 1 0 21326 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_208
timestamp 1607639953
transform 1 0 20222 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_232
timestamp 1607639953
transform 1 0 22430 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_260
timestamp 1607639953
transform 1 0 25006 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_248
timestamp 1607639953
transform 1 0 23902 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_247
timestamp 1607639953
transform 1 0 23534 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _068_
timestamp 1607639953
transform 1 0 23626 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_284
timestamp 1607639953
transform 1 0 27214 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_272
timestamp 1607639953
transform 1 0 26110 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_306
timestamp 1607639953
transform 1 0 29238 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_304
timestamp 1607639953
transform 1 0 29054 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_296
timestamp 1607639953
transform 1 0 28318 0 1 3808
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_248
timestamp 1607639953
transform 1 0 29146 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_330
timestamp 1607639953
transform 1 0 31446 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_318
timestamp 1607639953
transform 1 0 30342 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_342
timestamp 1607639953
transform 1 0 32550 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_367
timestamp 1607639953
transform 1 0 34850 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_354
timestamp 1607639953
transform 1 0 33654 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_249
timestamp 1607639953
transform 1 0 34758 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_391
timestamp 1607639953
transform 1 0 37058 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_379
timestamp 1607639953
transform 1 0 35954 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_415
timestamp 1607639953
transform 1 0 39266 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_403
timestamp 1607639953
transform 1 0 38162 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_440
timestamp 1607639953
transform 1 0 41566 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_428
timestamp 1607639953
transform 1 0 40462 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_250
timestamp 1607639953
transform 1 0 40370 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_452
timestamp 1607639953
transform 1 0 42670 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_476
timestamp 1607639953
transform 1 0 44878 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_464
timestamp 1607639953
transform 1 0 43774 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_501
timestamp 1607639953
transform 1 0 47178 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_489
timestamp 1607639953
transform 1 0 46074 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_251
timestamp 1607639953
transform 1 0 45982 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_525
timestamp 1607639953
transform 1 0 49386 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_513
timestamp 1607639953
transform 1 0 48282 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_550
timestamp 1607639953
transform 1 0 51686 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_537
timestamp 1607639953
transform 1 0 50490 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_252
timestamp 1607639953
transform 1 0 51594 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_562
timestamp 1607639953
transform 1 0 52790 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_586
timestamp 1607639953
transform 1 0 54998 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_574
timestamp 1607639953
transform 1 0 53894 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_611
timestamp 1607639953
transform 1 0 57298 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_598
timestamp 1607639953
transform 1 0 56102 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_253
timestamp 1607639953
transform 1 0 57206 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_623
timestamp 1607639953
transform 1 0 58402 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1607639953
transform -1 0 58862 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_15
timestamp 1607639953
transform 1 0 2466 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_3
timestamp 1607639953
transform 1 0 1362 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1607639953
transform 1 0 1086 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_44
timestamp 1607639953
transform 1 0 5134 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_32
timestamp 1607639953
transform 1 0 4030 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_27
timestamp 1607639953
transform 1 0 3570 0 -1 4896
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_254
timestamp 1607639953
transform 1 0 3938 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_56
timestamp 1607639953
transform 1 0 6238 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_80
timestamp 1607639953
transform 1 0 8446 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_68
timestamp 1607639953
transform 1 0 7342 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_105
timestamp 1607639953
transform 1 0 10746 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_93
timestamp 1607639953
transform 1 0 9642 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_255
timestamp 1607639953
transform 1 0 9550 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_129
timestamp 1607639953
transform 1 0 12954 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_117
timestamp 1607639953
transform 1 0 11850 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_154
timestamp 1607639953
transform 1 0 15254 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1607639953
transform 1 0 14058 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_256
timestamp 1607639953
transform 1 0 15162 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_166
timestamp 1607639953
transform 1 0 16358 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_190
timestamp 1607639953
transform 1 0 18566 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_178
timestamp 1607639953
transform 1 0 17462 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_215
timestamp 1607639953
transform 1 0 20866 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_202
timestamp 1607639953
transform 1 0 19670 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_257
timestamp 1607639953
transform 1 0 20774 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_239
timestamp 1607639953
transform 1 0 23074 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_227
timestamp 1607639953
transform 1 0 21970 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_263
timestamp 1607639953
transform 1 0 25282 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_251
timestamp 1607639953
transform 1 0 24178 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_276
timestamp 1607639953
transform 1 0 26478 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_258
timestamp 1607639953
transform 1 0 26386 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_300
timestamp 1607639953
transform 1 0 28686 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_288
timestamp 1607639953
transform 1 0 27582 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_324
timestamp 1607639953
transform 1 0 30894 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_312
timestamp 1607639953
transform 1 0 29790 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_349
timestamp 1607639953
transform 1 0 33194 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_337
timestamp 1607639953
transform 1 0 32090 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_259
timestamp 1607639953
transform 1 0 31998 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_373
timestamp 1607639953
transform 1 0 35402 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_361
timestamp 1607639953
transform 1 0 34298 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_385
timestamp 1607639953
transform 1 0 36506 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_410
timestamp 1607639953
transform 1 0 38806 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_398
timestamp 1607639953
transform 1 0 37702 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_260
timestamp 1607639953
transform 1 0 37610 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_434
timestamp 1607639953
transform 1 0 41014 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_422
timestamp 1607639953
transform 1 0 39910 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_459
timestamp 1607639953
transform 1 0 43314 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_446
timestamp 1607639953
transform 1 0 42118 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_261
timestamp 1607639953
transform 1 0 43222 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_483
timestamp 1607639953
transform 1 0 45522 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_471
timestamp 1607639953
transform 1 0 44418 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_495
timestamp 1607639953
transform 1 0 46626 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_520
timestamp 1607639953
transform 1 0 48926 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_507
timestamp 1607639953
transform 1 0 47730 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_262
timestamp 1607639953
transform 1 0 48834 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_544
timestamp 1607639953
transform 1 0 51134 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_532
timestamp 1607639953
transform 1 0 50030 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_568
timestamp 1607639953
transform 1 0 53342 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_556
timestamp 1607639953
transform 1 0 52238 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_593
timestamp 1607639953
transform 1 0 55642 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_581
timestamp 1607639953
transform 1 0 54538 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_263
timestamp 1607639953
transform 1 0 54446 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_605
timestamp 1607639953
transform 1 0 56746 0 -1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_617
timestamp 1607639953
transform 1 0 57850 0 -1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1607639953
transform -1 0 58862 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_15
timestamp 1607639953
transform 1 0 2466 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1607639953
transform 1 0 1362 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1607639953
transform 1 0 1086 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_39
timestamp 1607639953
transform 1 0 4674 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_27
timestamp 1607639953
transform 1 0 3570 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_62
timestamp 1607639953
transform 1 0 6790 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_59
timestamp 1607639953
transform 1 0 6514 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_51
timestamp 1607639953
transform 1 0 5778 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_264
timestamp 1607639953
transform 1 0 6698 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_84
timestamp 1607639953
transform 1 0 8814 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_74
timestamp 1607639953
transform 1 0 7894 0 1 4896
box -38 -48 222 592
use AOI21X1  AOI21X1
timestamp 1608117647
transform 1 0 8078 0 1 4896
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILLER_5_108
timestamp 1607639953
transform 1 0 11022 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_96
timestamp 1607639953
transform 1 0 9918 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_123
timestamp 1607639953
transform 1 0 12402 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_120
timestamp 1607639953
transform 1 0 12126 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_265
timestamp 1607639953
transform 1 0 12310 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_147
timestamp 1607639953
transform 1 0 14610 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_135
timestamp 1607639953
transform 1 0 13506 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_171
timestamp 1607639953
transform 1 0 16818 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_159
timestamp 1607639953
transform 1 0 15714 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_196
timestamp 1607639953
transform 1 0 19118 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_184
timestamp 1607639953
transform 1 0 18014 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_266
timestamp 1607639953
transform 1 0 17922 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_220
timestamp 1607639953
transform 1 0 21326 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_208
timestamp 1607639953
transform 1 0 20222 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_232
timestamp 1607639953
transform 1 0 22430 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_257
timestamp 1607639953
transform 1 0 24730 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_245
timestamp 1607639953
transform 1 0 23626 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_267
timestamp 1607639953
transform 1 0 23534 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_281
timestamp 1607639953
transform 1 0 26938 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_269
timestamp 1607639953
transform 1 0 25834 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_306
timestamp 1607639953
transform 1 0 29238 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_293
timestamp 1607639953
transform 1 0 28042 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_268
timestamp 1607639953
transform 1 0 29146 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_330
timestamp 1607639953
transform 1 0 31446 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_318
timestamp 1607639953
transform 1 0 30342 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_350
timestamp 1607639953
transform 1 0 33286 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_342
timestamp 1607639953
transform 1 0 32550 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_367
timestamp 1607639953
transform 1 0 34850 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_364
timestamp 1607639953
transform 1 0 34574 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_356
timestamp 1607639953
transform 1 0 33838 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_269
timestamp 1607639953
transform 1 0 34758 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _086_
timestamp 1607639953
transform 1 0 33562 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_391
timestamp 1607639953
transform 1 0 37058 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_379
timestamp 1607639953
transform 1 0 35954 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_415
timestamp 1607639953
transform 1 0 39266 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_403
timestamp 1607639953
transform 1 0 38162 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_440
timestamp 1607639953
transform 1 0 41566 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_428
timestamp 1607639953
transform 1 0 40462 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_270
timestamp 1607639953
transform 1 0 40370 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_452
timestamp 1607639953
transform 1 0 42670 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_476
timestamp 1607639953
transform 1 0 44878 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_464
timestamp 1607639953
transform 1 0 43774 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_505
timestamp 1607639953
transform 1 0 47546 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_493
timestamp 1607639953
transform 1 0 46442 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_489
timestamp 1607639953
transform 1 0 46074 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_271
timestamp 1607639953
transform 1 0 45982 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _012_
timestamp 1607639953
transform 1 0 46166 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_517
timestamp 1607639953
transform 1 0 48650 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_550
timestamp 1607639953
transform 1 0 51686 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_541
timestamp 1607639953
transform 1 0 50858 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_529
timestamp 1607639953
transform 1 0 49754 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_272
timestamp 1607639953
transform 1 0 51594 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_562
timestamp 1607639953
transform 1 0 52790 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_588
timestamp 1607639953
transform 1 0 55182 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_582
timestamp 1607639953
transform 1 0 54630 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_5_574
timestamp 1607639953
transform 1 0 53894 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _140_
timestamp 1607639953
transform 1 0 54906 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_611
timestamp 1607639953
transform 1 0 57298 0 1 4896
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_608
timestamp 1607639953
transform 1 0 57022 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_5_600
timestamp 1607639953
transform 1 0 56286 0 1 4896
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_273
timestamp 1607639953
transform 1 0 57206 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_623
timestamp 1607639953
transform 1 0 58402 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1607639953
transform -1 0 58862 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_15
timestamp 1607639953
transform 1 0 2466 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1607639953
transform 1 0 1362 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_15
timestamp 1607639953
transform 1 0 2466 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_3
timestamp 1607639953
transform 1 0 1362 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1607639953
transform 1 0 1086 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1607639953
transform 1 0 1086 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_39
timestamp 1607639953
transform 1 0 4674 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_27
timestamp 1607639953
transform 1 0 3570 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_44
timestamp 1607639953
transform 1 0 5134 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_32
timestamp 1607639953
transform 1 0 4030 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_27
timestamp 1607639953
transform 1 0 3570 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_274
timestamp 1607639953
transform 1 0 3938 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_62
timestamp 1607639953
transform 1 0 6790 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1607639953
transform 1 0 6514 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_51
timestamp 1607639953
transform 1 0 5778 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_63
timestamp 1607639953
transform 1 0 6882 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_51
timestamp 1607639953
transform 1 0 5778 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_284
timestamp 1607639953
transform 1 0 6698 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _120_
timestamp 1607639953
transform 1 0 5502 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_86
timestamp 1607639953
transform 1 0 8998 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_7_74
timestamp 1607639953
transform 1 0 7894 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_87
timestamp 1607639953
transform 1 0 9090 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_75
timestamp 1607639953
transform 1 0 7986 0 -1 5984
box -38 -48 1142 592
use AOI22X1  AOI22X1
timestamp 1608117647
transform 1 0 8078 0 1 5984
box 0 -48 920 592
use sky130_fd_sc_hd__decap_12  FILLER_7_110
timestamp 1607639953
transform 1 0 11206 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_98
timestamp 1607639953
transform 1 0 10102 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_103
timestamp 1607639953
transform 1 0 10562 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_99
timestamp 1607639953
transform 1 0 10194 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_93
timestamp 1607639953
transform 1 0 9642 0 -1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_91
timestamp 1607639953
transform 1 0 9458 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_275
timestamp 1607639953
transform 1 0 9550 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _011_
timestamp 1607639953
transform 1 0 10286 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_123
timestamp 1607639953
transform 1 0 12402 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_127
timestamp 1607639953
transform 1 0 12770 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_115
timestamp 1607639953
transform 1 0 11666 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_285
timestamp 1607639953
transform 1 0 12310 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_147
timestamp 1607639953
transform 1 0 14610 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_135
timestamp 1607639953
transform 1 0 13506 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_154
timestamp 1607639953
transform 1 0 15254 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_151
timestamp 1607639953
transform 1 0 14978 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_139
timestamp 1607639953
transform 1 0 13874 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_276
timestamp 1607639953
transform 1 0 15162 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_171
timestamp 1607639953
transform 1 0 16818 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_159
timestamp 1607639953
transform 1 0 15714 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_166
timestamp 1607639953
transform 1 0 16358 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_196
timestamp 1607639953
transform 1 0 19118 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_184
timestamp 1607639953
transform 1 0 18014 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_190
timestamp 1607639953
transform 1 0 18566 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_178
timestamp 1607639953
transform 1 0 17462 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_286
timestamp 1607639953
transform 1 0 17922 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_220
timestamp 1607639953
transform 1 0 21326 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_208
timestamp 1607639953
transform 1 0 20222 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_215
timestamp 1607639953
transform 1 0 20866 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_202
timestamp 1607639953
transform 1 0 19670 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_277
timestamp 1607639953
transform 1 0 20774 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_232
timestamp 1607639953
transform 1 0 22430 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_241
timestamp 1607639953
transform 1 0 23258 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_229
timestamp 1607639953
transform 1 0 22154 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_223
timestamp 1607639953
transform 1 0 21602 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _016_
timestamp 1607639953
transform 1 0 21878 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_257
timestamp 1607639953
transform 1 0 24730 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_245
timestamp 1607639953
transform 1 0 23626 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_253
timestamp 1607639953
transform 1 0 24362 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_287
timestamp 1607639953
transform 1 0 23534 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_281
timestamp 1607639953
transform 1 0 26938 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_269
timestamp 1607639953
transform 1 0 25834 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_276
timestamp 1607639953
transform 1 0 26478 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_273
timestamp 1607639953
transform 1 0 26202 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_265
timestamp 1607639953
transform 1 0 25466 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_278
timestamp 1607639953
transform 1 0 26386 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_306
timestamp 1607639953
transform 1 0 29238 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_293
timestamp 1607639953
transform 1 0 28042 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_307
timestamp 1607639953
transform 1 0 29330 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_295
timestamp 1607639953
transform 1 0 28226 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_288
timestamp 1607639953
transform 1 0 27582 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_288
timestamp 1607639953
transform 1 0 29146 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _039_
timestamp 1607639953
transform 1 0 27950 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_330
timestamp 1607639953
transform 1 0 31446 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_318
timestamp 1607639953
transform 1 0 30342 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_319
timestamp 1607639953
transform 1 0 30434 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_342
timestamp 1607639953
transform 1 0 32550 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_349
timestamp 1607639953
transform 1 0 33194 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_337
timestamp 1607639953
transform 1 0 32090 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_335
timestamp 1607639953
transform 1 0 31906 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_331
timestamp 1607639953
transform 1 0 31538 0 -1 5984
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_279
timestamp 1607639953
transform 1 0 31998 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_367
timestamp 1607639953
transform 1 0 34850 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_364
timestamp 1607639953
transform 1 0 34574 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_7_360
timestamp 1607639953
transform 1 0 34206 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_354
timestamp 1607639953
transform 1 0 33654 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_373
timestamp 1607639953
transform 1 0 35402 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_361
timestamp 1607639953
transform 1 0 34298 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_289
timestamp 1607639953
transform 1 0 34758 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _061_
timestamp 1607639953
transform 1 0 34298 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _035_
timestamp 1607639953
transform 1 0 35494 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_390
timestamp 1607639953
transform 1 0 36966 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_378
timestamp 1607639953
transform 1 0 35862 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_389
timestamp 1607639953
transform 1 0 36874 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_377
timestamp 1607639953
transform 1 0 35770 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _170_
timestamp 1607639953
transform 1 0 35586 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_7_414
timestamp 1607639953
transform 1 0 39174 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_402
timestamp 1607639953
transform 1 0 38070 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_410
timestamp 1607639953
transform 1 0 38806 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_398
timestamp 1607639953
transform 1 0 37702 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_280
timestamp 1607639953
transform 1 0 37610 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_440
timestamp 1607639953
transform 1 0 41566 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_428
timestamp 1607639953
transform 1 0 40462 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_426
timestamp 1607639953
transform 1 0 40278 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_434
timestamp 1607639953
transform 1 0 41014 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_422
timestamp 1607639953
transform 1 0 39910 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_290
timestamp 1607639953
transform 1 0 40370 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_458
timestamp 1607639953
transform 1 0 43222 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_454
timestamp 1607639953
transform 1 0 42854 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_448
timestamp 1607639953
transform 1 0 42302 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_6_459
timestamp 1607639953
transform 1 0 43314 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_446
timestamp 1607639953
transform 1 0 42118 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_281
timestamp 1607639953
transform 1 0 43222 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _115_
timestamp 1607639953
transform 1 0 42946 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _088_
timestamp 1607639953
transform 1 0 42578 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_7_482
timestamp 1607639953
transform 1 0 45430 0 1 5984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_7_470
timestamp 1607639953
transform 1 0 44326 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_483
timestamp 1607639953
transform 1 0 45522 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_471
timestamp 1607639953
transform 1 0 44418 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_501
timestamp 1607639953
transform 1 0 47178 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_489
timestamp 1607639953
transform 1 0 46074 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_495
timestamp 1607639953
transform 1 0 46626 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_291
timestamp 1607639953
transform 1 0 45982 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_525
timestamp 1607639953
transform 1 0 49386 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_513
timestamp 1607639953
transform 1 0 48282 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_520
timestamp 1607639953
transform 1 0 48926 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_507
timestamp 1607639953
transform 1 0 47730 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_282
timestamp 1607639953
transform 1 0 48834 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_550
timestamp 1607639953
transform 1 0 51686 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_537
timestamp 1607639953
transform 1 0 50490 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_544
timestamp 1607639953
transform 1 0 51134 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_532
timestamp 1607639953
transform 1 0 50030 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_292
timestamp 1607639953
transform 1 0 51594 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_562
timestamp 1607639953
transform 1 0 52790 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_568
timestamp 1607639953
transform 1 0 53342 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_556
timestamp 1607639953
transform 1 0 52238 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_586
timestamp 1607639953
transform 1 0 54998 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_574
timestamp 1607639953
transform 1 0 53894 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_593
timestamp 1607639953
transform 1 0 55642 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_581
timestamp 1607639953
transform 1 0 54538 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_283
timestamp 1607639953
transform 1 0 54446 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_611
timestamp 1607639953
transform 1 0 57298 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_598
timestamp 1607639953
transform 1 0 56102 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_605
timestamp 1607639953
transform 1 0 56746 0 -1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_293
timestamp 1607639953
transform 1 0 57206 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_7_623
timestamp 1607639953
transform 1 0 58402 0 1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_617
timestamp 1607639953
transform 1 0 57850 0 -1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1607639953
transform -1 0 58862 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1607639953
transform -1 0 58862 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1607639953
transform 1 0 2466 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1607639953
transform 1 0 1362 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1607639953
transform 1 0 1086 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_44
timestamp 1607639953
transform 1 0 5134 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_32
timestamp 1607639953
transform 1 0 4030 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_27
timestamp 1607639953
transform 1 0 3570 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_294
timestamp 1607639953
transform 1 0 3938 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_56
timestamp 1607639953
transform 1 0 6238 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_80
timestamp 1607639953
transform 1 0 8446 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_76
timestamp 1607639953
transform 1 0 8078 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_68
timestamp 1607639953
transform 1 0 7342 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _147_
timestamp 1607639953
transform 1 0 8170 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_105
timestamp 1607639953
transform 1 0 10746 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_93
timestamp 1607639953
transform 1 0 9642 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_295
timestamp 1607639953
transform 1 0 9550 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_129
timestamp 1607639953
transform 1 0 12954 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_117
timestamp 1607639953
transform 1 0 11850 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_154
timestamp 1607639953
transform 1 0 15254 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1607639953
transform 1 0 14058 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_296
timestamp 1607639953
transform 1 0 15162 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_166
timestamp 1607639953
transform 1 0 16358 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_190
timestamp 1607639953
transform 1 0 18566 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_178
timestamp 1607639953
transform 1 0 17462 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_215
timestamp 1607639953
transform 1 0 20866 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_202
timestamp 1607639953
transform 1 0 19670 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_297
timestamp 1607639953
transform 1 0 20774 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_239
timestamp 1607639953
transform 1 0 23074 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_227
timestamp 1607639953
transform 1 0 21970 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_263
timestamp 1607639953
transform 1 0 25282 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_251
timestamp 1607639953
transform 1 0 24178 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_276
timestamp 1607639953
transform 1 0 26478 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_298
timestamp 1607639953
transform 1 0 26386 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_300
timestamp 1607639953
transform 1 0 28686 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_288
timestamp 1607639953
transform 1 0 27582 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_324
timestamp 1607639953
transform 1 0 30894 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_312
timestamp 1607639953
transform 1 0 29790 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_349
timestamp 1607639953
transform 1 0 33194 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_337
timestamp 1607639953
transform 1 0 32090 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_299
timestamp 1607639953
transform 1 0 31998 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_373
timestamp 1607639953
transform 1 0 35402 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_361
timestamp 1607639953
transform 1 0 34298 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_385
timestamp 1607639953
transform 1 0 36506 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_410
timestamp 1607639953
transform 1 0 38806 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_398
timestamp 1607639953
transform 1 0 37702 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_300
timestamp 1607639953
transform 1 0 37610 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_434
timestamp 1607639953
transform 1 0 41014 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_422
timestamp 1607639953
transform 1 0 39910 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_459
timestamp 1607639953
transform 1 0 43314 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_446
timestamp 1607639953
transform 1 0 42118 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_301
timestamp 1607639953
transform 1 0 43222 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_483
timestamp 1607639953
transform 1 0 45522 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_471
timestamp 1607639953
transform 1 0 44418 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_495
timestamp 1607639953
transform 1 0 46626 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_520
timestamp 1607639953
transform 1 0 48926 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_507
timestamp 1607639953
transform 1 0 47730 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_302
timestamp 1607639953
transform 1 0 48834 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_548
timestamp 1607639953
transform 1 0 51502 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_544
timestamp 1607639953
transform 1 0 51134 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_532
timestamp 1607639953
transform 1 0 50030 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _038_
timestamp 1607639953
transform 1 0 51594 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_571
timestamp 1607639953
transform 1 0 53618 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_8_559
timestamp 1607639953
transform 1 0 52514 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_552
timestamp 1607639953
transform 1 0 51870 0 -1 7072
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _067_
timestamp 1607639953
transform 1 0 52238 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_593
timestamp 1607639953
transform 1 0 55642 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_581
timestamp 1607639953
transform 1 0 54538 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_579
timestamp 1607639953
transform 1 0 54354 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_303
timestamp 1607639953
transform 1 0 54446 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_605
timestamp 1607639953
transform 1 0 56746 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_617
timestamp 1607639953
transform 1 0 57850 0 -1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1607639953
transform -1 0 58862 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1607639953
transform 1 0 2466 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1607639953
transform 1 0 1362 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1607639953
transform 1 0 1086 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1607639953
transform 1 0 4674 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1607639953
transform 1 0 3570 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_62
timestamp 1607639953
transform 1 0 6790 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_59
timestamp 1607639953
transform 1 0 6514 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_9_51
timestamp 1607639953
transform 1 0 5778 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_304
timestamp 1607639953
transform 1 0 6698 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_82
timestamp 1607639953
transform 1 0 8630 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_74
timestamp 1607639953
transform 1 0 7894 0 1 7072
box -38 -48 222 592
use BUFX2  BUFX2
timestamp 1608117647
transform 1 0 8078 0 1 7072
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILLER_9_108
timestamp 1607639953
transform 1 0 11022 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_96
timestamp 1607639953
transform 1 0 9918 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_90
timestamp 1607639953
transform 1 0 9366 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _195_
timestamp 1607639953
transform 1 0 9642 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_123
timestamp 1607639953
transform 1 0 12402 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_120
timestamp 1607639953
transform 1 0 12126 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_305
timestamp 1607639953
transform 1 0 12310 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_147
timestamp 1607639953
transform 1 0 14610 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_135
timestamp 1607639953
transform 1 0 13506 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_171
timestamp 1607639953
transform 1 0 16818 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_9_159
timestamp 1607639953
transform 1 0 15714 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_196
timestamp 1607639953
transform 1 0 19118 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_184
timestamp 1607639953
transform 1 0 18014 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_180
timestamp 1607639953
transform 1 0 17646 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_306
timestamp 1607639953
transform 1 0 17922 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _023_
timestamp 1607639953
transform 1 0 17370 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_220
timestamp 1607639953
transform 1 0 21326 0 1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_9_208
timestamp 1607639953
transform 1 0 20222 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_241
timestamp 1607639953
transform 1 0 23258 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_229
timestamp 1607639953
transform 1 0 22154 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _154_
timestamp 1607639953
transform 1 0 21878 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_257
timestamp 1607639953
transform 1 0 24730 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_245
timestamp 1607639953
transform 1 0 23626 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_307
timestamp 1607639953
transform 1 0 23534 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_281
timestamp 1607639953
transform 1 0 26938 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_269
timestamp 1607639953
transform 1 0 25834 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_306
timestamp 1607639953
transform 1 0 29238 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_293
timestamp 1607639953
transform 1 0 28042 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_308
timestamp 1607639953
transform 1 0 29146 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_330
timestamp 1607639953
transform 1 0 31446 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_318
timestamp 1607639953
transform 1 0 30342 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_342
timestamp 1607639953
transform 1 0 32550 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_367
timestamp 1607639953
transform 1 0 34850 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_354
timestamp 1607639953
transform 1 0 33654 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_309
timestamp 1607639953
transform 1 0 34758 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_391
timestamp 1607639953
transform 1 0 37058 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_379
timestamp 1607639953
transform 1 0 35954 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_415
timestamp 1607639953
transform 1 0 39266 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_403
timestamp 1607639953
transform 1 0 38162 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_440
timestamp 1607639953
transform 1 0 41566 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_428
timestamp 1607639953
transform 1 0 40462 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_310
timestamp 1607639953
transform 1 0 40370 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_452
timestamp 1607639953
transform 1 0 42670 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_478
timestamp 1607639953
transform 1 0 45062 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_472
timestamp 1607639953
transform 1 0 44510 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_464
timestamp 1607639953
transform 1 0 43774 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _165_
timestamp 1607639953
transform 1 0 44786 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_501
timestamp 1607639953
transform 1 0 47178 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_489
timestamp 1607639953
transform 1 0 46074 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_486
timestamp 1607639953
transform 1 0 45798 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_311
timestamp 1607639953
transform 1 0 45982 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_9_525
timestamp 1607639953
transform 1 0 49386 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_513
timestamp 1607639953
transform 1 0 48282 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _054_
timestamp 1607639953
transform 1 0 49478 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_550
timestamp 1607639953
transform 1 0 51686 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_541
timestamp 1607639953
transform 1 0 50858 0 1 7072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_9_529
timestamp 1607639953
transform 1 0 49754 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_312
timestamp 1607639953
transform 1 0 51594 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_562
timestamp 1607639953
transform 1 0 52790 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_586
timestamp 1607639953
transform 1 0 54998 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_574
timestamp 1607639953
transform 1 0 53894 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_611
timestamp 1607639953
transform 1 0 57298 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_598
timestamp 1607639953
transform 1 0 56102 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_313
timestamp 1607639953
transform 1 0 57206 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_623
timestamp 1607639953
transform 1 0 58402 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1607639953
transform -1 0 58862 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1607639953
transform 1 0 2466 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1607639953
transform 1 0 1362 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1607639953
transform 1 0 1086 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_44
timestamp 1607639953
transform 1 0 5134 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_32
timestamp 1607639953
transform 1 0 4030 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_27
timestamp 1607639953
transform 1 0 3570 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_314
timestamp 1607639953
transform 1 0 3938 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_56
timestamp 1607639953
transform 1 0 6238 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_80
timestamp 1607639953
transform 1 0 8446 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_68
timestamp 1607639953
transform 1 0 7342 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_105
timestamp 1607639953
transform 1 0 10746 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_93
timestamp 1607639953
transform 1 0 9642 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_315
timestamp 1607639953
transform 1 0 9550 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _084_
timestamp 1607639953
transform 1 0 11022 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_123
timestamp 1607639953
transform 1 0 12402 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_111
timestamp 1607639953
transform 1 0 11298 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_154
timestamp 1607639953
transform 1 0 15254 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_147
timestamp 1607639953
transform 1 0 14610 0 -1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_10_135
timestamp 1607639953
transform 1 0 13506 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_316
timestamp 1607639953
transform 1 0 15162 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_166
timestamp 1607639953
transform 1 0 16358 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_190
timestamp 1607639953
transform 1 0 18566 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_178
timestamp 1607639953
transform 1 0 17462 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_215
timestamp 1607639953
transform 1 0 20866 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_202
timestamp 1607639953
transform 1 0 19670 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_317
timestamp 1607639953
transform 1 0 20774 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_239
timestamp 1607639953
transform 1 0 23074 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_227
timestamp 1607639953
transform 1 0 21970 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_263
timestamp 1607639953
transform 1 0 25282 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_251
timestamp 1607639953
transform 1 0 24178 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_276
timestamp 1607639953
transform 1 0 26478 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_318
timestamp 1607639953
transform 1 0 26386 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_300
timestamp 1607639953
transform 1 0 28686 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_288
timestamp 1607639953
transform 1 0 27582 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_324
timestamp 1607639953
transform 1 0 30894 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_312
timestamp 1607639953
transform 1 0 29790 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_349
timestamp 1607639953
transform 1 0 33194 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_337
timestamp 1607639953
transform 1 0 32090 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_319
timestamp 1607639953
transform 1 0 31998 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_373
timestamp 1607639953
transform 1 0 35402 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_361
timestamp 1607639953
transform 1 0 34298 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_385
timestamp 1607639953
transform 1 0 36506 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_410
timestamp 1607639953
transform 1 0 38806 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_398
timestamp 1607639953
transform 1 0 37702 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_320
timestamp 1607639953
transform 1 0 37610 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_434
timestamp 1607639953
transform 1 0 41014 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_422
timestamp 1607639953
transform 1 0 39910 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _071_
timestamp 1607639953
transform 1 0 41382 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_459
timestamp 1607639953
transform 1 0 43314 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_457
timestamp 1607639953
transform 1 0 43130 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_453
timestamp 1607639953
transform 1 0 42762 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_441
timestamp 1607639953
transform 1 0 41658 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_321
timestamp 1607639953
transform 1 0 43222 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_483
timestamp 1607639953
transform 1 0 45522 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_471
timestamp 1607639953
transform 1 0 44418 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_495
timestamp 1607639953
transform 1 0 46626 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_520
timestamp 1607639953
transform 1 0 48926 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_507
timestamp 1607639953
transform 1 0 47730 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_322
timestamp 1607639953
transform 1 0 48834 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_544
timestamp 1607639953
transform 1 0 51134 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_532
timestamp 1607639953
transform 1 0 50030 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_568
timestamp 1607639953
transform 1 0 53342 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_556
timestamp 1607639953
transform 1 0 52238 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_593
timestamp 1607639953
transform 1 0 55642 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_581
timestamp 1607639953
transform 1 0 54538 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_323
timestamp 1607639953
transform 1 0 54446 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_605
timestamp 1607639953
transform 1 0 56746 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_624
timestamp 1607639953
transform 1 0 58494 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_617
timestamp 1607639953
transform 1 0 57850 0 -1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1607639953
transform -1 0 58862 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _085_
timestamp 1607639953
transform 1 0 58218 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1607639953
transform 1 0 2466 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1607639953
transform 1 0 1362 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1607639953
transform 1 0 1086 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1607639953
transform 1 0 4674 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_27
timestamp 1607639953
transform 1 0 3570 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_62
timestamp 1607639953
transform 1 0 6790 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_59
timestamp 1607639953
transform 1 0 6514 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_11_51
timestamp 1607639953
transform 1 0 5778 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_324
timestamp 1607639953
transform 1 0 6698 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_84
timestamp 1607639953
transform 1 0 8814 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_74
timestamp 1607639953
transform 1 0 7894 0 1 8160
box -38 -48 222 592
use BUFX4  BUFX4
timestamp 1608117647
transform 1 0 8078 0 1 8160
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILLER_11_108
timestamp 1607639953
transform 1 0 11022 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_96
timestamp 1607639953
transform 1 0 9918 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_123
timestamp 1607639953
transform 1 0 12402 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_120
timestamp 1607639953
transform 1 0 12126 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_325
timestamp 1607639953
transform 1 0 12310 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_147
timestamp 1607639953
transform 1 0 14610 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_135
timestamp 1607639953
transform 1 0 13506 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_171
timestamp 1607639953
transform 1 0 16818 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_159
timestamp 1607639953
transform 1 0 15714 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_196
timestamp 1607639953
transform 1 0 19118 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_184
timestamp 1607639953
transform 1 0 18014 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_326
timestamp 1607639953
transform 1 0 17922 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_220
timestamp 1607639953
transform 1 0 21326 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_208
timestamp 1607639953
transform 1 0 20222 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_232
timestamp 1607639953
transform 1 0 22430 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_257
timestamp 1607639953
transform 1 0 24730 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_245
timestamp 1607639953
transform 1 0 23626 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_327
timestamp 1607639953
transform 1 0 23534 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_281
timestamp 1607639953
transform 1 0 26938 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_269
timestamp 1607639953
transform 1 0 25834 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_306
timestamp 1607639953
transform 1 0 29238 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_293
timestamp 1607639953
transform 1 0 28042 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_328
timestamp 1607639953
transform 1 0 29146 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_330
timestamp 1607639953
transform 1 0 31446 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_318
timestamp 1607639953
transform 1 0 30342 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_342
timestamp 1607639953
transform 1 0 32550 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_367
timestamp 1607639953
transform 1 0 34850 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_354
timestamp 1607639953
transform 1 0 33654 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_329
timestamp 1607639953
transform 1 0 34758 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_391
timestamp 1607639953
transform 1 0 37058 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_379
timestamp 1607639953
transform 1 0 35954 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_415
timestamp 1607639953
transform 1 0 39266 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_403
timestamp 1607639953
transform 1 0 38162 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _184_
timestamp 1607639953
transform 1 0 39542 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_440
timestamp 1607639953
transform 1 0 41566 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_428
timestamp 1607639953
transform 1 0 40462 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_421
timestamp 1607639953
transform 1 0 39818 0 1 8160
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_330
timestamp 1607639953
transform 1 0 40370 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_452
timestamp 1607639953
transform 1 0 42670 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_476
timestamp 1607639953
transform 1 0 44878 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_464
timestamp 1607639953
transform 1 0 43774 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_501
timestamp 1607639953
transform 1 0 47178 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_489
timestamp 1607639953
transform 1 0 46074 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_331
timestamp 1607639953
transform 1 0 45982 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_525
timestamp 1607639953
transform 1 0 49386 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_513
timestamp 1607639953
transform 1 0 48282 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_550
timestamp 1607639953
transform 1 0 51686 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_537
timestamp 1607639953
transform 1 0 50490 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_332
timestamp 1607639953
transform 1 0 51594 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_562
timestamp 1607639953
transform 1 0 52790 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_586
timestamp 1607639953
transform 1 0 54998 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_574
timestamp 1607639953
transform 1 0 53894 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_614
timestamp 1607639953
transform 1 0 57574 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_11_598
timestamp 1607639953
transform 1 0 56102 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_333
timestamp 1607639953
transform 1 0 57206 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _199_
timestamp 1607639953
transform 1 0 57298 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_11_622
timestamp 1607639953
transform 1 0 58310 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1607639953
transform -1 0 58862 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1607639953
transform 1 0 2466 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1607639953
transform 1 0 1362 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1607639953
transform 1 0 1086 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_44
timestamp 1607639953
transform 1 0 5134 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_32
timestamp 1607639953
transform 1 0 4030 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_27
timestamp 1607639953
transform 1 0 3570 0 -1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_334
timestamp 1607639953
transform 1 0 3938 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_56
timestamp 1607639953
transform 1 0 6238 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_80
timestamp 1607639953
transform 1 0 8446 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_68
timestamp 1607639953
transform 1 0 7342 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_105
timestamp 1607639953
transform 1 0 10746 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_93
timestamp 1607639953
transform 1 0 9642 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_335
timestamp 1607639953
transform 1 0 9550 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_129
timestamp 1607639953
transform 1 0 12954 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_117
timestamp 1607639953
transform 1 0 11850 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_154
timestamp 1607639953
transform 1 0 15254 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_141
timestamp 1607639953
transform 1 0 14058 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_336
timestamp 1607639953
transform 1 0 15162 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_166
timestamp 1607639953
transform 1 0 16358 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_198
timestamp 1607639953
transform 1 0 19302 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_190
timestamp 1607639953
transform 1 0 18566 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_178
timestamp 1607639953
transform 1 0 17462 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_215
timestamp 1607639953
transform 1 0 20866 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_211
timestamp 1607639953
transform 1 0 20498 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_12_203
timestamp 1607639953
transform 1 0 19762 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_337
timestamp 1607639953
transform 1 0 20774 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _022_
timestamp 1607639953
transform 1 0 19486 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_239
timestamp 1607639953
transform 1 0 23074 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_227
timestamp 1607639953
transform 1 0 21970 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_263
timestamp 1607639953
transform 1 0 25282 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_251
timestamp 1607639953
transform 1 0 24178 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_276
timestamp 1607639953
transform 1 0 26478 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_338
timestamp 1607639953
transform 1 0 26386 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_300
timestamp 1607639953
transform 1 0 28686 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_288
timestamp 1607639953
transform 1 0 27582 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_324
timestamp 1607639953
transform 1 0 30894 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_312
timestamp 1607639953
transform 1 0 29790 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_349
timestamp 1607639953
transform 1 0 33194 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_337
timestamp 1607639953
transform 1 0 32090 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_339
timestamp 1607639953
transform 1 0 31998 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_373
timestamp 1607639953
transform 1 0 35402 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_361
timestamp 1607639953
transform 1 0 34298 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_385
timestamp 1607639953
transform 1 0 36506 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_410
timestamp 1607639953
transform 1 0 38806 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_398
timestamp 1607639953
transform 1 0 37702 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_340
timestamp 1607639953
transform 1 0 37610 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_434
timestamp 1607639953
transform 1 0 41014 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_422
timestamp 1607639953
transform 1 0 39910 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_459
timestamp 1607639953
transform 1 0 43314 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_446
timestamp 1607639953
transform 1 0 42118 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_341
timestamp 1607639953
transform 1 0 43222 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_483
timestamp 1607639953
transform 1 0 45522 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_471
timestamp 1607639953
transform 1 0 44418 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_495
timestamp 1607639953
transform 1 0 46626 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_520
timestamp 1607639953
transform 1 0 48926 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_507
timestamp 1607639953
transform 1 0 47730 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_342
timestamp 1607639953
transform 1 0 48834 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_544
timestamp 1607639953
transform 1 0 51134 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_532
timestamp 1607639953
transform 1 0 50030 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_572
timestamp 1607639953
transform 1 0 53710 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_568
timestamp 1607639953
transform 1 0 53342 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_556
timestamp 1607639953
transform 1 0 52238 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _129_
timestamp 1607639953
transform 1 0 53434 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_593
timestamp 1607639953
transform 1 0 55642 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_581
timestamp 1607639953
transform 1 0 54538 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_343
timestamp 1607639953
transform 1 0 54446 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_605
timestamp 1607639953
transform 1 0 56746 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_617
timestamp 1607639953
transform 1 0 57850 0 -1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1607639953
transform -1 0 58862 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1607639953
transform 1 0 2466 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1607639953
transform 1 0 1362 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1607639953
transform 1 0 2466 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1607639953
transform 1 0 1362 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1607639953
transform 1 0 1086 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1607639953
transform 1 0 1086 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_44
timestamp 1607639953
transform 1 0 5134 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_32
timestamp 1607639953
transform 1 0 4030 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_27
timestamp 1607639953
transform 1 0 3570 0 -1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1607639953
transform 1 0 4674 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1607639953
transform 1 0 3570 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_354
timestamp 1607639953
transform 1 0 3938 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_56
timestamp 1607639953
transform 1 0 6238 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_62
timestamp 1607639953
transform 1 0 6790 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_59
timestamp 1607639953
transform 1 0 6514 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_51
timestamp 1607639953
transform 1 0 5778 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_344
timestamp 1607639953
transform 1 0 6698 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_80
timestamp 1607639953
transform 1 0 8446 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_68
timestamp 1607639953
transform 1 0 7342 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_74
timestamp 1607639953
transform 1 0 7894 0 1 9248
box -38 -48 222 592
use CLKBUF1  CLKBUF1
timestamp 1608117647
transform 1 0 8078 0 1 9248
box 0 -48 1656 592
use sky130_fd_sc_hd__decap_12  FILLER_14_105
timestamp 1607639953
transform 1 0 10746 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_93
timestamp 1607639953
transform 1 0 9642 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_106
timestamp 1607639953
transform 1 0 10838 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_94
timestamp 1607639953
transform 1 0 9734 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_355
timestamp 1607639953
transform 1 0 9550 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_129
timestamp 1607639953
transform 1 0 12954 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_117
timestamp 1607639953
transform 1 0 11850 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_123
timestamp 1607639953
transform 1 0 12402 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_118
timestamp 1607639953
transform 1 0 11942 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_345
timestamp 1607639953
transform 1 0 12310 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_154
timestamp 1607639953
transform 1 0 15254 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_141
timestamp 1607639953
transform 1 0 14058 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_147
timestamp 1607639953
transform 1 0 14610 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_135
timestamp 1607639953
transform 1 0 13506 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_356
timestamp 1607639953
transform 1 0 15162 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_166
timestamp 1607639953
transform 1 0 16358 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_171
timestamp 1607639953
transform 1 0 16818 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_159
timestamp 1607639953
transform 1 0 15714 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_190
timestamp 1607639953
transform 1 0 18566 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_178
timestamp 1607639953
transform 1 0 17462 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_196
timestamp 1607639953
transform 1 0 19118 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_184
timestamp 1607639953
transform 1 0 18014 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_346
timestamp 1607639953
transform 1 0 17922 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_215
timestamp 1607639953
transform 1 0 20866 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_202
timestamp 1607639953
transform 1 0 19670 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_220
timestamp 1607639953
transform 1 0 21326 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_208
timestamp 1607639953
transform 1 0 20222 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_357
timestamp 1607639953
transform 1 0 20774 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_239
timestamp 1607639953
transform 1 0 23074 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_227
timestamp 1607639953
transform 1 0 21970 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_232
timestamp 1607639953
transform 1 0 22430 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_263
timestamp 1607639953
transform 1 0 25282 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_251
timestamp 1607639953
transform 1 0 24178 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_257
timestamp 1607639953
transform 1 0 24730 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_245
timestamp 1607639953
transform 1 0 23626 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_347
timestamp 1607639953
transform 1 0 23534 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_284
timestamp 1607639953
transform 1 0 27214 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_276
timestamp 1607639953
transform 1 0 26478 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_281
timestamp 1607639953
transform 1 0 26938 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_269
timestamp 1607639953
transform 1 0 25834 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_358
timestamp 1607639953
transform 1 0 26386 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _100_
timestamp 1607639953
transform 1 0 27306 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_300
timestamp 1607639953
transform 1 0 28686 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_288
timestamp 1607639953
transform 1 0 27582 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_306
timestamp 1607639953
transform 1 0 29238 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_293
timestamp 1607639953
transform 1 0 28042 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_348
timestamp 1607639953
transform 1 0 29146 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_326
timestamp 1607639953
transform 1 0 31078 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_320
timestamp 1607639953
transform 1 0 30526 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_312
timestamp 1607639953
transform 1 0 29790 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_330
timestamp 1607639953
transform 1 0 31446 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_318
timestamp 1607639953
transform 1 0 30342 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _102_
timestamp 1607639953
transform 1 0 30802 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_349
timestamp 1607639953
transform 1 0 33194 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_337
timestamp 1607639953
transform 1 0 32090 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_334
timestamp 1607639953
transform 1 0 31814 0 -1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_350
timestamp 1607639953
transform 1 0 33286 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_338
timestamp 1607639953
transform 1 0 32182 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_334
timestamp 1607639953
transform 1 0 31814 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_359
timestamp 1607639953
transform 1 0 31998 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _141_
timestamp 1607639953
transform 1 0 31906 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_373
timestamp 1607639953
transform 1 0 35402 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_361
timestamp 1607639953
transform 1 0 34298 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_367
timestamp 1607639953
transform 1 0 34850 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_362
timestamp 1607639953
transform 1 0 34390 0 1 9248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_349
timestamp 1607639953
transform 1 0 34758 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_385
timestamp 1607639953
transform 1 0 36506 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_391
timestamp 1607639953
transform 1 0 37058 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_379
timestamp 1607639953
transform 1 0 35954 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_410
timestamp 1607639953
transform 1 0 38806 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_398
timestamp 1607639953
transform 1 0 37702 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_415
timestamp 1607639953
transform 1 0 39266 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_403
timestamp 1607639953
transform 1 0 38162 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_360
timestamp 1607639953
transform 1 0 37610 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_434
timestamp 1607639953
transform 1 0 41014 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_422
timestamp 1607639953
transform 1 0 39910 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_440
timestamp 1607639953
transform 1 0 41566 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_428
timestamp 1607639953
transform 1 0 40462 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_350
timestamp 1607639953
transform 1 0 40370 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_459
timestamp 1607639953
transform 1 0 43314 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_446
timestamp 1607639953
transform 1 0 42118 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_462
timestamp 1607639953
transform 1 0 43590 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_458
timestamp 1607639953
transform 1 0 43222 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_452
timestamp 1607639953
transform 1 0 42670 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_361
timestamp 1607639953
transform 1 0 43222 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _082_
timestamp 1607639953
transform 1 0 43314 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_483
timestamp 1607639953
transform 1 0 45522 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_471
timestamp 1607639953
transform 1 0 44418 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_474
timestamp 1607639953
transform 1 0 44694 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_495
timestamp 1607639953
transform 1 0 46626 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_505
timestamp 1607639953
transform 1 0 47546 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_501
timestamp 1607639953
transform 1 0 47178 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_489
timestamp 1607639953
transform 1 0 46074 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_486
timestamp 1607639953
transform 1 0 45798 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_351
timestamp 1607639953
transform 1 0 45982 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _206_
timestamp 1607639953
transform 1 0 47270 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_520
timestamp 1607639953
transform 1 0 48926 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_507
timestamp 1607639953
transform 1 0 47730 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_517
timestamp 1607639953
transform 1 0 48650 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_362
timestamp 1607639953
transform 1 0 48834 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_544
timestamp 1607639953
transform 1 0 51134 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_532
timestamp 1607639953
transform 1 0 50030 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_550
timestamp 1607639953
transform 1 0 51686 0 1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_13_541
timestamp 1607639953
transform 1 0 50858 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_529
timestamp 1607639953
transform 1 0 49754 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_352
timestamp 1607639953
transform 1 0 51594 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_568
timestamp 1607639953
transform 1 0 53342 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_556
timestamp 1607639953
transform 1 0 52238 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_571
timestamp 1607639953
transform 1 0 53618 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_559
timestamp 1607639953
transform 1 0 52514 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _159_
timestamp 1607639953
transform 1 0 52238 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_593
timestamp 1607639953
transform 1 0 55642 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_581
timestamp 1607639953
transform 1 0 54538 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_583
timestamp 1607639953
transform 1 0 54722 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_363
timestamp 1607639953
transform 1 0 54446 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_605
timestamp 1607639953
transform 1 0 56746 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_611
timestamp 1607639953
transform 1 0 57298 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_607
timestamp 1607639953
transform 1 0 56930 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_603
timestamp 1607639953
transform 1 0 56562 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_595
timestamp 1607639953
transform 1 0 55826 0 1 9248
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_353
timestamp 1607639953
transform 1 0 57206 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _020_
timestamp 1607639953
transform 1 0 56654 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_617
timestamp 1607639953
transform 1 0 57850 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_623
timestamp 1607639953
transform 1 0 58402 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1607639953
transform -1 0 58862 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1607639953
transform -1 0 58862 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1607639953
transform 1 0 2466 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1607639953
transform 1 0 1362 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1607639953
transform 1 0 1086 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1607639953
transform 1 0 4674 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1607639953
transform 1 0 3570 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_62
timestamp 1607639953
transform 1 0 6790 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_59
timestamp 1607639953
transform 1 0 6514 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_51
timestamp 1607639953
transform 1 0 5778 0 1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_364
timestamp 1607639953
transform 1 0 6698 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_74
timestamp 1607639953
transform 1 0 7894 0 1 10336
box -38 -48 222 592
use HAX1  HAX1
timestamp 1608117647
transform 1 0 8078 0 1 10336
box 0 -48 2024 592
use sky130_fd_sc_hd__decap_12  FILLER_15_110
timestamp 1607639953
transform 1 0 11206 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_98
timestamp 1607639953
transform 1 0 10102 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_123
timestamp 1607639953
transform 1 0 12402 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_365
timestamp 1607639953
transform 1 0 12310 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_147
timestamp 1607639953
transform 1 0 14610 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_135
timestamp 1607639953
transform 1 0 13506 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_171
timestamp 1607639953
transform 1 0 16818 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_159
timestamp 1607639953
transform 1 0 15714 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_196
timestamp 1607639953
transform 1 0 19118 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_184
timestamp 1607639953
transform 1 0 18014 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_366
timestamp 1607639953
transform 1 0 17922 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_220
timestamp 1607639953
transform 1 0 21326 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_208
timestamp 1607639953
transform 1 0 20222 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_232
timestamp 1607639953
transform 1 0 22430 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_257
timestamp 1607639953
transform 1 0 24730 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_245
timestamp 1607639953
transform 1 0 23626 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_367
timestamp 1607639953
transform 1 0 23534 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_281
timestamp 1607639953
transform 1 0 26938 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_269
timestamp 1607639953
transform 1 0 25834 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_306
timestamp 1607639953
transform 1 0 29238 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_293
timestamp 1607639953
transform 1 0 28042 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_368
timestamp 1607639953
transform 1 0 29146 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_330
timestamp 1607639953
transform 1 0 31446 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_318
timestamp 1607639953
transform 1 0 30342 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_342
timestamp 1607639953
transform 1 0 32550 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_367
timestamp 1607639953
transform 1 0 34850 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_354
timestamp 1607639953
transform 1 0 33654 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_369
timestamp 1607639953
transform 1 0 34758 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_391
timestamp 1607639953
transform 1 0 37058 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_379
timestamp 1607639953
transform 1 0 35954 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_415
timestamp 1607639953
transform 1 0 39266 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_403
timestamp 1607639953
transform 1 0 38162 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_440
timestamp 1607639953
transform 1 0 41566 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_428
timestamp 1607639953
transform 1 0 40462 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_370
timestamp 1607639953
transform 1 0 40370 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_459
timestamp 1607639953
transform 1 0 43314 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_447
timestamp 1607639953
transform 1 0 42210 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _171_
timestamp 1607639953
transform 1 0 41934 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_483
timestamp 1607639953
transform 1 0 45522 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_471
timestamp 1607639953
transform 1 0 44418 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_501
timestamp 1607639953
transform 1 0 47178 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_489
timestamp 1607639953
transform 1 0 46074 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_487
timestamp 1607639953
transform 1 0 45890 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_371
timestamp 1607639953
transform 1 0 45982 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_525
timestamp 1607639953
transform 1 0 49386 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_513
timestamp 1607639953
transform 1 0 48282 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_550
timestamp 1607639953
transform 1 0 51686 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_537
timestamp 1607639953
transform 1 0 50490 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_372
timestamp 1607639953
transform 1 0 51594 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_562
timestamp 1607639953
transform 1 0 52790 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_586
timestamp 1607639953
transform 1 0 54998 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_574
timestamp 1607639953
transform 1 0 53894 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_611
timestamp 1607639953
transform 1 0 57298 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_598
timestamp 1607639953
transform 1 0 56102 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_373
timestamp 1607639953
transform 1 0 57206 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_623
timestamp 1607639953
transform 1 0 58402 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1607639953
transform -1 0 58862 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1607639953
transform 1 0 2466 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1607639953
transform 1 0 1362 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1607639953
transform 1 0 1086 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_44
timestamp 1607639953
transform 1 0 5134 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_32
timestamp 1607639953
transform 1 0 4030 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_27
timestamp 1607639953
transform 1 0 3570 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_374
timestamp 1607639953
transform 1 0 3938 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_56
timestamp 1607639953
transform 1 0 6238 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_80
timestamp 1607639953
transform 1 0 8446 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_68
timestamp 1607639953
transform 1 0 7342 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_105
timestamp 1607639953
transform 1 0 10746 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_93
timestamp 1607639953
transform 1 0 9642 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_375
timestamp 1607639953
transform 1 0 9550 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_129
timestamp 1607639953
transform 1 0 12954 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_117
timestamp 1607639953
transform 1 0 11850 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_154
timestamp 1607639953
transform 1 0 15254 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_141
timestamp 1607639953
transform 1 0 14058 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_376
timestamp 1607639953
transform 1 0 15162 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_166
timestamp 1607639953
transform 1 0 16358 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_190
timestamp 1607639953
transform 1 0 18566 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_178
timestamp 1607639953
transform 1 0 17462 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_215
timestamp 1607639953
transform 1 0 20866 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_202
timestamp 1607639953
transform 1 0 19670 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_377
timestamp 1607639953
transform 1 0 20774 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_239
timestamp 1607639953
transform 1 0 23074 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_227
timestamp 1607639953
transform 1 0 21970 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_263
timestamp 1607639953
transform 1 0 25282 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_251
timestamp 1607639953
transform 1 0 24178 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_276
timestamp 1607639953
transform 1 0 26478 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_378
timestamp 1607639953
transform 1 0 26386 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_300
timestamp 1607639953
transform 1 0 28686 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_288
timestamp 1607639953
transform 1 0 27582 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_328
timestamp 1607639953
transform 1 0 31262 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_324
timestamp 1607639953
transform 1 0 30894 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_312
timestamp 1607639953
transform 1 0 29790 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _126_
timestamp 1607639953
transform 1 0 30986 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_349
timestamp 1607639953
transform 1 0 33194 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_337
timestamp 1607639953
transform 1 0 32090 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_379
timestamp 1607639953
transform 1 0 31998 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_373
timestamp 1607639953
transform 1 0 35402 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_361
timestamp 1607639953
transform 1 0 34298 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_385
timestamp 1607639953
transform 1 0 36506 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_410
timestamp 1607639953
transform 1 0 38806 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_398
timestamp 1607639953
transform 1 0 37702 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_380
timestamp 1607639953
transform 1 0 37610 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_434
timestamp 1607639953
transform 1 0 41014 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_422
timestamp 1607639953
transform 1 0 39910 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_459
timestamp 1607639953
transform 1 0 43314 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_446
timestamp 1607639953
transform 1 0 42118 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_381
timestamp 1607639953
transform 1 0 43222 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_483
timestamp 1607639953
transform 1 0 45522 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_471
timestamp 1607639953
transform 1 0 44418 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_495
timestamp 1607639953
transform 1 0 46626 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_520
timestamp 1607639953
transform 1 0 48926 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_507
timestamp 1607639953
transform 1 0 47730 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_382
timestamp 1607639953
transform 1 0 48834 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_544
timestamp 1607639953
transform 1 0 51134 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_532
timestamp 1607639953
transform 1 0 50030 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_568
timestamp 1607639953
transform 1 0 53342 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_556
timestamp 1607639953
transform 1 0 52238 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_593
timestamp 1607639953
transform 1 0 55642 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_581
timestamp 1607639953
transform 1 0 54538 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_383
timestamp 1607639953
transform 1 0 54446 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_605
timestamp 1607639953
transform 1 0 56746 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_617
timestamp 1607639953
transform 1 0 57850 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1607639953
transform -1 0 58862 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_15
timestamp 1607639953
transform 1 0 2466 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1607639953
transform 1 0 1362 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1607639953
transform 1 0 1086 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_39
timestamp 1607639953
transform 1 0 4674 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_27
timestamp 1607639953
transform 1 0 3570 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_62
timestamp 1607639953
transform 1 0 6790 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_59
timestamp 1607639953
transform 1 0 6514 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_17_51
timestamp 1607639953
transform 1 0 5778 0 1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_384
timestamp 1607639953
transform 1 0 6698 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_80
timestamp 1607639953
transform 1 0 8446 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_74
timestamp 1607639953
transform 1 0 7894 0 1 11424
box -38 -48 222 592
use INV  INV
timestamp 1608117647
transform 1 0 8078 0 1 11424
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_17_104
timestamp 1607639953
transform 1 0 10654 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_92
timestamp 1607639953
transform 1 0 9550 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_123
timestamp 1607639953
transform 1 0 12402 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_116
timestamp 1607639953
transform 1 0 11758 0 1 11424
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_385
timestamp 1607639953
transform 1 0 12310 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_147
timestamp 1607639953
transform 1 0 14610 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_135
timestamp 1607639953
transform 1 0 13506 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_171
timestamp 1607639953
transform 1 0 16818 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_159
timestamp 1607639953
transform 1 0 15714 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_196
timestamp 1607639953
transform 1 0 19118 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_184
timestamp 1607639953
transform 1 0 18014 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_386
timestamp 1607639953
transform 1 0 17922 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_220
timestamp 1607639953
transform 1 0 21326 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_208
timestamp 1607639953
transform 1 0 20222 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_232
timestamp 1607639953
transform 1 0 22430 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_257
timestamp 1607639953
transform 1 0 24730 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_245
timestamp 1607639953
transform 1 0 23626 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_387
timestamp 1607639953
transform 1 0 23534 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_281
timestamp 1607639953
transform 1 0 26938 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_269
timestamp 1607639953
transform 1 0 25834 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_306
timestamp 1607639953
transform 1 0 29238 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_293
timestamp 1607639953
transform 1 0 28042 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_388
timestamp 1607639953
transform 1 0 29146 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_330
timestamp 1607639953
transform 1 0 31446 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_318
timestamp 1607639953
transform 1 0 30342 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_342
timestamp 1607639953
transform 1 0 32550 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_367
timestamp 1607639953
transform 1 0 34850 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_354
timestamp 1607639953
transform 1 0 33654 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_389
timestamp 1607639953
transform 1 0 34758 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_391
timestamp 1607639953
transform 1 0 37058 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_379
timestamp 1607639953
transform 1 0 35954 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_415
timestamp 1607639953
transform 1 0 39266 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_403
timestamp 1607639953
transform 1 0 38162 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_440
timestamp 1607639953
transform 1 0 41566 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_428
timestamp 1607639953
transform 1 0 40462 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_390
timestamp 1607639953
transform 1 0 40370 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_452
timestamp 1607639953
transform 1 0 42670 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_476
timestamp 1607639953
transform 1 0 44878 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_464
timestamp 1607639953
transform 1 0 43774 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_501
timestamp 1607639953
transform 1 0 47178 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_489
timestamp 1607639953
transform 1 0 46074 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_391
timestamp 1607639953
transform 1 0 45982 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_525
timestamp 1607639953
transform 1 0 49386 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_513
timestamp 1607639953
transform 1 0 48282 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_550
timestamp 1607639953
transform 1 0 51686 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_537
timestamp 1607639953
transform 1 0 50490 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_392
timestamp 1607639953
transform 1 0 51594 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_562
timestamp 1607639953
transform 1 0 52790 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_586
timestamp 1607639953
transform 1 0 54998 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_574
timestamp 1607639953
transform 1 0 53894 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_611
timestamp 1607639953
transform 1 0 57298 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_598
timestamp 1607639953
transform 1 0 56102 0 1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_393
timestamp 1607639953
transform 1 0 57206 0 1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_623
timestamp 1607639953
transform 1 0 58402 0 1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1607639953
transform -1 0 58862 0 1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1607639953
transform 1 0 2466 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1607639953
transform 1 0 1362 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1607639953
transform 1 0 1086 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_44
timestamp 1607639953
transform 1 0 5134 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_32
timestamp 1607639953
transform 1 0 4030 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_27
timestamp 1607639953
transform 1 0 3570 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_394
timestamp 1607639953
transform 1 0 3938 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_56
timestamp 1607639953
transform 1 0 6238 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_80
timestamp 1607639953
transform 1 0 8446 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_68
timestamp 1607639953
transform 1 0 7342 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_105
timestamp 1607639953
transform 1 0 10746 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_93
timestamp 1607639953
transform 1 0 9642 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_395
timestamp 1607639953
transform 1 0 9550 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_129
timestamp 1607639953
transform 1 0 12954 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_117
timestamp 1607639953
transform 1 0 11850 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_154
timestamp 1607639953
transform 1 0 15254 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_141
timestamp 1607639953
transform 1 0 14058 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_396
timestamp 1607639953
transform 1 0 15162 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_166
timestamp 1607639953
transform 1 0 16358 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_190
timestamp 1607639953
transform 1 0 18566 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_178
timestamp 1607639953
transform 1 0 17462 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_215
timestamp 1607639953
transform 1 0 20866 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_202
timestamp 1607639953
transform 1 0 19670 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_397
timestamp 1607639953
transform 1 0 20774 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_239
timestamp 1607639953
transform 1 0 23074 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_227
timestamp 1607639953
transform 1 0 21970 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_263
timestamp 1607639953
transform 1 0 25282 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_251
timestamp 1607639953
transform 1 0 24178 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_276
timestamp 1607639953
transform 1 0 26478 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_398
timestamp 1607639953
transform 1 0 26386 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_300
timestamp 1607639953
transform 1 0 28686 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_288
timestamp 1607639953
transform 1 0 27582 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_324
timestamp 1607639953
transform 1 0 30894 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_312
timestamp 1607639953
transform 1 0 29790 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_349
timestamp 1607639953
transform 1 0 33194 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_337
timestamp 1607639953
transform 1 0 32090 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_399
timestamp 1607639953
transform 1 0 31998 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_373
timestamp 1607639953
transform 1 0 35402 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_361
timestamp 1607639953
transform 1 0 34298 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_385
timestamp 1607639953
transform 1 0 36506 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_413
timestamp 1607639953
transform 1 0 39082 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_401
timestamp 1607639953
transform 1 0 37978 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_400
timestamp 1607639953
transform 1 0 37610 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _186_
timestamp 1607639953
transform 1 0 37702 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_437
timestamp 1607639953
transform 1 0 41290 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_425
timestamp 1607639953
transform 1 0 40186 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_459
timestamp 1607639953
transform 1 0 43314 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_457
timestamp 1607639953
transform 1 0 43130 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_449
timestamp 1607639953
transform 1 0 42394 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_401
timestamp 1607639953
transform 1 0 43222 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_483
timestamp 1607639953
transform 1 0 45522 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_471
timestamp 1607639953
transform 1 0 44418 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_502
timestamp 1607639953
transform 1 0 47270 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_495
timestamp 1607639953
transform 1 0 46626 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _105_
timestamp 1607639953
transform 1 0 46994 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_18_520
timestamp 1607639953
transform 1 0 48926 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_518
timestamp 1607639953
transform 1 0 48742 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_514
timestamp 1607639953
transform 1 0 48374 0 -1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_402
timestamp 1607639953
transform 1 0 48834 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_544
timestamp 1607639953
transform 1 0 51134 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_532
timestamp 1607639953
transform 1 0 50030 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_568
timestamp 1607639953
transform 1 0 53342 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_556
timestamp 1607639953
transform 1 0 52238 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_593
timestamp 1607639953
transform 1 0 55642 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_581
timestamp 1607639953
transform 1 0 54538 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_403
timestamp 1607639953
transform 1 0 54446 0 -1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_605
timestamp 1607639953
transform 1 0 56746 0 -1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_617
timestamp 1607639953
transform 1 0 57850 0 -1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1607639953
transform -1 0 58862 0 -1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_15
timestamp 1607639953
transform 1 0 2466 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_3
timestamp 1607639953
transform 1 0 1362 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_15
timestamp 1607639953
transform 1 0 2466 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_3
timestamp 1607639953
transform 1 0 1362 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1607639953
transform 1 0 1086 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1607639953
transform 1 0 1086 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_44
timestamp 1607639953
transform 1 0 5134 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_32
timestamp 1607639953
transform 1 0 4030 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_27
timestamp 1607639953
transform 1 0 3570 0 -1 13600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_39
timestamp 1607639953
transform 1 0 4674 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_27
timestamp 1607639953
transform 1 0 3570 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_414
timestamp 1607639953
transform 1 0 3938 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_60
timestamp 1607639953
transform 1 0 6606 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_20_56
timestamp 1607639953
transform 1 0 6238 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_62
timestamp 1607639953
transform 1 0 6790 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_59
timestamp 1607639953
transform 1 0 6514 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_51
timestamp 1607639953
transform 1 0 5778 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_404
timestamp 1607639953
transform 1 0 6698 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _046_
timestamp 1607639953
transform 1 0 6330 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_84
timestamp 1607639953
transform 1 0 8814 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_20_72
timestamp 1607639953
transform 1 0 7710 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_80
timestamp 1607639953
transform 1 0 8446 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_74
timestamp 1607639953
transform 1 0 7894 0 1 12512
box -38 -48 222 592
use INVX1  INVX1
timestamp 1608117647
transform 1 0 8078 0 1 12512
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_20_105
timestamp 1607639953
transform 1 0 10746 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_93
timestamp 1607639953
transform 1 0 9642 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_108
timestamp 1607639953
transform 1 0 11022 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_96
timestamp 1607639953
transform 1 0 9918 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_92
timestamp 1607639953
transform 1 0 9550 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_415
timestamp 1607639953
transform 1 0 9550 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _070_
timestamp 1607639953
transform 1 0 9642 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_129
timestamp 1607639953
transform 1 0 12954 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_117
timestamp 1607639953
transform 1 0 11850 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_123
timestamp 1607639953
transform 1 0 12402 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_120
timestamp 1607639953
transform 1 0 12126 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_405
timestamp 1607639953
transform 1 0 12310 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_154
timestamp 1607639953
transform 1 0 15254 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_141
timestamp 1607639953
transform 1 0 14058 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_154
timestamp 1607639953
transform 1 0 15254 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_147
timestamp 1607639953
transform 1 0 14610 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_135
timestamp 1607639953
transform 1 0 13506 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_416
timestamp 1607639953
transform 1 0 15162 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _189_
timestamp 1607639953
transform 1 0 14978 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_166
timestamp 1607639953
transform 1 0 16358 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_166
timestamp 1607639953
transform 1 0 16358 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_190
timestamp 1607639953
transform 1 0 18566 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_178
timestamp 1607639953
transform 1 0 17462 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_196
timestamp 1607639953
transform 1 0 19118 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_184
timestamp 1607639953
transform 1 0 18014 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_182
timestamp 1607639953
transform 1 0 17830 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_178
timestamp 1607639953
transform 1 0 17462 0 1 12512
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_406
timestamp 1607639953
transform 1 0 17922 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_215
timestamp 1607639953
transform 1 0 20866 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_202
timestamp 1607639953
transform 1 0 19670 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_220
timestamp 1607639953
transform 1 0 21326 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_208
timestamp 1607639953
transform 1 0 20222 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_417
timestamp 1607639953
transform 1 0 20774 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_239
timestamp 1607639953
transform 1 0 23074 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_227
timestamp 1607639953
transform 1 0 21970 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_232
timestamp 1607639953
transform 1 0 22430 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_263
timestamp 1607639953
transform 1 0 25282 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_251
timestamp 1607639953
transform 1 0 24178 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_257
timestamp 1607639953
transform 1 0 24730 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_245
timestamp 1607639953
transform 1 0 23626 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_407
timestamp 1607639953
transform 1 0 23534 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_276
timestamp 1607639953
transform 1 0 26478 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_281
timestamp 1607639953
transform 1 0 26938 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_269
timestamp 1607639953
transform 1 0 25834 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_418
timestamp 1607639953
transform 1 0 26386 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_300
timestamp 1607639953
transform 1 0 28686 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_288
timestamp 1607639953
transform 1 0 27582 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_306
timestamp 1607639953
transform 1 0 29238 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_293
timestamp 1607639953
transform 1 0 28042 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_408
timestamp 1607639953
transform 1 0 29146 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_324
timestamp 1607639953
transform 1 0 30894 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_312
timestamp 1607639953
transform 1 0 29790 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_330
timestamp 1607639953
transform 1 0 31446 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_318
timestamp 1607639953
transform 1 0 30342 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_349
timestamp 1607639953
transform 1 0 33194 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_337
timestamp 1607639953
transform 1 0 32090 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_342
timestamp 1607639953
transform 1 0 32550 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_419
timestamp 1607639953
transform 1 0 31998 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_373
timestamp 1607639953
transform 1 0 35402 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_361
timestamp 1607639953
transform 1 0 34298 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_367
timestamp 1607639953
transform 1 0 34850 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_354
timestamp 1607639953
transform 1 0 33654 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_409
timestamp 1607639953
transform 1 0 34758 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_385
timestamp 1607639953
transform 1 0 36506 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_391
timestamp 1607639953
transform 1 0 37058 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_379
timestamp 1607639953
transform 1 0 35954 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_410
timestamp 1607639953
transform 1 0 38806 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_398
timestamp 1607639953
transform 1 0 37702 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_415
timestamp 1607639953
transform 1 0 39266 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_403
timestamp 1607639953
transform 1 0 38162 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_420
timestamp 1607639953
transform 1 0 37610 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_434
timestamp 1607639953
transform 1 0 41014 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_422
timestamp 1607639953
transform 1 0 39910 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_431
timestamp 1607639953
transform 1 0 40738 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_410
timestamp 1607639953
transform 1 0 40370 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _168_
timestamp 1607639953
transform 1 0 40462 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_459
timestamp 1607639953
transform 1 0 43314 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_446
timestamp 1607639953
transform 1 0 42118 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_455
timestamp 1607639953
transform 1 0 42946 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_443
timestamp 1607639953
transform 1 0 41842 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_421
timestamp 1607639953
transform 1 0 43222 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_483
timestamp 1607639953
transform 1 0 45522 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_471
timestamp 1607639953
transform 1 0 44418 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_479
timestamp 1607639953
transform 1 0 45154 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_19_467
timestamp 1607639953
transform 1 0 44050 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_495
timestamp 1607639953
transform 1 0 46626 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_504
timestamp 1607639953
transform 1 0 47454 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_492
timestamp 1607639953
transform 1 0 46350 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_487
timestamp 1607639953
transform 1 0 45890 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_411
timestamp 1607639953
transform 1 0 45982 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _001_
timestamp 1607639953
transform 1 0 46074 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_520
timestamp 1607639953
transform 1 0 48926 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_507
timestamp 1607639953
transform 1 0 47730 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_528
timestamp 1607639953
transform 1 0 49662 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_516
timestamp 1607639953
transform 1 0 48558 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_422
timestamp 1607639953
transform 1 0 48834 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_544
timestamp 1607639953
transform 1 0 51134 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_532
timestamp 1607639953
transform 1 0 50030 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_550
timestamp 1607639953
transform 1 0 51686 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_19_548
timestamp 1607639953
transform 1 0 51502 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_540
timestamp 1607639953
transform 1 0 50766 0 1 12512
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_412
timestamp 1607639953
transform 1 0 51594 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_568
timestamp 1607639953
transform 1 0 53342 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_556
timestamp 1607639953
transform 1 0 52238 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_562
timestamp 1607639953
transform 1 0 52790 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_593
timestamp 1607639953
transform 1 0 55642 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_581
timestamp 1607639953
transform 1 0 54538 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_586
timestamp 1607639953
transform 1 0 54998 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_574
timestamp 1607639953
transform 1 0 53894 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_423
timestamp 1607639953
transform 1 0 54446 0 -1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_605
timestamp 1607639953
transform 1 0 56746 0 -1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_611
timestamp 1607639953
transform 1 0 57298 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_598
timestamp 1607639953
transform 1 0 56102 0 1 12512
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_413
timestamp 1607639953
transform 1 0 57206 0 1 12512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_617
timestamp 1607639953
transform 1 0 57850 0 -1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_623
timestamp 1607639953
transform 1 0 58402 0 1 12512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1607639953
transform -1 0 58862 0 -1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1607639953
transform -1 0 58862 0 1 12512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_15
timestamp 1607639953
transform 1 0 2466 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1607639953
transform 1 0 1362 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1607639953
transform 1 0 1086 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_39
timestamp 1607639953
transform 1 0 4674 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_27
timestamp 1607639953
transform 1 0 3570 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_62
timestamp 1607639953
transform 1 0 6790 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_59
timestamp 1607639953
transform 1 0 6514 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_51
timestamp 1607639953
transform 1 0 5778 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_424
timestamp 1607639953
transform 1 0 6698 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_80
timestamp 1607639953
transform 1 0 8446 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_74
timestamp 1607639953
transform 1 0 7894 0 1 13600
box -38 -48 222 592
use INVX2  INVX2
timestamp 1608117647
transform 1 0 8078 0 1 13600
box 0 -48 368 592
use sky130_fd_sc_hd__decap_12  FILLER_21_104
timestamp 1607639953
transform 1 0 10654 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_92
timestamp 1607639953
transform 1 0 9550 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_126
timestamp 1607639953
transform 1 0 12678 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_116
timestamp 1607639953
transform 1 0 11758 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_425
timestamp 1607639953
transform 1 0 12310 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _081_
timestamp 1607639953
transform 1 0 12402 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_150
timestamp 1607639953
transform 1 0 14886 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_138
timestamp 1607639953
transform 1 0 13782 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_174
timestamp 1607639953
transform 1 0 17094 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_21_162
timestamp 1607639953
transform 1 0 15990 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_196
timestamp 1607639953
transform 1 0 19118 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_184
timestamp 1607639953
transform 1 0 18014 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_182
timestamp 1607639953
transform 1 0 17830 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_426
timestamp 1607639953
transform 1 0 17922 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_220
timestamp 1607639953
transform 1 0 21326 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_208
timestamp 1607639953
transform 1 0 20222 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_232
timestamp 1607639953
transform 1 0 22430 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_257
timestamp 1607639953
transform 1 0 24730 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_245
timestamp 1607639953
transform 1 0 23626 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_427
timestamp 1607639953
transform 1 0 23534 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_281
timestamp 1607639953
transform 1 0 26938 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_269
timestamp 1607639953
transform 1 0 25834 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_306
timestamp 1607639953
transform 1 0 29238 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_293
timestamp 1607639953
transform 1 0 28042 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_428
timestamp 1607639953
transform 1 0 29146 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_21_330
timestamp 1607639953
transform 1 0 31446 0 1 13600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_21_318
timestamp 1607639953
transform 1 0 30342 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_351
timestamp 1607639953
transform 1 0 33378 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_339
timestamp 1607639953
transform 1 0 32274 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _033_
timestamp 1607639953
transform 1 0 31998 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_367
timestamp 1607639953
transform 1 0 34850 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_363
timestamp 1607639953
transform 1 0 34482 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_429
timestamp 1607639953
transform 1 0 34758 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_391
timestamp 1607639953
transform 1 0 37058 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_379
timestamp 1607639953
transform 1 0 35954 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_415
timestamp 1607639953
transform 1 0 39266 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_403
timestamp 1607639953
transform 1 0 38162 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_440
timestamp 1607639953
transform 1 0 41566 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_428
timestamp 1607639953
transform 1 0 40462 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_430
timestamp 1607639953
transform 1 0 40370 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_452
timestamp 1607639953
transform 1 0 42670 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_476
timestamp 1607639953
transform 1 0 44878 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_464
timestamp 1607639953
transform 1 0 43774 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_504
timestamp 1607639953
transform 1 0 47454 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_492
timestamp 1607639953
transform 1 0 46350 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_431
timestamp 1607639953
transform 1 0 45982 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _205_
timestamp 1607639953
transform 1 0 46074 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_528
timestamp 1607639953
transform 1 0 49662 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_516
timestamp 1607639953
transform 1 0 48558 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_550
timestamp 1607639953
transform 1 0 51686 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_548
timestamp 1607639953
transform 1 0 51502 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_540
timestamp 1607639953
transform 1 0 50766 0 1 13600
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_432
timestamp 1607639953
transform 1 0 51594 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_562
timestamp 1607639953
transform 1 0 52790 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_586
timestamp 1607639953
transform 1 0 54998 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_574
timestamp 1607639953
transform 1 0 53894 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_611
timestamp 1607639953
transform 1 0 57298 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_598
timestamp 1607639953
transform 1 0 56102 0 1 13600
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_433
timestamp 1607639953
transform 1 0 57206 0 1 13600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_21_623
timestamp 1607639953
transform 1 0 58402 0 1 13600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1607639953
transform -1 0 58862 0 1 13600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_15
timestamp 1607639953
transform 1 0 2466 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_3
timestamp 1607639953
transform 1 0 1362 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1607639953
transform 1 0 1086 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_22_44
timestamp 1607639953
transform 1 0 5134 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_32
timestamp 1607639953
transform 1 0 4030 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_27
timestamp 1607639953
transform 1 0 3570 0 -1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_434
timestamp 1607639953
transform 1 0 3938 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_56
timestamp 1607639953
transform 1 0 6238 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_80
timestamp 1607639953
transform 1 0 8446 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_68
timestamp 1607639953
transform 1 0 7342 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_105
timestamp 1607639953
transform 1 0 10746 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_93
timestamp 1607639953
transform 1 0 9642 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_435
timestamp 1607639953
transform 1 0 9550 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_129
timestamp 1607639953
transform 1 0 12954 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_117
timestamp 1607639953
transform 1 0 11850 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_154
timestamp 1607639953
transform 1 0 15254 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_141
timestamp 1607639953
transform 1 0 14058 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_436
timestamp 1607639953
transform 1 0 15162 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_166
timestamp 1607639953
transform 1 0 16358 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_190
timestamp 1607639953
transform 1 0 18566 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_178
timestamp 1607639953
transform 1 0 17462 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_215
timestamp 1607639953
transform 1 0 20866 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_202
timestamp 1607639953
transform 1 0 19670 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_437
timestamp 1607639953
transform 1 0 20774 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_239
timestamp 1607639953
transform 1 0 23074 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_227
timestamp 1607639953
transform 1 0 21970 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_263
timestamp 1607639953
transform 1 0 25282 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_251
timestamp 1607639953
transform 1 0 24178 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_276
timestamp 1607639953
transform 1 0 26478 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_438
timestamp 1607639953
transform 1 0 26386 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_300
timestamp 1607639953
transform 1 0 28686 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_288
timestamp 1607639953
transform 1 0 27582 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_324
timestamp 1607639953
transform 1 0 30894 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_312
timestamp 1607639953
transform 1 0 29790 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_349
timestamp 1607639953
transform 1 0 33194 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_337
timestamp 1607639953
transform 1 0 32090 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_439
timestamp 1607639953
transform 1 0 31998 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_373
timestamp 1607639953
transform 1 0 35402 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_361
timestamp 1607639953
transform 1 0 34298 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_385
timestamp 1607639953
transform 1 0 36506 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_410
timestamp 1607639953
transform 1 0 38806 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_398
timestamp 1607639953
transform 1 0 37702 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_440
timestamp 1607639953
transform 1 0 37610 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_434
timestamp 1607639953
transform 1 0 41014 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_422
timestamp 1607639953
transform 1 0 39910 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_459
timestamp 1607639953
transform 1 0 43314 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_446
timestamp 1607639953
transform 1 0 42118 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_441
timestamp 1607639953
transform 1 0 43222 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_483
timestamp 1607639953
transform 1 0 45522 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_471
timestamp 1607639953
transform 1 0 44418 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_495
timestamp 1607639953
transform 1 0 46626 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_520
timestamp 1607639953
transform 1 0 48926 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_507
timestamp 1607639953
transform 1 0 47730 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_442
timestamp 1607639953
transform 1 0 48834 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_544
timestamp 1607639953
transform 1 0 51134 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_532
timestamp 1607639953
transform 1 0 50030 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_568
timestamp 1607639953
transform 1 0 53342 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_556
timestamp 1607639953
transform 1 0 52238 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_593
timestamp 1607639953
transform 1 0 55642 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_581
timestamp 1607639953
transform 1 0 54538 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_443
timestamp 1607639953
transform 1 0 54446 0 -1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_605
timestamp 1607639953
transform 1 0 56746 0 -1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_617
timestamp 1607639953
transform 1 0 57850 0 -1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1607639953
transform -1 0 58862 0 -1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1607639953
transform 1 0 2466 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1607639953
transform 1 0 1362 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1607639953
transform 1 0 1086 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_39
timestamp 1607639953
transform 1 0 4674 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1607639953
transform 1 0 3570 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_62
timestamp 1607639953
transform 1 0 6790 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_59
timestamp 1607639953
transform 1 0 6514 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_51
timestamp 1607639953
transform 1 0 5778 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_444
timestamp 1607639953
transform 1 0 6698 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_86
timestamp 1607639953
transform 1 0 8998 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_82
timestamp 1607639953
transform 1 0 8630 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_23_74
timestamp 1607639953
transform 1 0 7894 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _117_
timestamp 1607639953
transform 1 0 8722 0 1 14688
box -38 -48 314 592
use INVX4  INVX4
timestamp 1608117647
transform 1 0 8078 0 1 14688
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILLER_23_110
timestamp 1607639953
transform 1 0 11206 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_98
timestamp 1607639953
transform 1 0 10102 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_123
timestamp 1607639953
transform 1 0 12402 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_445
timestamp 1607639953
transform 1 0 12310 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_147
timestamp 1607639953
transform 1 0 14610 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_135
timestamp 1607639953
transform 1 0 13506 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_171
timestamp 1607639953
transform 1 0 16818 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_159
timestamp 1607639953
transform 1 0 15714 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_196
timestamp 1607639953
transform 1 0 19118 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_184
timestamp 1607639953
transform 1 0 18014 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_446
timestamp 1607639953
transform 1 0 17922 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_220
timestamp 1607639953
transform 1 0 21326 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_208
timestamp 1607639953
transform 1 0 20222 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_232
timestamp 1607639953
transform 1 0 22430 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_257
timestamp 1607639953
transform 1 0 24730 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_245
timestamp 1607639953
transform 1 0 23626 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_447
timestamp 1607639953
transform 1 0 23534 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_284
timestamp 1607639953
transform 1 0 27214 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_269
timestamp 1607639953
transform 1 0 25834 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _087_
timestamp 1607639953
transform 1 0 26938 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_23_306
timestamp 1607639953
transform 1 0 29238 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_304
timestamp 1607639953
transform 1 0 29054 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_296
timestamp 1607639953
transform 1 0 28318 0 1 14688
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_448
timestamp 1607639953
transform 1 0 29146 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_330
timestamp 1607639953
transform 1 0 31446 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_318
timestamp 1607639953
transform 1 0 30342 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_342
timestamp 1607639953
transform 1 0 32550 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_367
timestamp 1607639953
transform 1 0 34850 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_354
timestamp 1607639953
transform 1 0 33654 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_449
timestamp 1607639953
transform 1 0 34758 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_391
timestamp 1607639953
transform 1 0 37058 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_379
timestamp 1607639953
transform 1 0 35954 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_415
timestamp 1607639953
transform 1 0 39266 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_403
timestamp 1607639953
transform 1 0 38162 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_440
timestamp 1607639953
transform 1 0 41566 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_428
timestamp 1607639953
transform 1 0 40462 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_450
timestamp 1607639953
transform 1 0 40370 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_452
timestamp 1607639953
transform 1 0 42670 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_476
timestamp 1607639953
transform 1 0 44878 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_464
timestamp 1607639953
transform 1 0 43774 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_501
timestamp 1607639953
transform 1 0 47178 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_489
timestamp 1607639953
transform 1 0 46074 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_451
timestamp 1607639953
transform 1 0 45982 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_525
timestamp 1607639953
transform 1 0 49386 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_513
timestamp 1607639953
transform 1 0 48282 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_550
timestamp 1607639953
transform 1 0 51686 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_537
timestamp 1607639953
transform 1 0 50490 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_452
timestamp 1607639953
transform 1 0 51594 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_562
timestamp 1607639953
transform 1 0 52790 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_586
timestamp 1607639953
transform 1 0 54998 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_574
timestamp 1607639953
transform 1 0 53894 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_611
timestamp 1607639953
transform 1 0 57298 0 1 14688
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_609
timestamp 1607639953
transform 1 0 57114 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_605
timestamp 1607639953
transform 1 0 56746 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_598
timestamp 1607639953
transform 1 0 56102 0 1 14688
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_453
timestamp 1607639953
transform 1 0 57206 0 1 14688
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _094_
timestamp 1607639953
transform 1 0 56470 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_23_623
timestamp 1607639953
transform 1 0 58402 0 1 14688
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1607639953
transform -1 0 58862 0 1 14688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1607639953
transform 1 0 2466 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1607639953
transform 1 0 1362 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1607639953
transform 1 0 1086 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_35
timestamp 1607639953
transform 1 0 4306 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_27
timestamp 1607639953
transform 1 0 3570 0 -1 15776
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_454
timestamp 1607639953
transform 1 0 3938 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _152_
timestamp 1607639953
transform 1 0 4030 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_24_59
timestamp 1607639953
transform 1 0 6514 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_47
timestamp 1607639953
transform 1 0 5410 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_83
timestamp 1607639953
transform 1 0 8722 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_71
timestamp 1607639953
transform 1 0 7618 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_105
timestamp 1607639953
transform 1 0 10746 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_93
timestamp 1607639953
transform 1 0 9642 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_91
timestamp 1607639953
transform 1 0 9458 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_455
timestamp 1607639953
transform 1 0 9550 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_129
timestamp 1607639953
transform 1 0 12954 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_117
timestamp 1607639953
transform 1 0 11850 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_154
timestamp 1607639953
transform 1 0 15254 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_141
timestamp 1607639953
transform 1 0 14058 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_456
timestamp 1607639953
transform 1 0 15162 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_166
timestamp 1607639953
transform 1 0 16358 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_190
timestamp 1607639953
transform 1 0 18566 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_178
timestamp 1607639953
transform 1 0 17462 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_215
timestamp 1607639953
transform 1 0 20866 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_202
timestamp 1607639953
transform 1 0 19670 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_457
timestamp 1607639953
transform 1 0 20774 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_239
timestamp 1607639953
transform 1 0 23074 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_227
timestamp 1607639953
transform 1 0 21970 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_263
timestamp 1607639953
transform 1 0 25282 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_251
timestamp 1607639953
transform 1 0 24178 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_276
timestamp 1607639953
transform 1 0 26478 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_458
timestamp 1607639953
transform 1 0 26386 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_300
timestamp 1607639953
transform 1 0 28686 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_288
timestamp 1607639953
transform 1 0 27582 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_324
timestamp 1607639953
transform 1 0 30894 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_312
timestamp 1607639953
transform 1 0 29790 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_349
timestamp 1607639953
transform 1 0 33194 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_337
timestamp 1607639953
transform 1 0 32090 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_459
timestamp 1607639953
transform 1 0 31998 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_373
timestamp 1607639953
transform 1 0 35402 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_361
timestamp 1607639953
transform 1 0 34298 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_385
timestamp 1607639953
transform 1 0 36506 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_410
timestamp 1607639953
transform 1 0 38806 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_398
timestamp 1607639953
transform 1 0 37702 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_460
timestamp 1607639953
transform 1 0 37610 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_434
timestamp 1607639953
transform 1 0 41014 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_422
timestamp 1607639953
transform 1 0 39910 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_459
timestamp 1607639953
transform 1 0 43314 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_446
timestamp 1607639953
transform 1 0 42118 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_461
timestamp 1607639953
transform 1 0 43222 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_483
timestamp 1607639953
transform 1 0 45522 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_471
timestamp 1607639953
transform 1 0 44418 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_495
timestamp 1607639953
transform 1 0 46626 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_520
timestamp 1607639953
transform 1 0 48926 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_507
timestamp 1607639953
transform 1 0 47730 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_462
timestamp 1607639953
transform 1 0 48834 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_544
timestamp 1607639953
transform 1 0 51134 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_532
timestamp 1607639953
transform 1 0 50030 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_568
timestamp 1607639953
transform 1 0 53342 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_556
timestamp 1607639953
transform 1 0 52238 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_593
timestamp 1607639953
transform 1 0 55642 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_581
timestamp 1607639953
transform 1 0 54538 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_463
timestamp 1607639953
transform 1 0 54446 0 -1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_605
timestamp 1607639953
transform 1 0 56746 0 -1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_617
timestamp 1607639953
transform 1 0 57850 0 -1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1607639953
transform -1 0 58862 0 -1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1607639953
transform 1 0 2466 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1607639953
transform 1 0 1362 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1607639953
transform 1 0 1086 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_39
timestamp 1607639953
transform 1 0 4674 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1607639953
transform 1 0 3570 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_62
timestamp 1607639953
transform 1 0 6790 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_59
timestamp 1607639953
transform 1 0 6514 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_51
timestamp 1607639953
transform 1 0 5778 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_464
timestamp 1607639953
transform 1 0 6698 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_86
timestamp 1607639953
transform 1 0 8998 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_74
timestamp 1607639953
transform 1 0 7894 0 1 15776
box -38 -48 222 592
use INVX8  INVX8
timestamp 1608117647
transform 1 0 8078 0 1 15776
box 0 -48 920 592
use sky130_fd_sc_hd__decap_12  FILLER_25_110
timestamp 1607639953
transform 1 0 11206 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_98
timestamp 1607639953
transform 1 0 10102 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_123
timestamp 1607639953
transform 1 0 12402 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_465
timestamp 1607639953
transform 1 0 12310 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_147
timestamp 1607639953
transform 1 0 14610 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_135
timestamp 1607639953
transform 1 0 13506 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_170
timestamp 1607639953
transform 1 0 16726 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_159
timestamp 1607639953
transform 1 0 15714 0 1 15776
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _173_
timestamp 1607639953
transform 1 0 16450 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_25_196
timestamp 1607639953
transform 1 0 19118 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_184
timestamp 1607639953
transform 1 0 18014 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_182
timestamp 1607639953
transform 1 0 17830 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_466
timestamp 1607639953
transform 1 0 17922 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_220
timestamp 1607639953
transform 1 0 21326 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_208
timestamp 1607639953
transform 1 0 20222 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_232
timestamp 1607639953
transform 1 0 22430 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_257
timestamp 1607639953
transform 1 0 24730 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_245
timestamp 1607639953
transform 1 0 23626 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_467
timestamp 1607639953
transform 1 0 23534 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_281
timestamp 1607639953
transform 1 0 26938 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_269
timestamp 1607639953
transform 1 0 25834 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_306
timestamp 1607639953
transform 1 0 29238 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_293
timestamp 1607639953
transform 1 0 28042 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_468
timestamp 1607639953
transform 1 0 29146 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_330
timestamp 1607639953
transform 1 0 31446 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_318
timestamp 1607639953
transform 1 0 30342 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_342
timestamp 1607639953
transform 1 0 32550 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_367
timestamp 1607639953
transform 1 0 34850 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_354
timestamp 1607639953
transform 1 0 33654 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_469
timestamp 1607639953
transform 1 0 34758 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_391
timestamp 1607639953
transform 1 0 37058 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_379
timestamp 1607639953
transform 1 0 35954 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_415
timestamp 1607639953
transform 1 0 39266 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_403
timestamp 1607639953
transform 1 0 38162 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_440
timestamp 1607639953
transform 1 0 41566 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_428
timestamp 1607639953
transform 1 0 40462 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_470
timestamp 1607639953
transform 1 0 40370 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_452
timestamp 1607639953
transform 1 0 42670 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_476
timestamp 1607639953
transform 1 0 44878 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_464
timestamp 1607639953
transform 1 0 43774 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_501
timestamp 1607639953
transform 1 0 47178 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_489
timestamp 1607639953
transform 1 0 46074 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_471
timestamp 1607639953
transform 1 0 45982 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_525
timestamp 1607639953
transform 1 0 49386 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_513
timestamp 1607639953
transform 1 0 48282 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_550
timestamp 1607639953
transform 1 0 51686 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_537
timestamp 1607639953
transform 1 0 50490 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_472
timestamp 1607639953
transform 1 0 51594 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_562
timestamp 1607639953
transform 1 0 52790 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_586
timestamp 1607639953
transform 1 0 54998 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_574
timestamp 1607639953
transform 1 0 53894 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_611
timestamp 1607639953
transform 1 0 57298 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_598
timestamp 1607639953
transform 1 0 56102 0 1 15776
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_473
timestamp 1607639953
transform 1 0 57206 0 1 15776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_623
timestamp 1607639953
transform 1 0 58402 0 1 15776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1607639953
transform -1 0 58862 0 1 15776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_15
timestamp 1607639953
transform 1 0 2466 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_3
timestamp 1607639953
transform 1 0 1362 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_15
timestamp 1607639953
transform 1 0 2466 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_3
timestamp 1607639953
transform 1 0 1362 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1607639953
transform 1 0 1086 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1607639953
transform 1 0 1086 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_44
timestamp 1607639953
transform 1 0 5134 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_32
timestamp 1607639953
transform 1 0 4030 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_27
timestamp 1607639953
transform 1 0 3570 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_44
timestamp 1607639953
transform 1 0 5134 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_32
timestamp 1607639953
transform 1 0 4030 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_27
timestamp 1607639953
transform 1 0 3570 0 -1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_474
timestamp 1607639953
transform 1 0 3938 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _166_
timestamp 1607639953
transform 1 0 3754 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_62
timestamp 1607639953
transform 1 0 6790 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_60
timestamp 1607639953
transform 1 0 6606 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_56
timestamp 1607639953
transform 1 0 6238 0 1 16864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_56
timestamp 1607639953
transform 1 0 6238 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_484
timestamp 1607639953
transform 1 0 6698 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_74
timestamp 1607639953
transform 1 0 7894 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_80
timestamp 1607639953
transform 1 0 8446 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_68
timestamp 1607639953
transform 1 0 7342 0 -1 16864
box -38 -48 1142 592
use LATCH  LATCH
timestamp 1608117647
transform 1 0 8078 0 1 16864
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_12  FILLER_27_102
timestamp 1607639953
transform 1 0 10470 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_90
timestamp 1607639953
transform 1 0 9366 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_105
timestamp 1607639953
transform 1 0 10746 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_93
timestamp 1607639953
transform 1 0 9642 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_475
timestamp 1607639953
transform 1 0 9550 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_123
timestamp 1607639953
transform 1 0 12402 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_114
timestamp 1607639953
transform 1 0 11574 0 1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_26_129
timestamp 1607639953
transform 1 0 12954 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_117
timestamp 1607639953
transform 1 0 11850 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_485
timestamp 1607639953
transform 1 0 12310 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_147
timestamp 1607639953
transform 1 0 14610 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_135
timestamp 1607639953
transform 1 0 13506 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_154
timestamp 1607639953
transform 1 0 15254 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_141
timestamp 1607639953
transform 1 0 14058 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_476
timestamp 1607639953
transform 1 0 15162 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_171
timestamp 1607639953
transform 1 0 16818 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_159
timestamp 1607639953
transform 1 0 15714 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_166
timestamp 1607639953
transform 1 0 16358 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_196
timestamp 1607639953
transform 1 0 19118 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_184
timestamp 1607639953
transform 1 0 18014 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_190
timestamp 1607639953
transform 1 0 18566 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_178
timestamp 1607639953
transform 1 0 17462 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_486
timestamp 1607639953
transform 1 0 17922 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_220
timestamp 1607639953
transform 1 0 21326 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_208
timestamp 1607639953
transform 1 0 20222 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_215
timestamp 1607639953
transform 1 0 20866 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_202
timestamp 1607639953
transform 1 0 19670 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_477
timestamp 1607639953
transform 1 0 20774 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_232
timestamp 1607639953
transform 1 0 22430 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_239
timestamp 1607639953
transform 1 0 23074 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_227
timestamp 1607639953
transform 1 0 21970 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_257
timestamp 1607639953
transform 1 0 24730 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_245
timestamp 1607639953
transform 1 0 23626 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_263
timestamp 1607639953
transform 1 0 25282 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_251
timestamp 1607639953
transform 1 0 24178 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_487
timestamp 1607639953
transform 1 0 23534 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_281
timestamp 1607639953
transform 1 0 26938 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_269
timestamp 1607639953
transform 1 0 25834 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_276
timestamp 1607639953
transform 1 0 26478 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_478
timestamp 1607639953
transform 1 0 26386 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_306
timestamp 1607639953
transform 1 0 29238 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_293
timestamp 1607639953
transform 1 0 28042 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_300
timestamp 1607639953
transform 1 0 28686 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_288
timestamp 1607639953
transform 1 0 27582 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_488
timestamp 1607639953
transform 1 0 29146 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_330
timestamp 1607639953
transform 1 0 31446 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_318
timestamp 1607639953
transform 1 0 30342 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_324
timestamp 1607639953
transform 1 0 30894 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_312
timestamp 1607639953
transform 1 0 29790 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_342
timestamp 1607639953
transform 1 0 32550 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_349
timestamp 1607639953
transform 1 0 33194 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_337
timestamp 1607639953
transform 1 0 32090 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_479
timestamp 1607639953
transform 1 0 31998 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_367
timestamp 1607639953
transform 1 0 34850 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_354
timestamp 1607639953
transform 1 0 33654 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_373
timestamp 1607639953
transform 1 0 35402 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_361
timestamp 1607639953
transform 1 0 34298 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_489
timestamp 1607639953
transform 1 0 34758 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_391
timestamp 1607639953
transform 1 0 37058 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_379
timestamp 1607639953
transform 1 0 35954 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_385
timestamp 1607639953
transform 1 0 36506 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_415
timestamp 1607639953
transform 1 0 39266 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_403
timestamp 1607639953
transform 1 0 38162 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_410
timestamp 1607639953
transform 1 0 38806 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_398
timestamp 1607639953
transform 1 0 37702 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_480
timestamp 1607639953
transform 1 0 37610 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_440
timestamp 1607639953
transform 1 0 41566 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_428
timestamp 1607639953
transform 1 0 40462 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_434
timestamp 1607639953
transform 1 0 41014 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_422
timestamp 1607639953
transform 1 0 39910 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_490
timestamp 1607639953
transform 1 0 40370 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_452
timestamp 1607639953
transform 1 0 42670 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_459
timestamp 1607639953
transform 1 0 43314 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_446
timestamp 1607639953
transform 1 0 42118 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_481
timestamp 1607639953
transform 1 0 43222 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_476
timestamp 1607639953
transform 1 0 44878 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_464
timestamp 1607639953
transform 1 0 43774 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_483
timestamp 1607639953
transform 1 0 45522 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_471
timestamp 1607639953
transform 1 0 44418 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_501
timestamp 1607639953
transform 1 0 47178 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_489
timestamp 1607639953
transform 1 0 46074 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_495
timestamp 1607639953
transform 1 0 46626 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_491
timestamp 1607639953
transform 1 0 45982 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_525
timestamp 1607639953
transform 1 0 49386 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_513
timestamp 1607639953
transform 1 0 48282 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_520
timestamp 1607639953
transform 1 0 48926 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_507
timestamp 1607639953
transform 1 0 47730 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_482
timestamp 1607639953
transform 1 0 48834 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_550
timestamp 1607639953
transform 1 0 51686 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_537
timestamp 1607639953
transform 1 0 50490 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_544
timestamp 1607639953
transform 1 0 51134 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_532
timestamp 1607639953
transform 1 0 50030 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_492
timestamp 1607639953
transform 1 0 51594 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_562
timestamp 1607639953
transform 1 0 52790 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_568
timestamp 1607639953
transform 1 0 53342 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_556
timestamp 1607639953
transform 1 0 52238 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_586
timestamp 1607639953
transform 1 0 54998 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_574
timestamp 1607639953
transform 1 0 53894 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_593
timestamp 1607639953
transform 1 0 55642 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_581
timestamp 1607639953
transform 1 0 54538 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_483
timestamp 1607639953
transform 1 0 54446 0 -1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_611
timestamp 1607639953
transform 1 0 57298 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_598
timestamp 1607639953
transform 1 0 56102 0 1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_605
timestamp 1607639953
transform 1 0 56746 0 -1 16864
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_493
timestamp 1607639953
transform 1 0 57206 0 1 16864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_27_623
timestamp 1607639953
transform 1 0 58402 0 1 16864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_617
timestamp 1607639953
transform 1 0 57850 0 -1 16864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1607639953
transform -1 0 58862 0 1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1607639953
transform -1 0 58862 0 -1 16864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_15
timestamp 1607639953
transform 1 0 2466 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_3
timestamp 1607639953
transform 1 0 1362 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1607639953
transform 1 0 1086 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_44
timestamp 1607639953
transform 1 0 5134 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_32
timestamp 1607639953
transform 1 0 4030 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_27
timestamp 1607639953
transform 1 0 3570 0 -1 17952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_494
timestamp 1607639953
transform 1 0 3938 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_56
timestamp 1607639953
transform 1 0 6238 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_80
timestamp 1607639953
transform 1 0 8446 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_68
timestamp 1607639953
transform 1 0 7342 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_105
timestamp 1607639953
transform 1 0 10746 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_93
timestamp 1607639953
transform 1 0 9642 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_495
timestamp 1607639953
transform 1 0 9550 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_129
timestamp 1607639953
transform 1 0 12954 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_117
timestamp 1607639953
transform 1 0 11850 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_154
timestamp 1607639953
transform 1 0 15254 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_141
timestamp 1607639953
transform 1 0 14058 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_496
timestamp 1607639953
transform 1 0 15162 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_166
timestamp 1607639953
transform 1 0 16358 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_190
timestamp 1607639953
transform 1 0 18566 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_178
timestamp 1607639953
transform 1 0 17462 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_215
timestamp 1607639953
transform 1 0 20866 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_202
timestamp 1607639953
transform 1 0 19670 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_497
timestamp 1607639953
transform 1 0 20774 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_239
timestamp 1607639953
transform 1 0 23074 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_227
timestamp 1607639953
transform 1 0 21970 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_263
timestamp 1607639953
transform 1 0 25282 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_251
timestamp 1607639953
transform 1 0 24178 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_276
timestamp 1607639953
transform 1 0 26478 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_498
timestamp 1607639953
transform 1 0 26386 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_300
timestamp 1607639953
transform 1 0 28686 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_288
timestamp 1607639953
transform 1 0 27582 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_324
timestamp 1607639953
transform 1 0 30894 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_312
timestamp 1607639953
transform 1 0 29790 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_349
timestamp 1607639953
transform 1 0 33194 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_337
timestamp 1607639953
transform 1 0 32090 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_499
timestamp 1607639953
transform 1 0 31998 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_373
timestamp 1607639953
transform 1 0 35402 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_361
timestamp 1607639953
transform 1 0 34298 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_385
timestamp 1607639953
transform 1 0 36506 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_410
timestamp 1607639953
transform 1 0 38806 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_398
timestamp 1607639953
transform 1 0 37702 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_500
timestamp 1607639953
transform 1 0 37610 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_434
timestamp 1607639953
transform 1 0 41014 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_422
timestamp 1607639953
transform 1 0 39910 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_459
timestamp 1607639953
transform 1 0 43314 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_446
timestamp 1607639953
transform 1 0 42118 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_501
timestamp 1607639953
transform 1 0 43222 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_483
timestamp 1607639953
transform 1 0 45522 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_471
timestamp 1607639953
transform 1 0 44418 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_495
timestamp 1607639953
transform 1 0 46626 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_520
timestamp 1607639953
transform 1 0 48926 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_507
timestamp 1607639953
transform 1 0 47730 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_502
timestamp 1607639953
transform 1 0 48834 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_544
timestamp 1607639953
transform 1 0 51134 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_532
timestamp 1607639953
transform 1 0 50030 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_570
timestamp 1607639953
transform 1 0 53526 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_564
timestamp 1607639953
transform 1 0 52974 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_556
timestamp 1607639953
transform 1 0 52238 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _182_
timestamp 1607639953
transform 1 0 53250 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_593
timestamp 1607639953
transform 1 0 55642 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_581
timestamp 1607639953
transform 1 0 54538 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_578
timestamp 1607639953
transform 1 0 54262 0 -1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_503
timestamp 1607639953
transform 1 0 54446 0 -1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_605
timestamp 1607639953
transform 1 0 56746 0 -1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_617
timestamp 1607639953
transform 1 0 57850 0 -1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1607639953
transform -1 0 58862 0 -1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_15
timestamp 1607639953
transform 1 0 2466 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_3
timestamp 1607639953
transform 1 0 1362 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1607639953
transform 1 0 1086 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_39
timestamp 1607639953
transform 1 0 4674 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_27
timestamp 1607639953
transform 1 0 3570 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_62
timestamp 1607639953
transform 1 0 6790 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_59
timestamp 1607639953
transform 1 0 6514 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_51
timestamp 1607639953
transform 1 0 5778 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_504
timestamp 1607639953
transform 1 0 6698 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_88
timestamp 1607639953
transform 1 0 9182 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_74
timestamp 1607639953
transform 1 0 7894 0 1 17952
box -38 -48 222 592
use MUX2X1  MUX2X1
timestamp 1608117647
transform 1 0 8078 0 1 17952
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_29_100
timestamp 1607639953
transform 1 0 10286 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_123
timestamp 1607639953
transform 1 0 12402 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_120
timestamp 1607639953
transform 1 0 12126 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_29_112
timestamp 1607639953
transform 1 0 11390 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_505
timestamp 1607639953
transform 1 0 12310 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_147
timestamp 1607639953
transform 1 0 14610 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_135
timestamp 1607639953
transform 1 0 13506 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_171
timestamp 1607639953
transform 1 0 16818 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_159
timestamp 1607639953
transform 1 0 15714 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_196
timestamp 1607639953
transform 1 0 19118 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_184
timestamp 1607639953
transform 1 0 18014 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_506
timestamp 1607639953
transform 1 0 17922 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_220
timestamp 1607639953
transform 1 0 21326 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_208
timestamp 1607639953
transform 1 0 20222 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_232
timestamp 1607639953
transform 1 0 22430 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_257
timestamp 1607639953
transform 1 0 24730 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_245
timestamp 1607639953
transform 1 0 23626 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_507
timestamp 1607639953
transform 1 0 23534 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_281
timestamp 1607639953
transform 1 0 26938 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_269
timestamp 1607639953
transform 1 0 25834 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_306
timestamp 1607639953
transform 1 0 29238 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_293
timestamp 1607639953
transform 1 0 28042 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_508
timestamp 1607639953
transform 1 0 29146 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_330
timestamp 1607639953
transform 1 0 31446 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_318
timestamp 1607639953
transform 1 0 30342 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_341
timestamp 1607639953
transform 1 0 32458 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _017_
timestamp 1607639953
transform 1 0 32182 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_367
timestamp 1607639953
transform 1 0 34850 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_365
timestamp 1607639953
transform 1 0 34666 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_353
timestamp 1607639953
transform 1 0 33562 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_509
timestamp 1607639953
transform 1 0 34758 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_391
timestamp 1607639953
transform 1 0 37058 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_379
timestamp 1607639953
transform 1 0 35954 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_415
timestamp 1607639953
transform 1 0 39266 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_403
timestamp 1607639953
transform 1 0 38162 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_440
timestamp 1607639953
transform 1 0 41566 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_428
timestamp 1607639953
transform 1 0 40462 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_510
timestamp 1607639953
transform 1 0 40370 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_452
timestamp 1607639953
transform 1 0 42670 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_476
timestamp 1607639953
transform 1 0 44878 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_464
timestamp 1607639953
transform 1 0 43774 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_501
timestamp 1607639953
transform 1 0 47178 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_489
timestamp 1607639953
transform 1 0 46074 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_511
timestamp 1607639953
transform 1 0 45982 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_525
timestamp 1607639953
transform 1 0 49386 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_513
timestamp 1607639953
transform 1 0 48282 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_550
timestamp 1607639953
transform 1 0 51686 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_537
timestamp 1607639953
transform 1 0 50490 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_512
timestamp 1607639953
transform 1 0 51594 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_563
timestamp 1607639953
transform 1 0 52882 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_558
timestamp 1607639953
transform 1 0 52422 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _079_
timestamp 1607639953
transform 1 0 52606 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_587
timestamp 1607639953
transform 1 0 55090 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_575
timestamp 1607639953
transform 1 0 53986 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_611
timestamp 1607639953
transform 1 0 57298 0 1 17952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_607
timestamp 1607639953
transform 1 0 56930 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_599
timestamp 1607639953
transform 1 0 56194 0 1 17952
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_513
timestamp 1607639953
transform 1 0 57206 0 1 17952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_623
timestamp 1607639953
transform 1 0 58402 0 1 17952
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1607639953
transform -1 0 58862 0 1 17952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1607639953
transform 1 0 2466 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_3
timestamp 1607639953
transform 1 0 1362 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1607639953
transform 1 0 1086 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_44
timestamp 1607639953
transform 1 0 5134 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_32
timestamp 1607639953
transform 1 0 4030 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_27
timestamp 1607639953
transform 1 0 3570 0 -1 19040
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_514
timestamp 1607639953
transform 1 0 3938 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_56
timestamp 1607639953
transform 1 0 6238 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_80
timestamp 1607639953
transform 1 0 8446 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_68
timestamp 1607639953
transform 1 0 7342 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_105
timestamp 1607639953
transform 1 0 10746 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_93
timestamp 1607639953
transform 1 0 9642 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_515
timestamp 1607639953
transform 1 0 9550 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_129
timestamp 1607639953
transform 1 0 12954 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_117
timestamp 1607639953
transform 1 0 11850 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_154
timestamp 1607639953
transform 1 0 15254 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_141
timestamp 1607639953
transform 1 0 14058 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_516
timestamp 1607639953
transform 1 0 15162 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_166
timestamp 1607639953
transform 1 0 16358 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _108_
timestamp 1607639953
transform 1 0 17094 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_189
timestamp 1607639953
transform 1 0 18474 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_177
timestamp 1607639953
transform 1 0 17370 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_215
timestamp 1607639953
transform 1 0 20866 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_213
timestamp 1607639953
transform 1 0 20682 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_201
timestamp 1607639953
transform 1 0 19578 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_517
timestamp 1607639953
transform 1 0 20774 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_239
timestamp 1607639953
transform 1 0 23074 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_227
timestamp 1607639953
transform 1 0 21970 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_263
timestamp 1607639953
transform 1 0 25282 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_251
timestamp 1607639953
transform 1 0 24178 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_276
timestamp 1607639953
transform 1 0 26478 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_518
timestamp 1607639953
transform 1 0 26386 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_300
timestamp 1607639953
transform 1 0 28686 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_288
timestamp 1607639953
transform 1 0 27582 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_324
timestamp 1607639953
transform 1 0 30894 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_312
timestamp 1607639953
transform 1 0 29790 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_349
timestamp 1607639953
transform 1 0 33194 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_337
timestamp 1607639953
transform 1 0 32090 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_519
timestamp 1607639953
transform 1 0 31998 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_373
timestamp 1607639953
transform 1 0 35402 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_361
timestamp 1607639953
transform 1 0 34298 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_385
timestamp 1607639953
transform 1 0 36506 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_410
timestamp 1607639953
transform 1 0 38806 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_398
timestamp 1607639953
transform 1 0 37702 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_520
timestamp 1607639953
transform 1 0 37610 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_434
timestamp 1607639953
transform 1 0 41014 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_422
timestamp 1607639953
transform 1 0 39910 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_459
timestamp 1607639953
transform 1 0 43314 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_446
timestamp 1607639953
transform 1 0 42118 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_521
timestamp 1607639953
transform 1 0 43222 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_483
timestamp 1607639953
transform 1 0 45522 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_471
timestamp 1607639953
transform 1 0 44418 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_495
timestamp 1607639953
transform 1 0 46626 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_520
timestamp 1607639953
transform 1 0 48926 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_507
timestamp 1607639953
transform 1 0 47730 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_522
timestamp 1607639953
transform 1 0 48834 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_544
timestamp 1607639953
transform 1 0 51134 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_532
timestamp 1607639953
transform 1 0 50030 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_568
timestamp 1607639953
transform 1 0 53342 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_556
timestamp 1607639953
transform 1 0 52238 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_593
timestamp 1607639953
transform 1 0 55642 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_581
timestamp 1607639953
transform 1 0 54538 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_523
timestamp 1607639953
transform 1 0 54446 0 -1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_605
timestamp 1607639953
transform 1 0 56746 0 -1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_617
timestamp 1607639953
transform 1 0 57850 0 -1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1607639953
transform -1 0 58862 0 -1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1607639953
transform 1 0 2466 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1607639953
transform 1 0 1362 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1607639953
transform 1 0 1086 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_39
timestamp 1607639953
transform 1 0 4674 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_27
timestamp 1607639953
transform 1 0 3570 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_62
timestamp 1607639953
transform 1 0 6790 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_59
timestamp 1607639953
transform 1 0 6514 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_51
timestamp 1607639953
transform 1 0 5778 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_524
timestamp 1607639953
transform 1 0 6698 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_82
timestamp 1607639953
transform 1 0 8630 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_74
timestamp 1607639953
transform 1 0 7894 0 1 19040
box -38 -48 222 592
use NAND2X1  NAND2X1
timestamp 1608117647
transform 1 0 8078 0 1 19040
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILLER_31_108
timestamp 1607639953
transform 1 0 11022 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_96
timestamp 1607639953
transform 1 0 9918 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_90
timestamp 1607639953
transform 1 0 9366 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _024_
timestamp 1607639953
transform 1 0 9642 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_123
timestamp 1607639953
transform 1 0 12402 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_120
timestamp 1607639953
transform 1 0 12126 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_525
timestamp 1607639953
transform 1 0 12310 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _018_
timestamp 1607639953
transform 1 0 13138 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_146
timestamp 1607639953
transform 1 0 14518 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_134
timestamp 1607639953
transform 1 0 13414 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_170
timestamp 1607639953
transform 1 0 16726 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_158
timestamp 1607639953
transform 1 0 15622 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_196
timestamp 1607639953
transform 1 0 19118 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_184
timestamp 1607639953
transform 1 0 18014 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_182
timestamp 1607639953
transform 1 0 17830 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_526
timestamp 1607639953
transform 1 0 17922 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_220
timestamp 1607639953
transform 1 0 21326 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_208
timestamp 1607639953
transform 1 0 20222 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_232
timestamp 1607639953
transform 1 0 22430 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_257
timestamp 1607639953
transform 1 0 24730 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_245
timestamp 1607639953
transform 1 0 23626 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_527
timestamp 1607639953
transform 1 0 23534 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_281
timestamp 1607639953
transform 1 0 26938 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_269
timestamp 1607639953
transform 1 0 25834 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_293
timestamp 1607639953
transform 1 0 28042 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_528
timestamp 1607639953
transform 1 0 29146 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _122_
timestamp 1607639953
transform 1 0 29238 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_321
timestamp 1607639953
transform 1 0 30618 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_309
timestamp 1607639953
transform 1 0 29514 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_345
timestamp 1607639953
transform 1 0 32826 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_333
timestamp 1607639953
transform 1 0 31722 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_367
timestamp 1607639953
transform 1 0 34850 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_365
timestamp 1607639953
transform 1 0 34666 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_357
timestamp 1607639953
transform 1 0 33930 0 1 19040
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_529
timestamp 1607639953
transform 1 0 34758 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_391
timestamp 1607639953
transform 1 0 37058 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_379
timestamp 1607639953
transform 1 0 35954 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_415
timestamp 1607639953
transform 1 0 39266 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_403
timestamp 1607639953
transform 1 0 38162 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_440
timestamp 1607639953
transform 1 0 41566 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_428
timestamp 1607639953
transform 1 0 40462 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_530
timestamp 1607639953
transform 1 0 40370 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_452
timestamp 1607639953
transform 1 0 42670 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_476
timestamp 1607639953
transform 1 0 44878 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_464
timestamp 1607639953
transform 1 0 43774 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_501
timestamp 1607639953
transform 1 0 47178 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_489
timestamp 1607639953
transform 1 0 46074 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_531
timestamp 1607639953
transform 1 0 45982 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_525
timestamp 1607639953
transform 1 0 49386 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_513
timestamp 1607639953
transform 1 0 48282 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_550
timestamp 1607639953
transform 1 0 51686 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_537
timestamp 1607639953
transform 1 0 50490 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_532
timestamp 1607639953
transform 1 0 51594 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_562
timestamp 1607639953
transform 1 0 52790 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_586
timestamp 1607639953
transform 1 0 54998 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_574
timestamp 1607639953
transform 1 0 53894 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_611
timestamp 1607639953
transform 1 0 57298 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_598
timestamp 1607639953
transform 1 0 56102 0 1 19040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_533
timestamp 1607639953
transform 1 0 57206 0 1 19040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_31_623
timestamp 1607639953
transform 1 0 58402 0 1 19040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1607639953
transform -1 0 58862 0 1 19040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_15
timestamp 1607639953
transform 1 0 2466 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1607639953
transform 1 0 1362 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1607639953
transform 1 0 1086 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_44
timestamp 1607639953
transform 1 0 5134 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_32
timestamp 1607639953
transform 1 0 4030 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_27
timestamp 1607639953
transform 1 0 3570 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_534
timestamp 1607639953
transform 1 0 3938 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_56
timestamp 1607639953
transform 1 0 6238 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_80
timestamp 1607639953
transform 1 0 8446 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_68
timestamp 1607639953
transform 1 0 7342 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_105
timestamp 1607639953
transform 1 0 10746 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_93
timestamp 1607639953
transform 1 0 9642 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_535
timestamp 1607639953
transform 1 0 9550 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_129
timestamp 1607639953
transform 1 0 12954 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_117
timestamp 1607639953
transform 1 0 11850 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_154
timestamp 1607639953
transform 1 0 15254 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_141
timestamp 1607639953
transform 1 0 14058 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_536
timestamp 1607639953
transform 1 0 15162 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_166
timestamp 1607639953
transform 1 0 16358 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_190
timestamp 1607639953
transform 1 0 18566 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_178
timestamp 1607639953
transform 1 0 17462 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_215
timestamp 1607639953
transform 1 0 20866 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_202
timestamp 1607639953
transform 1 0 19670 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_537
timestamp 1607639953
transform 1 0 20774 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_239
timestamp 1607639953
transform 1 0 23074 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_227
timestamp 1607639953
transform 1 0 21970 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_263
timestamp 1607639953
transform 1 0 25282 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_251
timestamp 1607639953
transform 1 0 24178 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_276
timestamp 1607639953
transform 1 0 26478 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_538
timestamp 1607639953
transform 1 0 26386 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_300
timestamp 1607639953
transform 1 0 28686 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_288
timestamp 1607639953
transform 1 0 27582 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_324
timestamp 1607639953
transform 1 0 30894 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_312
timestamp 1607639953
transform 1 0 29790 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_349
timestamp 1607639953
transform 1 0 33194 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_337
timestamp 1607639953
transform 1 0 32090 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_539
timestamp 1607639953
transform 1 0 31998 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_373
timestamp 1607639953
transform 1 0 35402 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_361
timestamp 1607639953
transform 1 0 34298 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_385
timestamp 1607639953
transform 1 0 36506 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_410
timestamp 1607639953
transform 1 0 38806 0 -1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_398
timestamp 1607639953
transform 1 0 37702 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_540
timestamp 1607639953
transform 1 0 37610 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _009_
timestamp 1607639953
transform 1 0 39542 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_433
timestamp 1607639953
transform 1 0 40922 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_421
timestamp 1607639953
transform 1 0 39818 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_459
timestamp 1607639953
transform 1 0 43314 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_457
timestamp 1607639953
transform 1 0 43130 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_445
timestamp 1607639953
transform 1 0 42026 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_541
timestamp 1607639953
transform 1 0 43222 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_483
timestamp 1607639953
transform 1 0 45522 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_471
timestamp 1607639953
transform 1 0 44418 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_495
timestamp 1607639953
transform 1 0 46626 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_528
timestamp 1607639953
transform 1 0 49662 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_524
timestamp 1607639953
transform 1 0 49294 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_520
timestamp 1607639953
transform 1 0 48926 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_507
timestamp 1607639953
transform 1 0 47730 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_542
timestamp 1607639953
transform 1 0 48834 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _055_
timestamp 1607639953
transform 1 0 49386 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_540
timestamp 1607639953
transform 1 0 50766 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_564
timestamp 1607639953
transform 1 0 52974 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_552
timestamp 1607639953
transform 1 0 51870 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_593
timestamp 1607639953
transform 1 0 55642 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_581
timestamp 1607639953
transform 1 0 54538 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_576
timestamp 1607639953
transform 1 0 54078 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_543
timestamp 1607639953
transform 1 0 54446 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_605
timestamp 1607639953
transform 1 0 56746 0 -1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_621
timestamp 1607639953
transform 1 0 58218 0 -1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_617
timestamp 1607639953
transform 1 0 57850 0 -1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1607639953
transform -1 0 58862 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _063_
timestamp 1607639953
transform 1 0 57942 0 -1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1607639953
transform 1 0 2466 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1607639953
transform 1 0 1362 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1607639953
transform 1 0 2466 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1607639953
transform 1 0 1362 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1607639953
transform 1 0 1086 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1607639953
transform 1 0 1086 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_44
timestamp 1607639953
transform 1 0 5134 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_32
timestamp 1607639953
transform 1 0 4030 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_27
timestamp 1607639953
transform 1 0 3570 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_33
timestamp 1607639953
transform 1 0 4122 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_27
timestamp 1607639953
transform 1 0 3570 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_554
timestamp 1607639953
transform 1 0 3938 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _051_
timestamp 1607639953
transform 1 0 3846 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_56
timestamp 1607639953
transform 1 0 6238 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_62
timestamp 1607639953
transform 1 0 6790 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_57
timestamp 1607639953
transform 1 0 6330 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_45
timestamp 1607639953
transform 1 0 5226 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_544
timestamp 1607639953
transform 1 0 6698 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_80
timestamp 1607639953
transform 1 0 8446 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_68
timestamp 1607639953
transform 1 0 7342 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_84
timestamp 1607639953
transform 1 0 8814 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_74
timestamp 1607639953
transform 1 0 7894 0 1 20128
box -38 -48 222 592
use NAND3X1  NAND3X1
timestamp 1608117647
transform 1 0 8078 0 1 20128
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILLER_34_105
timestamp 1607639953
transform 1 0 10746 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_93
timestamp 1607639953
transform 1 0 9642 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_108
timestamp 1607639953
transform 1 0 11022 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_96
timestamp 1607639953
transform 1 0 9918 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_555
timestamp 1607639953
transform 1 0 9550 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_129
timestamp 1607639953
transform 1 0 12954 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_117
timestamp 1607639953
transform 1 0 11850 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_123
timestamp 1607639953
transform 1 0 12402 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_120
timestamp 1607639953
transform 1 0 12126 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_545
timestamp 1607639953
transform 1 0 12310 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_154
timestamp 1607639953
transform 1 0 15254 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_141
timestamp 1607639953
transform 1 0 14058 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_147
timestamp 1607639953
transform 1 0 14610 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_135
timestamp 1607639953
transform 1 0 13506 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_556
timestamp 1607639953
transform 1 0 15162 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_166
timestamp 1607639953
transform 1 0 16358 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_171
timestamp 1607639953
transform 1 0 16818 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_159
timestamp 1607639953
transform 1 0 15714 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_190
timestamp 1607639953
transform 1 0 18566 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_178
timestamp 1607639953
transform 1 0 17462 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_190
timestamp 1607639953
transform 1 0 18566 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_184
timestamp 1607639953
transform 1 0 18014 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_546
timestamp 1607639953
transform 1 0 17922 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _172_
timestamp 1607639953
transform 1 0 18290 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_215
timestamp 1607639953
transform 1 0 20866 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_202
timestamp 1607639953
transform 1 0 19670 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_214
timestamp 1607639953
transform 1 0 20774 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_202
timestamp 1607639953
transform 1 0 19670 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_557
timestamp 1607639953
transform 1 0 20774 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_239
timestamp 1607639953
transform 1 0 23074 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_227
timestamp 1607639953
transform 1 0 21970 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_238
timestamp 1607639953
transform 1 0 22982 0 1 20128
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_33_226
timestamp 1607639953
transform 1 0 21878 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_254
timestamp 1607639953
transform 1 0 24454 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_257
timestamp 1607639953
transform 1 0 24730 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_245
timestamp 1607639953
transform 1 0 23626 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_547
timestamp 1607639953
transform 1 0 23534 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _032_
timestamp 1607639953
transform 1 0 24178 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_276
timestamp 1607639953
transform 1 0 26478 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_274
timestamp 1607639953
transform 1 0 26294 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_266
timestamp 1607639953
transform 1 0 25558 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_281
timestamp 1607639953
transform 1 0 26938 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_269
timestamp 1607639953
transform 1 0 25834 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_558
timestamp 1607639953
transform 1 0 26386 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_300
timestamp 1607639953
transform 1 0 28686 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_288
timestamp 1607639953
transform 1 0 27582 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_306
timestamp 1607639953
transform 1 0 29238 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_304
timestamp 1607639953
transform 1 0 29054 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_300
timestamp 1607639953
transform 1 0 28686 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_293
timestamp 1607639953
transform 1 0 28042 0 1 20128
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_548
timestamp 1607639953
transform 1 0 29146 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _185_
timestamp 1607639953
transform 1 0 28410 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_34_328
timestamp 1607639953
transform 1 0 31262 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_324
timestamp 1607639953
transform 1 0 30894 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_312
timestamp 1607639953
transform 1 0 29790 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_330
timestamp 1607639953
transform 1 0 31446 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_318
timestamp 1607639953
transform 1 0 30342 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _151_
timestamp 1607639953
transform 1 0 31354 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_349
timestamp 1607639953
transform 1 0 33194 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_337
timestamp 1607639953
transform 1 0 32090 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_332
timestamp 1607639953
transform 1 0 31630 0 -1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_342
timestamp 1607639953
transform 1 0 32550 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_559
timestamp 1607639953
transform 1 0 31998 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_373
timestamp 1607639953
transform 1 0 35402 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_361
timestamp 1607639953
transform 1 0 34298 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_367
timestamp 1607639953
transform 1 0 34850 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_354
timestamp 1607639953
transform 1 0 33654 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_549
timestamp 1607639953
transform 1 0 34758 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_385
timestamp 1607639953
transform 1 0 36506 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_391
timestamp 1607639953
transform 1 0 37058 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_379
timestamp 1607639953
transform 1 0 35954 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_410
timestamp 1607639953
transform 1 0 38806 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_398
timestamp 1607639953
transform 1 0 37702 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_415
timestamp 1607639953
transform 1 0 39266 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_403
timestamp 1607639953
transform 1 0 38162 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_560
timestamp 1607639953
transform 1 0 37610 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_434
timestamp 1607639953
transform 1 0 41014 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_422
timestamp 1607639953
transform 1 0 39910 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_440
timestamp 1607639953
transform 1 0 41566 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_428
timestamp 1607639953
transform 1 0 40462 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_550
timestamp 1607639953
transform 1 0 40370 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_459
timestamp 1607639953
transform 1 0 43314 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_446
timestamp 1607639953
transform 1 0 42118 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_452
timestamp 1607639953
transform 1 0 42670 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_561
timestamp 1607639953
transform 1 0 43222 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_483
timestamp 1607639953
transform 1 0 45522 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_471
timestamp 1607639953
transform 1 0 44418 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_476
timestamp 1607639953
transform 1 0 44878 0 1 20128
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_464
timestamp 1607639953
transform 1 0 43774 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _114_
timestamp 1607639953
transform 1 0 45614 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_495
timestamp 1607639953
transform 1 0 46626 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_501
timestamp 1607639953
transform 1 0 47178 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_489
timestamp 1607639953
transform 1 0 46074 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_33_487
timestamp 1607639953
transform 1 0 45890 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_551
timestamp 1607639953
transform 1 0 45982 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_520
timestamp 1607639953
transform 1 0 48926 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_507
timestamp 1607639953
transform 1 0 47730 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_525
timestamp 1607639953
transform 1 0 49386 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_513
timestamp 1607639953
transform 1 0 48282 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_562
timestamp 1607639953
transform 1 0 48834 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_544
timestamp 1607639953
transform 1 0 51134 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_532
timestamp 1607639953
transform 1 0 50030 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_550
timestamp 1607639953
transform 1 0 51686 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_537
timestamp 1607639953
transform 1 0 50490 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_552
timestamp 1607639953
transform 1 0 51594 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_567
timestamp 1607639953
transform 1 0 53250 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_555
timestamp 1607639953
transform 1 0 52146 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_562
timestamp 1607639953
transform 1 0 52790 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _190_
timestamp 1607639953
transform 1 0 51870 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_593
timestamp 1607639953
transform 1 0 55642 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_581
timestamp 1607639953
transform 1 0 54538 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_579
timestamp 1607639953
transform 1 0 54354 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_586
timestamp 1607639953
transform 1 0 54998 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_574
timestamp 1607639953
transform 1 0 53894 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_563
timestamp 1607639953
transform 1 0 54446 0 -1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_605
timestamp 1607639953
transform 1 0 56746 0 -1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_611
timestamp 1607639953
transform 1 0 57298 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_598
timestamp 1607639953
transform 1 0 56102 0 1 20128
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_553
timestamp 1607639953
transform 1 0 57206 0 1 20128
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_617
timestamp 1607639953
transform 1 0 57850 0 -1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_623
timestamp 1607639953
transform 1 0 58402 0 1 20128
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1607639953
transform -1 0 58862 0 -1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1607639953
transform -1 0 58862 0 1 20128
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1607639953
transform 1 0 2466 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1607639953
transform 1 0 1362 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1607639953
transform 1 0 1086 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_39
timestamp 1607639953
transform 1 0 4674 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_27
timestamp 1607639953
transform 1 0 3570 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_62
timestamp 1607639953
transform 1 0 6790 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_59
timestamp 1607639953
transform 1 0 6514 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_51
timestamp 1607639953
transform 1 0 5778 0 1 21216
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_564
timestamp 1607639953
transform 1 0 6698 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_82
timestamp 1607639953
transform 1 0 8630 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_74
timestamp 1607639953
transform 1 0 7894 0 1 21216
box -38 -48 222 592
use NOR2X1  NOR2X1
timestamp 1608117647
transform 1 0 8078 0 1 21216
box 0 -48 552 592
use sky130_fd_sc_hd__decap_12  FILLER_35_106
timestamp 1607639953
transform 1 0 10838 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_94
timestamp 1607639953
transform 1 0 9734 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_123
timestamp 1607639953
transform 1 0 12402 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_118
timestamp 1607639953
transform 1 0 11942 0 1 21216
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_565
timestamp 1607639953
transform 1 0 12310 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_147
timestamp 1607639953
transform 1 0 14610 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_135
timestamp 1607639953
transform 1 0 13506 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_171
timestamp 1607639953
transform 1 0 16818 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_159
timestamp 1607639953
transform 1 0 15714 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_196
timestamp 1607639953
transform 1 0 19118 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_184
timestamp 1607639953
transform 1 0 18014 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_566
timestamp 1607639953
transform 1 0 17922 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_220
timestamp 1607639953
transform 1 0 21326 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_208
timestamp 1607639953
transform 1 0 20222 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_232
timestamp 1607639953
transform 1 0 22430 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_257
timestamp 1607639953
transform 1 0 24730 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_245
timestamp 1607639953
transform 1 0 23626 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_567
timestamp 1607639953
transform 1 0 23534 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_281
timestamp 1607639953
transform 1 0 26938 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_269
timestamp 1607639953
transform 1 0 25834 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_306
timestamp 1607639953
transform 1 0 29238 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_293
timestamp 1607639953
transform 1 0 28042 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_568
timestamp 1607639953
transform 1 0 29146 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_330
timestamp 1607639953
transform 1 0 31446 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_318
timestamp 1607639953
transform 1 0 30342 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_342
timestamp 1607639953
transform 1 0 32550 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_367
timestamp 1607639953
transform 1 0 34850 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_354
timestamp 1607639953
transform 1 0 33654 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_569
timestamp 1607639953
transform 1 0 34758 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_391
timestamp 1607639953
transform 1 0 37058 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_379
timestamp 1607639953
transform 1 0 35954 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_415
timestamp 1607639953
transform 1 0 39266 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_403
timestamp 1607639953
transform 1 0 38162 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_440
timestamp 1607639953
transform 1 0 41566 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_428
timestamp 1607639953
transform 1 0 40462 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_570
timestamp 1607639953
transform 1 0 40370 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_452
timestamp 1607639953
transform 1 0 42670 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_476
timestamp 1607639953
transform 1 0 44878 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_464
timestamp 1607639953
transform 1 0 43774 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_501
timestamp 1607639953
transform 1 0 47178 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_489
timestamp 1607639953
transform 1 0 46074 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_571
timestamp 1607639953
transform 1 0 45982 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_525
timestamp 1607639953
transform 1 0 49386 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_513
timestamp 1607639953
transform 1 0 48282 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_550
timestamp 1607639953
transform 1 0 51686 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_537
timestamp 1607639953
transform 1 0 50490 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_572
timestamp 1607639953
transform 1 0 51594 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_562
timestamp 1607639953
transform 1 0 52790 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_586
timestamp 1607639953
transform 1 0 54998 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_574
timestamp 1607639953
transform 1 0 53894 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_611
timestamp 1607639953
transform 1 0 57298 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_598
timestamp 1607639953
transform 1 0 56102 0 1 21216
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_573
timestamp 1607639953
transform 1 0 57206 0 1 21216
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_35_623
timestamp 1607639953
transform 1 0 58402 0 1 21216
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1607639953
transform -1 0 58862 0 1 21216
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1607639953
transform 1 0 2466 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1607639953
transform 1 0 1362 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1607639953
transform 1 0 1086 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_44
timestamp 1607639953
transform 1 0 5134 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_32
timestamp 1607639953
transform 1 0 4030 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_27
timestamp 1607639953
transform 1 0 3570 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_574
timestamp 1607639953
transform 1 0 3938 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_56
timestamp 1607639953
transform 1 0 6238 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_80
timestamp 1607639953
transform 1 0 8446 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_68
timestamp 1607639953
transform 1 0 7342 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_105
timestamp 1607639953
transform 1 0 10746 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_93
timestamp 1607639953
transform 1 0 9642 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_575
timestamp 1607639953
transform 1 0 9550 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_129
timestamp 1607639953
transform 1 0 12954 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_117
timestamp 1607639953
transform 1 0 11850 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_154
timestamp 1607639953
transform 1 0 15254 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_141
timestamp 1607639953
transform 1 0 14058 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_576
timestamp 1607639953
transform 1 0 15162 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_166
timestamp 1607639953
transform 1 0 16358 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_190
timestamp 1607639953
transform 1 0 18566 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_178
timestamp 1607639953
transform 1 0 17462 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_215
timestamp 1607639953
transform 1 0 20866 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_202
timestamp 1607639953
transform 1 0 19670 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_577
timestamp 1607639953
transform 1 0 20774 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_234
timestamp 1607639953
transform 1 0 22614 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_227
timestamp 1607639953
transform 1 0 21970 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _193_
timestamp 1607639953
transform 1 0 22338 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_258
timestamp 1607639953
transform 1 0 24822 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_246
timestamp 1607639953
transform 1 0 23718 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_276
timestamp 1607639953
transform 1 0 26478 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_274
timestamp 1607639953
transform 1 0 26294 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_270
timestamp 1607639953
transform 1 0 25926 0 -1 22304
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_578
timestamp 1607639953
transform 1 0 26386 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_300
timestamp 1607639953
transform 1 0 28686 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_288
timestamp 1607639953
transform 1 0 27582 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_324
timestamp 1607639953
transform 1 0 30894 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_312
timestamp 1607639953
transform 1 0 29790 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_349
timestamp 1607639953
transform 1 0 33194 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_337
timestamp 1607639953
transform 1 0 32090 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_579
timestamp 1607639953
transform 1 0 31998 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_363
timestamp 1607639953
transform 1 0 34482 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_357
timestamp 1607639953
transform 1 0 33930 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _056_
timestamp 1607639953
transform 1 0 34206 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_36_395
timestamp 1607639953
transform 1 0 37426 0 -1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_36_387
timestamp 1607639953
transform 1 0 36690 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_36_375
timestamp 1607639953
transform 1 0 35586 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_410
timestamp 1607639953
transform 1 0 38806 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_398
timestamp 1607639953
transform 1 0 37702 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_580
timestamp 1607639953
transform 1 0 37610 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_434
timestamp 1607639953
transform 1 0 41014 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_422
timestamp 1607639953
transform 1 0 39910 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_459
timestamp 1607639953
transform 1 0 43314 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_446
timestamp 1607639953
transform 1 0 42118 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_581
timestamp 1607639953
transform 1 0 43222 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_483
timestamp 1607639953
transform 1 0 45522 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_471
timestamp 1607639953
transform 1 0 44418 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_495
timestamp 1607639953
transform 1 0 46626 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_520
timestamp 1607639953
transform 1 0 48926 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_507
timestamp 1607639953
transform 1 0 47730 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_582
timestamp 1607639953
transform 1 0 48834 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_544
timestamp 1607639953
transform 1 0 51134 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_532
timestamp 1607639953
transform 1 0 50030 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_568
timestamp 1607639953
transform 1 0 53342 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_556
timestamp 1607639953
transform 1 0 52238 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_593
timestamp 1607639953
transform 1 0 55642 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_581
timestamp 1607639953
transform 1 0 54538 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_583
timestamp 1607639953
transform 1 0 54446 0 -1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_605
timestamp 1607639953
transform 1 0 56746 0 -1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_617
timestamp 1607639953
transform 1 0 57850 0 -1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1607639953
transform -1 0 58862 0 -1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_15
timestamp 1607639953
transform 1 0 2466 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_3
timestamp 1607639953
transform 1 0 1362 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1607639953
transform 1 0 1086 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_39
timestamp 1607639953
transform 1 0 4674 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_27
timestamp 1607639953
transform 1 0 3570 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_62
timestamp 1607639953
transform 1 0 6790 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_59
timestamp 1607639953
transform 1 0 6514 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_51
timestamp 1607639953
transform 1 0 5778 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_584
timestamp 1607639953
transform 1 0 6698 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_74
timestamp 1607639953
transform 1 0 7894 0 1 22304
box -38 -48 222 592
use NOR3X1  NOR3X1
timestamp 1608117647
transform 1 0 8078 0 1 22304
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_12  FILLER_37_102
timestamp 1607639953
transform 1 0 10470 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_90
timestamp 1607639953
transform 1 0 9366 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_123
timestamp 1607639953
transform 1 0 12402 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_114
timestamp 1607639953
transform 1 0 11574 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_585
timestamp 1607639953
transform 1 0 12310 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_147
timestamp 1607639953
transform 1 0 14610 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_135
timestamp 1607639953
transform 1 0 13506 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_171
timestamp 1607639953
transform 1 0 16818 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_159
timestamp 1607639953
transform 1 0 15714 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_196
timestamp 1607639953
transform 1 0 19118 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_184
timestamp 1607639953
transform 1 0 18014 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_586
timestamp 1607639953
transform 1 0 17922 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_220
timestamp 1607639953
transform 1 0 21326 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_208
timestamp 1607639953
transform 1 0 20222 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_232
timestamp 1607639953
transform 1 0 22430 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_257
timestamp 1607639953
transform 1 0 24730 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_245
timestamp 1607639953
transform 1 0 23626 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_587
timestamp 1607639953
transform 1 0 23534 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_281
timestamp 1607639953
transform 1 0 26938 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_269
timestamp 1607639953
transform 1 0 25834 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_306
timestamp 1607639953
transform 1 0 29238 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_293
timestamp 1607639953
transform 1 0 28042 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_588
timestamp 1607639953
transform 1 0 29146 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_330
timestamp 1607639953
transform 1 0 31446 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_318
timestamp 1607639953
transform 1 0 30342 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_342
timestamp 1607639953
transform 1 0 32550 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_367
timestamp 1607639953
transform 1 0 34850 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_354
timestamp 1607639953
transform 1 0 33654 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_589
timestamp 1607639953
transform 1 0 34758 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_391
timestamp 1607639953
transform 1 0 37058 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_379
timestamp 1607639953
transform 1 0 35954 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_415
timestamp 1607639953
transform 1 0 39266 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_403
timestamp 1607639953
transform 1 0 38162 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_440
timestamp 1607639953
transform 1 0 41566 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_436
timestamp 1607639953
transform 1 0 41198 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_428
timestamp 1607639953
transform 1 0 40462 0 1 22304
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_590
timestamp 1607639953
transform 1 0 40370 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _127_
timestamp 1607639953
transform 1 0 41290 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_452
timestamp 1607639953
transform 1 0 42670 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_476
timestamp 1607639953
transform 1 0 44878 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_464
timestamp 1607639953
transform 1 0 43774 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_501
timestamp 1607639953
transform 1 0 47178 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_489
timestamp 1607639953
transform 1 0 46074 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_591
timestamp 1607639953
transform 1 0 45982 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_525
timestamp 1607639953
transform 1 0 49386 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_513
timestamp 1607639953
transform 1 0 48282 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_550
timestamp 1607639953
transform 1 0 51686 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_537
timestamp 1607639953
transform 1 0 50490 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_592
timestamp 1607639953
transform 1 0 51594 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_562
timestamp 1607639953
transform 1 0 52790 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_586
timestamp 1607639953
transform 1 0 54998 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_574
timestamp 1607639953
transform 1 0 53894 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_611
timestamp 1607639953
transform 1 0 57298 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_598
timestamp 1607639953
transform 1 0 56102 0 1 22304
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_593
timestamp 1607639953
transform 1 0 57206 0 1 22304
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_623
timestamp 1607639953
transform 1 0 58402 0 1 22304
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1607639953
transform -1 0 58862 0 1 22304
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_15
timestamp 1607639953
transform 1 0 2466 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_3
timestamp 1607639953
transform 1 0 1362 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1607639953
transform 1 0 1086 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_44
timestamp 1607639953
transform 1 0 5134 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_32
timestamp 1607639953
transform 1 0 4030 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_27
timestamp 1607639953
transform 1 0 3570 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_594
timestamp 1607639953
transform 1 0 3938 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_64
timestamp 1607639953
transform 1 0 6974 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_60
timestamp 1607639953
transform 1 0 6606 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_56
timestamp 1607639953
transform 1 0 6238 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _113_
timestamp 1607639953
transform 1 0 6698 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_88
timestamp 1607639953
transform 1 0 9182 0 -1 23392
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_76
timestamp 1607639953
transform 1 0 8078 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_105
timestamp 1607639953
transform 1 0 10746 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_93
timestamp 1607639953
transform 1 0 9642 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_595
timestamp 1607639953
transform 1 0 9550 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_129
timestamp 1607639953
transform 1 0 12954 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_117
timestamp 1607639953
transform 1 0 11850 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_154
timestamp 1607639953
transform 1 0 15254 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_141
timestamp 1607639953
transform 1 0 14058 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_596
timestamp 1607639953
transform 1 0 15162 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_166
timestamp 1607639953
transform 1 0 16358 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_190
timestamp 1607639953
transform 1 0 18566 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_178
timestamp 1607639953
transform 1 0 17462 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_220
timestamp 1607639953
transform 1 0 21326 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_215
timestamp 1607639953
transform 1 0 20866 0 -1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_38_202
timestamp 1607639953
transform 1 0 19670 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_597
timestamp 1607639953
transform 1 0 20774 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _073_
timestamp 1607639953
transform 1 0 21050 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_38_232
timestamp 1607639953
transform 1 0 22430 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_256
timestamp 1607639953
transform 1 0 24638 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_244
timestamp 1607639953
transform 1 0 23534 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_276
timestamp 1607639953
transform 1 0 26478 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_274
timestamp 1607639953
transform 1 0 26294 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_38_268
timestamp 1607639953
transform 1 0 25742 0 -1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_598
timestamp 1607639953
transform 1 0 26386 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_300
timestamp 1607639953
transform 1 0 28686 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_288
timestamp 1607639953
transform 1 0 27582 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_324
timestamp 1607639953
transform 1 0 30894 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_312
timestamp 1607639953
transform 1 0 29790 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_349
timestamp 1607639953
transform 1 0 33194 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_337
timestamp 1607639953
transform 1 0 32090 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_599
timestamp 1607639953
transform 1 0 31998 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_373
timestamp 1607639953
transform 1 0 35402 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_361
timestamp 1607639953
transform 1 0 34298 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_385
timestamp 1607639953
transform 1 0 36506 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_410
timestamp 1607639953
transform 1 0 38806 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_398
timestamp 1607639953
transform 1 0 37702 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_600
timestamp 1607639953
transform 1 0 37610 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_434
timestamp 1607639953
transform 1 0 41014 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_422
timestamp 1607639953
transform 1 0 39910 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_459
timestamp 1607639953
transform 1 0 43314 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_446
timestamp 1607639953
transform 1 0 42118 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_601
timestamp 1607639953
transform 1 0 43222 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_483
timestamp 1607639953
transform 1 0 45522 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_471
timestamp 1607639953
transform 1 0 44418 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_495
timestamp 1607639953
transform 1 0 46626 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_520
timestamp 1607639953
transform 1 0 48926 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_507
timestamp 1607639953
transform 1 0 47730 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_602
timestamp 1607639953
transform 1 0 48834 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_544
timestamp 1607639953
transform 1 0 51134 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_532
timestamp 1607639953
transform 1 0 50030 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_568
timestamp 1607639953
transform 1 0 53342 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_556
timestamp 1607639953
transform 1 0 52238 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_593
timestamp 1607639953
transform 1 0 55642 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_581
timestamp 1607639953
transform 1 0 54538 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_603
timestamp 1607639953
transform 1 0 54446 0 -1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_605
timestamp 1607639953
transform 1 0 56746 0 -1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_617
timestamp 1607639953
transform 1 0 57850 0 -1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1607639953
transform -1 0 58862 0 -1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_40_15
timestamp 1607639953
transform 1 0 2466 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1607639953
transform 1 0 1362 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_15
timestamp 1607639953
transform 1 0 2466 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_3
timestamp 1607639953
transform 1 0 1362 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1607639953
transform 1 0 1086 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1607639953
transform 1 0 1086 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_40_44
timestamp 1607639953
transform 1 0 5134 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_32
timestamp 1607639953
transform 1 0 4030 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_27
timestamp 1607639953
transform 1 0 3570 0 -1 24480
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_39
timestamp 1607639953
transform 1 0 4674 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_27
timestamp 1607639953
transform 1 0 3570 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_614
timestamp 1607639953
transform 1 0 3938 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_56
timestamp 1607639953
transform 1 0 6238 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_62
timestamp 1607639953
transform 1 0 6790 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_59
timestamp 1607639953
transform 1 0 6514 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_39_51
timestamp 1607639953
transform 1 0 5778 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_604
timestamp 1607639953
transform 1 0 6698 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_80
timestamp 1607639953
transform 1 0 8446 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_68
timestamp 1607639953
transform 1 0 7342 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_84
timestamp 1607639953
transform 1 0 8814 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_74
timestamp 1607639953
transform 1 0 7894 0 1 23392
box -38 -48 222 592
use OAI21X1  OAI21X1
timestamp 1608117647
transform 1 0 8078 0 1 23392
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILLER_40_108
timestamp 1607639953
transform 1 0 11022 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_96
timestamp 1607639953
transform 1 0 9918 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_108
timestamp 1607639953
transform 1 0 11022 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_96
timestamp 1607639953
transform 1 0 9918 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_615
timestamp 1607639953
transform 1 0 9550 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _049_
timestamp 1607639953
transform 1 0 9642 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_40_132
timestamp 1607639953
transform 1 0 13230 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_120
timestamp 1607639953
transform 1 0 12126 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_123
timestamp 1607639953
transform 1 0 12402 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_120
timestamp 1607639953
transform 1 0 12126 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_605
timestamp 1607639953
transform 1 0 12310 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_154
timestamp 1607639953
transform 1 0 15254 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_152
timestamp 1607639953
transform 1 0 15070 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_144
timestamp 1607639953
transform 1 0 14334 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_39_147
timestamp 1607639953
transform 1 0 14610 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_135
timestamp 1607639953
transform 1 0 13506 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_616
timestamp 1607639953
transform 1 0 15162 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_166
timestamp 1607639953
transform 1 0 16358 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_171
timestamp 1607639953
transform 1 0 16818 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_159
timestamp 1607639953
transform 1 0 15714 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_198
timestamp 1607639953
transform 1 0 19302 0 -1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_190
timestamp 1607639953
transform 1 0 18566 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_178
timestamp 1607639953
transform 1 0 17462 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_196
timestamp 1607639953
transform 1 0 19118 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_184
timestamp 1607639953
transform 1 0 18014 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_606
timestamp 1607639953
transform 1 0 17922 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_215
timestamp 1607639953
transform 1 0 20866 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_211
timestamp 1607639953
transform 1 0 20498 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_40_203
timestamp 1607639953
transform 1 0 19762 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_39_220
timestamp 1607639953
transform 1 0 21326 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_208
timestamp 1607639953
transform 1 0 20222 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_617
timestamp 1607639953
transform 1 0 20774 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _064_
timestamp 1607639953
transform 1 0 19486 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_40_239
timestamp 1607639953
transform 1 0 23074 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_227
timestamp 1607639953
transform 1 0 21970 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_232
timestamp 1607639953
transform 1 0 22430 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_263
timestamp 1607639953
transform 1 0 25282 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_251
timestamp 1607639953
transform 1 0 24178 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_257
timestamp 1607639953
transform 1 0 24730 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_245
timestamp 1607639953
transform 1 0 23626 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_607
timestamp 1607639953
transform 1 0 23534 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_276
timestamp 1607639953
transform 1 0 26478 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_281
timestamp 1607639953
transform 1 0 26938 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_269
timestamp 1607639953
transform 1 0 25834 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_618
timestamp 1607639953
transform 1 0 26386 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_300
timestamp 1607639953
transform 1 0 28686 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_288
timestamp 1607639953
transform 1 0 27582 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_306
timestamp 1607639953
transform 1 0 29238 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_293
timestamp 1607639953
transform 1 0 28042 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_608
timestamp 1607639953
transform 1 0 29146 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_324
timestamp 1607639953
transform 1 0 30894 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_312
timestamp 1607639953
transform 1 0 29790 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_330
timestamp 1607639953
transform 1 0 31446 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_318
timestamp 1607639953
transform 1 0 30342 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_349
timestamp 1607639953
transform 1 0 33194 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_337
timestamp 1607639953
transform 1 0 32090 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_342
timestamp 1607639953
transform 1 0 32550 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_619
timestamp 1607639953
transform 1 0 31998 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_373
timestamp 1607639953
transform 1 0 35402 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_361
timestamp 1607639953
transform 1 0 34298 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_367
timestamp 1607639953
transform 1 0 34850 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_354
timestamp 1607639953
transform 1 0 33654 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_609
timestamp 1607639953
transform 1 0 34758 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_385
timestamp 1607639953
transform 1 0 36506 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_391
timestamp 1607639953
transform 1 0 37058 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_379
timestamp 1607639953
transform 1 0 35954 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_410
timestamp 1607639953
transform 1 0 38806 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_398
timestamp 1607639953
transform 1 0 37702 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_415
timestamp 1607639953
transform 1 0 39266 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_403
timestamp 1607639953
transform 1 0 38162 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_620
timestamp 1607639953
transform 1 0 37610 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_434
timestamp 1607639953
transform 1 0 41014 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_422
timestamp 1607639953
transform 1 0 39910 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_440
timestamp 1607639953
transform 1 0 41566 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_428
timestamp 1607639953
transform 1 0 40462 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_610
timestamp 1607639953
transform 1 0 40370 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_459
timestamp 1607639953
transform 1 0 43314 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_446
timestamp 1607639953
transform 1 0 42118 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_462
timestamp 1607639953
transform 1 0 43590 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_458
timestamp 1607639953
transform 1 0 43222 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_452
timestamp 1607639953
transform 1 0 42670 0 1 23392
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_621
timestamp 1607639953
transform 1 0 43222 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _180_
timestamp 1607639953
transform 1 0 43314 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_40_483
timestamp 1607639953
transform 1 0 45522 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_471
timestamp 1607639953
transform 1 0 44418 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_474
timestamp 1607639953
transform 1 0 44694 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_495
timestamp 1607639953
transform 1 0 46626 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_501
timestamp 1607639953
transform 1 0 47178 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_489
timestamp 1607639953
transform 1 0 46074 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_486
timestamp 1607639953
transform 1 0 45798 0 1 23392
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_611
timestamp 1607639953
transform 1 0 45982 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_524
timestamp 1607639953
transform 1 0 49294 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_520
timestamp 1607639953
transform 1 0 48926 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_507
timestamp 1607639953
transform 1 0 47730 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_528
timestamp 1607639953
transform 1 0 49662 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_513
timestamp 1607639953
transform 1 0 48282 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_622
timestamp 1607639953
transform 1 0 48834 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _093_
timestamp 1607639953
transform 1 0 49018 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _090_
timestamp 1607639953
transform 1 0 49386 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_40_548
timestamp 1607639953
transform 1 0 51502 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_536
timestamp 1607639953
transform 1 0 50398 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_550
timestamp 1607639953
transform 1 0 51686 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_39_548
timestamp 1607639953
transform 1 0 51502 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_540
timestamp 1607639953
transform 1 0 50766 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_612
timestamp 1607639953
transform 1 0 51594 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_572
timestamp 1607639953
transform 1 0 53710 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_40_560
timestamp 1607639953
transform 1 0 52606 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_562
timestamp 1607639953
transform 1 0 52790 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_593
timestamp 1607639953
transform 1 0 55642 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_581
timestamp 1607639953
transform 1 0 54538 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_586
timestamp 1607639953
transform 1 0 54998 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_574
timestamp 1607639953
transform 1 0 53894 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_623
timestamp 1607639953
transform 1 0 54446 0 -1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_605
timestamp 1607639953
transform 1 0 56746 0 -1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_614
timestamp 1607639953
transform 1 0 57574 0 1 23392
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_39_598
timestamp 1607639953
transform 1 0 56102 0 1 23392
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_613
timestamp 1607639953
transform 1 0 57206 0 1 23392
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _194_
timestamp 1607639953
transform 1 0 57298 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_40_617
timestamp 1607639953
transform 1 0 57850 0 -1 24480
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_622
timestamp 1607639953
transform 1 0 58310 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1607639953
transform -1 0 58862 0 -1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1607639953
transform -1 0 58862 0 1 23392
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_18
timestamp 1607639953
transform 1 0 2742 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_6
timestamp 1607639953
transform 1 0 1638 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1607639953
transform 1 0 1086 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _002_
timestamp 1607639953
transform 1 0 1362 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_42
timestamp 1607639953
transform 1 0 4950 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_30
timestamp 1607639953
transform 1 0 3846 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_62
timestamp 1607639953
transform 1 0 6790 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_60
timestamp 1607639953
transform 1 0 6606 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_54
timestamp 1607639953
transform 1 0 6054 0 1 24480
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_624
timestamp 1607639953
transform 1 0 6698 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_86
timestamp 1607639953
transform 1 0 8998 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_74
timestamp 1607639953
transform 1 0 7894 0 1 24480
box -38 -48 222 592
use OAI22X1  OAI22X1
timestamp 1608117647
transform 1 0 8078 0 1 24480
box 0 -48 920 592
use sky130_fd_sc_hd__decap_12  FILLER_41_110
timestamp 1607639953
transform 1 0 11206 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_98
timestamp 1607639953
transform 1 0 10102 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_123
timestamp 1607639953
transform 1 0 12402 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_625
timestamp 1607639953
transform 1 0 12310 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_147
timestamp 1607639953
transform 1 0 14610 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_135
timestamp 1607639953
transform 1 0 13506 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_171
timestamp 1607639953
transform 1 0 16818 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_159
timestamp 1607639953
transform 1 0 15714 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_196
timestamp 1607639953
transform 1 0 19118 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_184
timestamp 1607639953
transform 1 0 18014 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_626
timestamp 1607639953
transform 1 0 17922 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_220
timestamp 1607639953
transform 1 0 21326 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_208
timestamp 1607639953
transform 1 0 20222 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_232
timestamp 1607639953
transform 1 0 22430 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_257
timestamp 1607639953
transform 1 0 24730 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_245
timestamp 1607639953
transform 1 0 23626 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_627
timestamp 1607639953
transform 1 0 23534 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_281
timestamp 1607639953
transform 1 0 26938 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_269
timestamp 1607639953
transform 1 0 25834 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_306
timestamp 1607639953
transform 1 0 29238 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_293
timestamp 1607639953
transform 1 0 28042 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_628
timestamp 1607639953
transform 1 0 29146 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_330
timestamp 1607639953
transform 1 0 31446 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_318
timestamp 1607639953
transform 1 0 30342 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_342
timestamp 1607639953
transform 1 0 32550 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_367
timestamp 1607639953
transform 1 0 34850 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_354
timestamp 1607639953
transform 1 0 33654 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_629
timestamp 1607639953
transform 1 0 34758 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_391
timestamp 1607639953
transform 1 0 37058 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_379
timestamp 1607639953
transform 1 0 35954 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_415
timestamp 1607639953
transform 1 0 39266 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_403
timestamp 1607639953
transform 1 0 38162 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_440
timestamp 1607639953
transform 1 0 41566 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_428
timestamp 1607639953
transform 1 0 40462 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_630
timestamp 1607639953
transform 1 0 40370 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_452
timestamp 1607639953
transform 1 0 42670 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_476
timestamp 1607639953
transform 1 0 44878 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_464
timestamp 1607639953
transform 1 0 43774 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_501
timestamp 1607639953
transform 1 0 47178 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_489
timestamp 1607639953
transform 1 0 46074 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_631
timestamp 1607639953
transform 1 0 45982 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_525
timestamp 1607639953
transform 1 0 49386 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_513
timestamp 1607639953
transform 1 0 48282 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_550
timestamp 1607639953
transform 1 0 51686 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_537
timestamp 1607639953
transform 1 0 50490 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_632
timestamp 1607639953
transform 1 0 51594 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_562
timestamp 1607639953
transform 1 0 52790 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_586
timestamp 1607639953
transform 1 0 54998 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_574
timestamp 1607639953
transform 1 0 53894 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_611
timestamp 1607639953
transform 1 0 57298 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_598
timestamp 1607639953
transform 1 0 56102 0 1 24480
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_633
timestamp 1607639953
transform 1 0 57206 0 1 24480
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_623
timestamp 1607639953
transform 1 0 58402 0 1 24480
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1607639953
transform -1 0 58862 0 1 24480
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_15
timestamp 1607639953
transform 1 0 2466 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_3
timestamp 1607639953
transform 1 0 1362 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1607639953
transform 1 0 1086 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_44
timestamp 1607639953
transform 1 0 5134 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_32
timestamp 1607639953
transform 1 0 4030 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_27
timestamp 1607639953
transform 1 0 3570 0 -1 25568
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_634
timestamp 1607639953
transform 1 0 3938 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_56
timestamp 1607639953
transform 1 0 6238 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_80
timestamp 1607639953
transform 1 0 8446 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_68
timestamp 1607639953
transform 1 0 7342 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_105
timestamp 1607639953
transform 1 0 10746 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_93
timestamp 1607639953
transform 1 0 9642 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_635
timestamp 1607639953
transform 1 0 9550 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_129
timestamp 1607639953
transform 1 0 12954 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_117
timestamp 1607639953
transform 1 0 11850 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_154
timestamp 1607639953
transform 1 0 15254 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_141
timestamp 1607639953
transform 1 0 14058 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_636
timestamp 1607639953
transform 1 0 15162 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_166
timestamp 1607639953
transform 1 0 16358 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_190
timestamp 1607639953
transform 1 0 18566 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_178
timestamp 1607639953
transform 1 0 17462 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_215
timestamp 1607639953
transform 1 0 20866 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_202
timestamp 1607639953
transform 1 0 19670 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_637
timestamp 1607639953
transform 1 0 20774 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_239
timestamp 1607639953
transform 1 0 23074 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_227
timestamp 1607639953
transform 1 0 21970 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_263
timestamp 1607639953
transform 1 0 25282 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_251
timestamp 1607639953
transform 1 0 24178 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_276
timestamp 1607639953
transform 1 0 26478 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_638
timestamp 1607639953
transform 1 0 26386 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_300
timestamp 1607639953
transform 1 0 28686 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_288
timestamp 1607639953
transform 1 0 27582 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_324
timestamp 1607639953
transform 1 0 30894 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_312
timestamp 1607639953
transform 1 0 29790 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_349
timestamp 1607639953
transform 1 0 33194 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_337
timestamp 1607639953
transform 1 0 32090 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_639
timestamp 1607639953
transform 1 0 31998 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_373
timestamp 1607639953
transform 1 0 35402 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_361
timestamp 1607639953
transform 1 0 34298 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_385
timestamp 1607639953
transform 1 0 36506 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_410
timestamp 1607639953
transform 1 0 38806 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_398
timestamp 1607639953
transform 1 0 37702 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_640
timestamp 1607639953
transform 1 0 37610 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_434
timestamp 1607639953
transform 1 0 41014 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_422
timestamp 1607639953
transform 1 0 39910 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_459
timestamp 1607639953
transform 1 0 43314 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_446
timestamp 1607639953
transform 1 0 42118 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_641
timestamp 1607639953
transform 1 0 43222 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_483
timestamp 1607639953
transform 1 0 45522 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_471
timestamp 1607639953
transform 1 0 44418 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_495
timestamp 1607639953
transform 1 0 46626 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_520
timestamp 1607639953
transform 1 0 48926 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_507
timestamp 1607639953
transform 1 0 47730 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_642
timestamp 1607639953
transform 1 0 48834 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_544
timestamp 1607639953
transform 1 0 51134 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_532
timestamp 1607639953
transform 1 0 50030 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_568
timestamp 1607639953
transform 1 0 53342 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_556
timestamp 1607639953
transform 1 0 52238 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_593
timestamp 1607639953
transform 1 0 55642 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_581
timestamp 1607639953
transform 1 0 54538 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_643
timestamp 1607639953
transform 1 0 54446 0 -1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_605
timestamp 1607639953
transform 1 0 56746 0 -1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_617
timestamp 1607639953
transform 1 0 57850 0 -1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1607639953
transform -1 0 58862 0 -1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_15
timestamp 1607639953
transform 1 0 2466 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_3
timestamp 1607639953
transform 1 0 1362 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1607639953
transform 1 0 1086 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_39
timestamp 1607639953
transform 1 0 4674 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_27
timestamp 1607639953
transform 1 0 3570 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_62
timestamp 1607639953
transform 1 0 6790 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_59
timestamp 1607639953
transform 1 0 6514 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_51
timestamp 1607639953
transform 1 0 5778 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_644
timestamp 1607639953
transform 1 0 6698 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_84
timestamp 1607639953
transform 1 0 8814 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_75
timestamp 1607639953
transform 1 0 7986 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_70
timestamp 1607639953
transform 1 0 7526 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _121_
timestamp 1607639953
transform 1 0 7710 0 1 25568
box -38 -48 314 592
use OR2X1  OR2X1
timestamp 1608117647
transform 1 0 8078 0 1 25568
box 0 -48 736 592
use sky130_fd_sc_hd__fill_2  FILLER_43_108
timestamp 1607639953
transform 1 0 11022 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_43_96
timestamp 1607639953
transform 1 0 9918 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _031_
timestamp 1607639953
transform 1 0 11206 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_123
timestamp 1607639953
transform 1 0 12402 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_121
timestamp 1607639953
transform 1 0 12218 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_113
timestamp 1607639953
transform 1 0 11482 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_645
timestamp 1607639953
transform 1 0 12310 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_147
timestamp 1607639953
transform 1 0 14610 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_135
timestamp 1607639953
transform 1 0 13506 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_171
timestamp 1607639953
transform 1 0 16818 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_159
timestamp 1607639953
transform 1 0 15714 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_196
timestamp 1607639953
transform 1 0 19118 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_184
timestamp 1607639953
transform 1 0 18014 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_646
timestamp 1607639953
transform 1 0 17922 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_220
timestamp 1607639953
transform 1 0 21326 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_208
timestamp 1607639953
transform 1 0 20222 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_232
timestamp 1607639953
transform 1 0 22430 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_257
timestamp 1607639953
transform 1 0 24730 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_245
timestamp 1607639953
transform 1 0 23626 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_647
timestamp 1607639953
transform 1 0 23534 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_281
timestamp 1607639953
transform 1 0 26938 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_269
timestamp 1607639953
transform 1 0 25834 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_306
timestamp 1607639953
transform 1 0 29238 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_293
timestamp 1607639953
transform 1 0 28042 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_648
timestamp 1607639953
transform 1 0 29146 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_330
timestamp 1607639953
transform 1 0 31446 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_318
timestamp 1607639953
transform 1 0 30342 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_342
timestamp 1607639953
transform 1 0 32550 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_367
timestamp 1607639953
transform 1 0 34850 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_354
timestamp 1607639953
transform 1 0 33654 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_649
timestamp 1607639953
transform 1 0 34758 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_391
timestamp 1607639953
transform 1 0 37058 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_379
timestamp 1607639953
transform 1 0 35954 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_415
timestamp 1607639953
transform 1 0 39266 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_403
timestamp 1607639953
transform 1 0 38162 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_440
timestamp 1607639953
transform 1 0 41566 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_43_428
timestamp 1607639953
transform 1 0 40462 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_650
timestamp 1607639953
transform 1 0 40370 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_454
timestamp 1607639953
transform 1 0 42854 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_448
timestamp 1607639953
transform 1 0 42302 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _107_
timestamp 1607639953
transform 1 0 42578 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_43_478
timestamp 1607639953
transform 1 0 45062 0 1 25568
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_43_466
timestamp 1607639953
transform 1 0 43958 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_501
timestamp 1607639953
transform 1 0 47178 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_489
timestamp 1607639953
transform 1 0 46074 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_486
timestamp 1607639953
transform 1 0 45798 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_651
timestamp 1607639953
transform 1 0 45982 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_525
timestamp 1607639953
transform 1 0 49386 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_513
timestamp 1607639953
transform 1 0 48282 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_550
timestamp 1607639953
transform 1 0 51686 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_537
timestamp 1607639953
transform 1 0 50490 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_652
timestamp 1607639953
transform 1 0 51594 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_562
timestamp 1607639953
transform 1 0 52790 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_586
timestamp 1607639953
transform 1 0 54998 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_574
timestamp 1607639953
transform 1 0 53894 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_611
timestamp 1607639953
transform 1 0 57298 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_598
timestamp 1607639953
transform 1 0 56102 0 1 25568
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_653
timestamp 1607639953
transform 1 0 57206 0 1 25568
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_623
timestamp 1607639953
transform 1 0 58402 0 1 25568
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1607639953
transform -1 0 58862 0 1 25568
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_44_15
timestamp 1607639953
transform 1 0 2466 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_3
timestamp 1607639953
transform 1 0 1362 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1607639953
transform 1 0 1086 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_44_35
timestamp 1607639953
transform 1 0 4306 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_27
timestamp 1607639953
transform 1 0 3570 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_654
timestamp 1607639953
transform 1 0 3938 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _037_
timestamp 1607639953
transform 1 0 4030 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_44_59
timestamp 1607639953
transform 1 0 6514 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_47
timestamp 1607639953
transform 1 0 5410 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_83
timestamp 1607639953
transform 1 0 8722 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_71
timestamp 1607639953
transform 1 0 7618 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_105
timestamp 1607639953
transform 1 0 10746 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_93
timestamp 1607639953
transform 1 0 9642 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_91
timestamp 1607639953
transform 1 0 9458 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_655
timestamp 1607639953
transform 1 0 9550 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_129
timestamp 1607639953
transform 1 0 12954 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_117
timestamp 1607639953
transform 1 0 11850 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_154
timestamp 1607639953
transform 1 0 15254 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_141
timestamp 1607639953
transform 1 0 14058 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_656
timestamp 1607639953
transform 1 0 15162 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_166
timestamp 1607639953
transform 1 0 16358 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_190
timestamp 1607639953
transform 1 0 18566 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_178
timestamp 1607639953
transform 1 0 17462 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_215
timestamp 1607639953
transform 1 0 20866 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_202
timestamp 1607639953
transform 1 0 19670 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_657
timestamp 1607639953
transform 1 0 20774 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_239
timestamp 1607639953
transform 1 0 23074 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_227
timestamp 1607639953
transform 1 0 21970 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_263
timestamp 1607639953
transform 1 0 25282 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_251
timestamp 1607639953
transform 1 0 24178 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_276
timestamp 1607639953
transform 1 0 26478 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_658
timestamp 1607639953
transform 1 0 26386 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_300
timestamp 1607639953
transform 1 0 28686 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_288
timestamp 1607639953
transform 1 0 27582 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_324
timestamp 1607639953
transform 1 0 30894 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_312
timestamp 1607639953
transform 1 0 29790 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_349
timestamp 1607639953
transform 1 0 33194 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_337
timestamp 1607639953
transform 1 0 32090 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_659
timestamp 1607639953
transform 1 0 31998 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_373
timestamp 1607639953
transform 1 0 35402 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_361
timestamp 1607639953
transform 1 0 34298 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_385
timestamp 1607639953
transform 1 0 36506 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_408
timestamp 1607639953
transform 1 0 38622 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_404
timestamp 1607639953
transform 1 0 38254 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_398
timestamp 1607639953
transform 1 0 37702 0 -1 26656
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_660
timestamp 1607639953
transform 1 0 37610 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _027_
timestamp 1607639953
transform 1 0 38346 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_44_438
timestamp 1607639953
transform 1 0 41382 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_426
timestamp 1607639953
transform 1 0 40278 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_44_420
timestamp 1607639953
transform 1 0 39726 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _164_
timestamp 1607639953
transform 1 0 40002 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_44_459
timestamp 1607639953
transform 1 0 43314 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_450
timestamp 1607639953
transform 1 0 42486 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_661
timestamp 1607639953
transform 1 0 43222 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_483
timestamp 1607639953
transform 1 0 45522 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_471
timestamp 1607639953
transform 1 0 44418 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_495
timestamp 1607639953
transform 1 0 46626 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_520
timestamp 1607639953
transform 1 0 48926 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_507
timestamp 1607639953
transform 1 0 47730 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_662
timestamp 1607639953
transform 1 0 48834 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_548
timestamp 1607639953
transform 1 0 51502 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_536
timestamp 1607639953
transform 1 0 50398 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_532
timestamp 1607639953
transform 1 0 50030 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _188_
timestamp 1607639953
transform 1 0 50122 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_44_572
timestamp 1607639953
transform 1 0 53710 0 -1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_44_560
timestamp 1607639953
transform 1 0 52606 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_593
timestamp 1607639953
transform 1 0 55642 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_581
timestamp 1607639953
transform 1 0 54538 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_663
timestamp 1607639953
transform 1 0 54446 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_612
timestamp 1607639953
transform 1 0 57390 0 -1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_605
timestamp 1607639953
transform 1 0 56746 0 -1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _000_
timestamp 1607639953
transform 1 0 57114 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_44_624
timestamp 1607639953
transform 1 0 58494 0 -1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1607639953
transform -1 0 58862 0 -1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_15
timestamp 1607639953
transform 1 0 2466 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_3
timestamp 1607639953
transform 1 0 1362 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1607639953
transform 1 0 1086 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_39
timestamp 1607639953
transform 1 0 4674 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_27
timestamp 1607639953
transform 1 0 3570 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_62
timestamp 1607639953
transform 1 0 6790 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_59
timestamp 1607639953
transform 1 0 6514 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_45_51
timestamp 1607639953
transform 1 0 5778 0 1 26656
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_664
timestamp 1607639953
transform 1 0 6698 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_84
timestamp 1607639953
transform 1 0 8814 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_74
timestamp 1607639953
transform 1 0 7894 0 1 26656
box -38 -48 222 592
use OR2X2  OR2X2
timestamp 1608117647
transform 1 0 8078 0 1 26656
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILLER_45_108
timestamp 1607639953
transform 1 0 11022 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_96
timestamp 1607639953
transform 1 0 9918 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_123
timestamp 1607639953
transform 1 0 12402 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_120
timestamp 1607639953
transform 1 0 12126 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_665
timestamp 1607639953
transform 1 0 12310 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_147
timestamp 1607639953
transform 1 0 14610 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_135
timestamp 1607639953
transform 1 0 13506 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_171
timestamp 1607639953
transform 1 0 16818 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_159
timestamp 1607639953
transform 1 0 15714 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_196
timestamp 1607639953
transform 1 0 19118 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_184
timestamp 1607639953
transform 1 0 18014 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_666
timestamp 1607639953
transform 1 0 17922 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_220
timestamp 1607639953
transform 1 0 21326 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_208
timestamp 1607639953
transform 1 0 20222 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_232
timestamp 1607639953
transform 1 0 22430 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_257
timestamp 1607639953
transform 1 0 24730 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_245
timestamp 1607639953
transform 1 0 23626 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_667
timestamp 1607639953
transform 1 0 23534 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_281
timestamp 1607639953
transform 1 0 26938 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_269
timestamp 1607639953
transform 1 0 25834 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_306
timestamp 1607639953
transform 1 0 29238 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_293
timestamp 1607639953
transform 1 0 28042 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_668
timestamp 1607639953
transform 1 0 29146 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_330
timestamp 1607639953
transform 1 0 31446 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_318
timestamp 1607639953
transform 1 0 30342 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_342
timestamp 1607639953
transform 1 0 32550 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_367
timestamp 1607639953
transform 1 0 34850 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_354
timestamp 1607639953
transform 1 0 33654 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_669
timestamp 1607639953
transform 1 0 34758 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_391
timestamp 1607639953
transform 1 0 37058 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_379
timestamp 1607639953
transform 1 0 35954 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_415
timestamp 1607639953
transform 1 0 39266 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_403
timestamp 1607639953
transform 1 0 38162 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_440
timestamp 1607639953
transform 1 0 41566 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_428
timestamp 1607639953
transform 1 0 40462 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_670
timestamp 1607639953
transform 1 0 40370 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_452
timestamp 1607639953
transform 1 0 42670 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_476
timestamp 1607639953
transform 1 0 44878 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_464
timestamp 1607639953
transform 1 0 43774 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_501
timestamp 1607639953
transform 1 0 47178 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_489
timestamp 1607639953
transform 1 0 46074 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_671
timestamp 1607639953
transform 1 0 45982 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_525
timestamp 1607639953
transform 1 0 49386 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_513
timestamp 1607639953
transform 1 0 48282 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_537
timestamp 1607639953
transform 1 0 50490 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_672
timestamp 1607639953
transform 1 0 51594 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _167_
timestamp 1607639953
transform 1 0 51686 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_569
timestamp 1607639953
transform 1 0 53434 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_565
timestamp 1607639953
transform 1 0 53066 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_553
timestamp 1607639953
transform 1 0 51962 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _134_
timestamp 1607639953
transform 1 0 53158 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_593
timestamp 1607639953
transform 1 0 55642 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_581
timestamp 1607639953
transform 1 0 54538 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_611
timestamp 1607639953
transform 1 0 57298 0 1 26656
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_609
timestamp 1607639953
transform 1 0 57114 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_605
timestamp 1607639953
transform 1 0 56746 0 1 26656
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_673
timestamp 1607639953
transform 1 0 57206 0 1 26656
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_45_623
timestamp 1607639953
transform 1 0 58402 0 1 26656
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1607639953
transform -1 0 58862 0 1 26656
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_47_15
timestamp 1607639953
transform 1 0 2466 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_3
timestamp 1607639953
transform 1 0 1362 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_15
timestamp 1607639953
transform 1 0 2466 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_3
timestamp 1607639953
transform 1 0 1362 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1607639953
transform 1 0 1086 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1607639953
transform 1 0 1086 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_47_39
timestamp 1607639953
transform 1 0 4674 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_27
timestamp 1607639953
transform 1 0 3570 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_44
timestamp 1607639953
transform 1 0 5134 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_32
timestamp 1607639953
transform 1 0 4030 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_27
timestamp 1607639953
transform 1 0 3570 0 -1 27744
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_674
timestamp 1607639953
transform 1 0 3938 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_62
timestamp 1607639953
transform 1 0 6790 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_59
timestamp 1607639953
transform 1 0 6514 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_51
timestamp 1607639953
transform 1 0 5778 0 1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_46_56
timestamp 1607639953
transform 1 0 6238 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_684
timestamp 1607639953
transform 1 0 6698 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_84
timestamp 1607639953
transform 1 0 8814 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_74
timestamp 1607639953
transform 1 0 7894 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_46_80
timestamp 1607639953
transform 1 0 8446 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_68
timestamp 1607639953
transform 1 0 7342 0 -1 27744
box -38 -48 1142 592
use TBUFX1  TBUFX1
timestamp 1608117647
transform 1 0 8078 0 1 27744
box 0 -48 736 592
use sky130_fd_sc_hd__decap_12  FILLER_47_108
timestamp 1607639953
transform 1 0 11022 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_96
timestamp 1607639953
transform 1 0 9918 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_105
timestamp 1607639953
transform 1 0 10746 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_93
timestamp 1607639953
transform 1 0 9642 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_675
timestamp 1607639953
transform 1 0 9550 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_123
timestamp 1607639953
transform 1 0 12402 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_120
timestamp 1607639953
transform 1 0 12126 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_46_129
timestamp 1607639953
transform 1 0 12954 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_117
timestamp 1607639953
transform 1 0 11850 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_685
timestamp 1607639953
transform 1 0 12310 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_147
timestamp 1607639953
transform 1 0 14610 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_135
timestamp 1607639953
transform 1 0 13506 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_141
timestamp 1607639953
transform 1 0 14058 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_676
timestamp 1607639953
transform 1 0 15162 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _069_
timestamp 1607639953
transform 1 0 15254 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_47_171
timestamp 1607639953
transform 1 0 16818 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_159
timestamp 1607639953
transform 1 0 15714 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_169
timestamp 1607639953
transform 1 0 16634 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_157
timestamp 1607639953
transform 1 0 15530 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_196
timestamp 1607639953
transform 1 0 19118 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_184
timestamp 1607639953
transform 1 0 18014 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_193
timestamp 1607639953
transform 1 0 18842 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_181
timestamp 1607639953
transform 1 0 17738 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_686
timestamp 1607639953
transform 1 0 17922 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_220
timestamp 1607639953
transform 1 0 21326 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_208
timestamp 1607639953
transform 1 0 20222 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_215
timestamp 1607639953
transform 1 0 20866 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_213
timestamp 1607639953
transform 1 0 20682 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_205
timestamp 1607639953
transform 1 0 19946 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_677
timestamp 1607639953
transform 1 0 20774 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_232
timestamp 1607639953
transform 1 0 22430 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_239
timestamp 1607639953
transform 1 0 23074 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_227
timestamp 1607639953
transform 1 0 21970 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_257
timestamp 1607639953
transform 1 0 24730 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_245
timestamp 1607639953
transform 1 0 23626 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_263
timestamp 1607639953
transform 1 0 25282 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_251
timestamp 1607639953
transform 1 0 24178 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_687
timestamp 1607639953
transform 1 0 23534 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_281
timestamp 1607639953
transform 1 0 26938 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_269
timestamp 1607639953
transform 1 0 25834 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_276
timestamp 1607639953
transform 1 0 26478 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_678
timestamp 1607639953
transform 1 0 26386 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_306
timestamp 1607639953
transform 1 0 29238 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_293
timestamp 1607639953
transform 1 0 28042 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_300
timestamp 1607639953
transform 1 0 28686 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_288
timestamp 1607639953
transform 1 0 27582 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_688
timestamp 1607639953
transform 1 0 29146 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_330
timestamp 1607639953
transform 1 0 31446 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_318
timestamp 1607639953
transform 1 0 30342 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_324
timestamp 1607639953
transform 1 0 30894 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_312
timestamp 1607639953
transform 1 0 29790 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_342
timestamp 1607639953
transform 1 0 32550 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_349
timestamp 1607639953
transform 1 0 33194 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_337
timestamp 1607639953
transform 1 0 32090 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_679
timestamp 1607639953
transform 1 0 31998 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_367
timestamp 1607639953
transform 1 0 34850 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_354
timestamp 1607639953
transform 1 0 33654 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_373
timestamp 1607639953
transform 1 0 35402 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_361
timestamp 1607639953
transform 1 0 34298 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_689
timestamp 1607639953
transform 1 0 34758 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_391
timestamp 1607639953
transform 1 0 37058 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_379
timestamp 1607639953
transform 1 0 35954 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_385
timestamp 1607639953
transform 1 0 36506 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_415
timestamp 1607639953
transform 1 0 39266 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_403
timestamp 1607639953
transform 1 0 38162 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_410
timestamp 1607639953
transform 1 0 38806 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_398
timestamp 1607639953
transform 1 0 37702 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_680
timestamp 1607639953
transform 1 0 37610 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_440
timestamp 1607639953
transform 1 0 41566 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_428
timestamp 1607639953
transform 1 0 40462 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_434
timestamp 1607639953
transform 1 0 41014 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_422
timestamp 1607639953
transform 1 0 39910 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_690
timestamp 1607639953
transform 1 0 40370 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_452
timestamp 1607639953
transform 1 0 42670 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_459
timestamp 1607639953
transform 1 0 43314 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_446
timestamp 1607639953
transform 1 0 42118 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_681
timestamp 1607639953
transform 1 0 43222 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_476
timestamp 1607639953
transform 1 0 44878 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_464
timestamp 1607639953
transform 1 0 43774 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_483
timestamp 1607639953
transform 1 0 45522 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_471
timestamp 1607639953
transform 1 0 44418 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_501
timestamp 1607639953
transform 1 0 47178 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_489
timestamp 1607639953
transform 1 0 46074 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_495
timestamp 1607639953
transform 1 0 46626 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_691
timestamp 1607639953
transform 1 0 45982 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_525
timestamp 1607639953
transform 1 0 49386 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_513
timestamp 1607639953
transform 1 0 48282 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_520
timestamp 1607639953
transform 1 0 48926 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_507
timestamp 1607639953
transform 1 0 47730 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_682
timestamp 1607639953
transform 1 0 48834 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_550
timestamp 1607639953
transform 1 0 51686 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_537
timestamp 1607639953
transform 1 0 50490 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_544
timestamp 1607639953
transform 1 0 51134 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_532
timestamp 1607639953
transform 1 0 50030 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_692
timestamp 1607639953
transform 1 0 51594 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_562
timestamp 1607639953
transform 1 0 52790 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_568
timestamp 1607639953
transform 1 0 53342 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_556
timestamp 1607639953
transform 1 0 52238 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_586
timestamp 1607639953
transform 1 0 54998 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_574
timestamp 1607639953
transform 1 0 53894 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_593
timestamp 1607639953
transform 1 0 55642 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_581
timestamp 1607639953
transform 1 0 54538 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_683
timestamp 1607639953
transform 1 0 54446 0 -1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_611
timestamp 1607639953
transform 1 0 57298 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_598
timestamp 1607639953
transform 1 0 56102 0 1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_605
timestamp 1607639953
transform 1 0 56746 0 -1 27744
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_693
timestamp 1607639953
transform 1 0 57206 0 1 27744
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_623
timestamp 1607639953
transform 1 0 58402 0 1 27744
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_46_617
timestamp 1607639953
transform 1 0 57850 0 -1 27744
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1607639953
transform -1 0 58862 0 1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1607639953
transform -1 0 58862 0 -1 27744
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_48_15
timestamp 1607639953
transform 1 0 2466 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_3
timestamp 1607639953
transform 1 0 1362 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1607639953
transform 1 0 1086 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_48_44
timestamp 1607639953
transform 1 0 5134 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_32
timestamp 1607639953
transform 1 0 4030 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_30
timestamp 1607639953
transform 1 0 3846 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_694
timestamp 1607639953
transform 1 0 3938 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _050_
timestamp 1607639953
transform 1 0 3570 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_48_56
timestamp 1607639953
transform 1 0 6238 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_80
timestamp 1607639953
transform 1 0 8446 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_68
timestamp 1607639953
transform 1 0 7342 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_105
timestamp 1607639953
transform 1 0 10746 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_93
timestamp 1607639953
transform 1 0 9642 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_695
timestamp 1607639953
transform 1 0 9550 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_129
timestamp 1607639953
transform 1 0 12954 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_117
timestamp 1607639953
transform 1 0 11850 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_154
timestamp 1607639953
transform 1 0 15254 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_141
timestamp 1607639953
transform 1 0 14058 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_696
timestamp 1607639953
transform 1 0 15162 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_166
timestamp 1607639953
transform 1 0 16358 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_190
timestamp 1607639953
transform 1 0 18566 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_178
timestamp 1607639953
transform 1 0 17462 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_215
timestamp 1607639953
transform 1 0 20866 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_202
timestamp 1607639953
transform 1 0 19670 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_697
timestamp 1607639953
transform 1 0 20774 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_239
timestamp 1607639953
transform 1 0 23074 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_227
timestamp 1607639953
transform 1 0 21970 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_263
timestamp 1607639953
transform 1 0 25282 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_251
timestamp 1607639953
transform 1 0 24178 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_279
timestamp 1607639953
transform 1 0 26754 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_698
timestamp 1607639953
transform 1 0 26386 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _128_
timestamp 1607639953
transform 1 0 26478 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_48_303
timestamp 1607639953
transform 1 0 28962 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_291
timestamp 1607639953
transform 1 0 27858 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_327
timestamp 1607639953
transform 1 0 31170 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_315
timestamp 1607639953
transform 1 0 30066 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_349
timestamp 1607639953
transform 1 0 33194 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_337
timestamp 1607639953
transform 1 0 32090 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_335
timestamp 1607639953
transform 1 0 31906 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_699
timestamp 1607639953
transform 1 0 31998 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_373
timestamp 1607639953
transform 1 0 35402 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_361
timestamp 1607639953
transform 1 0 34298 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_385
timestamp 1607639953
transform 1 0 36506 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_410
timestamp 1607639953
transform 1 0 38806 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_398
timestamp 1607639953
transform 1 0 37702 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_700
timestamp 1607639953
transform 1 0 37610 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_434
timestamp 1607639953
transform 1 0 41014 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_422
timestamp 1607639953
transform 1 0 39910 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_459
timestamp 1607639953
transform 1 0 43314 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_446
timestamp 1607639953
transform 1 0 42118 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_701
timestamp 1607639953
transform 1 0 43222 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_483
timestamp 1607639953
transform 1 0 45522 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_471
timestamp 1607639953
transform 1 0 44418 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_495
timestamp 1607639953
transform 1 0 46626 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_520
timestamp 1607639953
transform 1 0 48926 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_507
timestamp 1607639953
transform 1 0 47730 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_702
timestamp 1607639953
transform 1 0 48834 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_544
timestamp 1607639953
transform 1 0 51134 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_532
timestamp 1607639953
transform 1 0 50030 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_568
timestamp 1607639953
transform 1 0 53342 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_556
timestamp 1607639953
transform 1 0 52238 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_593
timestamp 1607639953
transform 1 0 55642 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_581
timestamp 1607639953
transform 1 0 54538 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_703
timestamp 1607639953
transform 1 0 54446 0 -1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_605
timestamp 1607639953
transform 1 0 56746 0 -1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_617
timestamp 1607639953
transform 1 0 57850 0 -1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1607639953
transform -1 0 58862 0 -1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_49_15
timestamp 1607639953
transform 1 0 2466 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_3
timestamp 1607639953
transform 1 0 1362 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1607639953
transform 1 0 1086 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_49_39
timestamp 1607639953
transform 1 0 4674 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_27
timestamp 1607639953
transform 1 0 3570 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_62
timestamp 1607639953
transform 1 0 6790 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_59
timestamp 1607639953
transform 1 0 6514 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_51
timestamp 1607639953
transform 1 0 5778 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_704
timestamp 1607639953
transform 1 0 6698 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_88
timestamp 1607639953
transform 1 0 9182 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_74
timestamp 1607639953
transform 1 0 7894 0 1 28832
box -38 -48 222 592
use TBUFX2  TBUFX2
timestamp 1608117647
transform 1 0 8078 0 1 28832
box 0 -48 1104 592
use sky130_fd_sc_hd__decap_12  FILLER_49_100
timestamp 1607639953
transform 1 0 10286 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_123
timestamp 1607639953
transform 1 0 12402 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_120
timestamp 1607639953
transform 1 0 12126 0 1 28832
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_49_112
timestamp 1607639953
transform 1 0 11390 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_705
timestamp 1607639953
transform 1 0 12310 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_147
timestamp 1607639953
transform 1 0 14610 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_135
timestamp 1607639953
transform 1 0 13506 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_171
timestamp 1607639953
transform 1 0 16818 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_159
timestamp 1607639953
transform 1 0 15714 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_196
timestamp 1607639953
transform 1 0 19118 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_184
timestamp 1607639953
transform 1 0 18014 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_706
timestamp 1607639953
transform 1 0 17922 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_220
timestamp 1607639953
transform 1 0 21326 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_208
timestamp 1607639953
transform 1 0 20222 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_232
timestamp 1607639953
transform 1 0 22430 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_257
timestamp 1607639953
transform 1 0 24730 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_245
timestamp 1607639953
transform 1 0 23626 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_707
timestamp 1607639953
transform 1 0 23534 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_281
timestamp 1607639953
transform 1 0 26938 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_269
timestamp 1607639953
transform 1 0 25834 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_306
timestamp 1607639953
transform 1 0 29238 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_293
timestamp 1607639953
transform 1 0 28042 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_708
timestamp 1607639953
transform 1 0 29146 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_330
timestamp 1607639953
transform 1 0 31446 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_318
timestamp 1607639953
transform 1 0 30342 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_342
timestamp 1607639953
transform 1 0 32550 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_367
timestamp 1607639953
transform 1 0 34850 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_354
timestamp 1607639953
transform 1 0 33654 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_709
timestamp 1607639953
transform 1 0 34758 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_391
timestamp 1607639953
transform 1 0 37058 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_379
timestamp 1607639953
transform 1 0 35954 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_415
timestamp 1607639953
transform 1 0 39266 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_403
timestamp 1607639953
transform 1 0 38162 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_440
timestamp 1607639953
transform 1 0 41566 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_428
timestamp 1607639953
transform 1 0 40462 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_710
timestamp 1607639953
transform 1 0 40370 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_452
timestamp 1607639953
transform 1 0 42670 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_476
timestamp 1607639953
transform 1 0 44878 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_464
timestamp 1607639953
transform 1 0 43774 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_501
timestamp 1607639953
transform 1 0 47178 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_489
timestamp 1607639953
transform 1 0 46074 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_711
timestamp 1607639953
transform 1 0 45982 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_525
timestamp 1607639953
transform 1 0 49386 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_513
timestamp 1607639953
transform 1 0 48282 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_550
timestamp 1607639953
transform 1 0 51686 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_548
timestamp 1607639953
transform 1 0 51502 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_537
timestamp 1607639953
transform 1 0 50490 0 1 28832
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_712
timestamp 1607639953
transform 1 0 51594 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _101_
timestamp 1607639953
transform 1 0 51226 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_49_562
timestamp 1607639953
transform 1 0 52790 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_586
timestamp 1607639953
transform 1 0 54998 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_574
timestamp 1607639953
transform 1 0 53894 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_611
timestamp 1607639953
transform 1 0 57298 0 1 28832
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_598
timestamp 1607639953
transform 1 0 56102 0 1 28832
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_713
timestamp 1607639953
transform 1 0 57206 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _103_
timestamp 1607639953
transform 1 0 57666 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_49_624
timestamp 1607639953
transform 1 0 58494 0 1 28832
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_49_618
timestamp 1607639953
transform 1 0 57942 0 1 28832
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1607639953
transform -1 0 58862 0 1 28832
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_50_15
timestamp 1607639953
transform 1 0 2466 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_3
timestamp 1607639953
transform 1 0 1362 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1607639953
transform 1 0 1086 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_50_44
timestamp 1607639953
transform 1 0 5134 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_32
timestamp 1607639953
transform 1 0 4030 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_27
timestamp 1607639953
transform 1 0 3570 0 -1 29920
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_714
timestamp 1607639953
transform 1 0 3938 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_56
timestamp 1607639953
transform 1 0 6238 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_80
timestamp 1607639953
transform 1 0 8446 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_68
timestamp 1607639953
transform 1 0 7342 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_105
timestamp 1607639953
transform 1 0 10746 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_93
timestamp 1607639953
transform 1 0 9642 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_715
timestamp 1607639953
transform 1 0 9550 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_129
timestamp 1607639953
transform 1 0 12954 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_117
timestamp 1607639953
transform 1 0 11850 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_154
timestamp 1607639953
transform 1 0 15254 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_141
timestamp 1607639953
transform 1 0 14058 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_716
timestamp 1607639953
transform 1 0 15162 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_166
timestamp 1607639953
transform 1 0 16358 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_190
timestamp 1607639953
transform 1 0 18566 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_178
timestamp 1607639953
transform 1 0 17462 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_215
timestamp 1607639953
transform 1 0 20866 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_202
timestamp 1607639953
transform 1 0 19670 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_717
timestamp 1607639953
transform 1 0 20774 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_239
timestamp 1607639953
transform 1 0 23074 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_227
timestamp 1607639953
transform 1 0 21970 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_263
timestamp 1607639953
transform 1 0 25282 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_251
timestamp 1607639953
transform 1 0 24178 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_279
timestamp 1607639953
transform 1 0 26754 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_718
timestamp 1607639953
transform 1 0 26386 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _169_
timestamp 1607639953
transform 1 0 26478 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_50_303
timestamp 1607639953
transform 1 0 28962 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_291
timestamp 1607639953
transform 1 0 27858 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_327
timestamp 1607639953
transform 1 0 31170 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_50_315
timestamp 1607639953
transform 1 0 30066 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_349
timestamp 1607639953
transform 1 0 33194 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_337
timestamp 1607639953
transform 1 0 32090 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_335
timestamp 1607639953
transform 1 0 31906 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_719
timestamp 1607639953
transform 1 0 31998 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_373
timestamp 1607639953
transform 1 0 35402 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_361
timestamp 1607639953
transform 1 0 34298 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_385
timestamp 1607639953
transform 1 0 36506 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_410
timestamp 1607639953
transform 1 0 38806 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_398
timestamp 1607639953
transform 1 0 37702 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_720
timestamp 1607639953
transform 1 0 37610 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_434
timestamp 1607639953
transform 1 0 41014 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_422
timestamp 1607639953
transform 1 0 39910 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_459
timestamp 1607639953
transform 1 0 43314 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_446
timestamp 1607639953
transform 1 0 42118 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_721
timestamp 1607639953
transform 1 0 43222 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_471
timestamp 1607639953
transform 1 0 44418 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _153_
timestamp 1607639953
transform 1 0 45522 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_50_498
timestamp 1607639953
transform 1 0 46902 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_486
timestamp 1607639953
transform 1 0 45798 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_520
timestamp 1607639953
transform 1 0 48926 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_518
timestamp 1607639953
transform 1 0 48742 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_510
timestamp 1607639953
transform 1 0 48006 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_722
timestamp 1607639953
transform 1 0 48834 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_544
timestamp 1607639953
transform 1 0 51134 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_532
timestamp 1607639953
transform 1 0 50030 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_568
timestamp 1607639953
transform 1 0 53342 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_556
timestamp 1607639953
transform 1 0 52238 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_593
timestamp 1607639953
transform 1 0 55642 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_581
timestamp 1607639953
transform 1 0 54538 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_723
timestamp 1607639953
transform 1 0 54446 0 -1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_605
timestamp 1607639953
transform 1 0 56746 0 -1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_617
timestamp 1607639953
transform 1 0 57850 0 -1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1607639953
transform -1 0 58862 0 -1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_15
timestamp 1607639953
transform 1 0 2466 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_3
timestamp 1607639953
transform 1 0 1362 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1607639953
transform 1 0 1086 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_39
timestamp 1607639953
transform 1 0 4674 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_27
timestamp 1607639953
transform 1 0 3570 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_62
timestamp 1607639953
transform 1 0 6790 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_59
timestamp 1607639953
transform 1 0 6514 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_51_51
timestamp 1607639953
transform 1 0 5778 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_724
timestamp 1607639953
transform 1 0 6698 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_51_74
timestamp 1607639953
transform 1 0 7894 0 1 29920
box -38 -48 222 592
use XNOR2X1  XNOR2X1
timestamp 1608117647
transform 1 0 8078 0 1 29920
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_12  FILLER_51_102
timestamp 1607639953
transform 1 0 10470 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_90
timestamp 1607639953
transform 1 0 9366 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_131
timestamp 1607639953
transform 1 0 13138 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_123
timestamp 1607639953
transform 1 0 12402 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_51_114
timestamp 1607639953
transform 1 0 11574 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_725
timestamp 1607639953
transform 1 0 12310 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _010_
timestamp 1607639953
transform 1 0 13230 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_147
timestamp 1607639953
transform 1 0 14610 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_135
timestamp 1607639953
transform 1 0 13506 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_165
timestamp 1607639953
transform 1 0 16266 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_159
timestamp 1607639953
transform 1 0 15714 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _014_
timestamp 1607639953
transform 1 0 15990 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_196
timestamp 1607639953
transform 1 0 19118 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_184
timestamp 1607639953
transform 1 0 18014 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_177
timestamp 1607639953
transform 1 0 17370 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_726
timestamp 1607639953
transform 1 0 17922 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_220
timestamp 1607639953
transform 1 0 21326 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_208
timestamp 1607639953
transform 1 0 20222 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_232
timestamp 1607639953
transform 1 0 22430 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_257
timestamp 1607639953
transform 1 0 24730 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_245
timestamp 1607639953
transform 1 0 23626 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_727
timestamp 1607639953
transform 1 0 23534 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_281
timestamp 1607639953
transform 1 0 26938 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_269
timestamp 1607639953
transform 1 0 25834 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_306
timestamp 1607639953
transform 1 0 29238 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_293
timestamp 1607639953
transform 1 0 28042 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_728
timestamp 1607639953
transform 1 0 29146 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_330
timestamp 1607639953
transform 1 0 31446 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_51_318
timestamp 1607639953
transform 1 0 30342 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_343
timestamp 1607639953
transform 1 0 32642 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_338
timestamp 1607639953
transform 1 0 32182 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _208_
timestamp 1607639953
transform 1 0 32366 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_367
timestamp 1607639953
transform 1 0 34850 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_363
timestamp 1607639953
transform 1 0 34482 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_51_355
timestamp 1607639953
transform 1 0 33746 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_729
timestamp 1607639953
transform 1 0 34758 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_391
timestamp 1607639953
transform 1 0 37058 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_379
timestamp 1607639953
transform 1 0 35954 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_415
timestamp 1607639953
transform 1 0 39266 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_403
timestamp 1607639953
transform 1 0 38162 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_440
timestamp 1607639953
transform 1 0 41566 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_428
timestamp 1607639953
transform 1 0 40462 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_730
timestamp 1607639953
transform 1 0 40370 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_452
timestamp 1607639953
transform 1 0 42670 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_476
timestamp 1607639953
transform 1 0 44878 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_464
timestamp 1607639953
transform 1 0 43774 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_501
timestamp 1607639953
transform 1 0 47178 0 1 29920
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_51_489
timestamp 1607639953
transform 1 0 46074 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_731
timestamp 1607639953
transform 1 0 45982 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_525
timestamp 1607639953
transform 1 0 49386 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_513
timestamp 1607639953
transform 1 0 48282 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_509
timestamp 1607639953
transform 1 0 47914 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _083_
timestamp 1607639953
transform 1 0 48006 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_550
timestamp 1607639953
transform 1 0 51686 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_537
timestamp 1607639953
transform 1 0 50490 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_732
timestamp 1607639953
transform 1 0 51594 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_562
timestamp 1607639953
transform 1 0 52790 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_586
timestamp 1607639953
transform 1 0 54998 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_574
timestamp 1607639953
transform 1 0 53894 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_611
timestamp 1607639953
transform 1 0 57298 0 1 29920
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_608
timestamp 1607639953
transform 1 0 57022 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_51_604
timestamp 1607639953
transform 1 0 56654 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_598
timestamp 1607639953
transform 1 0 56102 0 1 29920
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_733
timestamp 1607639953
transform 1 0 57206 0 1 29920
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _201_
timestamp 1607639953
transform 1 0 56746 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_51_623
timestamp 1607639953
transform 1 0 58402 0 1 29920
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1607639953
transform -1 0 58862 0 1 29920
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_53_15
timestamp 1607639953
transform 1 0 2466 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_3
timestamp 1607639953
transform 1 0 1362 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_15
timestamp 1607639953
transform 1 0 2466 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_3
timestamp 1607639953
transform 1 0 1362 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1607639953
transform 1 0 1086 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1607639953
transform 1 0 1086 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_53_39
timestamp 1607639953
transform 1 0 4674 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_27
timestamp 1607639953
transform 1 0 3570 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_44
timestamp 1607639953
transform 1 0 5134 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_32
timestamp 1607639953
transform 1 0 4030 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_27
timestamp 1607639953
transform 1 0 3570 0 -1 31008
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_734
timestamp 1607639953
transform 1 0 3938 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_62
timestamp 1607639953
transform 1 0 6790 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_59
timestamp 1607639953
transform 1 0 6514 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_53_51
timestamp 1607639953
transform 1 0 5778 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_64
timestamp 1607639953
transform 1 0 6974 0 -1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_56
timestamp 1607639953
transform 1 0 6238 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_744
timestamp 1607639953
transform 1 0 6698 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _200_
timestamp 1607639953
transform 1 0 7158 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_53_74
timestamp 1607639953
transform 1 0 7894 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_81
timestamp 1607639953
transform 1 0 8538 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_52_69
timestamp 1607639953
transform 1 0 7434 0 -1 31008
box -38 -48 1142 592
use XOR2X1  XOR2X1
timestamp 1608117647
transform 1 0 8078 0 1 31008
box 0 -48 1288 592
use sky130_fd_sc_hd__decap_12  FILLER_53_102
timestamp 1607639953
transform 1 0 10470 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_90
timestamp 1607639953
transform 1 0 9366 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_105
timestamp 1607639953
transform 1 0 10746 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_93
timestamp 1607639953
transform 1 0 9642 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_89
timestamp 1607639953
transform 1 0 9274 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_735
timestamp 1607639953
transform 1 0 9550 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_123
timestamp 1607639953
transform 1 0 12402 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_114
timestamp 1607639953
transform 1 0 11574 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_52_129
timestamp 1607639953
transform 1 0 12954 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_117
timestamp 1607639953
transform 1 0 11850 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_745
timestamp 1607639953
transform 1 0 12310 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_147
timestamp 1607639953
transform 1 0 14610 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_135
timestamp 1607639953
transform 1 0 13506 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_154
timestamp 1607639953
transform 1 0 15254 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_141
timestamp 1607639953
transform 1 0 14058 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_736
timestamp 1607639953
transform 1 0 15162 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_171
timestamp 1607639953
transform 1 0 16818 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_159
timestamp 1607639953
transform 1 0 15714 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_166
timestamp 1607639953
transform 1 0 16358 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_196
timestamp 1607639953
transform 1 0 19118 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_184
timestamp 1607639953
transform 1 0 18014 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_190
timestamp 1607639953
transform 1 0 18566 0 -1 31008
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_52_178
timestamp 1607639953
transform 1 0 17462 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_746
timestamp 1607639953
transform 1 0 17922 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _047_
timestamp 1607639953
transform 1 0 19118 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_53_219
timestamp 1607639953
transform 1 0 21234 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_208
timestamp 1607639953
transform 1 0 20222 0 1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_52_215
timestamp 1607639953
transform 1 0 20866 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_211
timestamp 1607639953
transform 1 0 20498 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_52_203
timestamp 1607639953
transform 1 0 19762 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_199
timestamp 1607639953
transform 1 0 19394 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_737
timestamp 1607639953
transform 1 0 20774 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _130_
timestamp 1607639953
transform 1 0 20958 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _075_
timestamp 1607639953
transform 1 0 19486 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_53_231
timestamp 1607639953
transform 1 0 22338 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_239
timestamp 1607639953
transform 1 0 23074 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_227
timestamp 1607639953
transform 1 0 21970 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_257
timestamp 1607639953
transform 1 0 24730 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_245
timestamp 1607639953
transform 1 0 23626 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_243
timestamp 1607639953
transform 1 0 23442 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_263
timestamp 1607639953
transform 1 0 25282 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_251
timestamp 1607639953
transform 1 0 24178 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_747
timestamp 1607639953
transform 1 0 23534 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_281
timestamp 1607639953
transform 1 0 26938 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_269
timestamp 1607639953
transform 1 0 25834 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_276
timestamp 1607639953
transform 1 0 26478 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_738
timestamp 1607639953
transform 1 0 26386 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_306
timestamp 1607639953
transform 1 0 29238 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_293
timestamp 1607639953
transform 1 0 28042 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_300
timestamp 1607639953
transform 1 0 28686 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_288
timestamp 1607639953
transform 1 0 27582 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_748
timestamp 1607639953
transform 1 0 29146 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_330
timestamp 1607639953
transform 1 0 31446 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_318
timestamp 1607639953
transform 1 0 30342 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_324
timestamp 1607639953
transform 1 0 30894 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_312
timestamp 1607639953
transform 1 0 29790 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_342
timestamp 1607639953
transform 1 0 32550 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_349
timestamp 1607639953
transform 1 0 33194 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_337
timestamp 1607639953
transform 1 0 32090 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_739
timestamp 1607639953
transform 1 0 31998 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_367
timestamp 1607639953
transform 1 0 34850 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_354
timestamp 1607639953
transform 1 0 33654 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_373
timestamp 1607639953
transform 1 0 35402 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_361
timestamp 1607639953
transform 1 0 34298 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_749
timestamp 1607639953
transform 1 0 34758 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_391
timestamp 1607639953
transform 1 0 37058 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_379
timestamp 1607639953
transform 1 0 35954 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_385
timestamp 1607639953
transform 1 0 36506 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_415
timestamp 1607639953
transform 1 0 39266 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_403
timestamp 1607639953
transform 1 0 38162 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_410
timestamp 1607639953
transform 1 0 38806 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_398
timestamp 1607639953
transform 1 0 37702 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_740
timestamp 1607639953
transform 1 0 37610 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_440
timestamp 1607639953
transform 1 0 41566 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_428
timestamp 1607639953
transform 1 0 40462 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_434
timestamp 1607639953
transform 1 0 41014 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_422
timestamp 1607639953
transform 1 0 39910 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_750
timestamp 1607639953
transform 1 0 40370 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_452
timestamp 1607639953
transform 1 0 42670 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_459
timestamp 1607639953
transform 1 0 43314 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_446
timestamp 1607639953
transform 1 0 42118 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_741
timestamp 1607639953
transform 1 0 43222 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_476
timestamp 1607639953
transform 1 0 44878 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_464
timestamp 1607639953
transform 1 0 43774 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_483
timestamp 1607639953
transform 1 0 45522 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_471
timestamp 1607639953
transform 1 0 44418 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_501
timestamp 1607639953
transform 1 0 47178 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_489
timestamp 1607639953
transform 1 0 46074 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_495
timestamp 1607639953
transform 1 0 46626 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_751
timestamp 1607639953
transform 1 0 45982 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_525
timestamp 1607639953
transform 1 0 49386 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_513
timestamp 1607639953
transform 1 0 48282 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_520
timestamp 1607639953
transform 1 0 48926 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_507
timestamp 1607639953
transform 1 0 47730 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_742
timestamp 1607639953
transform 1 0 48834 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_550
timestamp 1607639953
transform 1 0 51686 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_537
timestamp 1607639953
transform 1 0 50490 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_544
timestamp 1607639953
transform 1 0 51134 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_532
timestamp 1607639953
transform 1 0 50030 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_752
timestamp 1607639953
transform 1 0 51594 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_562
timestamp 1607639953
transform 1 0 52790 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_568
timestamp 1607639953
transform 1 0 53342 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_556
timestamp 1607639953
transform 1 0 52238 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_586
timestamp 1607639953
transform 1 0 54998 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_574
timestamp 1607639953
transform 1 0 53894 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_593
timestamp 1607639953
transform 1 0 55642 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_581
timestamp 1607639953
transform 1 0 54538 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_743
timestamp 1607639953
transform 1 0 54446 0 -1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_611
timestamp 1607639953
transform 1 0 57298 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_598
timestamp 1607639953
transform 1 0 56102 0 1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_605
timestamp 1607639953
transform 1 0 56746 0 -1 31008
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_753
timestamp 1607639953
transform 1 0 57206 0 1 31008
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_53_623
timestamp 1607639953
transform 1 0 58402 0 1 31008
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_617
timestamp 1607639953
transform 1 0 57850 0 -1 31008
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1607639953
transform -1 0 58862 0 1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1607639953
transform -1 0 58862 0 -1 31008
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_15
timestamp 1607639953
transform 1 0 2466 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_3
timestamp 1607639953
transform 1 0 1362 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1607639953
transform 1 0 1086 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_44
timestamp 1607639953
transform 1 0 5134 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_40
timestamp 1607639953
transform 1 0 4766 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_32
timestamp 1607639953
transform 1 0 4030 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_54_27
timestamp 1607639953
transform 1 0 3570 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_754
timestamp 1607639953
transform 1 0 3938 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _131_
timestamp 1607639953
transform 1 0 4858 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_56
timestamp 1607639953
transform 1 0 6238 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_80
timestamp 1607639953
transform 1 0 8446 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_68
timestamp 1607639953
transform 1 0 7342 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_105
timestamp 1607639953
transform 1 0 10746 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_93
timestamp 1607639953
transform 1 0 9642 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_755
timestamp 1607639953
transform 1 0 9550 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_129
timestamp 1607639953
transform 1 0 12954 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_117
timestamp 1607639953
transform 1 0 11850 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_154
timestamp 1607639953
transform 1 0 15254 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_141
timestamp 1607639953
transform 1 0 14058 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_756
timestamp 1607639953
transform 1 0 15162 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_166
timestamp 1607639953
transform 1 0 16358 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_196
timestamp 1607639953
transform 1 0 19118 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_190
timestamp 1607639953
transform 1 0 18566 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_54_178
timestamp 1607639953
transform 1 0 17462 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _198_
timestamp 1607639953
transform 1 0 19210 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_54_215
timestamp 1607639953
transform 1 0 20866 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_212
timestamp 1607639953
transform 1 0 20590 0 -1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_54_200
timestamp 1607639953
transform 1 0 19486 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_757
timestamp 1607639953
transform 1 0 20774 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_239
timestamp 1607639953
transform 1 0 23074 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_227
timestamp 1607639953
transform 1 0 21970 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_223
timestamp 1607639953
transform 1 0 21602 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _026_
timestamp 1607639953
transform 1 0 21694 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_263
timestamp 1607639953
transform 1 0 25282 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_251
timestamp 1607639953
transform 1 0 24178 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_276
timestamp 1607639953
transform 1 0 26478 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_758
timestamp 1607639953
transform 1 0 26386 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_300
timestamp 1607639953
transform 1 0 28686 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_288
timestamp 1607639953
transform 1 0 27582 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_324
timestamp 1607639953
transform 1 0 30894 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_312
timestamp 1607639953
transform 1 0 29790 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_341
timestamp 1607639953
transform 1 0 32458 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_54_337
timestamp 1607639953
transform 1 0 32090 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_759
timestamp 1607639953
transform 1 0 31998 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _138_
timestamp 1607639953
transform 1 0 32182 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_365
timestamp 1607639953
transform 1 0 34666 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_353
timestamp 1607639953
transform 1 0 33562 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_393
timestamp 1607639953
transform 1 0 37242 0 -1 32096
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_389
timestamp 1607639953
transform 1 0 36874 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_377
timestamp 1607639953
transform 1 0 35770 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _196_
timestamp 1607639953
transform 1 0 36966 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_410
timestamp 1607639953
transform 1 0 38806 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_398
timestamp 1607639953
transform 1 0 37702 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_760
timestamp 1607639953
transform 1 0 37610 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_434
timestamp 1607639953
transform 1 0 41014 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_422
timestamp 1607639953
transform 1 0 39910 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_459
timestamp 1607639953
transform 1 0 43314 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_446
timestamp 1607639953
transform 1 0 42118 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_761
timestamp 1607639953
transform 1 0 43222 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_483
timestamp 1607639953
transform 1 0 45522 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_471
timestamp 1607639953
transform 1 0 44418 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_495
timestamp 1607639953
transform 1 0 46626 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_520
timestamp 1607639953
transform 1 0 48926 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_507
timestamp 1607639953
transform 1 0 47730 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_762
timestamp 1607639953
transform 1 0 48834 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_550
timestamp 1607639953
transform 1 0 51686 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_54_544
timestamp 1607639953
transform 1 0 51134 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_532
timestamp 1607639953
transform 1 0 50030 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _048_
timestamp 1607639953
transform 1 0 51410 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_562
timestamp 1607639953
transform 1 0 52790 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_593
timestamp 1607639953
transform 1 0 55642 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_581
timestamp 1607639953
transform 1 0 54538 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_574
timestamp 1607639953
transform 1 0 53894 0 -1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_763
timestamp 1607639953
transform 1 0 54446 0 -1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_605
timestamp 1607639953
transform 1 0 56746 0 -1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_617
timestamp 1607639953
transform 1 0 57850 0 -1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1607639953
transform -1 0 58862 0 -1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_55_15
timestamp 1607639953
transform 1 0 2466 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_3
timestamp 1607639953
transform 1 0 1362 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1607639953
transform 1 0 1086 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_55_39
timestamp 1607639953
transform 1 0 4674 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_27
timestamp 1607639953
transform 1 0 3570 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_62
timestamp 1607639953
transform 1 0 6790 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_59
timestamp 1607639953
transform 1 0 6514 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_55_51
timestamp 1607639953
transform 1 0 5778 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_764
timestamp 1607639953
transform 1 0 6698 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_86
timestamp 1607639953
transform 1 0 8998 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_74
timestamp 1607639953
transform 1 0 7894 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_102
timestamp 1607639953
transform 1 0 10470 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_98
timestamp 1607639953
transform 1 0 10102 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _098_
timestamp 1607639953
transform 1 0 10194 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_55_123
timestamp 1607639953
transform 1 0 12402 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_114
timestamp 1607639953
transform 1 0 11574 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_765
timestamp 1607639953
transform 1 0 12310 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_147
timestamp 1607639953
transform 1 0 14610 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_135
timestamp 1607639953
transform 1 0 13506 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_171
timestamp 1607639953
transform 1 0 16818 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_159
timestamp 1607639953
transform 1 0 15714 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_196
timestamp 1607639953
transform 1 0 19118 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_184
timestamp 1607639953
transform 1 0 18014 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_766
timestamp 1607639953
transform 1 0 17922 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_220
timestamp 1607639953
transform 1 0 21326 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_208
timestamp 1607639953
transform 1 0 20222 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_232
timestamp 1607639953
transform 1 0 22430 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_257
timestamp 1607639953
transform 1 0 24730 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_245
timestamp 1607639953
transform 1 0 23626 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_767
timestamp 1607639953
transform 1 0 23534 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_281
timestamp 1607639953
transform 1 0 26938 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_269
timestamp 1607639953
transform 1 0 25834 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_306
timestamp 1607639953
transform 1 0 29238 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_293
timestamp 1607639953
transform 1 0 28042 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_768
timestamp 1607639953
transform 1 0 29146 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_330
timestamp 1607639953
transform 1 0 31446 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_318
timestamp 1607639953
transform 1 0 30342 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_342
timestamp 1607639953
transform 1 0 32550 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_367
timestamp 1607639953
transform 1 0 34850 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_354
timestamp 1607639953
transform 1 0 33654 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_769
timestamp 1607639953
transform 1 0 34758 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_391
timestamp 1607639953
transform 1 0 37058 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_379
timestamp 1607639953
transform 1 0 35954 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_415
timestamp 1607639953
transform 1 0 39266 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_403
timestamp 1607639953
transform 1 0 38162 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_440
timestamp 1607639953
transform 1 0 41566 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_428
timestamp 1607639953
transform 1 0 40462 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_770
timestamp 1607639953
transform 1 0 40370 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_452
timestamp 1607639953
transform 1 0 42670 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_476
timestamp 1607639953
transform 1 0 44878 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_464
timestamp 1607639953
transform 1 0 43774 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_501
timestamp 1607639953
transform 1 0 47178 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_489
timestamp 1607639953
transform 1 0 46074 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_771
timestamp 1607639953
transform 1 0 45982 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_525
timestamp 1607639953
transform 1 0 49386 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_513
timestamp 1607639953
transform 1 0 48282 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_550
timestamp 1607639953
transform 1 0 51686 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_548
timestamp 1607639953
transform 1 0 51502 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_542
timestamp 1607639953
transform 1 0 50950 0 1 32096
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_55_537
timestamp 1607639953
transform 1 0 50490 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_772
timestamp 1607639953
transform 1 0 51594 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _158_
timestamp 1607639953
transform 1 0 50674 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_55_566
timestamp 1607639953
transform 1 0 53158 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_562
timestamp 1607639953
transform 1 0 52790 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _118_
timestamp 1607639953
transform 1 0 52882 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_55_590
timestamp 1607639953
transform 1 0 55366 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_578
timestamp 1607639953
transform 1 0 54262 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_611
timestamp 1607639953
transform 1 0 57298 0 1 32096
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_602
timestamp 1607639953
transform 1 0 56470 0 1 32096
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_773
timestamp 1607639953
transform 1 0 57206 0 1 32096
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_55_623
timestamp 1607639953
transform 1 0 58402 0 1 32096
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1607639953
transform -1 0 58862 0 1 32096
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_15
timestamp 1607639953
transform 1 0 2466 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_3
timestamp 1607639953
transform 1 0 1362 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1607639953
transform 1 0 1086 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_44
timestamp 1607639953
transform 1 0 5134 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_32
timestamp 1607639953
transform 1 0 4030 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_27
timestamp 1607639953
transform 1 0 3570 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_774
timestamp 1607639953
transform 1 0 3938 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_56
timestamp 1607639953
transform 1 0 6238 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_80
timestamp 1607639953
transform 1 0 8446 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_68
timestamp 1607639953
transform 1 0 7342 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_105
timestamp 1607639953
transform 1 0 10746 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_93
timestamp 1607639953
transform 1 0 9642 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_775
timestamp 1607639953
transform 1 0 9550 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_124
timestamp 1607639953
transform 1 0 12494 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_117
timestamp 1607639953
transform 1 0 11850 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _160_
timestamp 1607639953
transform 1 0 12218 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_154
timestamp 1607639953
transform 1 0 15254 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_56_152
timestamp 1607639953
transform 1 0 15070 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_148
timestamp 1607639953
transform 1 0 14702 0 -1 33184
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_136
timestamp 1607639953
transform 1 0 13598 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_776
timestamp 1607639953
transform 1 0 15162 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_166
timestamp 1607639953
transform 1 0 16358 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_190
timestamp 1607639953
transform 1 0 18566 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_178
timestamp 1607639953
transform 1 0 17462 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_215
timestamp 1607639953
transform 1 0 20866 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_202
timestamp 1607639953
transform 1 0 19670 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_777
timestamp 1607639953
transform 1 0 20774 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_239
timestamp 1607639953
transform 1 0 23074 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_227
timestamp 1607639953
transform 1 0 21970 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_263
timestamp 1607639953
transform 1 0 25282 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_251
timestamp 1607639953
transform 1 0 24178 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_276
timestamp 1607639953
transform 1 0 26478 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_778
timestamp 1607639953
transform 1 0 26386 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_300
timestamp 1607639953
transform 1 0 28686 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_288
timestamp 1607639953
transform 1 0 27582 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_324
timestamp 1607639953
transform 1 0 30894 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_312
timestamp 1607639953
transform 1 0 29790 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_349
timestamp 1607639953
transform 1 0 33194 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_337
timestamp 1607639953
transform 1 0 32090 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_779
timestamp 1607639953
transform 1 0 31998 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_373
timestamp 1607639953
transform 1 0 35402 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_361
timestamp 1607639953
transform 1 0 34298 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_385
timestamp 1607639953
transform 1 0 36506 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_410
timestamp 1607639953
transform 1 0 38806 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_398
timestamp 1607639953
transform 1 0 37702 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_780
timestamp 1607639953
transform 1 0 37610 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_434
timestamp 1607639953
transform 1 0 41014 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_422
timestamp 1607639953
transform 1 0 39910 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_459
timestamp 1607639953
transform 1 0 43314 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_446
timestamp 1607639953
transform 1 0 42118 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_781
timestamp 1607639953
transform 1 0 43222 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_483
timestamp 1607639953
transform 1 0 45522 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_471
timestamp 1607639953
transform 1 0 44418 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_495
timestamp 1607639953
transform 1 0 46626 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_520
timestamp 1607639953
transform 1 0 48926 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_507
timestamp 1607639953
transform 1 0 47730 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_782
timestamp 1607639953
transform 1 0 48834 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_544
timestamp 1607639953
transform 1 0 51134 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_532
timestamp 1607639953
transform 1 0 50030 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_568
timestamp 1607639953
transform 1 0 53342 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_556
timestamp 1607639953
transform 1 0 52238 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_593
timestamp 1607639953
transform 1 0 55642 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_581
timestamp 1607639953
transform 1 0 54538 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_783
timestamp 1607639953
transform 1 0 54446 0 -1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_605
timestamp 1607639953
transform 1 0 56746 0 -1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_617
timestamp 1607639953
transform 1 0 57850 0 -1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1607639953
transform -1 0 58862 0 -1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_57_15
timestamp 1607639953
transform 1 0 2466 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_3
timestamp 1607639953
transform 1 0 1362 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1607639953
transform 1 0 1086 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_57_39
timestamp 1607639953
transform 1 0 4674 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_27
timestamp 1607639953
transform 1 0 3570 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_62
timestamp 1607639953
transform 1 0 6790 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_60
timestamp 1607639953
transform 1 0 6606 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_51
timestamp 1607639953
transform 1 0 5778 0 1 33184
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_784
timestamp 1607639953
transform 1 0 6698 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _025_
timestamp 1607639953
transform 1 0 6330 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_57_86
timestamp 1607639953
transform 1 0 8998 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_74
timestamp 1607639953
transform 1 0 7894 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_110
timestamp 1607639953
transform 1 0 11206 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_98
timestamp 1607639953
transform 1 0 10102 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_123
timestamp 1607639953
transform 1 0 12402 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_785
timestamp 1607639953
transform 1 0 12310 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_147
timestamp 1607639953
transform 1 0 14610 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_135
timestamp 1607639953
transform 1 0 13506 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_171
timestamp 1607639953
transform 1 0 16818 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_159
timestamp 1607639953
transform 1 0 15714 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_196
timestamp 1607639953
transform 1 0 19118 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_184
timestamp 1607639953
transform 1 0 18014 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_786
timestamp 1607639953
transform 1 0 17922 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_220
timestamp 1607639953
transform 1 0 21326 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_208
timestamp 1607639953
transform 1 0 20222 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_232
timestamp 1607639953
transform 1 0 22430 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_257
timestamp 1607639953
transform 1 0 24730 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_245
timestamp 1607639953
transform 1 0 23626 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_787
timestamp 1607639953
transform 1 0 23534 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_281
timestamp 1607639953
transform 1 0 26938 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_269
timestamp 1607639953
transform 1 0 25834 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_306
timestamp 1607639953
transform 1 0 29238 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_293
timestamp 1607639953
transform 1 0 28042 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_788
timestamp 1607639953
transform 1 0 29146 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_330
timestamp 1607639953
transform 1 0 31446 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_318
timestamp 1607639953
transform 1 0 30342 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_342
timestamp 1607639953
transform 1 0 32550 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_367
timestamp 1607639953
transform 1 0 34850 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_354
timestamp 1607639953
transform 1 0 33654 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_789
timestamp 1607639953
transform 1 0 34758 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_391
timestamp 1607639953
transform 1 0 37058 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_379
timestamp 1607639953
transform 1 0 35954 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_415
timestamp 1607639953
transform 1 0 39266 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_403
timestamp 1607639953
transform 1 0 38162 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_440
timestamp 1607639953
transform 1 0 41566 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_428
timestamp 1607639953
transform 1 0 40462 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_790
timestamp 1607639953
transform 1 0 40370 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_452
timestamp 1607639953
transform 1 0 42670 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_476
timestamp 1607639953
transform 1 0 44878 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_464
timestamp 1607639953
transform 1 0 43774 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_504
timestamp 1607639953
transform 1 0 47454 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_492
timestamp 1607639953
transform 1 0 46350 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_791
timestamp 1607639953
transform 1 0 45982 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _177_
timestamp 1607639953
transform 1 0 46074 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_57_528
timestamp 1607639953
transform 1 0 49662 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_516
timestamp 1607639953
transform 1 0 48558 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_550
timestamp 1607639953
transform 1 0 51686 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_57_548
timestamp 1607639953
transform 1 0 51502 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_540
timestamp 1607639953
transform 1 0 50766 0 1 33184
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_792
timestamp 1607639953
transform 1 0 51594 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_562
timestamp 1607639953
transform 1 0 52790 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_586
timestamp 1607639953
transform 1 0 54998 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_574
timestamp 1607639953
transform 1 0 53894 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_611
timestamp 1607639953
transform 1 0 57298 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_598
timestamp 1607639953
transform 1 0 56102 0 1 33184
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_793
timestamp 1607639953
transform 1 0 57206 0 1 33184
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_623
timestamp 1607639953
transform 1 0 58402 0 1 33184
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1607639953
transform -1 0 58862 0 1 33184
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_58_15
timestamp 1607639953
transform 1 0 2466 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_3
timestamp 1607639953
transform 1 0 1362 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1607639953
transform 1 0 1086 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_58_44
timestamp 1607639953
transform 1 0 5134 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_32
timestamp 1607639953
transform 1 0 4030 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_27
timestamp 1607639953
transform 1 0 3570 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_794
timestamp 1607639953
transform 1 0 3938 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_56
timestamp 1607639953
transform 1 0 6238 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_80
timestamp 1607639953
transform 1 0 8446 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_68
timestamp 1607639953
transform 1 0 7342 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_105
timestamp 1607639953
transform 1 0 10746 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_93
timestamp 1607639953
transform 1 0 9642 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_795
timestamp 1607639953
transform 1 0 9550 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_129
timestamp 1607639953
transform 1 0 12954 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_117
timestamp 1607639953
transform 1 0 11850 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_154
timestamp 1607639953
transform 1 0 15254 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_141
timestamp 1607639953
transform 1 0 14058 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_796
timestamp 1607639953
transform 1 0 15162 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_166
timestamp 1607639953
transform 1 0 16358 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_190
timestamp 1607639953
transform 1 0 18566 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_178
timestamp 1607639953
transform 1 0 17462 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_215
timestamp 1607639953
transform 1 0 20866 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_202
timestamp 1607639953
transform 1 0 19670 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_797
timestamp 1607639953
transform 1 0 20774 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_239
timestamp 1607639953
transform 1 0 23074 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_227
timestamp 1607639953
transform 1 0 21970 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_263
timestamp 1607639953
transform 1 0 25282 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_251
timestamp 1607639953
transform 1 0 24178 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_276
timestamp 1607639953
transform 1 0 26478 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_798
timestamp 1607639953
transform 1 0 26386 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_300
timestamp 1607639953
transform 1 0 28686 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_288
timestamp 1607639953
transform 1 0 27582 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_324
timestamp 1607639953
transform 1 0 30894 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_312
timestamp 1607639953
transform 1 0 29790 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_349
timestamp 1607639953
transform 1 0 33194 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_337
timestamp 1607639953
transform 1 0 32090 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_799
timestamp 1607639953
transform 1 0 31998 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_373
timestamp 1607639953
transform 1 0 35402 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_58_361
timestamp 1607639953
transform 1 0 34298 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_58_394
timestamp 1607639953
transform 1 0 37334 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_58_386
timestamp 1607639953
transform 1 0 36598 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_381
timestamp 1607639953
transform 1 0 36138 0 -1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _074_
timestamp 1607639953
transform 1 0 36322 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_58_410
timestamp 1607639953
transform 1 0 38806 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_398
timestamp 1607639953
transform 1 0 37702 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_800
timestamp 1607639953
transform 1 0 37610 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_434
timestamp 1607639953
transform 1 0 41014 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_422
timestamp 1607639953
transform 1 0 39910 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_459
timestamp 1607639953
transform 1 0 43314 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_446
timestamp 1607639953
transform 1 0 42118 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_801
timestamp 1607639953
transform 1 0 43222 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _104_
timestamp 1607639953
transform 1 0 43406 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_58_475
timestamp 1607639953
transform 1 0 44786 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_463
timestamp 1607639953
transform 1 0 43682 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_499
timestamp 1607639953
transform 1 0 46994 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_487
timestamp 1607639953
transform 1 0 45890 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_520
timestamp 1607639953
transform 1 0 48926 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_511
timestamp 1607639953
transform 1 0 48098 0 -1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_802
timestamp 1607639953
transform 1 0 48834 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_544
timestamp 1607639953
transform 1 0 51134 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_532
timestamp 1607639953
transform 1 0 50030 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_568
timestamp 1607639953
transform 1 0 53342 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_556
timestamp 1607639953
transform 1 0 52238 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_593
timestamp 1607639953
transform 1 0 55642 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_581
timestamp 1607639953
transform 1 0 54538 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_803
timestamp 1607639953
transform 1 0 54446 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_605
timestamp 1607639953
transform 1 0 56746 0 -1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_624
timestamp 1607639953
transform 1 0 58494 0 -1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_617
timestamp 1607639953
transform 1 0 57850 0 -1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1607639953
transform -1 0 58862 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _097_
timestamp 1607639953
transform 1 0 58218 0 -1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_60_15
timestamp 1607639953
transform 1 0 2466 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_3
timestamp 1607639953
transform 1 0 1362 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_15
timestamp 1607639953
transform 1 0 2466 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_3
timestamp 1607639953
transform 1 0 1362 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1607639953
transform 1 0 1086 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1607639953
transform 1 0 1086 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_60_44
timestamp 1607639953
transform 1 0 5134 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_32
timestamp 1607639953
transform 1 0 4030 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_27
timestamp 1607639953
transform 1 0 3570 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_39
timestamp 1607639953
transform 1 0 4674 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_27
timestamp 1607639953
transform 1 0 3570 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_814
timestamp 1607639953
transform 1 0 3938 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_56
timestamp 1607639953
transform 1 0 6238 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_62
timestamp 1607639953
transform 1 0 6790 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_59
timestamp 1607639953
transform 1 0 6514 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_59_51
timestamp 1607639953
transform 1 0 5778 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_804
timestamp 1607639953
transform 1 0 6698 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_80
timestamp 1607639953
transform 1 0 8446 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_68
timestamp 1607639953
transform 1 0 7342 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_86
timestamp 1607639953
transform 1 0 8998 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_74
timestamp 1607639953
transform 1 0 7894 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_105
timestamp 1607639953
transform 1 0 10746 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_93
timestamp 1607639953
transform 1 0 9642 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_110
timestamp 1607639953
transform 1 0 11206 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_98
timestamp 1607639953
transform 1 0 10102 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_815
timestamp 1607639953
transform 1 0 9550 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_129
timestamp 1607639953
transform 1 0 12954 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_117
timestamp 1607639953
transform 1 0 11850 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_123
timestamp 1607639953
transform 1 0 12402 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_805
timestamp 1607639953
transform 1 0 12310 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_154
timestamp 1607639953
transform 1 0 15254 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_141
timestamp 1607639953
transform 1 0 14058 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_147
timestamp 1607639953
transform 1 0 14610 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_135
timestamp 1607639953
transform 1 0 13506 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_816
timestamp 1607639953
transform 1 0 15162 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_166
timestamp 1607639953
transform 1 0 16358 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_171
timestamp 1607639953
transform 1 0 16818 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_159
timestamp 1607639953
transform 1 0 15714 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_190
timestamp 1607639953
transform 1 0 18566 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_178
timestamp 1607639953
transform 1 0 17462 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_196
timestamp 1607639953
transform 1 0 19118 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_184
timestamp 1607639953
transform 1 0 18014 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_806
timestamp 1607639953
transform 1 0 17922 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_215
timestamp 1607639953
transform 1 0 20866 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_202
timestamp 1607639953
transform 1 0 19670 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_215
timestamp 1607639953
transform 1 0 20866 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_208
timestamp 1607639953
transform 1 0 20222 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_817
timestamp 1607639953
transform 1 0 20774 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _030_
timestamp 1607639953
transform 1 0 20590 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_60_239
timestamp 1607639953
transform 1 0 23074 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_227
timestamp 1607639953
transform 1 0 21970 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_239
timestamp 1607639953
transform 1 0 23074 0 1 34272
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_227
timestamp 1607639953
transform 1 0 21970 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_263
timestamp 1607639953
transform 1 0 25282 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_251
timestamp 1607639953
transform 1 0 24178 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_257
timestamp 1607639953
transform 1 0 24730 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_245
timestamp 1607639953
transform 1 0 23626 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_243
timestamp 1607639953
transform 1 0 23442 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_807
timestamp 1607639953
transform 1 0 23534 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_276
timestamp 1607639953
transform 1 0 26478 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_281
timestamp 1607639953
transform 1 0 26938 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_269
timestamp 1607639953
transform 1 0 25834 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_818
timestamp 1607639953
transform 1 0 26386 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_300
timestamp 1607639953
transform 1 0 28686 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_288
timestamp 1607639953
transform 1 0 27582 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_306
timestamp 1607639953
transform 1 0 29238 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_293
timestamp 1607639953
transform 1 0 28042 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_808
timestamp 1607639953
transform 1 0 29146 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_322
timestamp 1607639953
transform 1 0 30710 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_318
timestamp 1607639953
transform 1 0 30342 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_60_312
timestamp 1607639953
transform 1 0 29790 0 -1 35360
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_59_330
timestamp 1607639953
transform 1 0 31446 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_318
timestamp 1607639953
transform 1 0 30342 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _034_
timestamp 1607639953
transform 1 0 30434 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_60_349
timestamp 1607639953
transform 1 0 33194 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_337
timestamp 1607639953
transform 1 0 32090 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_334
timestamp 1607639953
transform 1 0 31814 0 -1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_59_342
timestamp 1607639953
transform 1 0 32550 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_819
timestamp 1607639953
transform 1 0 31998 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_373
timestamp 1607639953
transform 1 0 35402 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_361
timestamp 1607639953
transform 1 0 34298 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_367
timestamp 1607639953
transform 1 0 34850 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_354
timestamp 1607639953
transform 1 0 33654 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_809
timestamp 1607639953
transform 1 0 34758 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_385
timestamp 1607639953
transform 1 0 36506 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_391
timestamp 1607639953
transform 1 0 37058 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_379
timestamp 1607639953
transform 1 0 35954 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_410
timestamp 1607639953
transform 1 0 38806 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_398
timestamp 1607639953
transform 1 0 37702 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_415
timestamp 1607639953
transform 1 0 39266 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_403
timestamp 1607639953
transform 1 0 38162 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_820
timestamp 1607639953
transform 1 0 37610 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_434
timestamp 1607639953
transform 1 0 41014 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_422
timestamp 1607639953
transform 1 0 39910 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_440
timestamp 1607639953
transform 1 0 41566 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_428
timestamp 1607639953
transform 1 0 40462 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_810
timestamp 1607639953
transform 1 0 40370 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_459
timestamp 1607639953
transform 1 0 43314 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_446
timestamp 1607639953
transform 1 0 42118 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_452
timestamp 1607639953
transform 1 0 42670 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_821
timestamp 1607639953
transform 1 0 43222 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_483
timestamp 1607639953
transform 1 0 45522 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_471
timestamp 1607639953
transform 1 0 44418 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_476
timestamp 1607639953
transform 1 0 44878 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_464
timestamp 1607639953
transform 1 0 43774 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_495
timestamp 1607639953
transform 1 0 46626 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_501
timestamp 1607639953
transform 1 0 47178 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_489
timestamp 1607639953
transform 1 0 46074 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_811
timestamp 1607639953
transform 1 0 45982 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_520
timestamp 1607639953
transform 1 0 48926 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_507
timestamp 1607639953
transform 1 0 47730 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_525
timestamp 1607639953
transform 1 0 49386 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_513
timestamp 1607639953
transform 1 0 48282 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_822
timestamp 1607639953
transform 1 0 48834 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_544
timestamp 1607639953
transform 1 0 51134 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_532
timestamp 1607639953
transform 1 0 50030 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_550
timestamp 1607639953
transform 1 0 51686 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_541
timestamp 1607639953
transform 1 0 50858 0 1 34272
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_537
timestamp 1607639953
transform 1 0 50490 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_812
timestamp 1607639953
transform 1 0 51594 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _197_
timestamp 1607639953
transform 1 0 50582 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_60_564
timestamp 1607639953
transform 1 0 52974 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_560
timestamp 1607639953
transform 1 0 52606 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_556
timestamp 1607639953
transform 1 0 52238 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_562
timestamp 1607639953
transform 1 0 52790 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _176_
timestamp 1607639953
transform 1 0 52698 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_60_593
timestamp 1607639953
transform 1 0 55642 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_581
timestamp 1607639953
transform 1 0 54538 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_576
timestamp 1607639953
transform 1 0 54078 0 -1 35360
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_586
timestamp 1607639953
transform 1 0 54998 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_574
timestamp 1607639953
transform 1 0 53894 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_823
timestamp 1607639953
transform 1 0 54446 0 -1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_605
timestamp 1607639953
transform 1 0 56746 0 -1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_611
timestamp 1607639953
transform 1 0 57298 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_598
timestamp 1607639953
transform 1 0 56102 0 1 34272
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_813
timestamp 1607639953
transform 1 0 57206 0 1 34272
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_617
timestamp 1607639953
transform 1 0 57850 0 -1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_623
timestamp 1607639953
transform 1 0 58402 0 1 34272
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1607639953
transform -1 0 58862 0 -1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1607639953
transform -1 0 58862 0 1 34272
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_61_15
timestamp 1607639953
transform 1 0 2466 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_3
timestamp 1607639953
transform 1 0 1362 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1607639953
transform 1 0 1086 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_61_39
timestamp 1607639953
transform 1 0 4674 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_27
timestamp 1607639953
transform 1 0 3570 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_62
timestamp 1607639953
transform 1 0 6790 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_59
timestamp 1607639953
transform 1 0 6514 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_61_51
timestamp 1607639953
transform 1 0 5778 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_824
timestamp 1607639953
transform 1 0 6698 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_86
timestamp 1607639953
transform 1 0 8998 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_74
timestamp 1607639953
transform 1 0 7894 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_110
timestamp 1607639953
transform 1 0 11206 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_98
timestamp 1607639953
transform 1 0 10102 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_123
timestamp 1607639953
transform 1 0 12402 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_825
timestamp 1607639953
transform 1 0 12310 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_147
timestamp 1607639953
transform 1 0 14610 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_135
timestamp 1607639953
transform 1 0 13506 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_171
timestamp 1607639953
transform 1 0 16818 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_159
timestamp 1607639953
transform 1 0 15714 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_196
timestamp 1607639953
transform 1 0 19118 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_184
timestamp 1607639953
transform 1 0 18014 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_826
timestamp 1607639953
transform 1 0 17922 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_220
timestamp 1607639953
transform 1 0 21326 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_208
timestamp 1607639953
transform 1 0 20222 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_232
timestamp 1607639953
transform 1 0 22430 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_257
timestamp 1607639953
transform 1 0 24730 0 1 35360
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_61_245
timestamp 1607639953
transform 1 0 23626 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_827
timestamp 1607639953
transform 1 0 23534 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_281
timestamp 1607639953
transform 1 0 26938 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_269
timestamp 1607639953
transform 1 0 25834 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_265
timestamp 1607639953
transform 1 0 25466 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _040_
timestamp 1607639953
transform 1 0 25558 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_61_306
timestamp 1607639953
transform 1 0 29238 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_293
timestamp 1607639953
transform 1 0 28042 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_828
timestamp 1607639953
transform 1 0 29146 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_330
timestamp 1607639953
transform 1 0 31446 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_318
timestamp 1607639953
transform 1 0 30342 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_342
timestamp 1607639953
transform 1 0 32550 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_367
timestamp 1607639953
transform 1 0 34850 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_354
timestamp 1607639953
transform 1 0 33654 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_829
timestamp 1607639953
transform 1 0 34758 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_391
timestamp 1607639953
transform 1 0 37058 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_379
timestamp 1607639953
transform 1 0 35954 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_415
timestamp 1607639953
transform 1 0 39266 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_403
timestamp 1607639953
transform 1 0 38162 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_440
timestamp 1607639953
transform 1 0 41566 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_428
timestamp 1607639953
transform 1 0 40462 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_830
timestamp 1607639953
transform 1 0 40370 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_452
timestamp 1607639953
transform 1 0 42670 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_476
timestamp 1607639953
transform 1 0 44878 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_464
timestamp 1607639953
transform 1 0 43774 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_501
timestamp 1607639953
transform 1 0 47178 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_489
timestamp 1607639953
transform 1 0 46074 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_831
timestamp 1607639953
transform 1 0 45982 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_525
timestamp 1607639953
transform 1 0 49386 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_513
timestamp 1607639953
transform 1 0 48282 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_550
timestamp 1607639953
transform 1 0 51686 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_537
timestamp 1607639953
transform 1 0 50490 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_832
timestamp 1607639953
transform 1 0 51594 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_562
timestamp 1607639953
transform 1 0 52790 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_586
timestamp 1607639953
transform 1 0 54998 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_574
timestamp 1607639953
transform 1 0 53894 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_611
timestamp 1607639953
transform 1 0 57298 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_598
timestamp 1607639953
transform 1 0 56102 0 1 35360
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_833
timestamp 1607639953
transform 1 0 57206 0 1 35360
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_623
timestamp 1607639953
transform 1 0 58402 0 1 35360
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1607639953
transform -1 0 58862 0 1 35360
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_15
timestamp 1607639953
transform 1 0 2466 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_3
timestamp 1607639953
transform 1 0 1362 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1607639953
transform 1 0 1086 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_44
timestamp 1607639953
transform 1 0 5134 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_32
timestamp 1607639953
transform 1 0 4030 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_27
timestamp 1607639953
transform 1 0 3570 0 -1 36448
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_834
timestamp 1607639953
transform 1 0 3938 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_56
timestamp 1607639953
transform 1 0 6238 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_80
timestamp 1607639953
transform 1 0 8446 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_68
timestamp 1607639953
transform 1 0 7342 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_105
timestamp 1607639953
transform 1 0 10746 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_93
timestamp 1607639953
transform 1 0 9642 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_835
timestamp 1607639953
transform 1 0 9550 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_129
timestamp 1607639953
transform 1 0 12954 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_117
timestamp 1607639953
transform 1 0 11850 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_154
timestamp 1607639953
transform 1 0 15254 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_141
timestamp 1607639953
transform 1 0 14058 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_836
timestamp 1607639953
transform 1 0 15162 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_166
timestamp 1607639953
transform 1 0 16358 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_190
timestamp 1607639953
transform 1 0 18566 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_178
timestamp 1607639953
transform 1 0 17462 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_215
timestamp 1607639953
transform 1 0 20866 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_202
timestamp 1607639953
transform 1 0 19670 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_837
timestamp 1607639953
transform 1 0 20774 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_239
timestamp 1607639953
transform 1 0 23074 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_227
timestamp 1607639953
transform 1 0 21970 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_263
timestamp 1607639953
transform 1 0 25282 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_251
timestamp 1607639953
transform 1 0 24178 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_276
timestamp 1607639953
transform 1 0 26478 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_838
timestamp 1607639953
transform 1 0 26386 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_300
timestamp 1607639953
transform 1 0 28686 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_288
timestamp 1607639953
transform 1 0 27582 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_324
timestamp 1607639953
transform 1 0 30894 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_312
timestamp 1607639953
transform 1 0 29790 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_349
timestamp 1607639953
transform 1 0 33194 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_337
timestamp 1607639953
transform 1 0 32090 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_839
timestamp 1607639953
transform 1 0 31998 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_373
timestamp 1607639953
transform 1 0 35402 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_361
timestamp 1607639953
transform 1 0 34298 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_385
timestamp 1607639953
transform 1 0 36506 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_410
timestamp 1607639953
transform 1 0 38806 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_398
timestamp 1607639953
transform 1 0 37702 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_840
timestamp 1607639953
transform 1 0 37610 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_434
timestamp 1607639953
transform 1 0 41014 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_422
timestamp 1607639953
transform 1 0 39910 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_459
timestamp 1607639953
transform 1 0 43314 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_446
timestamp 1607639953
transform 1 0 42118 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_841
timestamp 1607639953
transform 1 0 43222 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_62_479
timestamp 1607639953
transform 1 0 45154 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_62_471
timestamp 1607639953
transform 1 0 44418 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _204_
timestamp 1607639953
transform 1 0 45430 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_497
timestamp 1607639953
transform 1 0 46810 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_485
timestamp 1607639953
transform 1 0 45706 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_520
timestamp 1607639953
transform 1 0 48926 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_517
timestamp 1607639953
transform 1 0 48650 0 -1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_62_509
timestamp 1607639953
transform 1 0 47914 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_842
timestamp 1607639953
transform 1 0 48834 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_544
timestamp 1607639953
transform 1 0 51134 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_532
timestamp 1607639953
transform 1 0 50030 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_568
timestamp 1607639953
transform 1 0 53342 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_556
timestamp 1607639953
transform 1 0 52238 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_593
timestamp 1607639953
transform 1 0 55642 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_581
timestamp 1607639953
transform 1 0 54538 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_843
timestamp 1607639953
transform 1 0 54446 0 -1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_605
timestamp 1607639953
transform 1 0 56746 0 -1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_617
timestamp 1607639953
transform 1 0 57850 0 -1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1607639953
transform -1 0 58862 0 -1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_15
timestamp 1607639953
transform 1 0 2466 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_3
timestamp 1607639953
transform 1 0 1362 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1607639953
transform 1 0 1086 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_39
timestamp 1607639953
transform 1 0 4674 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_27
timestamp 1607639953
transform 1 0 3570 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_62
timestamp 1607639953
transform 1 0 6790 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_63_59
timestamp 1607639953
transform 1 0 6514 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_51
timestamp 1607639953
transform 1 0 5778 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_844
timestamp 1607639953
transform 1 0 6698 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_86
timestamp 1607639953
transform 1 0 8998 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_74
timestamp 1607639953
transform 1 0 7894 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_110
timestamp 1607639953
transform 1 0 11206 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_98
timestamp 1607639953
transform 1 0 10102 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_123
timestamp 1607639953
transform 1 0 12402 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_845
timestamp 1607639953
transform 1 0 12310 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_147
timestamp 1607639953
transform 1 0 14610 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_135
timestamp 1607639953
transform 1 0 13506 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_171
timestamp 1607639953
transform 1 0 16818 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_159
timestamp 1607639953
transform 1 0 15714 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_196
timestamp 1607639953
transform 1 0 19118 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_184
timestamp 1607639953
transform 1 0 18014 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_846
timestamp 1607639953
transform 1 0 17922 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_220
timestamp 1607639953
transform 1 0 21326 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_208
timestamp 1607639953
transform 1 0 20222 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_232
timestamp 1607639953
transform 1 0 22430 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_257
timestamp 1607639953
transform 1 0 24730 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_245
timestamp 1607639953
transform 1 0 23626 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_847
timestamp 1607639953
transform 1 0 23534 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_281
timestamp 1607639953
transform 1 0 26938 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_269
timestamp 1607639953
transform 1 0 25834 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_306
timestamp 1607639953
transform 1 0 29238 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_293
timestamp 1607639953
transform 1 0 28042 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_848
timestamp 1607639953
transform 1 0 29146 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_318
timestamp 1607639953
transform 1 0 30342 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _162_
timestamp 1607639953
transform 1 0 31446 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_345
timestamp 1607639953
transform 1 0 32826 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_333
timestamp 1607639953
transform 1 0 31722 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_367
timestamp 1607639953
transform 1 0 34850 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_365
timestamp 1607639953
transform 1 0 34666 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_357
timestamp 1607639953
transform 1 0 33930 0 1 36448
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_849
timestamp 1607639953
transform 1 0 34758 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_391
timestamp 1607639953
transform 1 0 37058 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_379
timestamp 1607639953
transform 1 0 35954 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_415
timestamp 1607639953
transform 1 0 39266 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_403
timestamp 1607639953
transform 1 0 38162 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_440
timestamp 1607639953
transform 1 0 41566 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_428
timestamp 1607639953
transform 1 0 40462 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_850
timestamp 1607639953
transform 1 0 40370 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_452
timestamp 1607639953
transform 1 0 42670 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_481
timestamp 1607639953
transform 1 0 45338 0 1 36448
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_63_476
timestamp 1607639953
transform 1 0 44878 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_63_464
timestamp 1607639953
transform 1 0 43774 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _110_
timestamp 1607639953
transform 1 0 45062 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_501
timestamp 1607639953
transform 1 0 47178 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_489
timestamp 1607639953
transform 1 0 46074 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_487
timestamp 1607639953
transform 1 0 45890 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_851
timestamp 1607639953
transform 1 0 45982 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_525
timestamp 1607639953
transform 1 0 49386 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_513
timestamp 1607639953
transform 1 0 48282 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_550
timestamp 1607639953
transform 1 0 51686 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_537
timestamp 1607639953
transform 1 0 50490 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_852
timestamp 1607639953
transform 1 0 51594 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_562
timestamp 1607639953
transform 1 0 52790 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_586
timestamp 1607639953
transform 1 0 54998 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_574
timestamp 1607639953
transform 1 0 53894 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_611
timestamp 1607639953
transform 1 0 57298 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_598
timestamp 1607639953
transform 1 0 56102 0 1 36448
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_853
timestamp 1607639953
transform 1 0 57206 0 1 36448
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_63_623
timestamp 1607639953
transform 1 0 58402 0 1 36448
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1607639953
transform -1 0 58862 0 1 36448
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_15
timestamp 1607639953
transform 1 0 2466 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_3
timestamp 1607639953
transform 1 0 1362 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1607639953
transform 1 0 1086 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_44
timestamp 1607639953
transform 1 0 5134 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_32
timestamp 1607639953
transform 1 0 4030 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_27
timestamp 1607639953
transform 1 0 3570 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_854
timestamp 1607639953
transform 1 0 3938 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_56
timestamp 1607639953
transform 1 0 6238 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_80
timestamp 1607639953
transform 1 0 8446 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_68
timestamp 1607639953
transform 1 0 7342 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_105
timestamp 1607639953
transform 1 0 10746 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_93
timestamp 1607639953
transform 1 0 9642 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_855
timestamp 1607639953
transform 1 0 9550 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_130
timestamp 1607639953
transform 1 0 13046 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_125
timestamp 1607639953
transform 1 0 12586 0 -1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_117
timestamp 1607639953
transform 1 0 11850 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _059_
timestamp 1607639953
transform 1 0 12770 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_154
timestamp 1607639953
transform 1 0 15254 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_150
timestamp 1607639953
transform 1 0 14886 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_142
timestamp 1607639953
transform 1 0 14150 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_856
timestamp 1607639953
transform 1 0 15162 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_166
timestamp 1607639953
transform 1 0 16358 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_190
timestamp 1607639953
transform 1 0 18566 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_178
timestamp 1607639953
transform 1 0 17462 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_215
timestamp 1607639953
transform 1 0 20866 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_202
timestamp 1607639953
transform 1 0 19670 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_857
timestamp 1607639953
transform 1 0 20774 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_239
timestamp 1607639953
transform 1 0 23074 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_227
timestamp 1607639953
transform 1 0 21970 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_263
timestamp 1607639953
transform 1 0 25282 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_251
timestamp 1607639953
transform 1 0 24178 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_279
timestamp 1607639953
transform 1 0 26754 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_858
timestamp 1607639953
transform 1 0 26386 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _060_
timestamp 1607639953
transform 1 0 26478 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_307
timestamp 1607639953
transform 1 0 29330 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_303
timestamp 1607639953
transform 1 0 28962 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_291
timestamp 1607639953
transform 1 0 27858 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _155_
timestamp 1607639953
transform 1 0 29054 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_64_327
timestamp 1607639953
transform 1 0 31170 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_323
timestamp 1607639953
transform 1 0 30802 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_319
timestamp 1607639953
transform 1 0 30434 0 -1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _119_
timestamp 1607639953
transform 1 0 30894 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_349
timestamp 1607639953
transform 1 0 33194 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_337
timestamp 1607639953
transform 1 0 32090 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_335
timestamp 1607639953
transform 1 0 31906 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_859
timestamp 1607639953
transform 1 0 31998 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_373
timestamp 1607639953
transform 1 0 35402 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_361
timestamp 1607639953
transform 1 0 34298 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_385
timestamp 1607639953
transform 1 0 36506 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_410
timestamp 1607639953
transform 1 0 38806 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_398
timestamp 1607639953
transform 1 0 37702 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_860
timestamp 1607639953
transform 1 0 37610 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_434
timestamp 1607639953
transform 1 0 41014 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_422
timestamp 1607639953
transform 1 0 39910 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_459
timestamp 1607639953
transform 1 0 43314 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_446
timestamp 1607639953
transform 1 0 42118 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_861
timestamp 1607639953
transform 1 0 43222 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _003_
timestamp 1607639953
transform 1 0 43590 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_477
timestamp 1607639953
transform 1 0 44970 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_465
timestamp 1607639953
transform 1 0 43866 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_504
timestamp 1607639953
transform 1 0 47454 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_489
timestamp 1607639953
transform 1 0 46074 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _203_
timestamp 1607639953
transform 1 0 47178 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_520
timestamp 1607639953
transform 1 0 48926 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_516
timestamp 1607639953
transform 1 0 48558 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_862
timestamp 1607639953
transform 1 0 48834 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_544
timestamp 1607639953
transform 1 0 51134 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_532
timestamp 1607639953
transform 1 0 50030 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_568
timestamp 1607639953
transform 1 0 53342 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_556
timestamp 1607639953
transform 1 0 52238 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_593
timestamp 1607639953
transform 1 0 55642 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_581
timestamp 1607639953
transform 1 0 54538 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_863
timestamp 1607639953
transform 1 0 54446 0 -1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_605
timestamp 1607639953
transform 1 0 56746 0 -1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_617
timestamp 1607639953
transform 1 0 57850 0 -1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1607639953
transform -1 0 58862 0 -1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_65_15
timestamp 1607639953
transform 1 0 2466 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_3
timestamp 1607639953
transform 1 0 1362 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1607639953
transform 1 0 1086 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_65_39
timestamp 1607639953
transform 1 0 4674 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_27
timestamp 1607639953
transform 1 0 3570 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_62
timestamp 1607639953
transform 1 0 6790 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_65_59
timestamp 1607639953
transform 1 0 6514 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_65_51
timestamp 1607639953
transform 1 0 5778 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_864
timestamp 1607639953
transform 1 0 6698 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_86
timestamp 1607639953
transform 1 0 8998 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_74
timestamp 1607639953
transform 1 0 7894 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_110
timestamp 1607639953
transform 1 0 11206 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_98
timestamp 1607639953
transform 1 0 10102 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_123
timestamp 1607639953
transform 1 0 12402 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_865
timestamp 1607639953
transform 1 0 12310 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_147
timestamp 1607639953
transform 1 0 14610 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_135
timestamp 1607639953
transform 1 0 13506 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_171
timestamp 1607639953
transform 1 0 16818 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_159
timestamp 1607639953
transform 1 0 15714 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_196
timestamp 1607639953
transform 1 0 19118 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_184
timestamp 1607639953
transform 1 0 18014 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_866
timestamp 1607639953
transform 1 0 17922 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_220
timestamp 1607639953
transform 1 0 21326 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_208
timestamp 1607639953
transform 1 0 20222 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_232
timestamp 1607639953
transform 1 0 22430 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_257
timestamp 1607639953
transform 1 0 24730 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_245
timestamp 1607639953
transform 1 0 23626 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_867
timestamp 1607639953
transform 1 0 23534 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_281
timestamp 1607639953
transform 1 0 26938 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_269
timestamp 1607639953
transform 1 0 25834 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_306
timestamp 1607639953
transform 1 0 29238 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_293
timestamp 1607639953
transform 1 0 28042 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_868
timestamp 1607639953
transform 1 0 29146 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_330
timestamp 1607639953
transform 1 0 31446 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_318
timestamp 1607639953
transform 1 0 30342 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_342
timestamp 1607639953
transform 1 0 32550 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_367
timestamp 1607639953
transform 1 0 34850 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_354
timestamp 1607639953
transform 1 0 33654 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_869
timestamp 1607639953
transform 1 0 34758 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_391
timestamp 1607639953
transform 1 0 37058 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_379
timestamp 1607639953
transform 1 0 35954 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_415
timestamp 1607639953
transform 1 0 39266 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_403
timestamp 1607639953
transform 1 0 38162 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_440
timestamp 1607639953
transform 1 0 41566 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_428
timestamp 1607639953
transform 1 0 40462 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_870
timestamp 1607639953
transform 1 0 40370 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_452
timestamp 1607639953
transform 1 0 42670 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_476
timestamp 1607639953
transform 1 0 44878 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_464
timestamp 1607639953
transform 1 0 43774 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_501
timestamp 1607639953
transform 1 0 47178 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_489
timestamp 1607639953
transform 1 0 46074 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_871
timestamp 1607639953
transform 1 0 45982 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_525
timestamp 1607639953
transform 1 0 49386 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_65_513
timestamp 1607639953
transform 1 0 48282 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _144_
timestamp 1607639953
transform 1 0 49570 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_65_550
timestamp 1607639953
transform 1 0 51686 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_65_546
timestamp 1607639953
transform 1 0 51318 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_65_538
timestamp 1607639953
transform 1 0 50582 0 1 37536
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_534
timestamp 1607639953
transform 1 0 50214 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_530
timestamp 1607639953
transform 1 0 49846 0 1 37536
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_872
timestamp 1607639953
transform 1 0 51594 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _076_
timestamp 1607639953
transform 1 0 50306 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_65_567
timestamp 1607639953
transform 1 0 53250 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_555
timestamp 1607639953
transform 1 0 52146 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _191_
timestamp 1607639953
transform 1 0 51870 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_65_591
timestamp 1607639953
transform 1 0 55458 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_579
timestamp 1607639953
transform 1 0 54354 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_611
timestamp 1607639953
transform 1 0 57298 0 1 37536
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_65_609
timestamp 1607639953
transform 1 0 57114 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_65_603
timestamp 1607639953
transform 1 0 56562 0 1 37536
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_873
timestamp 1607639953
transform 1 0 57206 0 1 37536
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_65_623
timestamp 1607639953
transform 1 0 58402 0 1 37536
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1607639953
transform -1 0 58862 0 1 37536
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_67_3
timestamp 1607639953
transform 1 0 1362 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_66_3
timestamp 1607639953
transform 1 0 1362 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1607639953
transform 1 0 1086 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1607639953
transform 1 0 1086 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _106_
timestamp 1607639953
transform 1 0 1454 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _045_
timestamp 1607639953
transform 1 0 1638 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_67_21
timestamp 1607639953
transform 1 0 3018 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_9
timestamp 1607639953
transform 1 0 1914 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_19
timestamp 1607639953
transform 1 0 2834 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_7
timestamp 1607639953
transform 1 0 1730 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_33
timestamp 1607639953
transform 1 0 4122 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_44
timestamp 1607639953
transform 1 0 5134 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_32
timestamp 1607639953
transform 1 0 4030 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_874
timestamp 1607639953
transform 1 0 3938 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_62
timestamp 1607639953
transform 1 0 6790 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_57
timestamp 1607639953
transform 1 0 6330 0 1 38624
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_67_45
timestamp 1607639953
transform 1 0 5226 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_56
timestamp 1607639953
transform 1 0 6238 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_884
timestamp 1607639953
transform 1 0 6698 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_86
timestamp 1607639953
transform 1 0 8998 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_74
timestamp 1607639953
transform 1 0 7894 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_80
timestamp 1607639953
transform 1 0 8446 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_68
timestamp 1607639953
transform 1 0 7342 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_110
timestamp 1607639953
transform 1 0 11206 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_98
timestamp 1607639953
transform 1 0 10102 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_105
timestamp 1607639953
transform 1 0 10746 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_93
timestamp 1607639953
transform 1 0 9642 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_875
timestamp 1607639953
transform 1 0 9550 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_126
timestamp 1607639953
transform 1 0 12678 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_129
timestamp 1607639953
transform 1 0 12954 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_117
timestamp 1607639953
transform 1 0 11850 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_885
timestamp 1607639953
transform 1 0 12310 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _065_
timestamp 1607639953
transform 1 0 12402 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_67_150
timestamp 1607639953
transform 1 0 14886 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_138
timestamp 1607639953
transform 1 0 13782 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_154
timestamp 1607639953
transform 1 0 15254 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_141
timestamp 1607639953
transform 1 0 14058 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_876
timestamp 1607639953
transform 1 0 15162 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_174
timestamp 1607639953
transform 1 0 17094 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_67_162
timestamp 1607639953
transform 1 0 15990 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_166
timestamp 1607639953
transform 1 0 16358 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_196
timestamp 1607639953
transform 1 0 19118 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_184
timestamp 1607639953
transform 1 0 18014 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_67_182
timestamp 1607639953
transform 1 0 17830 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_190
timestamp 1607639953
transform 1 0 18566 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_178
timestamp 1607639953
transform 1 0 17462 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_886
timestamp 1607639953
transform 1 0 17922 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_67_216
timestamp 1607639953
transform 1 0 20958 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_67_208
timestamp 1607639953
transform 1 0 20222 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_66_215
timestamp 1607639953
transform 1 0 20866 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_202
timestamp 1607639953
transform 1 0 19670 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_877
timestamp 1607639953
transform 1 0 20774 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _179_
timestamp 1607639953
transform 1 0 21234 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_67_242
timestamp 1607639953
transform 1 0 23350 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_67_234
timestamp 1607639953
transform 1 0 22614 0 1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_67_222
timestamp 1607639953
transform 1 0 21510 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_239
timestamp 1607639953
transform 1 0 23074 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_227
timestamp 1607639953
transform 1 0 21970 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_257
timestamp 1607639953
transform 1 0 24730 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_245
timestamp 1607639953
transform 1 0 23626 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_263
timestamp 1607639953
transform 1 0 25282 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_251
timestamp 1607639953
transform 1 0 24178 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_887
timestamp 1607639953
transform 1 0 23534 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_281
timestamp 1607639953
transform 1 0 26938 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_269
timestamp 1607639953
transform 1 0 25834 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_276
timestamp 1607639953
transform 1 0 26478 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_878
timestamp 1607639953
transform 1 0 26386 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_306
timestamp 1607639953
transform 1 0 29238 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_293
timestamp 1607639953
transform 1 0 28042 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_300
timestamp 1607639953
transform 1 0 28686 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_288
timestamp 1607639953
transform 1 0 27582 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_888
timestamp 1607639953
transform 1 0 29146 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_330
timestamp 1607639953
transform 1 0 31446 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_318
timestamp 1607639953
transform 1 0 30342 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_324
timestamp 1607639953
transform 1 0 30894 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_312
timestamp 1607639953
transform 1 0 29790 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_342
timestamp 1607639953
transform 1 0 32550 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_349
timestamp 1607639953
transform 1 0 33194 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_337
timestamp 1607639953
transform 1 0 32090 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_879
timestamp 1607639953
transform 1 0 31998 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_367
timestamp 1607639953
transform 1 0 34850 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_354
timestamp 1607639953
transform 1 0 33654 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_373
timestamp 1607639953
transform 1 0 35402 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_361
timestamp 1607639953
transform 1 0 34298 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_889
timestamp 1607639953
transform 1 0 34758 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_391
timestamp 1607639953
transform 1 0 37058 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_379
timestamp 1607639953
transform 1 0 35954 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_385
timestamp 1607639953
transform 1 0 36506 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_415
timestamp 1607639953
transform 1 0 39266 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_403
timestamp 1607639953
transform 1 0 38162 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_410
timestamp 1607639953
transform 1 0 38806 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_398
timestamp 1607639953
transform 1 0 37702 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_880
timestamp 1607639953
transform 1 0 37610 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_440
timestamp 1607639953
transform 1 0 41566 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_428
timestamp 1607639953
transform 1 0 40462 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_434
timestamp 1607639953
transform 1 0 41014 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_422
timestamp 1607639953
transform 1 0 39910 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_890
timestamp 1607639953
transform 1 0 40370 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_452
timestamp 1607639953
transform 1 0 42670 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_459
timestamp 1607639953
transform 1 0 43314 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_446
timestamp 1607639953
transform 1 0 42118 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_881
timestamp 1607639953
transform 1 0 43222 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_476
timestamp 1607639953
transform 1 0 44878 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_464
timestamp 1607639953
transform 1 0 43774 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_483
timestamp 1607639953
transform 1 0 45522 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_471
timestamp 1607639953
transform 1 0 44418 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_501
timestamp 1607639953
transform 1 0 47178 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_489
timestamp 1607639953
transform 1 0 46074 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_66_503
timestamp 1607639953
transform 1 0 47362 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_66_495
timestamp 1607639953
transform 1 0 46626 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_891
timestamp 1607639953
transform 1 0 45982 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _139_
timestamp 1607639953
transform 1 0 47638 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_67_525
timestamp 1607639953
transform 1 0 49386 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_513
timestamp 1607639953
transform 1 0 48282 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_520
timestamp 1607639953
transform 1 0 48926 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_66_517
timestamp 1607639953
transform 1 0 48650 0 -1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_66_509
timestamp 1607639953
transform 1 0 47914 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_882
timestamp 1607639953
transform 1 0 48834 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_550
timestamp 1607639953
transform 1 0 51686 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_537
timestamp 1607639953
transform 1 0 50490 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_544
timestamp 1607639953
transform 1 0 51134 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_532
timestamp 1607639953
transform 1 0 50030 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_892
timestamp 1607639953
transform 1 0 51594 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_562
timestamp 1607639953
transform 1 0 52790 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_568
timestamp 1607639953
transform 1 0 53342 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_556
timestamp 1607639953
transform 1 0 52238 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_586
timestamp 1607639953
transform 1 0 54998 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_574
timestamp 1607639953
transform 1 0 53894 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_593
timestamp 1607639953
transform 1 0 55642 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_581
timestamp 1607639953
transform 1 0 54538 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_883
timestamp 1607639953
transform 1 0 54446 0 -1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_611
timestamp 1607639953
transform 1 0 57298 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_598
timestamp 1607639953
transform 1 0 56102 0 1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_605
timestamp 1607639953
transform 1 0 56746 0 -1 38624
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_893
timestamp 1607639953
transform 1 0 57206 0 1 38624
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_67_623
timestamp 1607639953
transform 1 0 58402 0 1 38624
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_66_617
timestamp 1607639953
transform 1 0 57850 0 -1 38624
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1607639953
transform -1 0 58862 0 1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1607639953
transform -1 0 58862 0 -1 38624
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_15
timestamp 1607639953
transform 1 0 2466 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_3
timestamp 1607639953
transform 1 0 1362 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1607639953
transform 1 0 1086 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_44
timestamp 1607639953
transform 1 0 5134 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_32
timestamp 1607639953
transform 1 0 4030 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_68_27
timestamp 1607639953
transform 1 0 3570 0 -1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_894
timestamp 1607639953
transform 1 0 3938 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_56
timestamp 1607639953
transform 1 0 6238 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_80
timestamp 1607639953
transform 1 0 8446 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_68
timestamp 1607639953
transform 1 0 7342 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_108
timestamp 1607639953
transform 1 0 11022 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_93
timestamp 1607639953
transform 1 0 9642 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_895
timestamp 1607639953
transform 1 0 9550 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _148_
timestamp 1607639953
transform 1 0 10746 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_132
timestamp 1607639953
transform 1 0 13230 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_120
timestamp 1607639953
transform 1 0 12126 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_154
timestamp 1607639953
transform 1 0 15254 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_152
timestamp 1607639953
transform 1 0 15070 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_144
timestamp 1607639953
transform 1 0 14334 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_896
timestamp 1607639953
transform 1 0 15162 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_166
timestamp 1607639953
transform 1 0 16358 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_190
timestamp 1607639953
transform 1 0 18566 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_178
timestamp 1607639953
transform 1 0 17462 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_215
timestamp 1607639953
transform 1 0 20866 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_202
timestamp 1607639953
transform 1 0 19670 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_897
timestamp 1607639953
transform 1 0 20774 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_239
timestamp 1607639953
transform 1 0 23074 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_227
timestamp 1607639953
transform 1 0 21970 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_263
timestamp 1607639953
transform 1 0 25282 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_251
timestamp 1607639953
transform 1 0 24178 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_276
timestamp 1607639953
transform 1 0 26478 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_898
timestamp 1607639953
transform 1 0 26386 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_300
timestamp 1607639953
transform 1 0 28686 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_288
timestamp 1607639953
transform 1 0 27582 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_324
timestamp 1607639953
transform 1 0 30894 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_312
timestamp 1607639953
transform 1 0 29790 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_349
timestamp 1607639953
transform 1 0 33194 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_337
timestamp 1607639953
transform 1 0 32090 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_899
timestamp 1607639953
transform 1 0 31998 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_373
timestamp 1607639953
transform 1 0 35402 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_361
timestamp 1607639953
transform 1 0 34298 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_385
timestamp 1607639953
transform 1 0 36506 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_410
timestamp 1607639953
transform 1 0 38806 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_398
timestamp 1607639953
transform 1 0 37702 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_900
timestamp 1607639953
transform 1 0 37610 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_434
timestamp 1607639953
transform 1 0 41014 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_422
timestamp 1607639953
transform 1 0 39910 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_459
timestamp 1607639953
transform 1 0 43314 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_446
timestamp 1607639953
transform 1 0 42118 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_901
timestamp 1607639953
transform 1 0 43222 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_483
timestamp 1607639953
transform 1 0 45522 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_471
timestamp 1607639953
transform 1 0 44418 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_495
timestamp 1607639953
transform 1 0 46626 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_520
timestamp 1607639953
transform 1 0 48926 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_507
timestamp 1607639953
transform 1 0 47730 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_902
timestamp 1607639953
transform 1 0 48834 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_544
timestamp 1607639953
transform 1 0 51134 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_532
timestamp 1607639953
transform 1 0 50030 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_568
timestamp 1607639953
transform 1 0 53342 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_556
timestamp 1607639953
transform 1 0 52238 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_593
timestamp 1607639953
transform 1 0 55642 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_581
timestamp 1607639953
transform 1 0 54538 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_903
timestamp 1607639953
transform 1 0 54446 0 -1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_605
timestamp 1607639953
transform 1 0 56746 0 -1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_617
timestamp 1607639953
transform 1 0 57850 0 -1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1607639953
transform -1 0 58862 0 -1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_69_15
timestamp 1607639953
transform 1 0 2466 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_3
timestamp 1607639953
transform 1 0 1362 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1607639953
transform 1 0 1086 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_69_39
timestamp 1607639953
transform 1 0 4674 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_27
timestamp 1607639953
transform 1 0 3570 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_62
timestamp 1607639953
transform 1 0 6790 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_69_59
timestamp 1607639953
transform 1 0 6514 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_69_51
timestamp 1607639953
transform 1 0 5778 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_904
timestamp 1607639953
transform 1 0 6698 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_86
timestamp 1607639953
transform 1 0 8998 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_74
timestamp 1607639953
transform 1 0 7894 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_110
timestamp 1607639953
transform 1 0 11206 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_98
timestamp 1607639953
transform 1 0 10102 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_123
timestamp 1607639953
transform 1 0 12402 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_905
timestamp 1607639953
transform 1 0 12310 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_147
timestamp 1607639953
transform 1 0 14610 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_135
timestamp 1607639953
transform 1 0 13506 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_171
timestamp 1607639953
transform 1 0 16818 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_159
timestamp 1607639953
transform 1 0 15714 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_196
timestamp 1607639953
transform 1 0 19118 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_184
timestamp 1607639953
transform 1 0 18014 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_906
timestamp 1607639953
transform 1 0 17922 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_220
timestamp 1607639953
transform 1 0 21326 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_208
timestamp 1607639953
transform 1 0 20222 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_232
timestamp 1607639953
transform 1 0 22430 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_257
timestamp 1607639953
transform 1 0 24730 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_245
timestamp 1607639953
transform 1 0 23626 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_907
timestamp 1607639953
transform 1 0 23534 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_284
timestamp 1607639953
transform 1 0 27214 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_269
timestamp 1607639953
transform 1 0 25834 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _007_
timestamp 1607639953
transform 1 0 26938 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_69_306
timestamp 1607639953
transform 1 0 29238 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_69_304
timestamp 1607639953
transform 1 0 29054 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_296
timestamp 1607639953
transform 1 0 28318 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_908
timestamp 1607639953
transform 1 0 29146 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_330
timestamp 1607639953
transform 1 0 31446 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_318
timestamp 1607639953
transform 1 0 30342 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_342
timestamp 1607639953
transform 1 0 32550 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_367
timestamp 1607639953
transform 1 0 34850 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_354
timestamp 1607639953
transform 1 0 33654 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_909
timestamp 1607639953
transform 1 0 34758 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_391
timestamp 1607639953
transform 1 0 37058 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_379
timestamp 1607639953
transform 1 0 35954 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_415
timestamp 1607639953
transform 1 0 39266 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_403
timestamp 1607639953
transform 1 0 38162 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_440
timestamp 1607639953
transform 1 0 41566 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_428
timestamp 1607639953
transform 1 0 40462 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_910
timestamp 1607639953
transform 1 0 40370 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_452
timestamp 1607639953
transform 1 0 42670 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_476
timestamp 1607639953
transform 1 0 44878 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_464
timestamp 1607639953
transform 1 0 43774 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_500
timestamp 1607639953
transform 1 0 47086 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_69_489
timestamp 1607639953
transform 1 0 46074 0 1 39712
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_911
timestamp 1607639953
transform 1 0 45982 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _111_
timestamp 1607639953
transform 1 0 46810 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_69_519
timestamp 1607639953
transform 1 0 48834 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_512
timestamp 1607639953
transform 1 0 48190 0 1 39712
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _078_
timestamp 1607639953
transform 1 0 48558 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_69_550
timestamp 1607639953
transform 1 0 51686 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_543
timestamp 1607639953
transform 1 0 51042 0 1 39712
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_69_531
timestamp 1607639953
transform 1 0 49938 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_912
timestamp 1607639953
transform 1 0 51594 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_562
timestamp 1607639953
transform 1 0 52790 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_586
timestamp 1607639953
transform 1 0 54998 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_574
timestamp 1607639953
transform 1 0 53894 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_611
timestamp 1607639953
transform 1 0 57298 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_598
timestamp 1607639953
transform 1 0 56102 0 1 39712
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_913
timestamp 1607639953
transform 1 0 57206 0 1 39712
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_69_623
timestamp 1607639953
transform 1 0 58402 0 1 39712
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1607639953
transform -1 0 58862 0 1 39712
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_70_15
timestamp 1607639953
transform 1 0 2466 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_3
timestamp 1607639953
transform 1 0 1362 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1607639953
transform 1 0 1086 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_70_44
timestamp 1607639953
transform 1 0 5134 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_32
timestamp 1607639953
transform 1 0 4030 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_70_27
timestamp 1607639953
transform 1 0 3570 0 -1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_914
timestamp 1607639953
transform 1 0 3938 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_56
timestamp 1607639953
transform 1 0 6238 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_80
timestamp 1607639953
transform 1 0 8446 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_68
timestamp 1607639953
transform 1 0 7342 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_105
timestamp 1607639953
transform 1 0 10746 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_70_93
timestamp 1607639953
transform 1 0 9642 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_915
timestamp 1607639953
transform 1 0 9550 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_130
timestamp 1607639953
transform 1 0 13046 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_118
timestamp 1607639953
transform 1 0 11942 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_70_113
timestamp 1607639953
transform 1 0 11482 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__conb_1  _089_
timestamp 1607639953
transform 1 0 11666 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_70_154
timestamp 1607639953
transform 1 0 15254 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_70_150
timestamp 1607639953
transform 1 0 14886 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_70_142
timestamp 1607639953
transform 1 0 14150 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_916
timestamp 1607639953
transform 1 0 15162 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_166
timestamp 1607639953
transform 1 0 16358 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_190
timestamp 1607639953
transform 1 0 18566 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_178
timestamp 1607639953
transform 1 0 17462 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_215
timestamp 1607639953
transform 1 0 20866 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_202
timestamp 1607639953
transform 1 0 19670 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_917
timestamp 1607639953
transform 1 0 20774 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_239
timestamp 1607639953
transform 1 0 23074 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_227
timestamp 1607639953
transform 1 0 21970 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_263
timestamp 1607639953
transform 1 0 25282 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_251
timestamp 1607639953
transform 1 0 24178 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_276
timestamp 1607639953
transform 1 0 26478 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_918
timestamp 1607639953
transform 1 0 26386 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_300
timestamp 1607639953
transform 1 0 28686 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_288
timestamp 1607639953
transform 1 0 27582 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_324
timestamp 1607639953
transform 1 0 30894 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_312
timestamp 1607639953
transform 1 0 29790 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_349
timestamp 1607639953
transform 1 0 33194 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_337
timestamp 1607639953
transform 1 0 32090 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_919
timestamp 1607639953
transform 1 0 31998 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_373
timestamp 1607639953
transform 1 0 35402 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_361
timestamp 1607639953
transform 1 0 34298 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_385
timestamp 1607639953
transform 1 0 36506 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_410
timestamp 1607639953
transform 1 0 38806 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_398
timestamp 1607639953
transform 1 0 37702 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_920
timestamp 1607639953
transform 1 0 37610 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_434
timestamp 1607639953
transform 1 0 41014 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_422
timestamp 1607639953
transform 1 0 39910 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_70_459
timestamp 1607639953
transform 1 0 43314 0 -1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_70_446
timestamp 1607639953
transform 1 0 42118 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_921
timestamp 1607639953
transform 1 0 43222 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _181_
timestamp 1607639953
transform 1 0 43498 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_70_476
timestamp 1607639953
transform 1 0 44878 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_464
timestamp 1607639953
transform 1 0 43774 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_500
timestamp 1607639953
transform 1 0 47086 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_488
timestamp 1607639953
transform 1 0 45982 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_520
timestamp 1607639953
transform 1 0 48926 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_518
timestamp 1607639953
transform 1 0 48742 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_70_512
timestamp 1607639953
transform 1 0 48190 0 -1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_922
timestamp 1607639953
transform 1 0 48834 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_544
timestamp 1607639953
transform 1 0 51134 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_532
timestamp 1607639953
transform 1 0 50030 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_568
timestamp 1607639953
transform 1 0 53342 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_556
timestamp 1607639953
transform 1 0 52238 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_593
timestamp 1607639953
transform 1 0 55642 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_581
timestamp 1607639953
transform 1 0 54538 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_923
timestamp 1607639953
transform 1 0 54446 0 -1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_605
timestamp 1607639953
transform 1 0 56746 0 -1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_617
timestamp 1607639953
transform 1 0 57850 0 -1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1607639953
transform -1 0 58862 0 -1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_71_15
timestamp 1607639953
transform 1 0 2466 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_3
timestamp 1607639953
transform 1 0 1362 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1607639953
transform 1 0 1086 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_71_39
timestamp 1607639953
transform 1 0 4674 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_27
timestamp 1607639953
transform 1 0 3570 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_62
timestamp 1607639953
transform 1 0 6790 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_71_59
timestamp 1607639953
transform 1 0 6514 0 1 40800
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_71_51
timestamp 1607639953
transform 1 0 5778 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_924
timestamp 1607639953
transform 1 0 6698 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_86
timestamp 1607639953
transform 1 0 8998 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_74
timestamp 1607639953
transform 1 0 7894 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_110
timestamp 1607639953
transform 1 0 11206 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_98
timestamp 1607639953
transform 1 0 10102 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_123
timestamp 1607639953
transform 1 0 12402 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_925
timestamp 1607639953
transform 1 0 12310 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_147
timestamp 1607639953
transform 1 0 14610 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_135
timestamp 1607639953
transform 1 0 13506 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_171
timestamp 1607639953
transform 1 0 16818 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_159
timestamp 1607639953
transform 1 0 15714 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_196
timestamp 1607639953
transform 1 0 19118 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_184
timestamp 1607639953
transform 1 0 18014 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_926
timestamp 1607639953
transform 1 0 17922 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_220
timestamp 1607639953
transform 1 0 21326 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_208
timestamp 1607639953
transform 1 0 20222 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_232
timestamp 1607639953
transform 1 0 22430 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_257
timestamp 1607639953
transform 1 0 24730 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_245
timestamp 1607639953
transform 1 0 23626 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_927
timestamp 1607639953
transform 1 0 23534 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_281
timestamp 1607639953
transform 1 0 26938 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_269
timestamp 1607639953
transform 1 0 25834 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_306
timestamp 1607639953
transform 1 0 29238 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_293
timestamp 1607639953
transform 1 0 28042 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_928
timestamp 1607639953
transform 1 0 29146 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_330
timestamp 1607639953
transform 1 0 31446 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_318
timestamp 1607639953
transform 1 0 30342 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_342
timestamp 1607639953
transform 1 0 32550 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_367
timestamp 1607639953
transform 1 0 34850 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_354
timestamp 1607639953
transform 1 0 33654 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_929
timestamp 1607639953
transform 1 0 34758 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_391
timestamp 1607639953
transform 1 0 37058 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_379
timestamp 1607639953
transform 1 0 35954 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_415
timestamp 1607639953
transform 1 0 39266 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_403
timestamp 1607639953
transform 1 0 38162 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_440
timestamp 1607639953
transform 1 0 41566 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_428
timestamp 1607639953
transform 1 0 40462 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_930
timestamp 1607639953
transform 1 0 40370 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_452
timestamp 1607639953
transform 1 0 42670 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_476
timestamp 1607639953
transform 1 0 44878 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_464
timestamp 1607639953
transform 1 0 43774 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_504
timestamp 1607639953
transform 1 0 47454 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_492
timestamp 1607639953
transform 1 0 46350 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_931
timestamp 1607639953
transform 1 0 45982 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _125_
timestamp 1607639953
transform 1 0 46074 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_71_528
timestamp 1607639953
transform 1 0 49662 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_516
timestamp 1607639953
transform 1 0 48558 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_550
timestamp 1607639953
transform 1 0 51686 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_71_548
timestamp 1607639953
transform 1 0 51502 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_71_540
timestamp 1607639953
transform 1 0 50766 0 1 40800
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_932
timestamp 1607639953
transform 1 0 51594 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_562
timestamp 1607639953
transform 1 0 52790 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_586
timestamp 1607639953
transform 1 0 54998 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_574
timestamp 1607639953
transform 1 0 53894 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_611
timestamp 1607639953
transform 1 0 57298 0 1 40800
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_71_598
timestamp 1607639953
transform 1 0 56102 0 1 40800
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_933
timestamp 1607639953
transform 1 0 57206 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _146_
timestamp 1607639953
transform 1 0 57666 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_71_624
timestamp 1607639953
transform 1 0 58494 0 1 40800
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_71_618
timestamp 1607639953
transform 1 0 57942 0 1 40800
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1607639953
transform -1 0 58862 0 1 40800
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_73_15
timestamp 1607639953
transform 1 0 2466 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_3
timestamp 1607639953
transform 1 0 1362 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_15
timestamp 1607639953
transform 1 0 2466 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_3
timestamp 1607639953
transform 1 0 1362 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1607639953
transform 1 0 1086 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1607639953
transform 1 0 1086 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_73_39
timestamp 1607639953
transform 1 0 4674 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_27
timestamp 1607639953
transform 1 0 3570 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_44
timestamp 1607639953
transform 1 0 5134 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_32
timestamp 1607639953
transform 1 0 4030 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_72_27
timestamp 1607639953
transform 1 0 3570 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_934
timestamp 1607639953
transform 1 0 3938 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_62
timestamp 1607639953
transform 1 0 6790 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_73_59
timestamp 1607639953
transform 1 0 6514 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_73_51
timestamp 1607639953
transform 1 0 5778 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_72_56
timestamp 1607639953
transform 1 0 6238 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_944
timestamp 1607639953
transform 1 0 6698 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_84
timestamp 1607639953
transform 1 0 8814 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_73_80
timestamp 1607639953
transform 1 0 8446 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_73_74
timestamp 1607639953
transform 1 0 7894 0 1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_72_80
timestamp 1607639953
transform 1 0 8446 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_68
timestamp 1607639953
transform 1 0 7342 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _092_
timestamp 1607639953
transform 1 0 8538 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_73_108
timestamp 1607639953
transform 1 0 11022 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_96
timestamp 1607639953
transform 1 0 9918 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_105
timestamp 1607639953
transform 1 0 10746 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_93
timestamp 1607639953
transform 1 0 9642 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_935
timestamp 1607639953
transform 1 0 9550 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_123
timestamp 1607639953
transform 1 0 12402 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_73_120
timestamp 1607639953
transform 1 0 12126 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_129
timestamp 1607639953
transform 1 0 12954 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_72_117
timestamp 1607639953
transform 1 0 11850 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_945
timestamp 1607639953
transform 1 0 12310 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_147
timestamp 1607639953
transform 1 0 14610 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_135
timestamp 1607639953
transform 1 0 13506 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_154
timestamp 1607639953
transform 1 0 15254 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_72_152
timestamp 1607639953
transform 1 0 15070 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_72_148
timestamp 1607639953
transform 1 0 14702 0 -1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_72_136
timestamp 1607639953
transform 1 0 13598 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_936
timestamp 1607639953
transform 1 0 15162 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _041_
timestamp 1607639953
transform 1 0 13322 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_73_171
timestamp 1607639953
transform 1 0 16818 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_159
timestamp 1607639953
transform 1 0 15714 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_166
timestamp 1607639953
transform 1 0 16358 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_187
timestamp 1607639953
transform 1 0 18290 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_190
timestamp 1607639953
transform 1 0 18566 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_178
timestamp 1607639953
transform 1 0 17462 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_946
timestamp 1607639953
transform 1 0 17922 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _132_
timestamp 1607639953
transform 1 0 18014 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_73_211
timestamp 1607639953
transform 1 0 20498 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_199
timestamp 1607639953
transform 1 0 19394 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_215
timestamp 1607639953
transform 1 0 20866 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_202
timestamp 1607639953
transform 1 0 19670 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_937
timestamp 1607639953
transform 1 0 20774 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_73_241
timestamp 1607639953
transform 1 0 23258 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_73_233
timestamp 1607639953
transform 1 0 22522 0 1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_73_229
timestamp 1607639953
transform 1 0 22154 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_73_223
timestamp 1607639953
transform 1 0 21602 0 1 41888
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_72_239
timestamp 1607639953
transform 1 0 23074 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_227
timestamp 1607639953
transform 1 0 21970 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _178_
timestamp 1607639953
transform 1 0 22246 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_73_257
timestamp 1607639953
transform 1 0 24730 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_245
timestamp 1607639953
transform 1 0 23626 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_263
timestamp 1607639953
transform 1 0 25282 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_251
timestamp 1607639953
transform 1 0 24178 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_947
timestamp 1607639953
transform 1 0 23534 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_281
timestamp 1607639953
transform 1 0 26938 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_269
timestamp 1607639953
transform 1 0 25834 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_276
timestamp 1607639953
transform 1 0 26478 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_938
timestamp 1607639953
transform 1 0 26386 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_306
timestamp 1607639953
transform 1 0 29238 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_73_293
timestamp 1607639953
transform 1 0 28042 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_300
timestamp 1607639953
transform 1 0 28686 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_288
timestamp 1607639953
transform 1 0 27582 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_948
timestamp 1607639953
transform 1 0 29146 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_325
timestamp 1607639953
transform 1 0 30986 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_313
timestamp 1607639953
transform 1 0 29882 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_324
timestamp 1607639953
transform 1 0 30894 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_312
timestamp 1607639953
transform 1 0 29790 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _005_
timestamp 1607639953
transform 1 0 29606 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_73_349
timestamp 1607639953
transform 1 0 33194 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_337
timestamp 1607639953
transform 1 0 32090 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_349
timestamp 1607639953
transform 1 0 33194 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_337
timestamp 1607639953
transform 1 0 32090 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_939
timestamp 1607639953
transform 1 0 31998 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_367
timestamp 1607639953
transform 1 0 34850 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_73_365
timestamp 1607639953
transform 1 0 34666 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_361
timestamp 1607639953
transform 1 0 34298 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_72_373
timestamp 1607639953
transform 1 0 35402 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_361
timestamp 1607639953
transform 1 0 34298 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_949
timestamp 1607639953
transform 1 0 34758 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_391
timestamp 1607639953
transform 1 0 37058 0 1 41888
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_73_379
timestamp 1607639953
transform 1 0 35954 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_385
timestamp 1607639953
transform 1 0 36506 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _058_
timestamp 1607639953
transform 1 0 37426 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_73_410
timestamp 1607639953
transform 1 0 38806 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_398
timestamp 1607639953
transform 1 0 37702 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_410
timestamp 1607639953
transform 1 0 38806 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_398
timestamp 1607639953
transform 1 0 37702 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_940
timestamp 1607639953
transform 1 0 37610 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_440
timestamp 1607639953
transform 1 0 41566 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_428
timestamp 1607639953
transform 1 0 40462 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_73_426
timestamp 1607639953
transform 1 0 40278 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_73_422
timestamp 1607639953
transform 1 0 39910 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_72_434
timestamp 1607639953
transform 1 0 41014 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_72_422
timestamp 1607639953
transform 1 0 39910 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_950
timestamp 1607639953
transform 1 0 40370 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _052_
timestamp 1607639953
transform 1 0 40002 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_73_452
timestamp 1607639953
transform 1 0 42670 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_459
timestamp 1607639953
transform 1 0 43314 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_72_456
timestamp 1607639953
transform 1 0 43038 0 -1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_72_448
timestamp 1607639953
transform 1 0 42302 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_72_442
timestamp 1607639953
transform 1 0 41750 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_941
timestamp 1607639953
transform 1 0 43222 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _143_
timestamp 1607639953
transform 1 0 42026 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_73_476
timestamp 1607639953
transform 1 0 44878 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_464
timestamp 1607639953
transform 1 0 43774 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_483
timestamp 1607639953
transform 1 0 45522 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_471
timestamp 1607639953
transform 1 0 44418 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_501
timestamp 1607639953
transform 1 0 47178 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_489
timestamp 1607639953
transform 1 0 46074 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_495
timestamp 1607639953
transform 1 0 46626 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_951
timestamp 1607639953
transform 1 0 45982 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_525
timestamp 1607639953
transform 1 0 49386 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_513
timestamp 1607639953
transform 1 0 48282 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_520
timestamp 1607639953
transform 1 0 48926 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_507
timestamp 1607639953
transform 1 0 47730 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_942
timestamp 1607639953
transform 1 0 48834 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_550
timestamp 1607639953
transform 1 0 51686 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_537
timestamp 1607639953
transform 1 0 50490 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_544
timestamp 1607639953
transform 1 0 51134 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_532
timestamp 1607639953
transform 1 0 50030 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_952
timestamp 1607639953
transform 1 0 51594 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_562
timestamp 1607639953
transform 1 0 52790 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_568
timestamp 1607639953
transform 1 0 53342 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_556
timestamp 1607639953
transform 1 0 52238 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_586
timestamp 1607639953
transform 1 0 54998 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_574
timestamp 1607639953
transform 1 0 53894 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_593
timestamp 1607639953
transform 1 0 55642 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_581
timestamp 1607639953
transform 1 0 54538 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_943
timestamp 1607639953
transform 1 0 54446 0 -1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_611
timestamp 1607639953
transform 1 0 57298 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_598
timestamp 1607639953
transform 1 0 56102 0 1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_605
timestamp 1607639953
transform 1 0 56746 0 -1 41888
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_953
timestamp 1607639953
transform 1 0 57206 0 1 41888
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_73_623
timestamp 1607639953
transform 1 0 58402 0 1 41888
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_72_617
timestamp 1607639953
transform 1 0 57850 0 -1 41888
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1607639953
transform -1 0 58862 0 1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1607639953
transform -1 0 58862 0 -1 41888
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_74_15
timestamp 1607639953
transform 1 0 2466 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_3
timestamp 1607639953
transform 1 0 1362 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1607639953
transform 1 0 1086 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_74_44
timestamp 1607639953
transform 1 0 5134 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_32
timestamp 1607639953
transform 1 0 4030 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_74_27
timestamp 1607639953
transform 1 0 3570 0 -1 42976
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_954
timestamp 1607639953
transform 1 0 3938 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_56
timestamp 1607639953
transform 1 0 6238 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_80
timestamp 1607639953
transform 1 0 8446 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_68
timestamp 1607639953
transform 1 0 7342 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_105
timestamp 1607639953
transform 1 0 10746 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_93
timestamp 1607639953
transform 1 0 9642 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_955
timestamp 1607639953
transform 1 0 9550 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_129
timestamp 1607639953
transform 1 0 12954 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_117
timestamp 1607639953
transform 1 0 11850 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_154
timestamp 1607639953
transform 1 0 15254 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_141
timestamp 1607639953
transform 1 0 14058 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_956
timestamp 1607639953
transform 1 0 15162 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_166
timestamp 1607639953
transform 1 0 16358 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_190
timestamp 1607639953
transform 1 0 18566 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_178
timestamp 1607639953
transform 1 0 17462 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_215
timestamp 1607639953
transform 1 0 20866 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_202
timestamp 1607639953
transform 1 0 19670 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_957
timestamp 1607639953
transform 1 0 20774 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_239
timestamp 1607639953
transform 1 0 23074 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_227
timestamp 1607639953
transform 1 0 21970 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_263
timestamp 1607639953
transform 1 0 25282 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_251
timestamp 1607639953
transform 1 0 24178 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_276
timestamp 1607639953
transform 1 0 26478 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_958
timestamp 1607639953
transform 1 0 26386 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_300
timestamp 1607639953
transform 1 0 28686 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_288
timestamp 1607639953
transform 1 0 27582 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_324
timestamp 1607639953
transform 1 0 30894 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_312
timestamp 1607639953
transform 1 0 29790 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_347
timestamp 1607639953
transform 1 0 33010 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_343
timestamp 1607639953
transform 1 0 32642 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_74_337
timestamp 1607639953
transform 1 0 32090 0 -1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_959
timestamp 1607639953
transform 1 0 31998 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _021_
timestamp 1607639953
transform 1 0 32734 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_74_371
timestamp 1607639953
transform 1 0 35218 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_359
timestamp 1607639953
transform 1 0 34114 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_74_395
timestamp 1607639953
transform 1 0 37426 0 -1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_74_383
timestamp 1607639953
transform 1 0 36322 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_410
timestamp 1607639953
transform 1 0 38806 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_398
timestamp 1607639953
transform 1 0 37702 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_960
timestamp 1607639953
transform 1 0 37610 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_434
timestamp 1607639953
transform 1 0 41014 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_422
timestamp 1607639953
transform 1 0 39910 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_459
timestamp 1607639953
transform 1 0 43314 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_446
timestamp 1607639953
transform 1 0 42118 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_961
timestamp 1607639953
transform 1 0 43222 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_483
timestamp 1607639953
transform 1 0 45522 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_471
timestamp 1607639953
transform 1 0 44418 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_495
timestamp 1607639953
transform 1 0 46626 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_520
timestamp 1607639953
transform 1 0 48926 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_507
timestamp 1607639953
transform 1 0 47730 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_962
timestamp 1607639953
transform 1 0 48834 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_544
timestamp 1607639953
transform 1 0 51134 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_532
timestamp 1607639953
transform 1 0 50030 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_568
timestamp 1607639953
transform 1 0 53342 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_556
timestamp 1607639953
transform 1 0 52238 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_593
timestamp 1607639953
transform 1 0 55642 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_581
timestamp 1607639953
transform 1 0 54538 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_963
timestamp 1607639953
transform 1 0 54446 0 -1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_605
timestamp 1607639953
transform 1 0 56746 0 -1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_74_617
timestamp 1607639953
transform 1 0 57850 0 -1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1607639953
transform -1 0 58862 0 -1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_75_15
timestamp 1607639953
transform 1 0 2466 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_3
timestamp 1607639953
transform 1 0 1362 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1607639953
transform 1 0 1086 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_75_39
timestamp 1607639953
transform 1 0 4674 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_75_27
timestamp 1607639953
transform 1 0 3570 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_62
timestamp 1607639953
transform 1 0 6790 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_75_59
timestamp 1607639953
transform 1 0 6514 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_75_51
timestamp 1607639953
transform 1 0 5778 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_75_47
timestamp 1607639953
transform 1 0 5410 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_964
timestamp 1607639953
transform 1 0 6698 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _137_
timestamp 1607639953
transform 1 0 5502 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_75_86
timestamp 1607639953
transform 1 0 8998 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_74
timestamp 1607639953
transform 1 0 7894 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_110
timestamp 1607639953
transform 1 0 11206 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_98
timestamp 1607639953
transform 1 0 10102 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_123
timestamp 1607639953
transform 1 0 12402 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_965
timestamp 1607639953
transform 1 0 12310 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_147
timestamp 1607639953
transform 1 0 14610 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_135
timestamp 1607639953
transform 1 0 13506 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_171
timestamp 1607639953
transform 1 0 16818 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_159
timestamp 1607639953
transform 1 0 15714 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_196
timestamp 1607639953
transform 1 0 19118 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_184
timestamp 1607639953
transform 1 0 18014 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_966
timestamp 1607639953
transform 1 0 17922 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_220
timestamp 1607639953
transform 1 0 21326 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_208
timestamp 1607639953
transform 1 0 20222 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_232
timestamp 1607639953
transform 1 0 22430 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_257
timestamp 1607639953
transform 1 0 24730 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_245
timestamp 1607639953
transform 1 0 23626 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_967
timestamp 1607639953
transform 1 0 23534 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_281
timestamp 1607639953
transform 1 0 26938 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_269
timestamp 1607639953
transform 1 0 25834 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_306
timestamp 1607639953
transform 1 0 29238 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_293
timestamp 1607639953
transform 1 0 28042 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_968
timestamp 1607639953
transform 1 0 29146 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_330
timestamp 1607639953
transform 1 0 31446 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_318
timestamp 1607639953
transform 1 0 30342 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_342
timestamp 1607639953
transform 1 0 32550 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_367
timestamp 1607639953
transform 1 0 34850 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_354
timestamp 1607639953
transform 1 0 33654 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_969
timestamp 1607639953
transform 1 0 34758 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_391
timestamp 1607639953
transform 1 0 37058 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_379
timestamp 1607639953
transform 1 0 35954 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_415
timestamp 1607639953
transform 1 0 39266 0 1 42976
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_75_403
timestamp 1607639953
transform 1 0 38162 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_431
timestamp 1607639953
transform 1 0 40738 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_75_425
timestamp 1607639953
transform 1 0 40186 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_75_421
timestamp 1607639953
transform 1 0 39818 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_970
timestamp 1607639953
transform 1 0 40370 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _175_
timestamp 1607639953
transform 1 0 40462 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _029_
timestamp 1607639953
transform 1 0 39910 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_75_455
timestamp 1607639953
transform 1 0 42946 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_443
timestamp 1607639953
transform 1 0 41842 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_75_479
timestamp 1607639953
transform 1 0 45154 0 1 42976
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_75_467
timestamp 1607639953
transform 1 0 44050 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_501
timestamp 1607639953
transform 1 0 47178 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_489
timestamp 1607639953
transform 1 0 46074 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_75_487
timestamp 1607639953
transform 1 0 45890 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_971
timestamp 1607639953
transform 1 0 45982 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_525
timestamp 1607639953
transform 1 0 49386 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_513
timestamp 1607639953
transform 1 0 48282 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_550
timestamp 1607639953
transform 1 0 51686 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_537
timestamp 1607639953
transform 1 0 50490 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_972
timestamp 1607639953
transform 1 0 51594 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_562
timestamp 1607639953
transform 1 0 52790 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_586
timestamp 1607639953
transform 1 0 54998 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_574
timestamp 1607639953
transform 1 0 53894 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_611
timestamp 1607639953
transform 1 0 57298 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_598
timestamp 1607639953
transform 1 0 56102 0 1 42976
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_973
timestamp 1607639953
transform 1 0 57206 0 1 42976
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_75_623
timestamp 1607639953
transform 1 0 58402 0 1 42976
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1607639953
transform -1 0 58862 0 1 42976
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_76_15
timestamp 1607639953
transform 1 0 2466 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_3
timestamp 1607639953
transform 1 0 1362 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1607639953
transform 1 0 1086 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_76_44
timestamp 1607639953
transform 1 0 5134 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_32
timestamp 1607639953
transform 1 0 4030 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_27
timestamp 1607639953
transform 1 0 3570 0 -1 44064
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_974
timestamp 1607639953
transform 1 0 3938 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_56
timestamp 1607639953
transform 1 0 6238 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_80
timestamp 1607639953
transform 1 0 8446 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_68
timestamp 1607639953
transform 1 0 7342 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_105
timestamp 1607639953
transform 1 0 10746 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_93
timestamp 1607639953
transform 1 0 9642 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_975
timestamp 1607639953
transform 1 0 9550 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_129
timestamp 1607639953
transform 1 0 12954 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_117
timestamp 1607639953
transform 1 0 11850 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_154
timestamp 1607639953
transform 1 0 15254 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_141
timestamp 1607639953
transform 1 0 14058 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_976
timestamp 1607639953
transform 1 0 15162 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_166
timestamp 1607639953
transform 1 0 16358 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_190
timestamp 1607639953
transform 1 0 18566 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_178
timestamp 1607639953
transform 1 0 17462 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_215
timestamp 1607639953
transform 1 0 20866 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_202
timestamp 1607639953
transform 1 0 19670 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_977
timestamp 1607639953
transform 1 0 20774 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_239
timestamp 1607639953
transform 1 0 23074 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_227
timestamp 1607639953
transform 1 0 21970 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_263
timestamp 1607639953
transform 1 0 25282 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_251
timestamp 1607639953
transform 1 0 24178 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_276
timestamp 1607639953
transform 1 0 26478 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_978
timestamp 1607639953
transform 1 0 26386 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_300
timestamp 1607639953
transform 1 0 28686 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_288
timestamp 1607639953
transform 1 0 27582 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_324
timestamp 1607639953
transform 1 0 30894 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_312
timestamp 1607639953
transform 1 0 29790 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_349
timestamp 1607639953
transform 1 0 33194 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_337
timestamp 1607639953
transform 1 0 32090 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_979
timestamp 1607639953
transform 1 0 31998 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_373
timestamp 1607639953
transform 1 0 35402 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_361
timestamp 1607639953
transform 1 0 34298 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_385
timestamp 1607639953
transform 1 0 36506 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_410
timestamp 1607639953
transform 1 0 38806 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_398
timestamp 1607639953
transform 1 0 37702 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_980
timestamp 1607639953
transform 1 0 37610 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_434
timestamp 1607639953
transform 1 0 41014 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_422
timestamp 1607639953
transform 1 0 39910 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_459
timestamp 1607639953
transform 1 0 43314 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_446
timestamp 1607639953
transform 1 0 42118 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_981
timestamp 1607639953
transform 1 0 43222 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_483
timestamp 1607639953
transform 1 0 45522 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_471
timestamp 1607639953
transform 1 0 44418 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_495
timestamp 1607639953
transform 1 0 46626 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_520
timestamp 1607639953
transform 1 0 48926 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_507
timestamp 1607639953
transform 1 0 47730 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_982
timestamp 1607639953
transform 1 0 48834 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_544
timestamp 1607639953
transform 1 0 51134 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_532
timestamp 1607639953
transform 1 0 50030 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_568
timestamp 1607639953
transform 1 0 53342 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_556
timestamp 1607639953
transform 1 0 52238 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_593
timestamp 1607639953
transform 1 0 55642 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_581
timestamp 1607639953
transform 1 0 54538 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_983
timestamp 1607639953
transform 1 0 54446 0 -1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_605
timestamp 1607639953
transform 1 0 56746 0 -1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_76_617
timestamp 1607639953
transform 1 0 57850 0 -1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1607639953
transform -1 0 58862 0 -1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_77_15
timestamp 1607639953
transform 1 0 2466 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_3
timestamp 1607639953
transform 1 0 1362 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1607639953
transform 1 0 1086 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_77_39
timestamp 1607639953
transform 1 0 4674 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_27
timestamp 1607639953
transform 1 0 3570 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_62
timestamp 1607639953
transform 1 0 6790 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_77_59
timestamp 1607639953
transform 1 0 6514 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_77_51
timestamp 1607639953
transform 1 0 5778 0 1 44064
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_984
timestamp 1607639953
transform 1 0 6698 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_86
timestamp 1607639953
transform 1 0 8998 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_74
timestamp 1607639953
transform 1 0 7894 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_110
timestamp 1607639953
transform 1 0 11206 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_98
timestamp 1607639953
transform 1 0 10102 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_123
timestamp 1607639953
transform 1 0 12402 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_985
timestamp 1607639953
transform 1 0 12310 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_147
timestamp 1607639953
transform 1 0 14610 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_135
timestamp 1607639953
transform 1 0 13506 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_171
timestamp 1607639953
transform 1 0 16818 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_159
timestamp 1607639953
transform 1 0 15714 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_196
timestamp 1607639953
transform 1 0 19118 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_184
timestamp 1607639953
transform 1 0 18014 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_986
timestamp 1607639953
transform 1 0 17922 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_220
timestamp 1607639953
transform 1 0 21326 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_208
timestamp 1607639953
transform 1 0 20222 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_232
timestamp 1607639953
transform 1 0 22430 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_257
timestamp 1607639953
transform 1 0 24730 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_245
timestamp 1607639953
transform 1 0 23626 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_987
timestamp 1607639953
transform 1 0 23534 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_281
timestamp 1607639953
transform 1 0 26938 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_269
timestamp 1607639953
transform 1 0 25834 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_306
timestamp 1607639953
transform 1 0 29238 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_293
timestamp 1607639953
transform 1 0 28042 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_988
timestamp 1607639953
transform 1 0 29146 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_330
timestamp 1607639953
transform 1 0 31446 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_318
timestamp 1607639953
transform 1 0 30342 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_342
timestamp 1607639953
transform 1 0 32550 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_367
timestamp 1607639953
transform 1 0 34850 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_354
timestamp 1607639953
transform 1 0 33654 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_989
timestamp 1607639953
transform 1 0 34758 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_391
timestamp 1607639953
transform 1 0 37058 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_379
timestamp 1607639953
transform 1 0 35954 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_415
timestamp 1607639953
transform 1 0 39266 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_403
timestamp 1607639953
transform 1 0 38162 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_440
timestamp 1607639953
transform 1 0 41566 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_428
timestamp 1607639953
transform 1 0 40462 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_990
timestamp 1607639953
transform 1 0 40370 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_452
timestamp 1607639953
transform 1 0 42670 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_476
timestamp 1607639953
transform 1 0 44878 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_464
timestamp 1607639953
transform 1 0 43774 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_501
timestamp 1607639953
transform 1 0 47178 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_489
timestamp 1607639953
transform 1 0 46074 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_991
timestamp 1607639953
transform 1 0 45982 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_525
timestamp 1607639953
transform 1 0 49386 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_513
timestamp 1607639953
transform 1 0 48282 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_550
timestamp 1607639953
transform 1 0 51686 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_537
timestamp 1607639953
transform 1 0 50490 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_992
timestamp 1607639953
transform 1 0 51594 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_562
timestamp 1607639953
transform 1 0 52790 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_586
timestamp 1607639953
transform 1 0 54998 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_574
timestamp 1607639953
transform 1 0 53894 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_611
timestamp 1607639953
transform 1 0 57298 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_598
timestamp 1607639953
transform 1 0 56102 0 1 44064
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_993
timestamp 1607639953
transform 1 0 57206 0 1 44064
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_77_623
timestamp 1607639953
transform 1 0 58402 0 1 44064
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1607639953
transform -1 0 58862 0 1 44064
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_78_14
timestamp 1607639953
transform 1 0 2374 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_3
timestamp 1607639953
transform 1 0 1362 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1607639953
transform 1 0 1086 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _133_
timestamp 1607639953
transform 1 0 2098 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_78_44
timestamp 1607639953
transform 1 0 5134 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_32
timestamp 1607639953
transform 1 0 4030 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_30
timestamp 1607639953
transform 1 0 3846 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_26
timestamp 1607639953
transform 1 0 3478 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_994
timestamp 1607639953
transform 1 0 3938 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_56
timestamp 1607639953
transform 1 0 6238 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_80
timestamp 1607639953
transform 1 0 8446 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_68
timestamp 1607639953
transform 1 0 7342 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_105
timestamp 1607639953
transform 1 0 10746 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_93
timestamp 1607639953
transform 1 0 9642 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_995
timestamp 1607639953
transform 1 0 9550 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_129
timestamp 1607639953
transform 1 0 12954 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_117
timestamp 1607639953
transform 1 0 11850 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_154
timestamp 1607639953
transform 1 0 15254 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_141
timestamp 1607639953
transform 1 0 14058 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_996
timestamp 1607639953
transform 1 0 15162 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_174
timestamp 1607639953
transform 1 0 17094 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_170
timestamp 1607639953
transform 1 0 16726 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_166
timestamp 1607639953
transform 1 0 16358 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__conb_1  _006_
timestamp 1607639953
transform 1 0 16818 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_78_198
timestamp 1607639953
transform 1 0 19302 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_186
timestamp 1607639953
transform 1 0 18198 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_215
timestamp 1607639953
transform 1 0 20866 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_78_210
timestamp 1607639953
transform 1 0 20406 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_997
timestamp 1607639953
transform 1 0 20774 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_239
timestamp 1607639953
transform 1 0 23074 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_227
timestamp 1607639953
transform 1 0 21970 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_255
timestamp 1607639953
transform 1 0 24546 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_251
timestamp 1607639953
transform 1 0 24178 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _099_
timestamp 1607639953
transform 1 0 24270 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_78_276
timestamp 1607639953
transform 1 0 26478 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_78_267
timestamp 1607639953
transform 1 0 25650 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_998
timestamp 1607639953
transform 1 0 26386 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_300
timestamp 1607639953
transform 1 0 28686 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_288
timestamp 1607639953
transform 1 0 27582 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_324
timestamp 1607639953
transform 1 0 30894 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_312
timestamp 1607639953
transform 1 0 29790 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_349
timestamp 1607639953
transform 1 0 33194 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_337
timestamp 1607639953
transform 1 0 32090 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_999
timestamp 1607639953
transform 1 0 31998 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_373
timestamp 1607639953
transform 1 0 35402 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_361
timestamp 1607639953
transform 1 0 34298 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_385
timestamp 1607639953
transform 1 0 36506 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_410
timestamp 1607639953
transform 1 0 38806 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_398
timestamp 1607639953
transform 1 0 37702 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1000
timestamp 1607639953
transform 1 0 37610 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_434
timestamp 1607639953
transform 1 0 41014 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_422
timestamp 1607639953
transform 1 0 39910 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_459
timestamp 1607639953
transform 1 0 43314 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_446
timestamp 1607639953
transform 1 0 42118 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1001
timestamp 1607639953
transform 1 0 43222 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_483
timestamp 1607639953
transform 1 0 45522 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_471
timestamp 1607639953
transform 1 0 44418 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_503
timestamp 1607639953
transform 1 0 47362 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_78_495
timestamp 1607639953
transform 1 0 46626 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _109_
timestamp 1607639953
transform 1 0 47454 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_78_520
timestamp 1607639953
transform 1 0 48926 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_507
timestamp 1607639953
transform 1 0 47730 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1002
timestamp 1607639953
transform 1 0 48834 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_544
timestamp 1607639953
transform 1 0 51134 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_532
timestamp 1607639953
transform 1 0 50030 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_568
timestamp 1607639953
transform 1 0 53342 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_556
timestamp 1607639953
transform 1 0 52238 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_581
timestamp 1607639953
transform 1 0 54538 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1003
timestamp 1607639953
transform 1 0 54446 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _145_
timestamp 1607639953
transform 1 0 55642 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_78_608
timestamp 1607639953
transform 1 0 57022 0 -1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_78_604
timestamp 1607639953
transform 1 0 56654 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_78_596
timestamp 1607639953
transform 1 0 55918 0 -1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _077_
timestamp 1607639953
transform 1 0 56746 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_78_624
timestamp 1607639953
transform 1 0 58494 0 -1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_620
timestamp 1607639953
transform 1 0 58126 0 -1 45152
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1607639953
transform -1 0 58862 0 -1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_80_15
timestamp 1607639953
transform 1 0 2466 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_3
timestamp 1607639953
transform 1 0 1362 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_15
timestamp 1607639953
transform 1 0 2466 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_3
timestamp 1607639953
transform 1 0 1362 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1607639953
transform 1 0 1086 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1607639953
transform 1 0 1086 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_80_44
timestamp 1607639953
transform 1 0 5134 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_32
timestamp 1607639953
transform 1 0 4030 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_27
timestamp 1607639953
transform 1 0 3570 0 -1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_79_39
timestamp 1607639953
transform 1 0 4674 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_27
timestamp 1607639953
transform 1 0 3570 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1014
timestamp 1607639953
transform 1 0 3938 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_56
timestamp 1607639953
transform 1 0 6238 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_62
timestamp 1607639953
transform 1 0 6790 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_79_59
timestamp 1607639953
transform 1 0 6514 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_79_51
timestamp 1607639953
transform 1 0 5778 0 1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1004
timestamp 1607639953
transform 1 0 6698 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_80
timestamp 1607639953
transform 1 0 8446 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_68
timestamp 1607639953
transform 1 0 7342 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_86
timestamp 1607639953
transform 1 0 8998 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_74
timestamp 1607639953
transform 1 0 7894 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_105
timestamp 1607639953
transform 1 0 10746 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_93
timestamp 1607639953
transform 1 0 9642 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_110
timestamp 1607639953
transform 1 0 11206 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_98
timestamp 1607639953
transform 1 0 10102 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1015
timestamp 1607639953
transform 1 0 9550 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_129
timestamp 1607639953
transform 1 0 12954 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_117
timestamp 1607639953
transform 1 0 11850 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_123
timestamp 1607639953
transform 1 0 12402 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1005
timestamp 1607639953
transform 1 0 12310 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_154
timestamp 1607639953
transform 1 0 15254 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_141
timestamp 1607639953
transform 1 0 14058 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_147
timestamp 1607639953
transform 1 0 14610 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_135
timestamp 1607639953
transform 1 0 13506 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1016
timestamp 1607639953
transform 1 0 15162 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_166
timestamp 1607639953
transform 1 0 16358 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_171
timestamp 1607639953
transform 1 0 16818 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_159
timestamp 1607639953
transform 1 0 15714 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_190
timestamp 1607639953
transform 1 0 18566 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_178
timestamp 1607639953
transform 1 0 17462 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_196
timestamp 1607639953
transform 1 0 19118 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_184
timestamp 1607639953
transform 1 0 18014 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1006
timestamp 1607639953
transform 1 0 17922 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_215
timestamp 1607639953
transform 1 0 20866 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_202
timestamp 1607639953
transform 1 0 19670 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_220
timestamp 1607639953
transform 1 0 21326 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_208
timestamp 1607639953
transform 1 0 20222 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1017
timestamp 1607639953
transform 1 0 20774 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_239
timestamp 1607639953
transform 1 0 23074 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_227
timestamp 1607639953
transform 1 0 21970 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_232
timestamp 1607639953
transform 1 0 22430 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_263
timestamp 1607639953
transform 1 0 25282 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_251
timestamp 1607639953
transform 1 0 24178 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_257
timestamp 1607639953
transform 1 0 24730 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_245
timestamp 1607639953
transform 1 0 23626 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1007
timestamp 1607639953
transform 1 0 23534 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_276
timestamp 1607639953
transform 1 0 26478 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_281
timestamp 1607639953
transform 1 0 26938 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_269
timestamp 1607639953
transform 1 0 25834 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1018
timestamp 1607639953
transform 1 0 26386 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_300
timestamp 1607639953
transform 1 0 28686 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_288
timestamp 1607639953
transform 1 0 27582 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_306
timestamp 1607639953
transform 1 0 29238 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_293
timestamp 1607639953
transform 1 0 28042 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1008
timestamp 1607639953
transform 1 0 29146 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_324
timestamp 1607639953
transform 1 0 30894 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_312
timestamp 1607639953
transform 1 0 29790 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_330
timestamp 1607639953
transform 1 0 31446 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_318
timestamp 1607639953
transform 1 0 30342 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_349
timestamp 1607639953
transform 1 0 33194 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_337
timestamp 1607639953
transform 1 0 32090 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_342
timestamp 1607639953
transform 1 0 32550 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1019
timestamp 1607639953
transform 1 0 31998 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_373
timestamp 1607639953
transform 1 0 35402 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_361
timestamp 1607639953
transform 1 0 34298 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_367
timestamp 1607639953
transform 1 0 34850 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_354
timestamp 1607639953
transform 1 0 33654 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1009
timestamp 1607639953
transform 1 0 34758 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_385
timestamp 1607639953
transform 1 0 36506 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_391
timestamp 1607639953
transform 1 0 37058 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_379
timestamp 1607639953
transform 1 0 35954 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_410
timestamp 1607639953
transform 1 0 38806 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_398
timestamp 1607639953
transform 1 0 37702 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_415
timestamp 1607639953
transform 1 0 39266 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_403
timestamp 1607639953
transform 1 0 38162 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1020
timestamp 1607639953
transform 1 0 37610 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_434
timestamp 1607639953
transform 1 0 41014 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_422
timestamp 1607639953
transform 1 0 39910 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_432
timestamp 1607639953
transform 1 0 40830 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_79_428
timestamp 1607639953
transform 1 0 40462 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1010
timestamp 1607639953
transform 1 0 40370 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _116_
timestamp 1607639953
transform 1 0 40554 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_80_459
timestamp 1607639953
transform 1 0 43314 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_446
timestamp 1607639953
transform 1 0 42118 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_456
timestamp 1607639953
transform 1 0 43038 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_444
timestamp 1607639953
transform 1 0 41934 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1021
timestamp 1607639953
transform 1 0 43222 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_483
timestamp 1607639953
transform 1 0 45522 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_471
timestamp 1607639953
transform 1 0 44418 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_79_480
timestamp 1607639953
transform 1 0 45246 0 1 45152
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_79_468
timestamp 1607639953
transform 1 0 44142 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_495
timestamp 1607639953
transform 1 0 46626 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_501
timestamp 1607639953
transform 1 0 47178 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_489
timestamp 1607639953
transform 1 0 46074 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1011
timestamp 1607639953
transform 1 0 45982 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_520
timestamp 1607639953
transform 1 0 48926 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_507
timestamp 1607639953
transform 1 0 47730 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_525
timestamp 1607639953
transform 1 0 49386 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_513
timestamp 1607639953
transform 1 0 48282 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1022
timestamp 1607639953
transform 1 0 48834 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_544
timestamp 1607639953
transform 1 0 51134 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_532
timestamp 1607639953
transform 1 0 50030 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_550
timestamp 1607639953
transform 1 0 51686 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_537
timestamp 1607639953
transform 1 0 50490 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1012
timestamp 1607639953
transform 1 0 51594 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_568
timestamp 1607639953
transform 1 0 53342 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_556
timestamp 1607639953
transform 1 0 52238 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_562
timestamp 1607639953
transform 1 0 52790 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_593
timestamp 1607639953
transform 1 0 55642 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_581
timestamp 1607639953
transform 1 0 54538 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_586
timestamp 1607639953
transform 1 0 54998 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_574
timestamp 1607639953
transform 1 0 53894 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1023
timestamp 1607639953
transform 1 0 54446 0 -1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_605
timestamp 1607639953
transform 1 0 56746 0 -1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_611
timestamp 1607639953
transform 1 0 57298 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_598
timestamp 1607639953
transform 1 0 56102 0 1 45152
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1013
timestamp 1607639953
transform 1 0 57206 0 1 45152
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_80_617
timestamp 1607639953
transform 1 0 57850 0 -1 46240
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_79_623
timestamp 1607639953
transform 1 0 58402 0 1 45152
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1607639953
transform -1 0 58862 0 -1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1607639953
transform -1 0 58862 0 1 45152
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_81_15
timestamp 1607639953
transform 1 0 2466 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_3
timestamp 1607639953
transform 1 0 1362 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1607639953
transform 1 0 1086 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_81_43
timestamp 1607639953
transform 1 0 5042 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_39
timestamp 1607639953
transform 1 0 4674 0 1 46240
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_81_27
timestamp 1607639953
transform 1 0 3570 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _161_
timestamp 1607639953
transform 1 0 5134 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_81_62
timestamp 1607639953
transform 1 0 6790 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_81_59
timestamp 1607639953
transform 1 0 6514 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_81_47
timestamp 1607639953
transform 1 0 5410 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1024
timestamp 1607639953
transform 1 0 6698 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_86
timestamp 1607639953
transform 1 0 8998 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_74
timestamp 1607639953
transform 1 0 7894 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_110
timestamp 1607639953
transform 1 0 11206 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_98
timestamp 1607639953
transform 1 0 10102 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_123
timestamp 1607639953
transform 1 0 12402 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1025
timestamp 1607639953
transform 1 0 12310 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_147
timestamp 1607639953
transform 1 0 14610 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_135
timestamp 1607639953
transform 1 0 13506 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_171
timestamp 1607639953
transform 1 0 16818 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_159
timestamp 1607639953
transform 1 0 15714 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_196
timestamp 1607639953
transform 1 0 19118 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_184
timestamp 1607639953
transform 1 0 18014 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1026
timestamp 1607639953
transform 1 0 17922 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_220
timestamp 1607639953
transform 1 0 21326 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_208
timestamp 1607639953
transform 1 0 20222 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_232
timestamp 1607639953
transform 1 0 22430 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_257
timestamp 1607639953
transform 1 0 24730 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_245
timestamp 1607639953
transform 1 0 23626 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1027
timestamp 1607639953
transform 1 0 23534 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_281
timestamp 1607639953
transform 1 0 26938 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_269
timestamp 1607639953
transform 1 0 25834 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_306
timestamp 1607639953
transform 1 0 29238 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_293
timestamp 1607639953
transform 1 0 28042 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1028
timestamp 1607639953
transform 1 0 29146 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_330
timestamp 1607639953
transform 1 0 31446 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_318
timestamp 1607639953
transform 1 0 30342 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_342
timestamp 1607639953
transform 1 0 32550 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_367
timestamp 1607639953
transform 1 0 34850 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_354
timestamp 1607639953
transform 1 0 33654 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1029
timestamp 1607639953
transform 1 0 34758 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_391
timestamp 1607639953
transform 1 0 37058 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_379
timestamp 1607639953
transform 1 0 35954 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_415
timestamp 1607639953
transform 1 0 39266 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_403
timestamp 1607639953
transform 1 0 38162 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_440
timestamp 1607639953
transform 1 0 41566 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_428
timestamp 1607639953
transform 1 0 40462 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1030
timestamp 1607639953
transform 1 0 40370 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_452
timestamp 1607639953
transform 1 0 42670 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_476
timestamp 1607639953
transform 1 0 44878 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_464
timestamp 1607639953
transform 1 0 43774 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_501
timestamp 1607639953
transform 1 0 47178 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_489
timestamp 1607639953
transform 1 0 46074 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1031
timestamp 1607639953
transform 1 0 45982 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_525
timestamp 1607639953
transform 1 0 49386 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_513
timestamp 1607639953
transform 1 0 48282 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_81_550
timestamp 1607639953
transform 1 0 51686 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_81_537
timestamp 1607639953
transform 1 0 50490 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1032
timestamp 1607639953
transform 1 0 51594 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_567
timestamp 1607639953
transform 1 0 53250 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_555
timestamp 1607639953
transform 1 0 52146 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _135_
timestamp 1607639953
transform 1 0 51870 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_81_591
timestamp 1607639953
transform 1 0 55458 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_579
timestamp 1607639953
transform 1 0 54354 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_611
timestamp 1607639953
transform 1 0 57298 0 1 46240
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_81_609
timestamp 1607639953
transform 1 0 57114 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_81_603
timestamp 1607639953
transform 1 0 56562 0 1 46240
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1033
timestamp 1607639953
transform 1 0 57206 0 1 46240
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_81_623
timestamp 1607639953
transform 1 0 58402 0 1 46240
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1607639953
transform -1 0 58862 0 1 46240
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_15
timestamp 1607639953
transform 1 0 2466 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_3
timestamp 1607639953
transform 1 0 1362 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1607639953
transform 1 0 1086 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_44
timestamp 1607639953
transform 1 0 5134 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_32
timestamp 1607639953
transform 1 0 4030 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_27
timestamp 1607639953
transform 1 0 3570 0 -1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1034
timestamp 1607639953
transform 1 0 3938 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_56
timestamp 1607639953
transform 1 0 6238 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_80
timestamp 1607639953
transform 1 0 8446 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_68
timestamp 1607639953
transform 1 0 7342 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_105
timestamp 1607639953
transform 1 0 10746 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_93
timestamp 1607639953
transform 1 0 9642 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1035
timestamp 1607639953
transform 1 0 9550 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_129
timestamp 1607639953
transform 1 0 12954 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_117
timestamp 1607639953
transform 1 0 11850 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_154
timestamp 1607639953
transform 1 0 15254 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_141
timestamp 1607639953
transform 1 0 14058 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1036
timestamp 1607639953
transform 1 0 15162 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_166
timestamp 1607639953
transform 1 0 16358 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_190
timestamp 1607639953
transform 1 0 18566 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_178
timestamp 1607639953
transform 1 0 17462 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_215
timestamp 1607639953
transform 1 0 20866 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_202
timestamp 1607639953
transform 1 0 19670 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1037
timestamp 1607639953
transform 1 0 20774 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_239
timestamp 1607639953
transform 1 0 23074 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_227
timestamp 1607639953
transform 1 0 21970 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_263
timestamp 1607639953
transform 1 0 25282 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_251
timestamp 1607639953
transform 1 0 24178 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_280
timestamp 1607639953
transform 1 0 26846 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_276
timestamp 1607639953
transform 1 0 26478 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1038
timestamp 1607639953
transform 1 0 26386 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _080_
timestamp 1607639953
transform 1 0 26570 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_304
timestamp 1607639953
transform 1 0 29054 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_292
timestamp 1607639953
transform 1 0 27950 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_328
timestamp 1607639953
transform 1 0 31262 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_82_316
timestamp 1607639953
transform 1 0 30158 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_349
timestamp 1607639953
transform 1 0 33194 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_337
timestamp 1607639953
transform 1 0 32090 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1039
timestamp 1607639953
transform 1 0 31998 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_373
timestamp 1607639953
transform 1 0 35402 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_361
timestamp 1607639953
transform 1 0 34298 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_385
timestamp 1607639953
transform 1 0 36506 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_410
timestamp 1607639953
transform 1 0 38806 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_398
timestamp 1607639953
transform 1 0 37702 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1040
timestamp 1607639953
transform 1 0 37610 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_434
timestamp 1607639953
transform 1 0 41014 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_422
timestamp 1607639953
transform 1 0 39910 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_459
timestamp 1607639953
transform 1 0 43314 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_446
timestamp 1607639953
transform 1 0 42118 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1041
timestamp 1607639953
transform 1 0 43222 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_483
timestamp 1607639953
transform 1 0 45522 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_471
timestamp 1607639953
transform 1 0 44418 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_495
timestamp 1607639953
transform 1 0 46626 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_520
timestamp 1607639953
transform 1 0 48926 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_507
timestamp 1607639953
transform 1 0 47730 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1042
timestamp 1607639953
transform 1 0 48834 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_544
timestamp 1607639953
transform 1 0 51134 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_532
timestamp 1607639953
transform 1 0 50030 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_568
timestamp 1607639953
transform 1 0 53342 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_556
timestamp 1607639953
transform 1 0 52238 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_593
timestamp 1607639953
transform 1 0 55642 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_581
timestamp 1607639953
transform 1 0 54538 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1043
timestamp 1607639953
transform 1 0 54446 0 -1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_605
timestamp 1607639953
transform 1 0 56746 0 -1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_617
timestamp 1607639953
transform 1 0 57850 0 -1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1607639953
transform -1 0 58862 0 -1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_83_15
timestamp 1607639953
transform 1 0 2466 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_3
timestamp 1607639953
transform 1 0 1362 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1607639953
transform 1 0 1086 0 1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_83_39
timestamp 1607639953
transform 1 0 4674 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_27
timestamp 1607639953
transform 1 0 3570 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_62
timestamp 1607639953
transform 1 0 6790 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_83_59
timestamp 1607639953
transform 1 0 6514 0 1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_83_51
timestamp 1607639953
transform 1 0 5778 0 1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1044
timestamp 1607639953
transform 1 0 6698 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_83_86
timestamp 1607639953
transform 1 0 8998 0 1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_83_74
timestamp 1607639953
transform 1 0 7894 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_109
timestamp 1607639953
transform 1 0 11114 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_97
timestamp 1607639953
transform 1 0 10010 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _044_
timestamp 1607639953
transform 1 0 9734 0 1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_83_123
timestamp 1607639953
transform 1 0 12402 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_83_121
timestamp 1607639953
transform 1 0 12218 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1045
timestamp 1607639953
transform 1 0 12310 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_150
timestamp 1607639953
transform 1 0 14886 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_135
timestamp 1607639953
transform 1 0 13506 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _004_
timestamp 1607639953
transform 1 0 14610 0 1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_83_174
timestamp 1607639953
transform 1 0 17094 0 1 47328
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_83_162
timestamp 1607639953
transform 1 0 15990 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_196
timestamp 1607639953
transform 1 0 19118 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_184
timestamp 1607639953
transform 1 0 18014 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_83_182
timestamp 1607639953
transform 1 0 17830 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1046
timestamp 1607639953
transform 1 0 17922 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_220
timestamp 1607639953
transform 1 0 21326 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_208
timestamp 1607639953
transform 1 0 20222 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_232
timestamp 1607639953
transform 1 0 22430 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_257
timestamp 1607639953
transform 1 0 24730 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_245
timestamp 1607639953
transform 1 0 23626 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1047
timestamp 1607639953
transform 1 0 23534 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_281
timestamp 1607639953
transform 1 0 26938 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_269
timestamp 1607639953
transform 1 0 25834 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_306
timestamp 1607639953
transform 1 0 29238 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_293
timestamp 1607639953
transform 1 0 28042 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1048
timestamp 1607639953
transform 1 0 29146 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_330
timestamp 1607639953
transform 1 0 31446 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_318
timestamp 1607639953
transform 1 0 30342 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_342
timestamp 1607639953
transform 1 0 32550 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_367
timestamp 1607639953
transform 1 0 34850 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_354
timestamp 1607639953
transform 1 0 33654 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1049
timestamp 1607639953
transform 1 0 34758 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_391
timestamp 1607639953
transform 1 0 37058 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_379
timestamp 1607639953
transform 1 0 35954 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_415
timestamp 1607639953
transform 1 0 39266 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_403
timestamp 1607639953
transform 1 0 38162 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_440
timestamp 1607639953
transform 1 0 41566 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_428
timestamp 1607639953
transform 1 0 40462 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1050
timestamp 1607639953
transform 1 0 40370 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_452
timestamp 1607639953
transform 1 0 42670 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_83_482
timestamp 1607639953
transform 1 0 45430 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_83_476
timestamp 1607639953
transform 1 0 44878 0 1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_83_464
timestamp 1607639953
transform 1 0 43774 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _036_
timestamp 1607639953
transform 1 0 45522 0 1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_83_501
timestamp 1607639953
transform 1 0 47178 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_489
timestamp 1607639953
transform 1 0 46074 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_83_486
timestamp 1607639953
transform 1 0 45798 0 1 47328
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1051
timestamp 1607639953
transform 1 0 45982 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_525
timestamp 1607639953
transform 1 0 49386 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_513
timestamp 1607639953
transform 1 0 48282 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_550
timestamp 1607639953
transform 1 0 51686 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_537
timestamp 1607639953
transform 1 0 50490 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1052
timestamp 1607639953
transform 1 0 51594 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_83_562
timestamp 1607639953
transform 1 0 52790 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_586
timestamp 1607639953
transform 1 0 54998 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_574
timestamp 1607639953
transform 1 0 53894 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_611
timestamp 1607639953
transform 1 0 57298 0 1 47328
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_83_598
timestamp 1607639953
transform 1 0 56102 0 1 47328
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1053
timestamp 1607639953
transform 1 0 57206 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _008_
timestamp 1607639953
transform 1 0 57666 0 1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_83_624
timestamp 1607639953
transform 1 0 58494 0 1 47328
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_83_618
timestamp 1607639953
transform 1 0 57942 0 1 47328
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1607639953
transform -1 0 58862 0 1 47328
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_84_15
timestamp 1607639953
transform 1 0 2466 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_3
timestamp 1607639953
transform 1 0 1362 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1607639953
transform 1 0 1086 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_84_44
timestamp 1607639953
transform 1 0 5134 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_32
timestamp 1607639953
transform 1 0 4030 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_84_27
timestamp 1607639953
transform 1 0 3570 0 -1 48416
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1054
timestamp 1607639953
transform 1 0 3938 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_56
timestamp 1607639953
transform 1 0 6238 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_80
timestamp 1607639953
transform 1 0 8446 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_68
timestamp 1607639953
transform 1 0 7342 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_105
timestamp 1607639953
transform 1 0 10746 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_93
timestamp 1607639953
transform 1 0 9642 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1055
timestamp 1607639953
transform 1 0 9550 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_129
timestamp 1607639953
transform 1 0 12954 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_117
timestamp 1607639953
transform 1 0 11850 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_154
timestamp 1607639953
transform 1 0 15254 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_141
timestamp 1607639953
transform 1 0 14058 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1056
timestamp 1607639953
transform 1 0 15162 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_172
timestamp 1607639953
transform 1 0 16910 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_84_166
timestamp 1607639953
transform 1 0 16358 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _187_
timestamp 1607639953
transform 1 0 16634 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_84_196
timestamp 1607639953
transform 1 0 19118 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_184
timestamp 1607639953
transform 1 0 18014 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_215
timestamp 1607639953
transform 1 0 20866 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_84_208
timestamp 1607639953
transform 1 0 20222 0 -1 48416
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1057
timestamp 1607639953
transform 1 0 20774 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_239
timestamp 1607639953
transform 1 0 23074 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_227
timestamp 1607639953
transform 1 0 21970 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_263
timestamp 1607639953
transform 1 0 25282 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_251
timestamp 1607639953
transform 1 0 24178 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_276
timestamp 1607639953
transform 1 0 26478 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1058
timestamp 1607639953
transform 1 0 26386 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_300
timestamp 1607639953
transform 1 0 28686 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_288
timestamp 1607639953
transform 1 0 27582 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_324
timestamp 1607639953
transform 1 0 30894 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_312
timestamp 1607639953
transform 1 0 29790 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_349
timestamp 1607639953
transform 1 0 33194 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_337
timestamp 1607639953
transform 1 0 32090 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1059
timestamp 1607639953
transform 1 0 31998 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_373
timestamp 1607639953
transform 1 0 35402 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_361
timestamp 1607639953
transform 1 0 34298 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_385
timestamp 1607639953
transform 1 0 36506 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_410
timestamp 1607639953
transform 1 0 38806 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_398
timestamp 1607639953
transform 1 0 37702 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1060
timestamp 1607639953
transform 1 0 37610 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_434
timestamp 1607639953
transform 1 0 41014 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_422
timestamp 1607639953
transform 1 0 39910 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_459
timestamp 1607639953
transform 1 0 43314 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_446
timestamp 1607639953
transform 1 0 42118 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1061
timestamp 1607639953
transform 1 0 43222 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_483
timestamp 1607639953
transform 1 0 45522 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_471
timestamp 1607639953
transform 1 0 44418 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_495
timestamp 1607639953
transform 1 0 46626 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_520
timestamp 1607639953
transform 1 0 48926 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_507
timestamp 1607639953
transform 1 0 47730 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1062
timestamp 1607639953
transform 1 0 48834 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_544
timestamp 1607639953
transform 1 0 51134 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_532
timestamp 1607639953
transform 1 0 50030 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_568
timestamp 1607639953
transform 1 0 53342 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_556
timestamp 1607639953
transform 1 0 52238 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_593
timestamp 1607639953
transform 1 0 55642 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_581
timestamp 1607639953
transform 1 0 54538 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1063
timestamp 1607639953
transform 1 0 54446 0 -1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_605
timestamp 1607639953
transform 1 0 56746 0 -1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_84_617
timestamp 1607639953
transform 1 0 57850 0 -1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1607639953
transform -1 0 58862 0 -1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_86_15
timestamp 1607639953
transform 1 0 2466 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_3
timestamp 1607639953
transform 1 0 1362 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_15
timestamp 1607639953
transform 1 0 2466 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_3
timestamp 1607639953
transform 1 0 1362 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1607639953
transform 1 0 1086 0 -1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1607639953
transform 1 0 1086 0 1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_86_44
timestamp 1607639953
transform 1 0 5134 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_32
timestamp 1607639953
transform 1 0 4030 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_27
timestamp 1607639953
transform 1 0 3570 0 -1 49504
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_85_39
timestamp 1607639953
transform 1 0 4674 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_27
timestamp 1607639953
transform 1 0 3570 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1074
timestamp 1607639953
transform 1 0 3938 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_56
timestamp 1607639953
transform 1 0 6238 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_62
timestamp 1607639953
transform 1 0 6790 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_85_59
timestamp 1607639953
transform 1 0 6514 0 1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_85_51
timestamp 1607639953
transform 1 0 5778 0 1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1064
timestamp 1607639953
transform 1 0 6698 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_80
timestamp 1607639953
transform 1 0 8446 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_68
timestamp 1607639953
transform 1 0 7342 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_86
timestamp 1607639953
transform 1 0 8998 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_74
timestamp 1607639953
transform 1 0 7894 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_105
timestamp 1607639953
transform 1 0 10746 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_93
timestamp 1607639953
transform 1 0 9642 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_110
timestamp 1607639953
transform 1 0 11206 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_98
timestamp 1607639953
transform 1 0 10102 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1075
timestamp 1607639953
transform 1 0 9550 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_129
timestamp 1607639953
transform 1 0 12954 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_117
timestamp 1607639953
transform 1 0 11850 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_123
timestamp 1607639953
transform 1 0 12402 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1065
timestamp 1607639953
transform 1 0 12310 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_154
timestamp 1607639953
transform 1 0 15254 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_141
timestamp 1607639953
transform 1 0 14058 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_147
timestamp 1607639953
transform 1 0 14610 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_135
timestamp 1607639953
transform 1 0 13506 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1076
timestamp 1607639953
transform 1 0 15162 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_166
timestamp 1607639953
transform 1 0 16358 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_171
timestamp 1607639953
transform 1 0 16818 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_159
timestamp 1607639953
transform 1 0 15714 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_188
timestamp 1607639953
transform 1 0 18382 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_86_184
timestamp 1607639953
transform 1 0 18014 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_86_178
timestamp 1607639953
transform 1 0 17462 0 -1 49504
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_85_196
timestamp 1607639953
transform 1 0 19118 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_184
timestamp 1607639953
transform 1 0 18014 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1066
timestamp 1607639953
transform 1 0 17922 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _202_
timestamp 1607639953
transform 1 0 18106 0 -1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_86_215
timestamp 1607639953
transform 1 0 20866 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_86_212
timestamp 1607639953
transform 1 0 20590 0 -1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_86_200
timestamp 1607639953
transform 1 0 19486 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_220
timestamp 1607639953
transform 1 0 21326 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_208
timestamp 1607639953
transform 1 0 20222 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1077
timestamp 1607639953
transform 1 0 20774 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_239
timestamp 1607639953
transform 1 0 23074 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_227
timestamp 1607639953
transform 1 0 21970 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_232
timestamp 1607639953
transform 1 0 22430 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_263
timestamp 1607639953
transform 1 0 25282 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_251
timestamp 1607639953
transform 1 0 24178 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_257
timestamp 1607639953
transform 1 0 24730 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_245
timestamp 1607639953
transform 1 0 23626 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1067
timestamp 1607639953
transform 1 0 23534 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_276
timestamp 1607639953
transform 1 0 26478 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_281
timestamp 1607639953
transform 1 0 26938 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_269
timestamp 1607639953
transform 1 0 25834 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1078
timestamp 1607639953
transform 1 0 26386 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_300
timestamp 1607639953
transform 1 0 28686 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_288
timestamp 1607639953
transform 1 0 27582 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_306
timestamp 1607639953
transform 1 0 29238 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_293
timestamp 1607639953
transform 1 0 28042 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1068
timestamp 1607639953
transform 1 0 29146 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_324
timestamp 1607639953
transform 1 0 30894 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_312
timestamp 1607639953
transform 1 0 29790 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_330
timestamp 1607639953
transform 1 0 31446 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_318
timestamp 1607639953
transform 1 0 30342 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_86_349
timestamp 1607639953
transform 1 0 33194 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_337
timestamp 1607639953
transform 1 0 32090 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_342
timestamp 1607639953
transform 1 0 32550 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1079
timestamp 1607639953
transform 1 0 31998 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _136_
timestamp 1607639953
transform 1 0 33286 0 -1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_86_365
timestamp 1607639953
transform 1 0 34666 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_353
timestamp 1607639953
transform 1 0 33562 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_367
timestamp 1607639953
transform 1 0 34850 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_354
timestamp 1607639953
transform 1 0 33654 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1069
timestamp 1607639953
transform 1 0 34758 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_86_389
timestamp 1607639953
transform 1 0 36874 0 -1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_86_377
timestamp 1607639953
transform 1 0 35770 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_391
timestamp 1607639953
transform 1 0 37058 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_379
timestamp 1607639953
transform 1 0 35954 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_410
timestamp 1607639953
transform 1 0 38806 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_398
timestamp 1607639953
transform 1 0 37702 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_415
timestamp 1607639953
transform 1 0 39266 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_403
timestamp 1607639953
transform 1 0 38162 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1080
timestamp 1607639953
transform 1 0 37610 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_434
timestamp 1607639953
transform 1 0 41014 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_422
timestamp 1607639953
transform 1 0 39910 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_440
timestamp 1607639953
transform 1 0 41566 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_428
timestamp 1607639953
transform 1 0 40462 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1070
timestamp 1607639953
transform 1 0 40370 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_459
timestamp 1607639953
transform 1 0 43314 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_446
timestamp 1607639953
transform 1 0 42118 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_452
timestamp 1607639953
transform 1 0 42670 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1081
timestamp 1607639953
transform 1 0 43222 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_483
timestamp 1607639953
transform 1 0 45522 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_471
timestamp 1607639953
transform 1 0 44418 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_474
timestamp 1607639953
transform 1 0 44694 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_85_470
timestamp 1607639953
transform 1 0 44326 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_85_464
timestamp 1607639953
transform 1 0 43774 0 1 48416
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  _192_
timestamp 1607639953
transform 1 0 44418 0 1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_86_495
timestamp 1607639953
transform 1 0 46626 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_501
timestamp 1607639953
transform 1 0 47178 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_489
timestamp 1607639953
transform 1 0 46074 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_85_486
timestamp 1607639953
transform 1 0 45798 0 1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1071
timestamp 1607639953
transform 1 0 45982 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_520
timestamp 1607639953
transform 1 0 48926 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_507
timestamp 1607639953
transform 1 0 47730 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_524
timestamp 1607639953
transform 1 0 49294 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_85_513
timestamp 1607639953
transform 1 0 48282 0 1 48416
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1082
timestamp 1607639953
transform 1 0 48834 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _156_
timestamp 1607639953
transform 1 0 49018 0 1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_86_544
timestamp 1607639953
transform 1 0 51134 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_532
timestamp 1607639953
transform 1 0 50030 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_550
timestamp 1607639953
transform 1 0 51686 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_85_548
timestamp 1607639953
transform 1 0 51502 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_85_536
timestamp 1607639953
transform 1 0 50398 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1072
timestamp 1607639953
transform 1 0 51594 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_568
timestamp 1607639953
transform 1 0 53342 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_556
timestamp 1607639953
transform 1 0 52238 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_562
timestamp 1607639953
transform 1 0 52790 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_593
timestamp 1607639953
transform 1 0 55642 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_86_581
timestamp 1607639953
transform 1 0 54538 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_586
timestamp 1607639953
transform 1 0 54998 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_574
timestamp 1607639953
transform 1 0 53894 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1083
timestamp 1607639953
transform 1 0 54446 0 -1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_605
timestamp 1607639953
transform 1 0 56746 0 -1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_611
timestamp 1607639953
transform 1 0 57298 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_85_598
timestamp 1607639953
transform 1 0 56102 0 1 48416
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1073
timestamp 1607639953
transform 1 0 57206 0 1 48416
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_86_617
timestamp 1607639953
transform 1 0 57850 0 -1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_85_623
timestamp 1607639953
transform 1 0 58402 0 1 48416
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1607639953
transform -1 0 58862 0 -1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1607639953
transform -1 0 58862 0 1 48416
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_87_15
timestamp 1607639953
transform 1 0 2466 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_3
timestamp 1607639953
transform 1 0 1362 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_174
timestamp 1607639953
transform 1 0 1086 0 1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_87_39
timestamp 1607639953
transform 1 0 4674 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_27
timestamp 1607639953
transform 1 0 3570 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_62
timestamp 1607639953
transform 1 0 6790 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_87_59
timestamp 1607639953
transform 1 0 6514 0 1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_87_51
timestamp 1607639953
transform 1 0 5778 0 1 49504
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1084
timestamp 1607639953
transform 1 0 6698 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_86
timestamp 1607639953
transform 1 0 8998 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_74
timestamp 1607639953
transform 1 0 7894 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_110
timestamp 1607639953
transform 1 0 11206 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_98
timestamp 1607639953
transform 1 0 10102 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_123
timestamp 1607639953
transform 1 0 12402 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1085
timestamp 1607639953
transform 1 0 12310 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_147
timestamp 1607639953
transform 1 0 14610 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_135
timestamp 1607639953
transform 1 0 13506 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_171
timestamp 1607639953
transform 1 0 16818 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_159
timestamp 1607639953
transform 1 0 15714 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_196
timestamp 1607639953
transform 1 0 19118 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_184
timestamp 1607639953
transform 1 0 18014 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1086
timestamp 1607639953
transform 1 0 17922 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_220
timestamp 1607639953
transform 1 0 21326 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_208
timestamp 1607639953
transform 1 0 20222 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_232
timestamp 1607639953
transform 1 0 22430 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_257
timestamp 1607639953
transform 1 0 24730 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_245
timestamp 1607639953
transform 1 0 23626 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1087
timestamp 1607639953
transform 1 0 23534 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_281
timestamp 1607639953
transform 1 0 26938 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_269
timestamp 1607639953
transform 1 0 25834 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_306
timestamp 1607639953
transform 1 0 29238 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_293
timestamp 1607639953
transform 1 0 28042 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1088
timestamp 1607639953
transform 1 0 29146 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_330
timestamp 1607639953
transform 1 0 31446 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_318
timestamp 1607639953
transform 1 0 30342 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_342
timestamp 1607639953
transform 1 0 32550 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_367
timestamp 1607639953
transform 1 0 34850 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_354
timestamp 1607639953
transform 1 0 33654 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1089
timestamp 1607639953
transform 1 0 34758 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_391
timestamp 1607639953
transform 1 0 37058 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_379
timestamp 1607639953
transform 1 0 35954 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_415
timestamp 1607639953
transform 1 0 39266 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_403
timestamp 1607639953
transform 1 0 38162 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_440
timestamp 1607639953
transform 1 0 41566 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_428
timestamp 1607639953
transform 1 0 40462 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1090
timestamp 1607639953
transform 1 0 40370 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_452
timestamp 1607639953
transform 1 0 42670 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_476
timestamp 1607639953
transform 1 0 44878 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_464
timestamp 1607639953
transform 1 0 43774 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_501
timestamp 1607639953
transform 1 0 47178 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_489
timestamp 1607639953
transform 1 0 46074 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1091
timestamp 1607639953
transform 1 0 45982 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_525
timestamp 1607639953
transform 1 0 49386 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_513
timestamp 1607639953
transform 1 0 48282 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_550
timestamp 1607639953
transform 1 0 51686 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_537
timestamp 1607639953
transform 1 0 50490 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1092
timestamp 1607639953
transform 1 0 51594 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_87_562
timestamp 1607639953
transform 1 0 52790 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_586
timestamp 1607639953
transform 1 0 54998 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_574
timestamp 1607639953
transform 1 0 53894 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_611
timestamp 1607639953
transform 1 0 57298 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_87_598
timestamp 1607639953
transform 1 0 56102 0 1 49504
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1093
timestamp 1607639953
transform 1 0 57206 0 1 49504
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_87_623
timestamp 1607639953
transform 1 0 58402 0 1 49504
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_175
timestamp 1607639953
transform -1 0 58862 0 1 49504
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_88_15
timestamp 1607639953
transform 1 0 2466 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_3
timestamp 1607639953
transform 1 0 1362 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_176
timestamp 1607639953
transform 1 0 1086 0 -1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_88_44
timestamp 1607639953
transform 1 0 5134 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_32
timestamp 1607639953
transform 1 0 4030 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_88_27
timestamp 1607639953
transform 1 0 3570 0 -1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1094
timestamp 1607639953
transform 1 0 3938 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_56
timestamp 1607639953
transform 1 0 6238 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_80
timestamp 1607639953
transform 1 0 8446 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_68
timestamp 1607639953
transform 1 0 7342 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_105
timestamp 1607639953
transform 1 0 10746 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_93
timestamp 1607639953
transform 1 0 9642 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1095
timestamp 1607639953
transform 1 0 9550 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_129
timestamp 1607639953
transform 1 0 12954 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_117
timestamp 1607639953
transform 1 0 11850 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_88_154
timestamp 1607639953
transform 1 0 15254 0 -1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_88_141
timestamp 1607639953
transform 1 0 14058 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1096
timestamp 1607639953
transform 1 0 15162 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_168
timestamp 1607639953
transform 1 0 16542 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_88_162
timestamp 1607639953
transform 1 0 15990 0 -1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _142_
timestamp 1607639953
transform 1 0 16266 0 -1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_88_192
timestamp 1607639953
transform 1 0 18750 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_180
timestamp 1607639953
transform 1 0 17646 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_215
timestamp 1607639953
transform 1 0 20866 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_88_212
timestamp 1607639953
transform 1 0 20590 0 -1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_88_204
timestamp 1607639953
transform 1 0 19854 0 -1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1097
timestamp 1607639953
transform 1 0 20774 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_239
timestamp 1607639953
transform 1 0 23074 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_227
timestamp 1607639953
transform 1 0 21970 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_263
timestamp 1607639953
transform 1 0 25282 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_251
timestamp 1607639953
transform 1 0 24178 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_276
timestamp 1607639953
transform 1 0 26478 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1098
timestamp 1607639953
transform 1 0 26386 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_300
timestamp 1607639953
transform 1 0 28686 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_288
timestamp 1607639953
transform 1 0 27582 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_324
timestamp 1607639953
transform 1 0 30894 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_312
timestamp 1607639953
transform 1 0 29790 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_349
timestamp 1607639953
transform 1 0 33194 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_337
timestamp 1607639953
transform 1 0 32090 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1099
timestamp 1607639953
transform 1 0 31998 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_373
timestamp 1607639953
transform 1 0 35402 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_361
timestamp 1607639953
transform 1 0 34298 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_385
timestamp 1607639953
transform 1 0 36506 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_410
timestamp 1607639953
transform 1 0 38806 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_398
timestamp 1607639953
transform 1 0 37702 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1100
timestamp 1607639953
transform 1 0 37610 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_434
timestamp 1607639953
transform 1 0 41014 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_422
timestamp 1607639953
transform 1 0 39910 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_459
timestamp 1607639953
transform 1 0 43314 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_446
timestamp 1607639953
transform 1 0 42118 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1101
timestamp 1607639953
transform 1 0 43222 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_483
timestamp 1607639953
transform 1 0 45522 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_471
timestamp 1607639953
transform 1 0 44418 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_495
timestamp 1607639953
transform 1 0 46626 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_520
timestamp 1607639953
transform 1 0 48926 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_507
timestamp 1607639953
transform 1 0 47730 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1102
timestamp 1607639953
transform 1 0 48834 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_544
timestamp 1607639953
transform 1 0 51134 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_532
timestamp 1607639953
transform 1 0 50030 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_568
timestamp 1607639953
transform 1 0 53342 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_556
timestamp 1607639953
transform 1 0 52238 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_593
timestamp 1607639953
transform 1 0 55642 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_88_581
timestamp 1607639953
transform 1 0 54538 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1103
timestamp 1607639953
transform 1 0 54446 0 -1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_88_605
timestamp 1607639953
transform 1 0 56746 0 -1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_88_617
timestamp 1607639953
transform 1 0 57850 0 -1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_177
timestamp 1607639953
transform -1 0 58862 0 -1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_89_15
timestamp 1607639953
transform 1 0 2466 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_3
timestamp 1607639953
transform 1 0 1362 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_178
timestamp 1607639953
transform 1 0 1086 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_89_39
timestamp 1607639953
transform 1 0 4674 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_27
timestamp 1607639953
transform 1 0 3570 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_62
timestamp 1607639953
transform 1 0 6790 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_89_59
timestamp 1607639953
transform 1 0 6514 0 1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_89_51
timestamp 1607639953
transform 1 0 5778 0 1 50592
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1104
timestamp 1607639953
transform 1 0 6698 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_86
timestamp 1607639953
transform 1 0 8998 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_74
timestamp 1607639953
transform 1 0 7894 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_110
timestamp 1607639953
transform 1 0 11206 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_98
timestamp 1607639953
transform 1 0 10102 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_123
timestamp 1607639953
transform 1 0 12402 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1105
timestamp 1607639953
transform 1 0 12310 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_147
timestamp 1607639953
transform 1 0 14610 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_135
timestamp 1607639953
transform 1 0 13506 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_171
timestamp 1607639953
transform 1 0 16818 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_159
timestamp 1607639953
transform 1 0 15714 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_196
timestamp 1607639953
transform 1 0 19118 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_184
timestamp 1607639953
transform 1 0 18014 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1106
timestamp 1607639953
transform 1 0 17922 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_220
timestamp 1607639953
transform 1 0 21326 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_208
timestamp 1607639953
transform 1 0 20222 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_232
timestamp 1607639953
transform 1 0 22430 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_257
timestamp 1607639953
transform 1 0 24730 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_245
timestamp 1607639953
transform 1 0 23626 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1107
timestamp 1607639953
transform 1 0 23534 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_281
timestamp 1607639953
transform 1 0 26938 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_269
timestamp 1607639953
transform 1 0 25834 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_306
timestamp 1607639953
transform 1 0 29238 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_293
timestamp 1607639953
transform 1 0 28042 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1108
timestamp 1607639953
transform 1 0 29146 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_330
timestamp 1607639953
transform 1 0 31446 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_318
timestamp 1607639953
transform 1 0 30342 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_342
timestamp 1607639953
transform 1 0 32550 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_367
timestamp 1607639953
transform 1 0 34850 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_354
timestamp 1607639953
transform 1 0 33654 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1109
timestamp 1607639953
transform 1 0 34758 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_391
timestamp 1607639953
transform 1 0 37058 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_379
timestamp 1607639953
transform 1 0 35954 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_415
timestamp 1607639953
transform 1 0 39266 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_403
timestamp 1607639953
transform 1 0 38162 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_440
timestamp 1607639953
transform 1 0 41566 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_428
timestamp 1607639953
transform 1 0 40462 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1110
timestamp 1607639953
transform 1 0 40370 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_452
timestamp 1607639953
transform 1 0 42670 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_476
timestamp 1607639953
transform 1 0 44878 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_464
timestamp 1607639953
transform 1 0 43774 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_89_505
timestamp 1607639953
transform 1 0 47546 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_89_501
timestamp 1607639953
transform 1 0 47178 0 1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_89_489
timestamp 1607639953
transform 1 0 46074 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1111
timestamp 1607639953
transform 1 0 45982 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _015_
timestamp 1607639953
transform 1 0 47638 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_89_521
timestamp 1607639953
transform 1 0 49018 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_509
timestamp 1607639953
transform 1 0 47914 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_550
timestamp 1607639953
transform 1 0 51686 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_89_545
timestamp 1607639953
transform 1 0 51226 0 1 50592
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_89_533
timestamp 1607639953
transform 1 0 50122 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1112
timestamp 1607639953
transform 1 0 51594 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_89_562
timestamp 1607639953
transform 1 0 52790 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_586
timestamp 1607639953
transform 1 0 54998 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_574
timestamp 1607639953
transform 1 0 53894 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_611
timestamp 1607639953
transform 1 0 57298 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_89_598
timestamp 1607639953
transform 1 0 56102 0 1 50592
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1113
timestamp 1607639953
transform 1 0 57206 0 1 50592
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_89_623
timestamp 1607639953
transform 1 0 58402 0 1 50592
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_179
timestamp 1607639953
transform -1 0 58862 0 1 50592
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_90_15
timestamp 1607639953
transform 1 0 2466 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_3
timestamp 1607639953
transform 1 0 1362 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_180
timestamp 1607639953
transform 1 0 1086 0 -1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_90_44
timestamp 1607639953
transform 1 0 5134 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_32
timestamp 1607639953
transform 1 0 4030 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_90_27
timestamp 1607639953
transform 1 0 3570 0 -1 51680
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1114
timestamp 1607639953
transform 1 0 3938 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_56
timestamp 1607639953
transform 1 0 6238 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_90_84
timestamp 1607639953
transform 1 0 8814 0 -1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_90_80
timestamp 1607639953
transform 1 0 8446 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_68
timestamp 1607639953
transform 1 0 7342 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _124_
timestamp 1607639953
transform 1 0 8538 0 -1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_90_105
timestamp 1607639953
transform 1 0 10746 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_93
timestamp 1607639953
transform 1 0 9642 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1115
timestamp 1607639953
transform 1 0 9550 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_129
timestamp 1607639953
transform 1 0 12954 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_117
timestamp 1607639953
transform 1 0 11850 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_154
timestamp 1607639953
transform 1 0 15254 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_141
timestamp 1607639953
transform 1 0 14058 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1116
timestamp 1607639953
transform 1 0 15162 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_166
timestamp 1607639953
transform 1 0 16358 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_190
timestamp 1607639953
transform 1 0 18566 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_178
timestamp 1607639953
transform 1 0 17462 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_215
timestamp 1607639953
transform 1 0 20866 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_202
timestamp 1607639953
transform 1 0 19670 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1117
timestamp 1607639953
transform 1 0 20774 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_239
timestamp 1607639953
transform 1 0 23074 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_227
timestamp 1607639953
transform 1 0 21970 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_263
timestamp 1607639953
transform 1 0 25282 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_251
timestamp 1607639953
transform 1 0 24178 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_276
timestamp 1607639953
transform 1 0 26478 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1118
timestamp 1607639953
transform 1 0 26386 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_300
timestamp 1607639953
transform 1 0 28686 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_288
timestamp 1607639953
transform 1 0 27582 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_324
timestamp 1607639953
transform 1 0 30894 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_312
timestamp 1607639953
transform 1 0 29790 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_349
timestamp 1607639953
transform 1 0 33194 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_337
timestamp 1607639953
transform 1 0 32090 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1119
timestamp 1607639953
transform 1 0 31998 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_373
timestamp 1607639953
transform 1 0 35402 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_361
timestamp 1607639953
transform 1 0 34298 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_385
timestamp 1607639953
transform 1 0 36506 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_410
timestamp 1607639953
transform 1 0 38806 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_398
timestamp 1607639953
transform 1 0 37702 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1120
timestamp 1607639953
transform 1 0 37610 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_434
timestamp 1607639953
transform 1 0 41014 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_422
timestamp 1607639953
transform 1 0 39910 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_459
timestamp 1607639953
transform 1 0 43314 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_446
timestamp 1607639953
transform 1 0 42118 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1121
timestamp 1607639953
transform 1 0 43222 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_483
timestamp 1607639953
transform 1 0 45522 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_471
timestamp 1607639953
transform 1 0 44418 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_495
timestamp 1607639953
transform 1 0 46626 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_520
timestamp 1607639953
transform 1 0 48926 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_507
timestamp 1607639953
transform 1 0 47730 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1122
timestamp 1607639953
transform 1 0 48834 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_544
timestamp 1607639953
transform 1 0 51134 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_532
timestamp 1607639953
transform 1 0 50030 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_568
timestamp 1607639953
transform 1 0 53342 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_556
timestamp 1607639953
transform 1 0 52238 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_593
timestamp 1607639953
transform 1 0 55642 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_90_581
timestamp 1607639953
transform 1 0 54538 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1123
timestamp 1607639953
transform 1 0 54446 0 -1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_90_605
timestamp 1607639953
transform 1 0 56746 0 -1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_90_617
timestamp 1607639953
transform 1 0 57850 0 -1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_181
timestamp 1607639953
transform -1 0 58862 0 -1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_91_15
timestamp 1607639953
transform 1 0 2466 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_3
timestamp 1607639953
transform 1 0 1362 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_182
timestamp 1607639953
transform 1 0 1086 0 1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_91_39
timestamp 1607639953
transform 1 0 4674 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_27
timestamp 1607639953
transform 1 0 3570 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_62
timestamp 1607639953
transform 1 0 6790 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_91_59
timestamp 1607639953
transform 1 0 6514 0 1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_91_51
timestamp 1607639953
transform 1 0 5778 0 1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1124
timestamp 1607639953
transform 1 0 6698 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_86
timestamp 1607639953
transform 1 0 8998 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_74
timestamp 1607639953
transform 1 0 7894 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_110
timestamp 1607639953
transform 1 0 11206 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_98
timestamp 1607639953
transform 1 0 10102 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_123
timestamp 1607639953
transform 1 0 12402 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1125
timestamp 1607639953
transform 1 0 12310 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_147
timestamp 1607639953
transform 1 0 14610 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_135
timestamp 1607639953
transform 1 0 13506 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_171
timestamp 1607639953
transform 1 0 16818 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_159
timestamp 1607639953
transform 1 0 15714 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_196
timestamp 1607639953
transform 1 0 19118 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_184
timestamp 1607639953
transform 1 0 18014 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1126
timestamp 1607639953
transform 1 0 17922 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_220
timestamp 1607639953
transform 1 0 21326 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_208
timestamp 1607639953
transform 1 0 20222 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_232
timestamp 1607639953
transform 1 0 22430 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_257
timestamp 1607639953
transform 1 0 24730 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_245
timestamp 1607639953
transform 1 0 23626 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1127
timestamp 1607639953
transform 1 0 23534 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_281
timestamp 1607639953
transform 1 0 26938 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_269
timestamp 1607639953
transform 1 0 25834 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_306
timestamp 1607639953
transform 1 0 29238 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_293
timestamp 1607639953
transform 1 0 28042 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1128
timestamp 1607639953
transform 1 0 29146 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_330
timestamp 1607639953
transform 1 0 31446 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_318
timestamp 1607639953
transform 1 0 30342 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_342
timestamp 1607639953
transform 1 0 32550 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_367
timestamp 1607639953
transform 1 0 34850 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_354
timestamp 1607639953
transform 1 0 33654 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1129
timestamp 1607639953
transform 1 0 34758 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_391
timestamp 1607639953
transform 1 0 37058 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_379
timestamp 1607639953
transform 1 0 35954 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_415
timestamp 1607639953
transform 1 0 39266 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_403
timestamp 1607639953
transform 1 0 38162 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_440
timestamp 1607639953
transform 1 0 41566 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_428
timestamp 1607639953
transform 1 0 40462 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1130
timestamp 1607639953
transform 1 0 40370 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_452
timestamp 1607639953
transform 1 0 42670 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_476
timestamp 1607639953
transform 1 0 44878 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_464
timestamp 1607639953
transform 1 0 43774 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_501
timestamp 1607639953
transform 1 0 47178 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_489
timestamp 1607639953
transform 1 0 46074 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1131
timestamp 1607639953
transform 1 0 45982 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_525
timestamp 1607639953
transform 1 0 49386 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_513
timestamp 1607639953
transform 1 0 48282 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_550
timestamp 1607639953
transform 1 0 51686 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_537
timestamp 1607639953
transform 1 0 50490 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1132
timestamp 1607639953
transform 1 0 51594 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_91_562
timestamp 1607639953
transform 1 0 52790 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_586
timestamp 1607639953
transform 1 0 54998 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_91_574
timestamp 1607639953
transform 1 0 53894 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_91_611
timestamp 1607639953
transform 1 0 57298 0 1 51680
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_91_598
timestamp 1607639953
transform 1 0 56102 0 1 51680
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1133
timestamp 1607639953
transform 1 0 57206 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_91_624
timestamp 1607639953
transform 1 0 58494 0 1 51680
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_91_619
timestamp 1607639953
transform 1 0 58034 0 1 51680
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_183
timestamp 1607639953
transform -1 0 58862 0 1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _112_
timestamp 1607639953
transform 1 0 58218 0 1 51680
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_93_15
timestamp 1607639953
transform 1 0 2466 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_3
timestamp 1607639953
transform 1 0 1362 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_15
timestamp 1607639953
transform 1 0 2466 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_3
timestamp 1607639953
transform 1 0 1362 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_186
timestamp 1607639953
transform 1 0 1086 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_184
timestamp 1607639953
transform 1 0 1086 0 -1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_93_39
timestamp 1607639953
transform 1 0 4674 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_27
timestamp 1607639953
transform 1 0 3570 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_44
timestamp 1607639953
transform 1 0 5134 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_32
timestamp 1607639953
transform 1 0 4030 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_92_27
timestamp 1607639953
transform 1 0 3570 0 -1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1134
timestamp 1607639953
transform 1 0 3938 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_62
timestamp 1607639953
transform 1 0 6790 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_93_59
timestamp 1607639953
transform 1 0 6514 0 1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_93_51
timestamp 1607639953
transform 1 0 5778 0 1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_92_56
timestamp 1607639953
transform 1 0 6238 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1144
timestamp 1607639953
transform 1 0 6698 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_86
timestamp 1607639953
transform 1 0 8998 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_74
timestamp 1607639953
transform 1 0 7894 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_80
timestamp 1607639953
transform 1 0 8446 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_68
timestamp 1607639953
transform 1 0 7342 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_110
timestamp 1607639953
transform 1 0 11206 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_98
timestamp 1607639953
transform 1 0 10102 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_105
timestamp 1607639953
transform 1 0 10746 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_93
timestamp 1607639953
transform 1 0 9642 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1135
timestamp 1607639953
transform 1 0 9550 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_123
timestamp 1607639953
transform 1 0 12402 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_129
timestamp 1607639953
transform 1 0 12954 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_117
timestamp 1607639953
transform 1 0 11850 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1145
timestamp 1607639953
transform 1 0 12310 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_147
timestamp 1607639953
transform 1 0 14610 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_135
timestamp 1607639953
transform 1 0 13506 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_154
timestamp 1607639953
transform 1 0 15254 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_141
timestamp 1607639953
transform 1 0 14058 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1136
timestamp 1607639953
transform 1 0 15162 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_93_174
timestamp 1607639953
transform 1 0 17094 0 1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_93_159
timestamp 1607639953
transform 1 0 15714 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_166
timestamp 1607639953
transform 1 0 16358 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _042_
timestamp 1607639953
transform 1 0 16818 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_93_196
timestamp 1607639953
transform 1 0 19118 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_184
timestamp 1607639953
transform 1 0 18014 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_93_182
timestamp 1607639953
transform 1 0 17830 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_92_198
timestamp 1607639953
transform 1 0 19302 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_92_194
timestamp 1607639953
transform 1 0 18934 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_92_190
timestamp 1607639953
transform 1 0 18566 0 -1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_92_178
timestamp 1607639953
transform 1 0 17462 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1146
timestamp 1607639953
transform 1 0 17922 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _072_
timestamp 1607639953
transform 1 0 19026 0 -1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_93_220
timestamp 1607639953
transform 1 0 21326 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_208
timestamp 1607639953
transform 1 0 20222 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_215
timestamp 1607639953
transform 1 0 20866 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_92_210
timestamp 1607639953
transform 1 0 20406 0 -1 52768
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1137
timestamp 1607639953
transform 1 0 20774 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_232
timestamp 1607639953
transform 1 0 22430 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_239
timestamp 1607639953
transform 1 0 23074 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_227
timestamp 1607639953
transform 1 0 21970 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_257
timestamp 1607639953
transform 1 0 24730 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_245
timestamp 1607639953
transform 1 0 23626 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_263
timestamp 1607639953
transform 1 0 25282 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_251
timestamp 1607639953
transform 1 0 24178 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1147
timestamp 1607639953
transform 1 0 23534 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_281
timestamp 1607639953
transform 1 0 26938 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_269
timestamp 1607639953
transform 1 0 25834 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_276
timestamp 1607639953
transform 1 0 26478 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1138
timestamp 1607639953
transform 1 0 26386 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_306
timestamp 1607639953
transform 1 0 29238 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_293
timestamp 1607639953
transform 1 0 28042 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_300
timestamp 1607639953
transform 1 0 28686 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_288
timestamp 1607639953
transform 1 0 27582 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1148
timestamp 1607639953
transform 1 0 29146 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_330
timestamp 1607639953
transform 1 0 31446 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_318
timestamp 1607639953
transform 1 0 30342 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_324
timestamp 1607639953
transform 1 0 30894 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_312
timestamp 1607639953
transform 1 0 29790 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_342
timestamp 1607639953
transform 1 0 32550 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_349
timestamp 1607639953
transform 1 0 33194 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_337
timestamp 1607639953
transform 1 0 32090 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1139
timestamp 1607639953
transform 1 0 31998 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_367
timestamp 1607639953
transform 1 0 34850 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_354
timestamp 1607639953
transform 1 0 33654 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_373
timestamp 1607639953
transform 1 0 35402 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_361
timestamp 1607639953
transform 1 0 34298 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1149
timestamp 1607639953
transform 1 0 34758 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_93_391
timestamp 1607639953
transform 1 0 37058 0 1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_93_379
timestamp 1607639953
transform 1 0 35954 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_385
timestamp 1607639953
transform 1 0 36506 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_93_417
timestamp 1607639953
transform 1 0 39450 0 1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_93_405
timestamp 1607639953
transform 1 0 38346 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_93_399
timestamp 1607639953
transform 1 0 37794 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_92_410
timestamp 1607639953
transform 1 0 38806 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_398
timestamp 1607639953
transform 1 0 37702 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1140
timestamp 1607639953
transform 1 0 37610 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _043_
timestamp 1607639953
transform 1 0 38070 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_93_440
timestamp 1607639953
transform 1 0 41566 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_428
timestamp 1607639953
transform 1 0 40462 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_93_425
timestamp 1607639953
transform 1 0 40186 0 1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_92_434
timestamp 1607639953
transform 1 0 41014 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_422
timestamp 1607639953
transform 1 0 39910 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1150
timestamp 1607639953
transform 1 0 40370 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_452
timestamp 1607639953
transform 1 0 42670 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_459
timestamp 1607639953
transform 1 0 43314 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_446
timestamp 1607639953
transform 1 0 42118 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1141
timestamp 1607639953
transform 1 0 43222 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_476
timestamp 1607639953
transform 1 0 44878 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_464
timestamp 1607639953
transform 1 0 43774 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_483
timestamp 1607639953
transform 1 0 45522 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_471
timestamp 1607639953
transform 1 0 44418 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_506
timestamp 1607639953
transform 1 0 47638 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_93_501
timestamp 1607639953
transform 1 0 47178 0 1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_93_489
timestamp 1607639953
transform 1 0 46074 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_495
timestamp 1607639953
transform 1 0 46626 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1151
timestamp 1607639953
transform 1 0 45982 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _096_
timestamp 1607639953
transform 1 0 47362 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_93_518
timestamp 1607639953
transform 1 0 48742 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_520
timestamp 1607639953
transform 1 0 48926 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_507
timestamp 1607639953
transform 1 0 47730 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1142
timestamp 1607639953
transform 1 0 48834 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_550
timestamp 1607639953
transform 1 0 51686 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_93_548
timestamp 1607639953
transform 1 0 51502 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_93_542
timestamp 1607639953
transform 1 0 50950 0 1 52768
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_93_530
timestamp 1607639953
transform 1 0 49846 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_544
timestamp 1607639953
transform 1 0 51134 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_532
timestamp 1607639953
transform 1 0 50030 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1152
timestamp 1607639953
transform 1 0 51594 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_562
timestamp 1607639953
transform 1 0 52790 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_568
timestamp 1607639953
transform 1 0 53342 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_556
timestamp 1607639953
transform 1 0 52238 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_586
timestamp 1607639953
transform 1 0 54998 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_574
timestamp 1607639953
transform 1 0 53894 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_593
timestamp 1607639953
transform 1 0 55642 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_581
timestamp 1607639953
transform 1 0 54538 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1143
timestamp 1607639953
transform 1 0 54446 0 -1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_93_611
timestamp 1607639953
transform 1 0 57298 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_93_598
timestamp 1607639953
transform 1 0 56102 0 1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_92_605
timestamp 1607639953
transform 1 0 56746 0 -1 52768
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1153
timestamp 1607639953
transform 1 0 57206 0 1 52768
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_93_623
timestamp 1607639953
transform 1 0 58402 0 1 52768
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_92_617
timestamp 1607639953
transform 1 0 57850 0 -1 52768
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_187
timestamp 1607639953
transform -1 0 58862 0 1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_185
timestamp 1607639953
transform -1 0 58862 0 -1 52768
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_94_15
timestamp 1607639953
transform 1 0 2466 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_3
timestamp 1607639953
transform 1 0 1362 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_188
timestamp 1607639953
transform 1 0 1086 0 -1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_94_44
timestamp 1607639953
transform 1 0 5134 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_32
timestamp 1607639953
transform 1 0 4030 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_94_27
timestamp 1607639953
transform 1 0 3570 0 -1 53856
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1154
timestamp 1607639953
transform 1 0 3938 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_56
timestamp 1607639953
transform 1 0 6238 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_80
timestamp 1607639953
transform 1 0 8446 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_68
timestamp 1607639953
transform 1 0 7342 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_105
timestamp 1607639953
transform 1 0 10746 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_93
timestamp 1607639953
transform 1 0 9642 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1155
timestamp 1607639953
transform 1 0 9550 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_129
timestamp 1607639953
transform 1 0 12954 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_117
timestamp 1607639953
transform 1 0 11850 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_154
timestamp 1607639953
transform 1 0 15254 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_141
timestamp 1607639953
transform 1 0 14058 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1156
timestamp 1607639953
transform 1 0 15162 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_166
timestamp 1607639953
transform 1 0 16358 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_190
timestamp 1607639953
transform 1 0 18566 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_178
timestamp 1607639953
transform 1 0 17462 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_215
timestamp 1607639953
transform 1 0 20866 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_202
timestamp 1607639953
transform 1 0 19670 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1157
timestamp 1607639953
transform 1 0 20774 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_239
timestamp 1607639953
transform 1 0 23074 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_227
timestamp 1607639953
transform 1 0 21970 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_263
timestamp 1607639953
transform 1 0 25282 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_251
timestamp 1607639953
transform 1 0 24178 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_276
timestamp 1607639953
transform 1 0 26478 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1158
timestamp 1607639953
transform 1 0 26386 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_300
timestamp 1607639953
transform 1 0 28686 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_288
timestamp 1607639953
transform 1 0 27582 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_324
timestamp 1607639953
transform 1 0 30894 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_312
timestamp 1607639953
transform 1 0 29790 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_349
timestamp 1607639953
transform 1 0 33194 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_337
timestamp 1607639953
transform 1 0 32090 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1159
timestamp 1607639953
transform 1 0 31998 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_373
timestamp 1607639953
transform 1 0 35402 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_361
timestamp 1607639953
transform 1 0 34298 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_385
timestamp 1607639953
transform 1 0 36506 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_410
timestamp 1607639953
transform 1 0 38806 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_398
timestamp 1607639953
transform 1 0 37702 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1160
timestamp 1607639953
transform 1 0 37610 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_434
timestamp 1607639953
transform 1 0 41014 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_422
timestamp 1607639953
transform 1 0 39910 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_459
timestamp 1607639953
transform 1 0 43314 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_446
timestamp 1607639953
transform 1 0 42118 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1161
timestamp 1607639953
transform 1 0 43222 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_483
timestamp 1607639953
transform 1 0 45522 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_471
timestamp 1607639953
transform 1 0 44418 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_495
timestamp 1607639953
transform 1 0 46626 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_520
timestamp 1607639953
transform 1 0 48926 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_507
timestamp 1607639953
transform 1 0 47730 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1162
timestamp 1607639953
transform 1 0 48834 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_544
timestamp 1607639953
transform 1 0 51134 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_532
timestamp 1607639953
transform 1 0 50030 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_568
timestamp 1607639953
transform 1 0 53342 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_556
timestamp 1607639953
transform 1 0 52238 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_593
timestamp 1607639953
transform 1 0 55642 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_94_581
timestamp 1607639953
transform 1 0 54538 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1163
timestamp 1607639953
transform 1 0 54446 0 -1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_94_605
timestamp 1607639953
transform 1 0 56746 0 -1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_94_623
timestamp 1607639953
transform 1 0 58402 0 -1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_94_617
timestamp 1607639953
transform 1 0 57850 0 -1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_189
timestamp 1607639953
transform -1 0 58862 0 -1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _057_
timestamp 1607639953
transform 1 0 58126 0 -1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_95_15
timestamp 1607639953
transform 1 0 2466 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_3
timestamp 1607639953
transform 1 0 1362 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_190
timestamp 1607639953
transform 1 0 1086 0 1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_95_39
timestamp 1607639953
transform 1 0 4674 0 1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_95_27
timestamp 1607639953
transform 1 0 3570 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_62
timestamp 1607639953
transform 1 0 6790 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_95_59
timestamp 1607639953
transform 1 0 6514 0 1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_95_51
timestamp 1607639953
transform 1 0 5778 0 1 53856
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_95_47
timestamp 1607639953
transform 1 0 5410 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1164
timestamp 1607639953
transform 1 0 6698 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _157_
timestamp 1607639953
transform 1 0 5502 0 1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_95_86
timestamp 1607639953
transform 1 0 8998 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_74
timestamp 1607639953
transform 1 0 7894 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_110
timestamp 1607639953
transform 1 0 11206 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_98
timestamp 1607639953
transform 1 0 10102 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_123
timestamp 1607639953
transform 1 0 12402 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1165
timestamp 1607639953
transform 1 0 12310 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_147
timestamp 1607639953
transform 1 0 14610 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_135
timestamp 1607639953
transform 1 0 13506 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_171
timestamp 1607639953
transform 1 0 16818 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_159
timestamp 1607639953
transform 1 0 15714 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_196
timestamp 1607639953
transform 1 0 19118 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_184
timestamp 1607639953
transform 1 0 18014 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1166
timestamp 1607639953
transform 1 0 17922 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_220
timestamp 1607639953
transform 1 0 21326 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_208
timestamp 1607639953
transform 1 0 20222 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_232
timestamp 1607639953
transform 1 0 22430 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_257
timestamp 1607639953
transform 1 0 24730 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_245
timestamp 1607639953
transform 1 0 23626 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1167
timestamp 1607639953
transform 1 0 23534 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_281
timestamp 1607639953
transform 1 0 26938 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_269
timestamp 1607639953
transform 1 0 25834 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_306
timestamp 1607639953
transform 1 0 29238 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_293
timestamp 1607639953
transform 1 0 28042 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1168
timestamp 1607639953
transform 1 0 29146 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_330
timestamp 1607639953
transform 1 0 31446 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_318
timestamp 1607639953
transform 1 0 30342 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_342
timestamp 1607639953
transform 1 0 32550 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_367
timestamp 1607639953
transform 1 0 34850 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_354
timestamp 1607639953
transform 1 0 33654 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1169
timestamp 1607639953
transform 1 0 34758 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_391
timestamp 1607639953
transform 1 0 37058 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_379
timestamp 1607639953
transform 1 0 35954 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_415
timestamp 1607639953
transform 1 0 39266 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_403
timestamp 1607639953
transform 1 0 38162 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_440
timestamp 1607639953
transform 1 0 41566 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_428
timestamp 1607639953
transform 1 0 40462 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1170
timestamp 1607639953
transform 1 0 40370 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_452
timestamp 1607639953
transform 1 0 42670 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_476
timestamp 1607639953
transform 1 0 44878 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_464
timestamp 1607639953
transform 1 0 43774 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_501
timestamp 1607639953
transform 1 0 47178 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_489
timestamp 1607639953
transform 1 0 46074 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1171
timestamp 1607639953
transform 1 0 45982 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_525
timestamp 1607639953
transform 1 0 49386 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_513
timestamp 1607639953
transform 1 0 48282 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_550
timestamp 1607639953
transform 1 0 51686 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_537
timestamp 1607639953
transform 1 0 50490 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1172
timestamp 1607639953
transform 1 0 51594 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_95_562
timestamp 1607639953
transform 1 0 52790 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_586
timestamp 1607639953
transform 1 0 54998 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_574
timestamp 1607639953
transform 1 0 53894 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_611
timestamp 1607639953
transform 1 0 57298 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_95_598
timestamp 1607639953
transform 1 0 56102 0 1 53856
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1173
timestamp 1607639953
transform 1 0 57206 0 1 53856
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_95_623
timestamp 1607639953
transform 1 0 58402 0 1 53856
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_191
timestamp 1607639953
transform -1 0 58862 0 1 53856
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_96_15
timestamp 1607639953
transform 1 0 2466 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_3
timestamp 1607639953
transform 1 0 1362 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_192
timestamp 1607639953
transform 1 0 1086 0 -1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_96_44
timestamp 1607639953
transform 1 0 5134 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_32
timestamp 1607639953
transform 1 0 4030 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_96_27
timestamp 1607639953
transform 1 0 3570 0 -1 54944
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1174
timestamp 1607639953
transform 1 0 3938 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_56
timestamp 1607639953
transform 1 0 6238 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_80
timestamp 1607639953
transform 1 0 8446 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_68
timestamp 1607639953
transform 1 0 7342 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_105
timestamp 1607639953
transform 1 0 10746 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_93
timestamp 1607639953
transform 1 0 9642 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1175
timestamp 1607639953
transform 1 0 9550 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_129
timestamp 1607639953
transform 1 0 12954 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_117
timestamp 1607639953
transform 1 0 11850 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_154
timestamp 1607639953
transform 1 0 15254 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_141
timestamp 1607639953
transform 1 0 14058 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1176
timestamp 1607639953
transform 1 0 15162 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_96_174
timestamp 1607639953
transform 1 0 17094 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_96_166
timestamp 1607639953
transform 1 0 16358 0 -1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _163_
timestamp 1607639953
transform 1 0 17186 0 -1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_96_190
timestamp 1607639953
transform 1 0 18566 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_178
timestamp 1607639953
transform 1 0 17462 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_96_215
timestamp 1607639953
transform 1 0 20866 0 -1 54944
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_96_202
timestamp 1607639953
transform 1 0 19670 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1177
timestamp 1607639953
transform 1 0 20774 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_236
timestamp 1607639953
transform 1 0 22798 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_224
timestamp 1607639953
transform 1 0 21694 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _149_
timestamp 1607639953
transform 1 0 21418 0 -1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_96_264
timestamp 1607639953
transform 1 0 25374 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_96_260
timestamp 1607639953
transform 1 0 25006 0 -1 54944
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_96_248
timestamp 1607639953
transform 1 0 23902 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_276
timestamp 1607639953
transform 1 0 26478 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_96_274
timestamp 1607639953
transform 1 0 26294 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_96_268
timestamp 1607639953
transform 1 0 25742 0 -1 54944
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1178
timestamp 1607639953
transform 1 0 26386 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _019_
timestamp 1607639953
transform 1 0 25466 0 -1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_96_300
timestamp 1607639953
transform 1 0 28686 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_288
timestamp 1607639953
transform 1 0 27582 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_324
timestamp 1607639953
transform 1 0 30894 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_312
timestamp 1607639953
transform 1 0 29790 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_349
timestamp 1607639953
transform 1 0 33194 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_337
timestamp 1607639953
transform 1 0 32090 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1179
timestamp 1607639953
transform 1 0 31998 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_373
timestamp 1607639953
transform 1 0 35402 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_361
timestamp 1607639953
transform 1 0 34298 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_385
timestamp 1607639953
transform 1 0 36506 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_410
timestamp 1607639953
transform 1 0 38806 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_398
timestamp 1607639953
transform 1 0 37702 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1180
timestamp 1607639953
transform 1 0 37610 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_434
timestamp 1607639953
transform 1 0 41014 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_422
timestamp 1607639953
transform 1 0 39910 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_459
timestamp 1607639953
transform 1 0 43314 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_96_450
timestamp 1607639953
transform 1 0 42486 0 -1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_96_446
timestamp 1607639953
transform 1 0 42118 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1181
timestamp 1607639953
transform 1 0 43222 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _062_
timestamp 1607639953
transform 1 0 42210 0 -1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_96_483
timestamp 1607639953
transform 1 0 45522 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_471
timestamp 1607639953
transform 1 0 44418 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_96_503
timestamp 1607639953
transform 1 0 47362 0 -1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_96_495
timestamp 1607639953
transform 1 0 46626 0 -1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  _207_
timestamp 1607639953
transform 1 0 47638 0 -1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_96_520
timestamp 1607639953
transform 1 0 48926 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_96_517
timestamp 1607639953
transform 1 0 48650 0 -1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_96_509
timestamp 1607639953
transform 1 0 47914 0 -1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1182
timestamp 1607639953
transform 1 0 48834 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_544
timestamp 1607639953
transform 1 0 51134 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_532
timestamp 1607639953
transform 1 0 50030 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_568
timestamp 1607639953
transform 1 0 53342 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_556
timestamp 1607639953
transform 1 0 52238 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_593
timestamp 1607639953
transform 1 0 55642 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_96_581
timestamp 1607639953
transform 1 0 54538 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1183
timestamp 1607639953
transform 1 0 54446 0 -1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_96_605
timestamp 1607639953
transform 1 0 56746 0 -1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_96_617
timestamp 1607639953
transform 1 0 57850 0 -1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_193
timestamp 1607639953
transform -1 0 58862 0 -1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_97_15
timestamp 1607639953
transform 1 0 2466 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_3
timestamp 1607639953
transform 1 0 1362 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_194
timestamp 1607639953
transform 1 0 1086 0 1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_97_39
timestamp 1607639953
transform 1 0 4674 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_27
timestamp 1607639953
transform 1 0 3570 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_62
timestamp 1607639953
transform 1 0 6790 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_97_59
timestamp 1607639953
transform 1 0 6514 0 1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_97_51
timestamp 1607639953
transform 1 0 5778 0 1 54944
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1184
timestamp 1607639953
transform 1 0 6698 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_86
timestamp 1607639953
transform 1 0 8998 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_74
timestamp 1607639953
transform 1 0 7894 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_110
timestamp 1607639953
transform 1 0 11206 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_98
timestamp 1607639953
transform 1 0 10102 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_123
timestamp 1607639953
transform 1 0 12402 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1185
timestamp 1607639953
transform 1 0 12310 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_147
timestamp 1607639953
transform 1 0 14610 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_135
timestamp 1607639953
transform 1 0 13506 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_171
timestamp 1607639953
transform 1 0 16818 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_159
timestamp 1607639953
transform 1 0 15714 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_196
timestamp 1607639953
transform 1 0 19118 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_184
timestamp 1607639953
transform 1 0 18014 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1186
timestamp 1607639953
transform 1 0 17922 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_220
timestamp 1607639953
transform 1 0 21326 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_208
timestamp 1607639953
transform 1 0 20222 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_232
timestamp 1607639953
transform 1 0 22430 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_257
timestamp 1607639953
transform 1 0 24730 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_245
timestamp 1607639953
transform 1 0 23626 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1187
timestamp 1607639953
transform 1 0 23534 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_281
timestamp 1607639953
transform 1 0 26938 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_269
timestamp 1607639953
transform 1 0 25834 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_306
timestamp 1607639953
transform 1 0 29238 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_293
timestamp 1607639953
transform 1 0 28042 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1188
timestamp 1607639953
transform 1 0 29146 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_330
timestamp 1607639953
transform 1 0 31446 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_318
timestamp 1607639953
transform 1 0 30342 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_342
timestamp 1607639953
transform 1 0 32550 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_367
timestamp 1607639953
transform 1 0 34850 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_354
timestamp 1607639953
transform 1 0 33654 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1189
timestamp 1607639953
transform 1 0 34758 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_391
timestamp 1607639953
transform 1 0 37058 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_379
timestamp 1607639953
transform 1 0 35954 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_415
timestamp 1607639953
transform 1 0 39266 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_403
timestamp 1607639953
transform 1 0 38162 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_440
timestamp 1607639953
transform 1 0 41566 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_428
timestamp 1607639953
transform 1 0 40462 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1190
timestamp 1607639953
transform 1 0 40370 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_452
timestamp 1607639953
transform 1 0 42670 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_476
timestamp 1607639953
transform 1 0 44878 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_464
timestamp 1607639953
transform 1 0 43774 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_501
timestamp 1607639953
transform 1 0 47178 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_489
timestamp 1607639953
transform 1 0 46074 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1191
timestamp 1607639953
transform 1 0 45982 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_525
timestamp 1607639953
transform 1 0 49386 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_513
timestamp 1607639953
transform 1 0 48282 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_550
timestamp 1607639953
transform 1 0 51686 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_537
timestamp 1607639953
transform 1 0 50490 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1192
timestamp 1607639953
transform 1 0 51594 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_97_562
timestamp 1607639953
transform 1 0 52790 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_586
timestamp 1607639953
transform 1 0 54998 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_574
timestamp 1607639953
transform 1 0 53894 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_611
timestamp 1607639953
transform 1 0 57298 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_97_598
timestamp 1607639953
transform 1 0 56102 0 1 54944
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1193
timestamp 1607639953
transform 1 0 57206 0 1 54944
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_97_623
timestamp 1607639953
transform 1 0 58402 0 1 54944
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_195
timestamp 1607639953
transform -1 0 58862 0 1 54944
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_98_15
timestamp 1607639953
transform 1 0 2466 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_3
timestamp 1607639953
transform 1 0 1362 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_196
timestamp 1607639953
transform 1 0 1086 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_98_44
timestamp 1607639953
transform 1 0 5134 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_98_40
timestamp 1607639953
transform 1 0 4766 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_98_32
timestamp 1607639953
transform 1 0 4030 0 -1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_98_27
timestamp 1607639953
transform 1 0 3570 0 -1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1194
timestamp 1607639953
transform 1 0 3938 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _123_
timestamp 1607639953
transform 1 0 4858 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_98_56
timestamp 1607639953
transform 1 0 6238 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_80
timestamp 1607639953
transform 1 0 8446 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_68
timestamp 1607639953
transform 1 0 7342 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_105
timestamp 1607639953
transform 1 0 10746 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_93
timestamp 1607639953
transform 1 0 9642 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1195
timestamp 1607639953
transform 1 0 9550 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_129
timestamp 1607639953
transform 1 0 12954 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_117
timestamp 1607639953
transform 1 0 11850 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_154
timestamp 1607639953
transform 1 0 15254 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_141
timestamp 1607639953
transform 1 0 14058 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1196
timestamp 1607639953
transform 1 0 15162 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_166
timestamp 1607639953
transform 1 0 16358 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_190
timestamp 1607639953
transform 1 0 18566 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_178
timestamp 1607639953
transform 1 0 17462 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_215
timestamp 1607639953
transform 1 0 20866 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_202
timestamp 1607639953
transform 1 0 19670 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1197
timestamp 1607639953
transform 1 0 20774 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_239
timestamp 1607639953
transform 1 0 23074 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_227
timestamp 1607639953
transform 1 0 21970 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_263
timestamp 1607639953
transform 1 0 25282 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_251
timestamp 1607639953
transform 1 0 24178 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_276
timestamp 1607639953
transform 1 0 26478 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1198
timestamp 1607639953
transform 1 0 26386 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_300
timestamp 1607639953
transform 1 0 28686 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_288
timestamp 1607639953
transform 1 0 27582 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_324
timestamp 1607639953
transform 1 0 30894 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_312
timestamp 1607639953
transform 1 0 29790 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_349
timestamp 1607639953
transform 1 0 33194 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_337
timestamp 1607639953
transform 1 0 32090 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1199
timestamp 1607639953
transform 1 0 31998 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_373
timestamp 1607639953
transform 1 0 35402 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_361
timestamp 1607639953
transform 1 0 34298 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_385
timestamp 1607639953
transform 1 0 36506 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_410
timestamp 1607639953
transform 1 0 38806 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_398
timestamp 1607639953
transform 1 0 37702 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1200
timestamp 1607639953
transform 1 0 37610 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_434
timestamp 1607639953
transform 1 0 41014 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_422
timestamp 1607639953
transform 1 0 39910 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_459
timestamp 1607639953
transform 1 0 43314 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_446
timestamp 1607639953
transform 1 0 42118 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1201
timestamp 1607639953
transform 1 0 43222 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_483
timestamp 1607639953
transform 1 0 45522 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_471
timestamp 1607639953
transform 1 0 44418 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_495
timestamp 1607639953
transform 1 0 46626 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_520
timestamp 1607639953
transform 1 0 48926 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_507
timestamp 1607639953
transform 1 0 47730 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1202
timestamp 1607639953
transform 1 0 48834 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_544
timestamp 1607639953
transform 1 0 51134 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_532
timestamp 1607639953
transform 1 0 50030 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_568
timestamp 1607639953
transform 1 0 53342 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_556
timestamp 1607639953
transform 1 0 52238 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_593
timestamp 1607639953
transform 1 0 55642 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_98_581
timestamp 1607639953
transform 1 0 54538 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1203
timestamp 1607639953
transform 1 0 54446 0 -1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_98_605
timestamp 1607639953
transform 1 0 56746 0 -1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_98_617
timestamp 1607639953
transform 1 0 57850 0 -1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_197
timestamp 1607639953
transform -1 0 58862 0 -1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_100_15
timestamp 1607639953
transform 1 0 2466 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_3
timestamp 1607639953
transform 1 0 1362 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_15
timestamp 1607639953
transform 1 0 2466 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_3
timestamp 1607639953
transform 1 0 1362 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_200
timestamp 1607639953
transform 1 0 1086 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_198
timestamp 1607639953
transform 1 0 1086 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_100_44
timestamp 1607639953
transform 1 0 5134 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_32
timestamp 1607639953
transform 1 0 4030 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_100_27
timestamp 1607639953
transform 1 0 3570 0 -1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_99_39
timestamp 1607639953
transform 1 0 4674 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_27
timestamp 1607639953
transform 1 0 3570 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1214
timestamp 1607639953
transform 1 0 3938 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_56
timestamp 1607639953
transform 1 0 6238 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_62
timestamp 1607639953
transform 1 0 6790 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_99_59
timestamp 1607639953
transform 1 0 6514 0 1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_99_51
timestamp 1607639953
transform 1 0 5778 0 1 56032
box -38 -48 774 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1204
timestamp 1607639953
transform 1 0 6698 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_80
timestamp 1607639953
transform 1 0 8446 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_68
timestamp 1607639953
transform 1 0 7342 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_86
timestamp 1607639953
transform 1 0 8998 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_74
timestamp 1607639953
transform 1 0 7894 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_105
timestamp 1607639953
transform 1 0 10746 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_93
timestamp 1607639953
transform 1 0 9642 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_110
timestamp 1607639953
transform 1 0 11206 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_98
timestamp 1607639953
transform 1 0 10102 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1215
timestamp 1607639953
transform 1 0 9550 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_129
timestamp 1607639953
transform 1 0 12954 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_117
timestamp 1607639953
transform 1 0 11850 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_123
timestamp 1607639953
transform 1 0 12402 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1205
timestamp 1607639953
transform 1 0 12310 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_154
timestamp 1607639953
transform 1 0 15254 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_141
timestamp 1607639953
transform 1 0 14058 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_147
timestamp 1607639953
transform 1 0 14610 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_135
timestamp 1607639953
transform 1 0 13506 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1216
timestamp 1607639953
transform 1 0 15162 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_166
timestamp 1607639953
transform 1 0 16358 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_171
timestamp 1607639953
transform 1 0 16818 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_159
timestamp 1607639953
transform 1 0 15714 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_190
timestamp 1607639953
transform 1 0 18566 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_178
timestamp 1607639953
transform 1 0 17462 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_196
timestamp 1607639953
transform 1 0 19118 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_184
timestamp 1607639953
transform 1 0 18014 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1206
timestamp 1607639953
transform 1 0 17922 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_215
timestamp 1607639953
transform 1 0 20866 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_202
timestamp 1607639953
transform 1 0 19670 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_220
timestamp 1607639953
transform 1 0 21326 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_208
timestamp 1607639953
transform 1 0 20222 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1217
timestamp 1607639953
transform 1 0 20774 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_239
timestamp 1607639953
transform 1 0 23074 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_227
timestamp 1607639953
transform 1 0 21970 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_232
timestamp 1607639953
transform 1 0 22430 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_262
timestamp 1607639953
transform 1 0 25190 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_100_251
timestamp 1607639953
transform 1 0 24178 0 -1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_99_257
timestamp 1607639953
transform 1 0 24730 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_245
timestamp 1607639953
transform 1 0 23626 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1207
timestamp 1607639953
transform 1 0 23534 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _066_
timestamp 1607639953
transform 1 0 24914 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_100_276
timestamp 1607639953
transform 1 0 26478 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_100_274
timestamp 1607639953
transform 1 0 26294 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_281
timestamp 1607639953
transform 1 0 26938 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_269
timestamp 1607639953
transform 1 0 25834 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1218
timestamp 1607639953
transform 1 0 26386 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_300
timestamp 1607639953
transform 1 0 28686 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_288
timestamp 1607639953
transform 1 0 27582 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_306
timestamp 1607639953
transform 1 0 29238 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_293
timestamp 1607639953
transform 1 0 28042 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1208
timestamp 1607639953
transform 1 0 29146 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_324
timestamp 1607639953
transform 1 0 30894 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_312
timestamp 1607639953
transform 1 0 29790 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_330
timestamp 1607639953
transform 1 0 31446 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_318
timestamp 1607639953
transform 1 0 30342 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_342
timestamp 1607639953
transform 1 0 32550 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_100_337
timestamp 1607639953
transform 1 0 32090 0 -1 57120
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_99_342
timestamp 1607639953
transform 1 0 32550 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1219
timestamp 1607639953
transform 1 0 31998 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _183_
timestamp 1607639953
transform 1 0 32274 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_100_366
timestamp 1607639953
transform 1 0 34758 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_354
timestamp 1607639953
transform 1 0 33654 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_367
timestamp 1607639953
transform 1 0 34850 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_354
timestamp 1607639953
transform 1 0 33654 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1209
timestamp 1607639953
transform 1 0 34758 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_100_396
timestamp 1607639953
transform 1 0 37518 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_100_390
timestamp 1607639953
transform 1 0 36966 0 -1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_100_378
timestamp 1607639953
transform 1 0 35862 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_391
timestamp 1607639953
transform 1 0 37058 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_379
timestamp 1607639953
transform 1 0 35954 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_410
timestamp 1607639953
transform 1 0 38806 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_398
timestamp 1607639953
transform 1 0 37702 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_415
timestamp 1607639953
transform 1 0 39266 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_403
timestamp 1607639953
transform 1 0 38162 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1220
timestamp 1607639953
transform 1 0 37610 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_434
timestamp 1607639953
transform 1 0 41014 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_422
timestamp 1607639953
transform 1 0 39910 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_440
timestamp 1607639953
transform 1 0 41566 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_428
timestamp 1607639953
transform 1 0 40462 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1210
timestamp 1607639953
transform 1 0 40370 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_459
timestamp 1607639953
transform 1 0 43314 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_446
timestamp 1607639953
transform 1 0 42118 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_452
timestamp 1607639953
transform 1 0 42670 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1221
timestamp 1607639953
transform 1 0 43222 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_483
timestamp 1607639953
transform 1 0 45522 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_471
timestamp 1607639953
transform 1 0 44418 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_476
timestamp 1607639953
transform 1 0 44878 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_464
timestamp 1607639953
transform 1 0 43774 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_495
timestamp 1607639953
transform 1 0 46626 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_501
timestamp 1607639953
transform 1 0 47178 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_489
timestamp 1607639953
transform 1 0 46074 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1211
timestamp 1607639953
transform 1 0 45982 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_520
timestamp 1607639953
transform 1 0 48926 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_507
timestamp 1607639953
transform 1 0 47730 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_520
timestamp 1607639953
transform 1 0 48926 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_99_513
timestamp 1607639953
transform 1 0 48282 0 1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1222
timestamp 1607639953
transform 1 0 48834 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__conb_1  _013_
timestamp 1607639953
transform 1 0 48650 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_100_544
timestamp 1607639953
transform 1 0 51134 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_532
timestamp 1607639953
transform 1 0 50030 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_550
timestamp 1607639953
transform 1 0 51686 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_99_548
timestamp 1607639953
transform 1 0 51502 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_99_544
timestamp 1607639953
transform 1 0 51134 0 1 56032
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_99_532
timestamp 1607639953
transform 1 0 50030 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1212
timestamp 1607639953
transform 1 0 51594 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_100_571
timestamp 1607639953
transform 1 0 53618 0 -1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_100_559
timestamp 1607639953
transform 1 0 52514 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_562
timestamp 1607639953
transform 1 0 52790 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__conb_1  _095_
timestamp 1607639953
transform 1 0 52238 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_100_593
timestamp 1607639953
transform 1 0 55642 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_100_581
timestamp 1607639953
transform 1 0 54538 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_100_579
timestamp 1607639953
transform 1 0 54354 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_99_586
timestamp 1607639953
transform 1 0 54998 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_574
timestamp 1607639953
transform 1 0 53894 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1223
timestamp 1607639953
transform 1 0 54446 0 -1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_100_605
timestamp 1607639953
transform 1 0 56746 0 -1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_611
timestamp 1607639953
transform 1 0 57298 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_99_598
timestamp 1607639953
transform 1 0 56102 0 1 56032
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1213
timestamp 1607639953
transform 1 0 57206 0 1 56032
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_100_617
timestamp 1607639953
transform 1 0 57850 0 -1 57120
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_99_623
timestamp 1607639953
transform 1 0 58402 0 1 56032
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_201
timestamp 1607639953
transform -1 0 58862 0 -1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_199
timestamp 1607639953
transform -1 0 58862 0 1 56032
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_101_15
timestamp 1607639953
transform 1 0 2466 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_3
timestamp 1607639953
transform 1 0 1362 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_202
timestamp 1607639953
transform 1 0 1086 0 1 57120
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_101_44
timestamp 1607639953
transform 1 0 5134 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_32
timestamp 1607639953
transform 1 0 4030 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_101_27
timestamp 1607639953
transform 1 0 3570 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1224
timestamp 1607639953
transform 1 0 3938 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_63
timestamp 1607639953
transform 1 0 6882 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_56
timestamp 1607639953
transform 1 0 6238 0 1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1225
timestamp 1607639953
transform 1 0 6790 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_101_87
timestamp 1607639953
transform 1 0 9090 0 1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_101_75
timestamp 1607639953
transform 1 0 7986 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_106
timestamp 1607639953
transform 1 0 10838 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_94
timestamp 1607639953
transform 1 0 9734 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1226
timestamp 1607639953
transform 1 0 9642 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_125
timestamp 1607639953
transform 1 0 12586 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_118
timestamp 1607639953
transform 1 0 11942 0 1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1227
timestamp 1607639953
transform 1 0 12494 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_101_149
timestamp 1607639953
transform 1 0 14794 0 1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_101_137
timestamp 1607639953
transform 1 0 13690 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_168
timestamp 1607639953
transform 1 0 16542 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_156
timestamp 1607639953
transform 1 0 15438 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1228
timestamp 1607639953
transform 1 0 15346 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_187
timestamp 1607639953
transform 1 0 18290 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_180
timestamp 1607639953
transform 1 0 17646 0 1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1229
timestamp 1607639953
transform 1 0 18198 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_218
timestamp 1607639953
transform 1 0 21142 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_211
timestamp 1607639953
transform 1 0 20498 0 1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_101_199
timestamp 1607639953
transform 1 0 19394 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1230
timestamp 1607639953
transform 1 0 21050 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_101_242
timestamp 1607639953
transform 1 0 23350 0 1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_101_230
timestamp 1607639953
transform 1 0 22246 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_261
timestamp 1607639953
transform 1 0 25098 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_249
timestamp 1607639953
transform 1 0 23994 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1231
timestamp 1607639953
transform 1 0 23902 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_280
timestamp 1607639953
transform 1 0 26846 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_273
timestamp 1607639953
transform 1 0 26202 0 1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1232
timestamp 1607639953
transform 1 0 26754 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_101_304
timestamp 1607639953
transform 1 0 29054 0 1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_101_292
timestamp 1607639953
transform 1 0 27950 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_323
timestamp 1607639953
transform 1 0 30802 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_311
timestamp 1607639953
transform 1 0 29698 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1233
timestamp 1607639953
transform 1 0 29606 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_342
timestamp 1607639953
transform 1 0 32550 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_335
timestamp 1607639953
transform 1 0 31906 0 1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1234
timestamp 1607639953
transform 1 0 32458 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_373
timestamp 1607639953
transform 1 0 35402 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_366
timestamp 1607639953
transform 1 0 34758 0 1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_101_354
timestamp 1607639953
transform 1 0 33654 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1235
timestamp 1607639953
transform 1 0 35310 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_385
timestamp 1607639953
transform 1 0 36506 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_416
timestamp 1607639953
transform 1 0 39358 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_404
timestamp 1607639953
transform 1 0 38254 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_397
timestamp 1607639953
transform 1 0 37610 0 1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1236
timestamp 1607639953
transform 1 0 38162 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_435
timestamp 1607639953
transform 1 0 41106 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_428
timestamp 1607639953
transform 1 0 40462 0 1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1237
timestamp 1607639953
transform 1 0 41014 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_101_459
timestamp 1607639953
transform 1 0 43314 0 1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_101_447
timestamp 1607639953
transform 1 0 42210 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_478
timestamp 1607639953
transform 1 0 45062 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_466
timestamp 1607639953
transform 1 0 43958 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1238
timestamp 1607639953
transform 1 0 43866 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_497
timestamp 1607639953
transform 1 0 46810 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_490
timestamp 1607639953
transform 1 0 46166 0 1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1239
timestamp 1607639953
transform 1 0 46718 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_528
timestamp 1607639953
transform 1 0 49662 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_521
timestamp 1607639953
transform 1 0 49018 0 1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_101_509
timestamp 1607639953
transform 1 0 47914 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1240
timestamp 1607639953
transform 1 0 49570 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_540
timestamp 1607639953
transform 1 0 50766 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_571
timestamp 1607639953
transform 1 0 53618 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_101_559
timestamp 1607639953
transform 1 0 52514 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_552
timestamp 1607639953
transform 1 0 51870 0 1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1241
timestamp 1607639953
transform 1 0 52422 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_101_590
timestamp 1607639953
transform 1 0 55366 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_101_583
timestamp 1607639953
transform 1 0 54722 0 1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1242
timestamp 1607639953
transform 1 0 55274 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_101_614
timestamp 1607639953
transform 1 0 57574 0 1 57120
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_101_602
timestamp 1607639953
transform 1 0 56470 0 1 57120
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_101_621
timestamp 1607639953
transform 1 0 58218 0 1 57120
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_1243
timestamp 1607639953
transform 1 0 58126 0 1 57120
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_203
timestamp 1607639953
transform -1 0 58862 0 1 57120
box -38 -48 314 592
<< labels >>
rlabel metal2 s 184 59200 240 60000 6 io_in[0]
port 0 nsew default input
rlabel metal2 s 15916 59200 15972 60000 6 io_in[10]
port 1 nsew default input
rlabel metal2 s 17480 59200 17536 60000 6 io_in[11]
port 2 nsew default input
rlabel metal2 s 19044 59200 19100 60000 6 io_in[12]
port 3 nsew default input
rlabel metal2 s 20700 59200 20756 60000 6 io_in[13]
port 4 nsew default input
rlabel metal2 s 22264 59200 22320 60000 6 io_in[14]
port 5 nsew default input
rlabel metal2 s 23828 59200 23884 60000 6 io_in[15]
port 6 nsew default input
rlabel metal2 s 25392 59200 25448 60000 6 io_in[16]
port 7 nsew default input
rlabel metal2 s 26956 59200 27012 60000 6 io_in[17]
port 8 nsew default input
rlabel metal2 s 28520 59200 28576 60000 6 io_in[18]
port 9 nsew default input
rlabel metal2 s 30176 59200 30232 60000 6 io_in[19]
port 10 nsew default input
rlabel metal2 s 1748 59200 1804 60000 6 io_in[1]
port 11 nsew default input
rlabel metal2 s 31740 59200 31796 60000 6 io_in[20]
port 12 nsew default input
rlabel metal2 s 33304 59200 33360 60000 6 io_in[21]
port 13 nsew default input
rlabel metal2 s 34868 59200 34924 60000 6 io_in[22]
port 14 nsew default input
rlabel metal2 s 36432 59200 36488 60000 6 io_in[23]
port 15 nsew default input
rlabel metal2 s 37996 59200 38052 60000 6 io_in[24]
port 16 nsew default input
rlabel metal2 s 39560 59200 39616 60000 6 io_in[25]
port 17 nsew default input
rlabel metal2 s 41216 59200 41272 60000 6 io_in[26]
port 18 nsew default input
rlabel metal2 s 42780 59200 42836 60000 6 io_in[27]
port 19 nsew default input
rlabel metal2 s 44344 59200 44400 60000 6 io_in[28]
port 20 nsew default input
rlabel metal2 s 45908 59200 45964 60000 6 io_in[29]
port 21 nsew default input
rlabel metal2 s 3312 59200 3368 60000 6 io_in[2]
port 22 nsew default input
rlabel metal2 s 47472 59200 47528 60000 6 io_in[30]
port 23 nsew default input
rlabel metal2 s 49036 59200 49092 60000 6 io_in[31]
port 24 nsew default input
rlabel metal2 s 50692 59200 50748 60000 6 io_in[32]
port 25 nsew default input
rlabel metal2 s 52256 59200 52312 60000 6 io_in[33]
port 26 nsew default input
rlabel metal2 s 53820 59200 53876 60000 6 io_in[34]
port 27 nsew default input
rlabel metal2 s 55384 59200 55440 60000 6 io_in[35]
port 28 nsew default input
rlabel metal2 s 56948 59200 57004 60000 6 io_in[36]
port 29 nsew default input
rlabel metal2 s 58512 59200 58568 60000 6 io_in[37]
port 30 nsew default input
rlabel metal2 s 4876 59200 4932 60000 6 io_in[3]
port 31 nsew default input
rlabel metal2 s 6440 59200 6496 60000 6 io_in[4]
port 32 nsew default input
rlabel metal2 s 8004 59200 8060 60000 6 io_in[5]
port 33 nsew default input
rlabel metal2 s 9568 59200 9624 60000 6 io_in[6]
port 34 nsew default input
rlabel metal2 s 11224 59200 11280 60000 6 io_in[7]
port 35 nsew default input
rlabel metal2 s 12788 59200 12844 60000 6 io_in[8]
port 36 nsew default input
rlabel metal2 s 14352 59200 14408 60000 6 io_in[9]
port 37 nsew default input
rlabel metal2 s 644 59200 700 60000 6 io_oeb[0]
port 38 nsew default tristate
rlabel metal2 s 16468 59200 16524 60000 6 io_oeb[10]
port 39 nsew default tristate
rlabel metal2 s 18032 59200 18088 60000 6 io_oeb[11]
port 40 nsew default tristate
rlabel metal2 s 19596 59200 19652 60000 6 io_oeb[12]
port 41 nsew default tristate
rlabel metal2 s 21160 59200 21216 60000 6 io_oeb[13]
port 42 nsew default tristate
rlabel metal2 s 22724 59200 22780 60000 6 io_oeb[14]
port 43 nsew default tristate
rlabel metal2 s 24380 59200 24436 60000 6 io_oeb[15]
port 44 nsew default tristate
rlabel metal2 s 25944 59200 26000 60000 6 io_oeb[16]
port 45 nsew default tristate
rlabel metal2 s 27508 59200 27564 60000 6 io_oeb[17]
port 46 nsew default tristate
rlabel metal2 s 29072 59200 29128 60000 6 io_oeb[18]
port 47 nsew default tristate
rlabel metal2 s 30636 59200 30692 60000 6 io_oeb[19]
port 48 nsew default tristate
rlabel metal2 s 2208 59200 2264 60000 6 io_oeb[1]
port 49 nsew default tristate
rlabel metal2 s 32200 59200 32256 60000 6 io_oeb[20]
port 50 nsew default tristate
rlabel metal2 s 33856 59200 33912 60000 6 io_oeb[21]
port 51 nsew default tristate
rlabel metal2 s 35420 59200 35476 60000 6 io_oeb[22]
port 52 nsew default tristate
rlabel metal2 s 36984 59200 37040 60000 6 io_oeb[23]
port 53 nsew default tristate
rlabel metal2 s 38548 59200 38604 60000 6 io_oeb[24]
port 54 nsew default tristate
rlabel metal2 s 40112 59200 40168 60000 6 io_oeb[25]
port 55 nsew default tristate
rlabel metal2 s 41676 59200 41732 60000 6 io_oeb[26]
port 56 nsew default tristate
rlabel metal2 s 43240 59200 43296 60000 6 io_oeb[27]
port 57 nsew default tristate
rlabel metal2 s 44896 59200 44952 60000 6 io_oeb[28]
port 58 nsew default tristate
rlabel metal2 s 46460 59200 46516 60000 6 io_oeb[29]
port 59 nsew default tristate
rlabel metal2 s 3864 59200 3920 60000 6 io_oeb[2]
port 60 nsew default tristate
rlabel metal2 s 48024 59200 48080 60000 6 io_oeb[30]
port 61 nsew default tristate
rlabel metal2 s 49588 59200 49644 60000 6 io_oeb[31]
port 62 nsew default tristate
rlabel metal2 s 51152 59200 51208 60000 6 io_oeb[32]
port 63 nsew default tristate
rlabel metal2 s 52716 59200 52772 60000 6 io_oeb[33]
port 64 nsew default tristate
rlabel metal2 s 54372 59200 54428 60000 6 io_oeb[34]
port 65 nsew default tristate
rlabel metal2 s 55936 59200 55992 60000 6 io_oeb[35]
port 66 nsew default tristate
rlabel metal2 s 57500 59200 57556 60000 6 io_oeb[36]
port 67 nsew default tristate
rlabel metal2 s 59064 59200 59120 60000 6 io_oeb[37]
port 68 nsew default tristate
rlabel metal2 s 5428 59200 5484 60000 6 io_oeb[3]
port 69 nsew default tristate
rlabel metal2 s 6992 59200 7048 60000 6 io_oeb[4]
port 70 nsew default tristate
rlabel metal2 s 8556 59200 8612 60000 6 io_oeb[5]
port 71 nsew default tristate
rlabel metal2 s 10120 59200 10176 60000 6 io_oeb[6]
port 72 nsew default tristate
rlabel metal2 s 11684 59200 11740 60000 6 io_oeb[7]
port 73 nsew default tristate
rlabel metal2 s 13248 59200 13304 60000 6 io_oeb[8]
port 74 nsew default tristate
rlabel metal2 s 14904 59200 14960 60000 6 io_oeb[9]
port 75 nsew default tristate
rlabel metal2 s 1196 59200 1252 60000 6 io_out[0]
port 76 nsew default tristate
rlabel metal2 s 17020 59200 17076 60000 6 io_out[10]
port 77 nsew default tristate
rlabel metal2 s 18584 59200 18640 60000 6 io_out[11]
port 78 nsew default tristate
rlabel metal2 s 20148 59200 20204 60000 6 io_out[12]
port 79 nsew default tristate
rlabel metal2 s 21712 59200 21768 60000 6 io_out[13]
port 80 nsew default tristate
rlabel metal2 s 23276 59200 23332 60000 6 io_out[14]
port 81 nsew default tristate
rlabel metal2 s 24840 59200 24896 60000 6 io_out[15]
port 82 nsew default tristate
rlabel metal2 s 26404 59200 26460 60000 6 io_out[16]
port 83 nsew default tristate
rlabel metal2 s 28060 59200 28116 60000 6 io_out[17]
port 84 nsew default tristate
rlabel metal2 s 29624 59200 29680 60000 6 io_out[18]
port 85 nsew default tristate
rlabel metal2 s 31188 59200 31244 60000 6 io_out[19]
port 86 nsew default tristate
rlabel metal2 s 2760 59200 2816 60000 6 io_out[1]
port 87 nsew default tristate
rlabel metal2 s 32752 59200 32808 60000 6 io_out[20]
port 88 nsew default tristate
rlabel metal2 s 34316 59200 34372 60000 6 io_out[21]
port 89 nsew default tristate
rlabel metal2 s 35880 59200 35936 60000 6 io_out[22]
port 90 nsew default tristate
rlabel metal2 s 37536 59200 37592 60000 6 io_out[23]
port 91 nsew default tristate
rlabel metal2 s 39100 59200 39156 60000 6 io_out[24]
port 92 nsew default tristate
rlabel metal2 s 40664 59200 40720 60000 6 io_out[25]
port 93 nsew default tristate
rlabel metal2 s 42228 59200 42284 60000 6 io_out[26]
port 94 nsew default tristate
rlabel metal2 s 43792 59200 43848 60000 6 io_out[27]
port 95 nsew default tristate
rlabel metal2 s 45356 59200 45412 60000 6 io_out[28]
port 96 nsew default tristate
rlabel metal2 s 47012 59200 47068 60000 6 io_out[29]
port 97 nsew default tristate
rlabel metal2 s 4324 59200 4380 60000 6 io_out[2]
port 98 nsew default tristate
rlabel metal2 s 48576 59200 48632 60000 6 io_out[30]
port 99 nsew default tristate
rlabel metal2 s 50140 59200 50196 60000 6 io_out[31]
port 100 nsew default tristate
rlabel metal2 s 51704 59200 51760 60000 6 io_out[32]
port 101 nsew default tristate
rlabel metal2 s 53268 59200 53324 60000 6 io_out[33]
port 102 nsew default tristate
rlabel metal2 s 54832 59200 54888 60000 6 io_out[34]
port 103 nsew default tristate
rlabel metal2 s 56396 59200 56452 60000 6 io_out[35]
port 104 nsew default tristate
rlabel metal2 s 58052 59200 58108 60000 6 io_out[36]
port 105 nsew default tristate
rlabel metal2 s 59616 59200 59672 60000 6 io_out[37]
port 106 nsew default tristate
rlabel metal2 s 5888 59200 5944 60000 6 io_out[3]
port 107 nsew default tristate
rlabel metal2 s 7544 59200 7600 60000 6 io_out[4]
port 108 nsew default tristate
rlabel metal2 s 9108 59200 9164 60000 6 io_out[5]
port 109 nsew default tristate
rlabel metal2 s 10672 59200 10728 60000 6 io_out[6]
port 110 nsew default tristate
rlabel metal2 s 12236 59200 12292 60000 6 io_out[7]
port 111 nsew default tristate
rlabel metal2 s 13800 59200 13856 60000 6 io_out[8]
port 112 nsew default tristate
rlabel metal2 s 15364 59200 15420 60000 6 io_out[9]
port 113 nsew default tristate
rlabel metal2 s 12972 0 13028 800 6 la_data_in[0]
port 114 nsew default input
rlabel metal2 s 49680 0 49736 800 6 la_data_in[100]
port 115 nsew default input
rlabel metal2 s 50048 0 50104 800 6 la_data_in[101]
port 116 nsew default input
rlabel metal2 s 50416 0 50472 800 6 la_data_in[102]
port 117 nsew default input
rlabel metal2 s 50784 0 50840 800 6 la_data_in[103]
port 118 nsew default input
rlabel metal2 s 51152 0 51208 800 6 la_data_in[104]
port 119 nsew default input
rlabel metal2 s 51520 0 51576 800 6 la_data_in[105]
port 120 nsew default input
rlabel metal2 s 51888 0 51944 800 6 la_data_in[106]
port 121 nsew default input
rlabel metal2 s 52256 0 52312 800 6 la_data_in[107]
port 122 nsew default input
rlabel metal2 s 52624 0 52680 800 6 la_data_in[108]
port 123 nsew default input
rlabel metal2 s 52992 0 53048 800 6 la_data_in[109]
port 124 nsew default input
rlabel metal2 s 16560 0 16616 800 6 la_data_in[10]
port 125 nsew default input
rlabel metal2 s 53360 0 53416 800 6 la_data_in[110]
port 126 nsew default input
rlabel metal2 s 53728 0 53784 800 6 la_data_in[111]
port 127 nsew default input
rlabel metal2 s 54096 0 54152 800 6 la_data_in[112]
port 128 nsew default input
rlabel metal2 s 54464 0 54520 800 6 la_data_in[113]
port 129 nsew default input
rlabel metal2 s 54832 0 54888 800 6 la_data_in[114]
port 130 nsew default input
rlabel metal2 s 55200 0 55256 800 6 la_data_in[115]
port 131 nsew default input
rlabel metal2 s 55568 0 55624 800 6 la_data_in[116]
port 132 nsew default input
rlabel metal2 s 55936 0 55992 800 6 la_data_in[117]
port 133 nsew default input
rlabel metal2 s 56304 0 56360 800 6 la_data_in[118]
port 134 nsew default input
rlabel metal2 s 56672 0 56728 800 6 la_data_in[119]
port 135 nsew default input
rlabel metal2 s 16928 0 16984 800 6 la_data_in[11]
port 136 nsew default input
rlabel metal2 s 57040 0 57096 800 6 la_data_in[120]
port 137 nsew default input
rlabel metal2 s 57408 0 57464 800 6 la_data_in[121]
port 138 nsew default input
rlabel metal2 s 57776 0 57832 800 6 la_data_in[122]
port 139 nsew default input
rlabel metal2 s 58144 0 58200 800 6 la_data_in[123]
port 140 nsew default input
rlabel metal2 s 58512 0 58568 800 6 la_data_in[124]
port 141 nsew default input
rlabel metal2 s 58880 0 58936 800 6 la_data_in[125]
port 142 nsew default input
rlabel metal2 s 59248 0 59304 800 6 la_data_in[126]
port 143 nsew default input
rlabel metal2 s 59616 0 59672 800 6 la_data_in[127]
port 144 nsew default input
rlabel metal2 s 17296 0 17352 800 6 la_data_in[12]
port 145 nsew default input
rlabel metal2 s 17664 0 17720 800 6 la_data_in[13]
port 146 nsew default input
rlabel metal2 s 18032 0 18088 800 6 la_data_in[14]
port 147 nsew default input
rlabel metal2 s 18400 0 18456 800 6 la_data_in[15]
port 148 nsew default input
rlabel metal2 s 18768 0 18824 800 6 la_data_in[16]
port 149 nsew default input
rlabel metal2 s 19136 0 19192 800 6 la_data_in[17]
port 150 nsew default input
rlabel metal2 s 19504 0 19560 800 6 la_data_in[18]
port 151 nsew default input
rlabel metal2 s 19872 0 19928 800 6 la_data_in[19]
port 152 nsew default input
rlabel metal2 s 13340 0 13396 800 6 la_data_in[1]
port 153 nsew default input
rlabel metal2 s 20240 0 20296 800 6 la_data_in[20]
port 154 nsew default input
rlabel metal2 s 20608 0 20664 800 6 la_data_in[21]
port 155 nsew default input
rlabel metal2 s 20976 0 21032 800 6 la_data_in[22]
port 156 nsew default input
rlabel metal2 s 21344 0 21400 800 6 la_data_in[23]
port 157 nsew default input
rlabel metal2 s 21712 0 21768 800 6 la_data_in[24]
port 158 nsew default input
rlabel metal2 s 22080 0 22136 800 6 la_data_in[25]
port 159 nsew default input
rlabel metal2 s 22448 0 22504 800 6 la_data_in[26]
port 160 nsew default input
rlabel metal2 s 22816 0 22872 800 6 la_data_in[27]
port 161 nsew default input
rlabel metal2 s 23184 0 23240 800 6 la_data_in[28]
port 162 nsew default input
rlabel metal2 s 23552 0 23608 800 6 la_data_in[29]
port 163 nsew default input
rlabel metal2 s 13708 0 13764 800 6 la_data_in[2]
port 164 nsew default input
rlabel metal2 s 23920 0 23976 800 6 la_data_in[30]
port 165 nsew default input
rlabel metal2 s 24288 0 24344 800 6 la_data_in[31]
port 166 nsew default input
rlabel metal2 s 24656 0 24712 800 6 la_data_in[32]
port 167 nsew default input
rlabel metal2 s 25024 0 25080 800 6 la_data_in[33]
port 168 nsew default input
rlabel metal2 s 25392 0 25448 800 6 la_data_in[34]
port 169 nsew default input
rlabel metal2 s 25760 0 25816 800 6 la_data_in[35]
port 170 nsew default input
rlabel metal2 s 26128 0 26184 800 6 la_data_in[36]
port 171 nsew default input
rlabel metal2 s 26496 0 26552 800 6 la_data_in[37]
port 172 nsew default input
rlabel metal2 s 26864 0 26920 800 6 la_data_in[38]
port 173 nsew default input
rlabel metal2 s 27232 0 27288 800 6 la_data_in[39]
port 174 nsew default input
rlabel metal2 s 14076 0 14132 800 6 la_data_in[3]
port 175 nsew default input
rlabel metal2 s 27600 0 27656 800 6 la_data_in[40]
port 176 nsew default input
rlabel metal2 s 27968 0 28024 800 6 la_data_in[41]
port 177 nsew default input
rlabel metal2 s 28336 0 28392 800 6 la_data_in[42]
port 178 nsew default input
rlabel metal2 s 28704 0 28760 800 6 la_data_in[43]
port 179 nsew default input
rlabel metal2 s 29072 0 29128 800 6 la_data_in[44]
port 180 nsew default input
rlabel metal2 s 29440 0 29496 800 6 la_data_in[45]
port 181 nsew default input
rlabel metal2 s 29808 0 29864 800 6 la_data_in[46]
port 182 nsew default input
rlabel metal2 s 30176 0 30232 800 6 la_data_in[47]
port 183 nsew default input
rlabel metal2 s 30544 0 30600 800 6 la_data_in[48]
port 184 nsew default input
rlabel metal2 s 30912 0 30968 800 6 la_data_in[49]
port 185 nsew default input
rlabel metal2 s 14444 0 14500 800 6 la_data_in[4]
port 186 nsew default input
rlabel metal2 s 31280 0 31336 800 6 la_data_in[50]
port 187 nsew default input
rlabel metal2 s 31648 0 31704 800 6 la_data_in[51]
port 188 nsew default input
rlabel metal2 s 32016 0 32072 800 6 la_data_in[52]
port 189 nsew default input
rlabel metal2 s 32384 0 32440 800 6 la_data_in[53]
port 190 nsew default input
rlabel metal2 s 32752 0 32808 800 6 la_data_in[54]
port 191 nsew default input
rlabel metal2 s 33120 0 33176 800 6 la_data_in[55]
port 192 nsew default input
rlabel metal2 s 33488 0 33544 800 6 la_data_in[56]
port 193 nsew default input
rlabel metal2 s 33856 0 33912 800 6 la_data_in[57]
port 194 nsew default input
rlabel metal2 s 34224 0 34280 800 6 la_data_in[58]
port 195 nsew default input
rlabel metal2 s 34592 0 34648 800 6 la_data_in[59]
port 196 nsew default input
rlabel metal2 s 14812 0 14868 800 6 la_data_in[5]
port 197 nsew default input
rlabel metal2 s 34960 0 35016 800 6 la_data_in[60]
port 198 nsew default input
rlabel metal2 s 35328 0 35384 800 6 la_data_in[61]
port 199 nsew default input
rlabel metal2 s 35696 0 35752 800 6 la_data_in[62]
port 200 nsew default input
rlabel metal2 s 36064 0 36120 800 6 la_data_in[63]
port 201 nsew default input
rlabel metal2 s 36432 0 36488 800 6 la_data_in[64]
port 202 nsew default input
rlabel metal2 s 36800 0 36856 800 6 la_data_in[65]
port 203 nsew default input
rlabel metal2 s 37168 0 37224 800 6 la_data_in[66]
port 204 nsew default input
rlabel metal2 s 37536 0 37592 800 6 la_data_in[67]
port 205 nsew default input
rlabel metal2 s 37904 0 37960 800 6 la_data_in[68]
port 206 nsew default input
rlabel metal2 s 38272 0 38328 800 6 la_data_in[69]
port 207 nsew default input
rlabel metal2 s 15088 0 15144 800 6 la_data_in[6]
port 208 nsew default input
rlabel metal2 s 38640 0 38696 800 6 la_data_in[70]
port 209 nsew default input
rlabel metal2 s 39008 0 39064 800 6 la_data_in[71]
port 210 nsew default input
rlabel metal2 s 39376 0 39432 800 6 la_data_in[72]
port 211 nsew default input
rlabel metal2 s 39744 0 39800 800 6 la_data_in[73]
port 212 nsew default input
rlabel metal2 s 40112 0 40168 800 6 la_data_in[74]
port 213 nsew default input
rlabel metal2 s 40480 0 40536 800 6 la_data_in[75]
port 214 nsew default input
rlabel metal2 s 40848 0 40904 800 6 la_data_in[76]
port 215 nsew default input
rlabel metal2 s 41216 0 41272 800 6 la_data_in[77]
port 216 nsew default input
rlabel metal2 s 41584 0 41640 800 6 la_data_in[78]
port 217 nsew default input
rlabel metal2 s 41952 0 42008 800 6 la_data_in[79]
port 218 nsew default input
rlabel metal2 s 15456 0 15512 800 6 la_data_in[7]
port 219 nsew default input
rlabel metal2 s 42320 0 42376 800 6 la_data_in[80]
port 220 nsew default input
rlabel metal2 s 42688 0 42744 800 6 la_data_in[81]
port 221 nsew default input
rlabel metal2 s 43056 0 43112 800 6 la_data_in[82]
port 222 nsew default input
rlabel metal2 s 43424 0 43480 800 6 la_data_in[83]
port 223 nsew default input
rlabel metal2 s 43792 0 43848 800 6 la_data_in[84]
port 224 nsew default input
rlabel metal2 s 44160 0 44216 800 6 la_data_in[85]
port 225 nsew default input
rlabel metal2 s 44528 0 44584 800 6 la_data_in[86]
port 226 nsew default input
rlabel metal2 s 44896 0 44952 800 6 la_data_in[87]
port 227 nsew default input
rlabel metal2 s 45264 0 45320 800 6 la_data_in[88]
port 228 nsew default input
rlabel metal2 s 45632 0 45688 800 6 la_data_in[89]
port 229 nsew default input
rlabel metal2 s 15824 0 15880 800 6 la_data_in[8]
port 230 nsew default input
rlabel metal2 s 46000 0 46056 800 6 la_data_in[90]
port 231 nsew default input
rlabel metal2 s 46368 0 46424 800 6 la_data_in[91]
port 232 nsew default input
rlabel metal2 s 46736 0 46792 800 6 la_data_in[92]
port 233 nsew default input
rlabel metal2 s 47104 0 47160 800 6 la_data_in[93]
port 234 nsew default input
rlabel metal2 s 47472 0 47528 800 6 la_data_in[94]
port 235 nsew default input
rlabel metal2 s 47840 0 47896 800 6 la_data_in[95]
port 236 nsew default input
rlabel metal2 s 48208 0 48264 800 6 la_data_in[96]
port 237 nsew default input
rlabel metal2 s 48576 0 48632 800 6 la_data_in[97]
port 238 nsew default input
rlabel metal2 s 48944 0 49000 800 6 la_data_in[98]
port 239 nsew default input
rlabel metal2 s 49312 0 49368 800 6 la_data_in[99]
port 240 nsew default input
rlabel metal2 s 16192 0 16248 800 6 la_data_in[9]
port 241 nsew default input
rlabel metal2 s 13064 0 13120 800 6 la_data_out[0]
port 242 nsew default tristate
rlabel metal2 s 49772 0 49828 800 6 la_data_out[100]
port 243 nsew default tristate
rlabel metal2 s 50140 0 50196 800 6 la_data_out[101]
port 244 nsew default tristate
rlabel metal2 s 50508 0 50564 800 6 la_data_out[102]
port 245 nsew default tristate
rlabel metal2 s 50876 0 50932 800 6 la_data_out[103]
port 246 nsew default tristate
rlabel metal2 s 51244 0 51300 800 6 la_data_out[104]
port 247 nsew default tristate
rlabel metal2 s 51612 0 51668 800 6 la_data_out[105]
port 248 nsew default tristate
rlabel metal2 s 51980 0 52036 800 6 la_data_out[106]
port 249 nsew default tristate
rlabel metal2 s 52348 0 52404 800 6 la_data_out[107]
port 250 nsew default tristate
rlabel metal2 s 52716 0 52772 800 6 la_data_out[108]
port 251 nsew default tristate
rlabel metal2 s 53084 0 53140 800 6 la_data_out[109]
port 252 nsew default tristate
rlabel metal2 s 16744 0 16800 800 6 la_data_out[10]
port 253 nsew default tristate
rlabel metal2 s 53452 0 53508 800 6 la_data_out[110]
port 254 nsew default tristate
rlabel metal2 s 53820 0 53876 800 6 la_data_out[111]
port 255 nsew default tristate
rlabel metal2 s 54188 0 54244 800 6 la_data_out[112]
port 256 nsew default tristate
rlabel metal2 s 54556 0 54612 800 6 la_data_out[113]
port 257 nsew default tristate
rlabel metal2 s 54924 0 54980 800 6 la_data_out[114]
port 258 nsew default tristate
rlabel metal2 s 55292 0 55348 800 6 la_data_out[115]
port 259 nsew default tristate
rlabel metal2 s 55660 0 55716 800 6 la_data_out[116]
port 260 nsew default tristate
rlabel metal2 s 56028 0 56084 800 6 la_data_out[117]
port 261 nsew default tristate
rlabel metal2 s 56396 0 56452 800 6 la_data_out[118]
port 262 nsew default tristate
rlabel metal2 s 56764 0 56820 800 6 la_data_out[119]
port 263 nsew default tristate
rlabel metal2 s 17112 0 17168 800 6 la_data_out[11]
port 264 nsew default tristate
rlabel metal2 s 57132 0 57188 800 6 la_data_out[120]
port 265 nsew default tristate
rlabel metal2 s 57500 0 57556 800 6 la_data_out[121]
port 266 nsew default tristate
rlabel metal2 s 57868 0 57924 800 6 la_data_out[122]
port 267 nsew default tristate
rlabel metal2 s 58236 0 58292 800 6 la_data_out[123]
port 268 nsew default tristate
rlabel metal2 s 58604 0 58660 800 6 la_data_out[124]
port 269 nsew default tristate
rlabel metal2 s 58972 0 59028 800 6 la_data_out[125]
port 270 nsew default tristate
rlabel metal2 s 59340 0 59396 800 6 la_data_out[126]
port 271 nsew default tristate
rlabel metal2 s 59708 0 59764 800 6 la_data_out[127]
port 272 nsew default tristate
rlabel metal2 s 17480 0 17536 800 6 la_data_out[12]
port 273 nsew default tristate
rlabel metal2 s 17848 0 17904 800 6 la_data_out[13]
port 274 nsew default tristate
rlabel metal2 s 18216 0 18272 800 6 la_data_out[14]
port 275 nsew default tristate
rlabel metal2 s 18584 0 18640 800 6 la_data_out[15]
port 276 nsew default tristate
rlabel metal2 s 18952 0 19008 800 6 la_data_out[16]
port 277 nsew default tristate
rlabel metal2 s 19320 0 19376 800 6 la_data_out[17]
port 278 nsew default tristate
rlabel metal2 s 19688 0 19744 800 6 la_data_out[18]
port 279 nsew default tristate
rlabel metal2 s 20056 0 20112 800 6 la_data_out[19]
port 280 nsew default tristate
rlabel metal2 s 13432 0 13488 800 6 la_data_out[1]
port 281 nsew default tristate
rlabel metal2 s 20424 0 20480 800 6 la_data_out[20]
port 282 nsew default tristate
rlabel metal2 s 20792 0 20848 800 6 la_data_out[21]
port 283 nsew default tristate
rlabel metal2 s 21160 0 21216 800 6 la_data_out[22]
port 284 nsew default tristate
rlabel metal2 s 21528 0 21584 800 6 la_data_out[23]
port 285 nsew default tristate
rlabel metal2 s 21896 0 21952 800 6 la_data_out[24]
port 286 nsew default tristate
rlabel metal2 s 22264 0 22320 800 6 la_data_out[25]
port 287 nsew default tristate
rlabel metal2 s 22632 0 22688 800 6 la_data_out[26]
port 288 nsew default tristate
rlabel metal2 s 23000 0 23056 800 6 la_data_out[27]
port 289 nsew default tristate
rlabel metal2 s 23368 0 23424 800 6 la_data_out[28]
port 290 nsew default tristate
rlabel metal2 s 23736 0 23792 800 6 la_data_out[29]
port 291 nsew default tristate
rlabel metal2 s 13800 0 13856 800 6 la_data_out[2]
port 292 nsew default tristate
rlabel metal2 s 24104 0 24160 800 6 la_data_out[30]
port 293 nsew default tristate
rlabel metal2 s 24472 0 24528 800 6 la_data_out[31]
port 294 nsew default tristate
rlabel metal2 s 24840 0 24896 800 6 la_data_out[32]
port 295 nsew default tristate
rlabel metal2 s 25208 0 25264 800 6 la_data_out[33]
port 296 nsew default tristate
rlabel metal2 s 25576 0 25632 800 6 la_data_out[34]
port 297 nsew default tristate
rlabel metal2 s 25944 0 26000 800 6 la_data_out[35]
port 298 nsew default tristate
rlabel metal2 s 26312 0 26368 800 6 la_data_out[36]
port 299 nsew default tristate
rlabel metal2 s 26680 0 26736 800 6 la_data_out[37]
port 300 nsew default tristate
rlabel metal2 s 27048 0 27104 800 6 la_data_out[38]
port 301 nsew default tristate
rlabel metal2 s 27416 0 27472 800 6 la_data_out[39]
port 302 nsew default tristate
rlabel metal2 s 14168 0 14224 800 6 la_data_out[3]
port 303 nsew default tristate
rlabel metal2 s 27784 0 27840 800 6 la_data_out[40]
port 304 nsew default tristate
rlabel metal2 s 28152 0 28208 800 6 la_data_out[41]
port 305 nsew default tristate
rlabel metal2 s 28520 0 28576 800 6 la_data_out[42]
port 306 nsew default tristate
rlabel metal2 s 28888 0 28944 800 6 la_data_out[43]
port 307 nsew default tristate
rlabel metal2 s 29256 0 29312 800 6 la_data_out[44]
port 308 nsew default tristate
rlabel metal2 s 29624 0 29680 800 6 la_data_out[45]
port 309 nsew default tristate
rlabel metal2 s 29992 0 30048 800 6 la_data_out[46]
port 310 nsew default tristate
rlabel metal2 s 30268 0 30324 800 6 la_data_out[47]
port 311 nsew default tristate
rlabel metal2 s 30636 0 30692 800 6 la_data_out[48]
port 312 nsew default tristate
rlabel metal2 s 31004 0 31060 800 6 la_data_out[49]
port 313 nsew default tristate
rlabel metal2 s 14536 0 14592 800 6 la_data_out[4]
port 314 nsew default tristate
rlabel metal2 s 31372 0 31428 800 6 la_data_out[50]
port 315 nsew default tristate
rlabel metal2 s 31740 0 31796 800 6 la_data_out[51]
port 316 nsew default tristate
rlabel metal2 s 32108 0 32164 800 6 la_data_out[52]
port 317 nsew default tristate
rlabel metal2 s 32476 0 32532 800 6 la_data_out[53]
port 318 nsew default tristate
rlabel metal2 s 32844 0 32900 800 6 la_data_out[54]
port 319 nsew default tristate
rlabel metal2 s 33212 0 33268 800 6 la_data_out[55]
port 320 nsew default tristate
rlabel metal2 s 33580 0 33636 800 6 la_data_out[56]
port 321 nsew default tristate
rlabel metal2 s 33948 0 34004 800 6 la_data_out[57]
port 322 nsew default tristate
rlabel metal2 s 34316 0 34372 800 6 la_data_out[58]
port 323 nsew default tristate
rlabel metal2 s 34684 0 34740 800 6 la_data_out[59]
port 324 nsew default tristate
rlabel metal2 s 14904 0 14960 800 6 la_data_out[5]
port 325 nsew default tristate
rlabel metal2 s 35052 0 35108 800 6 la_data_out[60]
port 326 nsew default tristate
rlabel metal2 s 35420 0 35476 800 6 la_data_out[61]
port 327 nsew default tristate
rlabel metal2 s 35788 0 35844 800 6 la_data_out[62]
port 328 nsew default tristate
rlabel metal2 s 36156 0 36212 800 6 la_data_out[63]
port 329 nsew default tristate
rlabel metal2 s 36524 0 36580 800 6 la_data_out[64]
port 330 nsew default tristate
rlabel metal2 s 36892 0 36948 800 6 la_data_out[65]
port 331 nsew default tristate
rlabel metal2 s 37260 0 37316 800 6 la_data_out[66]
port 332 nsew default tristate
rlabel metal2 s 37628 0 37684 800 6 la_data_out[67]
port 333 nsew default tristate
rlabel metal2 s 37996 0 38052 800 6 la_data_out[68]
port 334 nsew default tristate
rlabel metal2 s 38364 0 38420 800 6 la_data_out[69]
port 335 nsew default tristate
rlabel metal2 s 15272 0 15328 800 6 la_data_out[6]
port 336 nsew default tristate
rlabel metal2 s 38732 0 38788 800 6 la_data_out[70]
port 337 nsew default tristate
rlabel metal2 s 39100 0 39156 800 6 la_data_out[71]
port 338 nsew default tristate
rlabel metal2 s 39468 0 39524 800 6 la_data_out[72]
port 339 nsew default tristate
rlabel metal2 s 39836 0 39892 800 6 la_data_out[73]
port 340 nsew default tristate
rlabel metal2 s 40204 0 40260 800 6 la_data_out[74]
port 341 nsew default tristate
rlabel metal2 s 40572 0 40628 800 6 la_data_out[75]
port 342 nsew default tristate
rlabel metal2 s 40940 0 40996 800 6 la_data_out[76]
port 343 nsew default tristate
rlabel metal2 s 41308 0 41364 800 6 la_data_out[77]
port 344 nsew default tristate
rlabel metal2 s 41676 0 41732 800 6 la_data_out[78]
port 345 nsew default tristate
rlabel metal2 s 42044 0 42100 800 6 la_data_out[79]
port 346 nsew default tristate
rlabel metal2 s 15640 0 15696 800 6 la_data_out[7]
port 347 nsew default tristate
rlabel metal2 s 42412 0 42468 800 6 la_data_out[80]
port 348 nsew default tristate
rlabel metal2 s 42780 0 42836 800 6 la_data_out[81]
port 349 nsew default tristate
rlabel metal2 s 43148 0 43204 800 6 la_data_out[82]
port 350 nsew default tristate
rlabel metal2 s 43516 0 43572 800 6 la_data_out[83]
port 351 nsew default tristate
rlabel metal2 s 43884 0 43940 800 6 la_data_out[84]
port 352 nsew default tristate
rlabel metal2 s 44252 0 44308 800 6 la_data_out[85]
port 353 nsew default tristate
rlabel metal2 s 44620 0 44676 800 6 la_data_out[86]
port 354 nsew default tristate
rlabel metal2 s 44988 0 45044 800 6 la_data_out[87]
port 355 nsew default tristate
rlabel metal2 s 45356 0 45412 800 6 la_data_out[88]
port 356 nsew default tristate
rlabel metal2 s 45724 0 45780 800 6 la_data_out[89]
port 357 nsew default tristate
rlabel metal2 s 16008 0 16064 800 6 la_data_out[8]
port 358 nsew default tristate
rlabel metal2 s 46092 0 46148 800 6 la_data_out[90]
port 359 nsew default tristate
rlabel metal2 s 46460 0 46516 800 6 la_data_out[91]
port 360 nsew default tristate
rlabel metal2 s 46828 0 46884 800 6 la_data_out[92]
port 361 nsew default tristate
rlabel metal2 s 47196 0 47252 800 6 la_data_out[93]
port 362 nsew default tristate
rlabel metal2 s 47564 0 47620 800 6 la_data_out[94]
port 363 nsew default tristate
rlabel metal2 s 47932 0 47988 800 6 la_data_out[95]
port 364 nsew default tristate
rlabel metal2 s 48300 0 48356 800 6 la_data_out[96]
port 365 nsew default tristate
rlabel metal2 s 48668 0 48724 800 6 la_data_out[97]
port 366 nsew default tristate
rlabel metal2 s 49036 0 49092 800 6 la_data_out[98]
port 367 nsew default tristate
rlabel metal2 s 49404 0 49460 800 6 la_data_out[99]
port 368 nsew default tristate
rlabel metal2 s 16376 0 16432 800 6 la_data_out[9]
port 369 nsew default tristate
rlabel metal2 s 13156 0 13212 800 6 la_oen[0]
port 370 nsew default input
rlabel metal2 s 49864 0 49920 800 6 la_oen[100]
port 371 nsew default input
rlabel metal2 s 50232 0 50288 800 6 la_oen[101]
port 372 nsew default input
rlabel metal2 s 50600 0 50656 800 6 la_oen[102]
port 373 nsew default input
rlabel metal2 s 50968 0 51024 800 6 la_oen[103]
port 374 nsew default input
rlabel metal2 s 51336 0 51392 800 6 la_oen[104]
port 375 nsew default input
rlabel metal2 s 51704 0 51760 800 6 la_oen[105]
port 376 nsew default input
rlabel metal2 s 52072 0 52128 800 6 la_oen[106]
port 377 nsew default input
rlabel metal2 s 52440 0 52496 800 6 la_oen[107]
port 378 nsew default input
rlabel metal2 s 52808 0 52864 800 6 la_oen[108]
port 379 nsew default input
rlabel metal2 s 53176 0 53232 800 6 la_oen[109]
port 380 nsew default input
rlabel metal2 s 16836 0 16892 800 6 la_oen[10]
port 381 nsew default input
rlabel metal2 s 53544 0 53600 800 6 la_oen[110]
port 382 nsew default input
rlabel metal2 s 53912 0 53968 800 6 la_oen[111]
port 383 nsew default input
rlabel metal2 s 54280 0 54336 800 6 la_oen[112]
port 384 nsew default input
rlabel metal2 s 54648 0 54704 800 6 la_oen[113]
port 385 nsew default input
rlabel metal2 s 55016 0 55072 800 6 la_oen[114]
port 386 nsew default input
rlabel metal2 s 55384 0 55440 800 6 la_oen[115]
port 387 nsew default input
rlabel metal2 s 55752 0 55808 800 6 la_oen[116]
port 388 nsew default input
rlabel metal2 s 56120 0 56176 800 6 la_oen[117]
port 389 nsew default input
rlabel metal2 s 56488 0 56544 800 6 la_oen[118]
port 390 nsew default input
rlabel metal2 s 56856 0 56912 800 6 la_oen[119]
port 391 nsew default input
rlabel metal2 s 17204 0 17260 800 6 la_oen[11]
port 392 nsew default input
rlabel metal2 s 57224 0 57280 800 6 la_oen[120]
port 393 nsew default input
rlabel metal2 s 57592 0 57648 800 6 la_oen[121]
port 394 nsew default input
rlabel metal2 s 57960 0 58016 800 6 la_oen[122]
port 395 nsew default input
rlabel metal2 s 58328 0 58384 800 6 la_oen[123]
port 396 nsew default input
rlabel metal2 s 58696 0 58752 800 6 la_oen[124]
port 397 nsew default input
rlabel metal2 s 59064 0 59120 800 6 la_oen[125]
port 398 nsew default input
rlabel metal2 s 59432 0 59488 800 6 la_oen[126]
port 399 nsew default input
rlabel metal2 s 59800 0 59856 800 6 la_oen[127]
port 400 nsew default input
rlabel metal2 s 17572 0 17628 800 6 la_oen[12]
port 401 nsew default input
rlabel metal2 s 17940 0 17996 800 6 la_oen[13]
port 402 nsew default input
rlabel metal2 s 18308 0 18364 800 6 la_oen[14]
port 403 nsew default input
rlabel metal2 s 18676 0 18732 800 6 la_oen[15]
port 404 nsew default input
rlabel metal2 s 19044 0 19100 800 6 la_oen[16]
port 405 nsew default input
rlabel metal2 s 19412 0 19468 800 6 la_oen[17]
port 406 nsew default input
rlabel metal2 s 19780 0 19836 800 6 la_oen[18]
port 407 nsew default input
rlabel metal2 s 20148 0 20204 800 6 la_oen[19]
port 408 nsew default input
rlabel metal2 s 13524 0 13580 800 6 la_oen[1]
port 409 nsew default input
rlabel metal2 s 20516 0 20572 800 6 la_oen[20]
port 410 nsew default input
rlabel metal2 s 20884 0 20940 800 6 la_oen[21]
port 411 nsew default input
rlabel metal2 s 21252 0 21308 800 6 la_oen[22]
port 412 nsew default input
rlabel metal2 s 21620 0 21676 800 6 la_oen[23]
port 413 nsew default input
rlabel metal2 s 21988 0 22044 800 6 la_oen[24]
port 414 nsew default input
rlabel metal2 s 22356 0 22412 800 6 la_oen[25]
port 415 nsew default input
rlabel metal2 s 22724 0 22780 800 6 la_oen[26]
port 416 nsew default input
rlabel metal2 s 23092 0 23148 800 6 la_oen[27]
port 417 nsew default input
rlabel metal2 s 23460 0 23516 800 6 la_oen[28]
port 418 nsew default input
rlabel metal2 s 23828 0 23884 800 6 la_oen[29]
port 419 nsew default input
rlabel metal2 s 13892 0 13948 800 6 la_oen[2]
port 420 nsew default input
rlabel metal2 s 24196 0 24252 800 6 la_oen[30]
port 421 nsew default input
rlabel metal2 s 24564 0 24620 800 6 la_oen[31]
port 422 nsew default input
rlabel metal2 s 24932 0 24988 800 6 la_oen[32]
port 423 nsew default input
rlabel metal2 s 25300 0 25356 800 6 la_oen[33]
port 424 nsew default input
rlabel metal2 s 25668 0 25724 800 6 la_oen[34]
port 425 nsew default input
rlabel metal2 s 26036 0 26092 800 6 la_oen[35]
port 426 nsew default input
rlabel metal2 s 26404 0 26460 800 6 la_oen[36]
port 427 nsew default input
rlabel metal2 s 26772 0 26828 800 6 la_oen[37]
port 428 nsew default input
rlabel metal2 s 27140 0 27196 800 6 la_oen[38]
port 429 nsew default input
rlabel metal2 s 27508 0 27564 800 6 la_oen[39]
port 430 nsew default input
rlabel metal2 s 14260 0 14316 800 6 la_oen[3]
port 431 nsew default input
rlabel metal2 s 27876 0 27932 800 6 la_oen[40]
port 432 nsew default input
rlabel metal2 s 28244 0 28300 800 6 la_oen[41]
port 433 nsew default input
rlabel metal2 s 28612 0 28668 800 6 la_oen[42]
port 434 nsew default input
rlabel metal2 s 28980 0 29036 800 6 la_oen[43]
port 435 nsew default input
rlabel metal2 s 29348 0 29404 800 6 la_oen[44]
port 436 nsew default input
rlabel metal2 s 29716 0 29772 800 6 la_oen[45]
port 437 nsew default input
rlabel metal2 s 30084 0 30140 800 6 la_oen[46]
port 438 nsew default input
rlabel metal2 s 30452 0 30508 800 6 la_oen[47]
port 439 nsew default input
rlabel metal2 s 30820 0 30876 800 6 la_oen[48]
port 440 nsew default input
rlabel metal2 s 31188 0 31244 800 6 la_oen[49]
port 441 nsew default input
rlabel metal2 s 14628 0 14684 800 6 la_oen[4]
port 442 nsew default input
rlabel metal2 s 31556 0 31612 800 6 la_oen[50]
port 443 nsew default input
rlabel metal2 s 31924 0 31980 800 6 la_oen[51]
port 444 nsew default input
rlabel metal2 s 32292 0 32348 800 6 la_oen[52]
port 445 nsew default input
rlabel metal2 s 32660 0 32716 800 6 la_oen[53]
port 446 nsew default input
rlabel metal2 s 33028 0 33084 800 6 la_oen[54]
port 447 nsew default input
rlabel metal2 s 33396 0 33452 800 6 la_oen[55]
port 448 nsew default input
rlabel metal2 s 33764 0 33820 800 6 la_oen[56]
port 449 nsew default input
rlabel metal2 s 34132 0 34188 800 6 la_oen[57]
port 450 nsew default input
rlabel metal2 s 34500 0 34556 800 6 la_oen[58]
port 451 nsew default input
rlabel metal2 s 34868 0 34924 800 6 la_oen[59]
port 452 nsew default input
rlabel metal2 s 14996 0 15052 800 6 la_oen[5]
port 453 nsew default input
rlabel metal2 s 35236 0 35292 800 6 la_oen[60]
port 454 nsew default input
rlabel metal2 s 35604 0 35660 800 6 la_oen[61]
port 455 nsew default input
rlabel metal2 s 35972 0 36028 800 6 la_oen[62]
port 456 nsew default input
rlabel metal2 s 36340 0 36396 800 6 la_oen[63]
port 457 nsew default input
rlabel metal2 s 36708 0 36764 800 6 la_oen[64]
port 458 nsew default input
rlabel metal2 s 37076 0 37132 800 6 la_oen[65]
port 459 nsew default input
rlabel metal2 s 37444 0 37500 800 6 la_oen[66]
port 460 nsew default input
rlabel metal2 s 37812 0 37868 800 6 la_oen[67]
port 461 nsew default input
rlabel metal2 s 38180 0 38236 800 6 la_oen[68]
port 462 nsew default input
rlabel metal2 s 38548 0 38604 800 6 la_oen[69]
port 463 nsew default input
rlabel metal2 s 15364 0 15420 800 6 la_oen[6]
port 464 nsew default input
rlabel metal2 s 38916 0 38972 800 6 la_oen[70]
port 465 nsew default input
rlabel metal2 s 39284 0 39340 800 6 la_oen[71]
port 466 nsew default input
rlabel metal2 s 39652 0 39708 800 6 la_oen[72]
port 467 nsew default input
rlabel metal2 s 40020 0 40076 800 6 la_oen[73]
port 468 nsew default input
rlabel metal2 s 40388 0 40444 800 6 la_oen[74]
port 469 nsew default input
rlabel metal2 s 40756 0 40812 800 6 la_oen[75]
port 470 nsew default input
rlabel metal2 s 41124 0 41180 800 6 la_oen[76]
port 471 nsew default input
rlabel metal2 s 41492 0 41548 800 6 la_oen[77]
port 472 nsew default input
rlabel metal2 s 41860 0 41916 800 6 la_oen[78]
port 473 nsew default input
rlabel metal2 s 42228 0 42284 800 6 la_oen[79]
port 474 nsew default input
rlabel metal2 s 15732 0 15788 800 6 la_oen[7]
port 475 nsew default input
rlabel metal2 s 42596 0 42652 800 6 la_oen[80]
port 476 nsew default input
rlabel metal2 s 42964 0 43020 800 6 la_oen[81]
port 477 nsew default input
rlabel metal2 s 43332 0 43388 800 6 la_oen[82]
port 478 nsew default input
rlabel metal2 s 43700 0 43756 800 6 la_oen[83]
port 479 nsew default input
rlabel metal2 s 44068 0 44124 800 6 la_oen[84]
port 480 nsew default input
rlabel metal2 s 44436 0 44492 800 6 la_oen[85]
port 481 nsew default input
rlabel metal2 s 44804 0 44860 800 6 la_oen[86]
port 482 nsew default input
rlabel metal2 s 45080 0 45136 800 6 la_oen[87]
port 483 nsew default input
rlabel metal2 s 45448 0 45504 800 6 la_oen[88]
port 484 nsew default input
rlabel metal2 s 45816 0 45872 800 6 la_oen[89]
port 485 nsew default input
rlabel metal2 s 16100 0 16156 800 6 la_oen[8]
port 486 nsew default input
rlabel metal2 s 46184 0 46240 800 6 la_oen[90]
port 487 nsew default input
rlabel metal2 s 46552 0 46608 800 6 la_oen[91]
port 488 nsew default input
rlabel metal2 s 46920 0 46976 800 6 la_oen[92]
port 489 nsew default input
rlabel metal2 s 47288 0 47344 800 6 la_oen[93]
port 490 nsew default input
rlabel metal2 s 47656 0 47712 800 6 la_oen[94]
port 491 nsew default input
rlabel metal2 s 48024 0 48080 800 6 la_oen[95]
port 492 nsew default input
rlabel metal2 s 48392 0 48448 800 6 la_oen[96]
port 493 nsew default input
rlabel metal2 s 48760 0 48816 800 6 la_oen[97]
port 494 nsew default input
rlabel metal2 s 49128 0 49184 800 6 la_oen[98]
port 495 nsew default input
rlabel metal2 s 49496 0 49552 800 6 la_oen[99]
port 496 nsew default input
rlabel metal2 s 16468 0 16524 800 6 la_oen[9]
port 497 nsew default input
rlabel metal2 s 0 0 56 800 6 wb_clk_i
port 498 nsew default input
rlabel metal2 s 92 0 148 800 6 wb_rst_i
port 499 nsew default input
rlabel metal2 s 184 0 240 800 6 wbs_ack_o
port 500 nsew default tristate
rlabel metal2 s 644 0 700 800 6 wbs_adr_i[0]
port 501 nsew default input
rlabel metal2 s 4876 0 4932 800 6 wbs_adr_i[10]
port 502 nsew default input
rlabel metal2 s 5244 0 5300 800 6 wbs_adr_i[11]
port 503 nsew default input
rlabel metal2 s 5612 0 5668 800 6 wbs_adr_i[12]
port 504 nsew default input
rlabel metal2 s 5980 0 6036 800 6 wbs_adr_i[13]
port 505 nsew default input
rlabel metal2 s 6348 0 6404 800 6 wbs_adr_i[14]
port 506 nsew default input
rlabel metal2 s 6716 0 6772 800 6 wbs_adr_i[15]
port 507 nsew default input
rlabel metal2 s 7084 0 7140 800 6 wbs_adr_i[16]
port 508 nsew default input
rlabel metal2 s 7452 0 7508 800 6 wbs_adr_i[17]
port 509 nsew default input
rlabel metal2 s 7820 0 7876 800 6 wbs_adr_i[18]
port 510 nsew default input
rlabel metal2 s 8188 0 8244 800 6 wbs_adr_i[19]
port 511 nsew default input
rlabel metal2 s 1196 0 1252 800 6 wbs_adr_i[1]
port 512 nsew default input
rlabel metal2 s 8556 0 8612 800 6 wbs_adr_i[20]
port 513 nsew default input
rlabel metal2 s 8924 0 8980 800 6 wbs_adr_i[21]
port 514 nsew default input
rlabel metal2 s 9292 0 9348 800 6 wbs_adr_i[22]
port 515 nsew default input
rlabel metal2 s 9660 0 9716 800 6 wbs_adr_i[23]
port 516 nsew default input
rlabel metal2 s 10028 0 10084 800 6 wbs_adr_i[24]
port 517 nsew default input
rlabel metal2 s 10396 0 10452 800 6 wbs_adr_i[25]
port 518 nsew default input
rlabel metal2 s 10764 0 10820 800 6 wbs_adr_i[26]
port 519 nsew default input
rlabel metal2 s 11132 0 11188 800 6 wbs_adr_i[27]
port 520 nsew default input
rlabel metal2 s 11500 0 11556 800 6 wbs_adr_i[28]
port 521 nsew default input
rlabel metal2 s 11868 0 11924 800 6 wbs_adr_i[29]
port 522 nsew default input
rlabel metal2 s 1656 0 1712 800 6 wbs_adr_i[2]
port 523 nsew default input
rlabel metal2 s 12236 0 12292 800 6 wbs_adr_i[30]
port 524 nsew default input
rlabel metal2 s 12604 0 12660 800 6 wbs_adr_i[31]
port 525 nsew default input
rlabel metal2 s 2116 0 2172 800 6 wbs_adr_i[3]
port 526 nsew default input
rlabel metal2 s 2668 0 2724 800 6 wbs_adr_i[4]
port 527 nsew default input
rlabel metal2 s 3036 0 3092 800 6 wbs_adr_i[5]
port 528 nsew default input
rlabel metal2 s 3404 0 3460 800 6 wbs_adr_i[6]
port 529 nsew default input
rlabel metal2 s 3772 0 3828 800 6 wbs_adr_i[7]
port 530 nsew default input
rlabel metal2 s 4140 0 4196 800 6 wbs_adr_i[8]
port 531 nsew default input
rlabel metal2 s 4508 0 4564 800 6 wbs_adr_i[9]
port 532 nsew default input
rlabel metal2 s 276 0 332 800 6 wbs_cyc_i
port 533 nsew default input
rlabel metal2 s 828 0 884 800 6 wbs_dat_i[0]
port 534 nsew default input
rlabel metal2 s 4968 0 5024 800 6 wbs_dat_i[10]
port 535 nsew default input
rlabel metal2 s 5336 0 5392 800 6 wbs_dat_i[11]
port 536 nsew default input
rlabel metal2 s 5704 0 5760 800 6 wbs_dat_i[12]
port 537 nsew default input
rlabel metal2 s 6072 0 6128 800 6 wbs_dat_i[13]
port 538 nsew default input
rlabel metal2 s 6440 0 6496 800 6 wbs_dat_i[14]
port 539 nsew default input
rlabel metal2 s 6808 0 6864 800 6 wbs_dat_i[15]
port 540 nsew default input
rlabel metal2 s 7176 0 7232 800 6 wbs_dat_i[16]
port 541 nsew default input
rlabel metal2 s 7544 0 7600 800 6 wbs_dat_i[17]
port 542 nsew default input
rlabel metal2 s 7912 0 7968 800 6 wbs_dat_i[18]
port 543 nsew default input
rlabel metal2 s 8280 0 8336 800 6 wbs_dat_i[19]
port 544 nsew default input
rlabel metal2 s 1288 0 1344 800 6 wbs_dat_i[1]
port 545 nsew default input
rlabel metal2 s 8648 0 8704 800 6 wbs_dat_i[20]
port 546 nsew default input
rlabel metal2 s 9016 0 9072 800 6 wbs_dat_i[21]
port 547 nsew default input
rlabel metal2 s 9384 0 9440 800 6 wbs_dat_i[22]
port 548 nsew default input
rlabel metal2 s 9752 0 9808 800 6 wbs_dat_i[23]
port 549 nsew default input
rlabel metal2 s 10120 0 10176 800 6 wbs_dat_i[24]
port 550 nsew default input
rlabel metal2 s 10488 0 10544 800 6 wbs_dat_i[25]
port 551 nsew default input
rlabel metal2 s 10856 0 10912 800 6 wbs_dat_i[26]
port 552 nsew default input
rlabel metal2 s 11224 0 11280 800 6 wbs_dat_i[27]
port 553 nsew default input
rlabel metal2 s 11592 0 11648 800 6 wbs_dat_i[28]
port 554 nsew default input
rlabel metal2 s 11960 0 12016 800 6 wbs_dat_i[29]
port 555 nsew default input
rlabel metal2 s 1748 0 1804 800 6 wbs_dat_i[2]
port 556 nsew default input
rlabel metal2 s 12328 0 12384 800 6 wbs_dat_i[30]
port 557 nsew default input
rlabel metal2 s 12696 0 12752 800 6 wbs_dat_i[31]
port 558 nsew default input
rlabel metal2 s 2300 0 2356 800 6 wbs_dat_i[3]
port 559 nsew default input
rlabel metal2 s 2760 0 2816 800 6 wbs_dat_i[4]
port 560 nsew default input
rlabel metal2 s 3128 0 3184 800 6 wbs_dat_i[5]
port 561 nsew default input
rlabel metal2 s 3496 0 3552 800 6 wbs_dat_i[6]
port 562 nsew default input
rlabel metal2 s 3864 0 3920 800 6 wbs_dat_i[7]
port 563 nsew default input
rlabel metal2 s 4232 0 4288 800 6 wbs_dat_i[8]
port 564 nsew default input
rlabel metal2 s 4600 0 4656 800 6 wbs_dat_i[9]
port 565 nsew default input
rlabel metal2 s 920 0 976 800 6 wbs_dat_o[0]
port 566 nsew default tristate
rlabel metal2 s 5060 0 5116 800 6 wbs_dat_o[10]
port 567 nsew default tristate
rlabel metal2 s 5428 0 5484 800 6 wbs_dat_o[11]
port 568 nsew default tristate
rlabel metal2 s 5796 0 5852 800 6 wbs_dat_o[12]
port 569 nsew default tristate
rlabel metal2 s 6164 0 6220 800 6 wbs_dat_o[13]
port 570 nsew default tristate
rlabel metal2 s 6532 0 6588 800 6 wbs_dat_o[14]
port 571 nsew default tristate
rlabel metal2 s 6900 0 6956 800 6 wbs_dat_o[15]
port 572 nsew default tristate
rlabel metal2 s 7268 0 7324 800 6 wbs_dat_o[16]
port 573 nsew default tristate
rlabel metal2 s 7636 0 7692 800 6 wbs_dat_o[17]
port 574 nsew default tristate
rlabel metal2 s 8004 0 8060 800 6 wbs_dat_o[18]
port 575 nsew default tristate
rlabel metal2 s 8372 0 8428 800 6 wbs_dat_o[19]
port 576 nsew default tristate
rlabel metal2 s 1380 0 1436 800 6 wbs_dat_o[1]
port 577 nsew default tristate
rlabel metal2 s 8740 0 8796 800 6 wbs_dat_o[20]
port 578 nsew default tristate
rlabel metal2 s 9108 0 9164 800 6 wbs_dat_o[21]
port 579 nsew default tristate
rlabel metal2 s 9476 0 9532 800 6 wbs_dat_o[22]
port 580 nsew default tristate
rlabel metal2 s 9844 0 9900 800 6 wbs_dat_o[23]
port 581 nsew default tristate
rlabel metal2 s 10212 0 10268 800 6 wbs_dat_o[24]
port 582 nsew default tristate
rlabel metal2 s 10580 0 10636 800 6 wbs_dat_o[25]
port 583 nsew default tristate
rlabel metal2 s 10948 0 11004 800 6 wbs_dat_o[26]
port 584 nsew default tristate
rlabel metal2 s 11316 0 11372 800 6 wbs_dat_o[27]
port 585 nsew default tristate
rlabel metal2 s 11684 0 11740 800 6 wbs_dat_o[28]
port 586 nsew default tristate
rlabel metal2 s 12052 0 12108 800 6 wbs_dat_o[29]
port 587 nsew default tristate
rlabel metal2 s 1932 0 1988 800 6 wbs_dat_o[2]
port 588 nsew default tristate
rlabel metal2 s 12420 0 12476 800 6 wbs_dat_o[30]
port 589 nsew default tristate
rlabel metal2 s 12788 0 12844 800 6 wbs_dat_o[31]
port 590 nsew default tristate
rlabel metal2 s 2392 0 2448 800 6 wbs_dat_o[3]
port 591 nsew default tristate
rlabel metal2 s 2852 0 2908 800 6 wbs_dat_o[4]
port 592 nsew default tristate
rlabel metal2 s 3220 0 3276 800 6 wbs_dat_o[5]
port 593 nsew default tristate
rlabel metal2 s 3588 0 3644 800 6 wbs_dat_o[6]
port 594 nsew default tristate
rlabel metal2 s 3956 0 4012 800 6 wbs_dat_o[7]
port 595 nsew default tristate
rlabel metal2 s 4324 0 4380 800 6 wbs_dat_o[8]
port 596 nsew default tristate
rlabel metal2 s 4692 0 4748 800 6 wbs_dat_o[9]
port 597 nsew default tristate
rlabel metal2 s 1012 0 1068 800 6 wbs_sel_i[0]
port 598 nsew default input
rlabel metal2 s 1564 0 1620 800 6 wbs_sel_i[1]
port 599 nsew default input
rlabel metal2 s 2024 0 2080 800 6 wbs_sel_i[2]
port 600 nsew default input
rlabel metal2 s 2484 0 2540 800 6 wbs_sel_i[3]
port 601 nsew default input
rlabel metal2 s 460 0 516 800 6 wbs_stb_i
port 602 nsew default input
rlabel metal2 s 552 0 608 800 6 wbs_we_i
port 603 nsew default input
rlabel metal4 s 4190 2128 4510 57712 6 VPWR
port 604 nsew default input
rlabel metal4 s 19550 2128 19870 57712 6 VGND
port 605 nsew default input
<< properties >>
string FIXED_BBOX 0 0 59856 60000
<< end >>
