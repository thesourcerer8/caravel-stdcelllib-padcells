VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO NOR3X1
  CLASS CORE ;
  FOREIGN NOR3X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.440 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
        RECT 0.000 2.480 6.440 2.960 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
        RECT 0.000 -0.240 6.440 0.240 ;
    END
  END gnd
  PIN Y
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
        RECT 0.320 1.740 0.610 2.030 ;
        RECT 5.840 1.740 6.130 2.030 ;
        RECT 0.390 0.920 0.530 1.740 ;
        RECT 5.910 0.920 6.050 1.740 ;
        RECT 0.390 0.780 6.050 0.920 ;
        RECT 1.240 0.570 1.530 0.780 ;
        RECT 3.080 0.570 3.370 0.780 ;
    END
  END Y
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
        RECT 2.620 1.310 2.910 1.380 ;
        RECT 3.540 1.310 3.830 1.510 ;
        RECT 2.620 1.220 3.830 1.310 ;
        RECT 2.620 1.170 3.750 1.220 ;
        RECT 2.620 1.090 2.910 1.170 ;
    END
  END A
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
        RECT 4.460 1.350 4.750 1.640 ;
    END
    PORT
      LAYER met2 ;
        RECT 1.700 1.090 1.990 1.640 ;
    END
  END B
  PIN C
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
        RECT 5.380 1.350 5.670 1.640 ;
    END
    PORT
      LAYER met2 ;
        RECT 0.780 1.090 1.070 1.640 ;
    END
  END C
END NOR3X1
END LIBRARY

