magic
tech sky130A
timestamp 1607791616
<< end >>
