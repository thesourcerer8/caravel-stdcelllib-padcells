VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_project_wrapper
  CLASS BLOCK ;
  FOREIGN user_project_wrapper ;
  ORIGIN 0.000 0.000 ;
  SIZE 2920.000 BY 3520.000 ;
  PIN analog_io[0]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 28.980 2924.800 30.180 ;
    END
  END analog_io[0]
  PIN analog_io[10]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2374.980 2924.800 2376.180 ;
    END
  END analog_io[10]
  PIN analog_io[11]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2609.580 2924.800 2610.780 ;
    END
  END analog_io[11]
  PIN analog_io[12]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2844.180 2924.800 2845.380 ;
    END
  END analog_io[12]
  PIN analog_io[13]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3078.780 2924.800 3079.980 ;
    END
  END analog_io[13]
  PIN analog_io[14]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 3313.380 2924.800 3314.580 ;
    END
  END analog_io[14]
  PIN analog_io[15]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2879.090 3517.600 2879.650 3524.800 ;
    END
  END analog_io[15]
  PIN analog_io[16]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2554.790 3517.600 2555.350 3524.800 ;
    END
  END analog_io[16]
  PIN analog_io[17]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 2230.490 3517.600 2231.050 3524.800 ;
    END
  END analog_io[17]
  PIN analog_io[18]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1905.730 3517.600 1906.290 3524.800 ;
    END
  END analog_io[18]
  PIN analog_io[19]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1581.430 3517.600 1581.990 3524.800 ;
    END
  END analog_io[19]
  PIN analog_io[1]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 263.580 2924.800 264.780 ;
    END
  END analog_io[1]
  PIN analog_io[20]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 1257.130 3517.600 1257.690 3524.800 ;
    END
  END analog_io[20]
  PIN analog_io[21]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 932.370 3517.600 932.930 3524.800 ;
    END
  END analog_io[21]
  PIN analog_io[22]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 608.070 3517.600 608.630 3524.800 ;
    END
  END analog_io[22]
  PIN analog_io[23]
    DIRECTION INOUT ;
    PORT
      LAYER met2 ;
        RECT 283.770 3517.600 284.330 3524.800 ;
    END
  END analog_io[23]
  PIN analog_io[24]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3482.700 2.400 3483.900 ;
    END
  END analog_io[24]
  PIN analog_io[25]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 3195.060 2.400 3196.260 ;
    END
  END analog_io[25]
  PIN analog_io[26]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2908.100 2.400 2909.300 ;
    END
  END analog_io[26]
  PIN analog_io[27]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2620.460 2.400 2621.660 ;
    END
  END analog_io[27]
  PIN analog_io[28]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2333.500 2.400 2334.700 ;
    END
  END analog_io[28]
  PIN analog_io[29]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 2045.860 2.400 2047.060 ;
    END
  END analog_io[29]
  PIN analog_io[2]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 498.180 2924.800 499.380 ;
    END
  END analog_io[2]
  PIN analog_io[30]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT -4.800 1758.900 2.400 1760.100 ;
    END
  END analog_io[30]
  PIN analog_io[3]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 732.780 2924.800 733.980 ;
    END
  END analog_io[3]
  PIN analog_io[4]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 967.380 2924.800 968.580 ;
    END
  END analog_io[4]
  PIN analog_io[5]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1201.980 2924.800 1203.180 ;
    END
  END analog_io[5]
  PIN analog_io[6]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1436.580 2924.800 1437.780 ;
    END
  END analog_io[6]
  PIN analog_io[7]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1671.180 2924.800 1672.380 ;
    END
  END analog_io[7]
  PIN analog_io[8]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 1905.780 2924.800 1906.980 ;
    END
  END analog_io[8]
  PIN analog_io[9]
    DIRECTION INOUT ;
    PORT
      LAYER met3 ;
        RECT 2917.600 2140.380 2924.800 2141.580 ;
    END
  END analog_io[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1145.470 89.660 1145.790 89.720 ;
        RECT 2898.990 89.660 2899.310 89.720 ;
        RECT 1145.470 89.520 2899.310 89.660 ;
        RECT 1145.470 89.460 1145.790 89.520 ;
        RECT 2898.990 89.460 2899.310 89.520 ;
      LAYER via ;
        RECT 1145.500 89.460 1145.760 89.720 ;
        RECT 2899.020 89.460 2899.280 89.720 ;
      LAYER met2 ;
        RECT 1150.920 1996.210 1151.200 2000.000 ;
        RECT 1145.560 1996.070 1151.200 1996.210 ;
        RECT 1145.560 89.750 1145.700 1996.070 ;
        RECT 1150.920 1996.000 1151.200 1996.070 ;
        RECT 1145.500 89.430 1145.760 89.750 ;
        RECT 2899.020 89.430 2899.280 89.750 ;
        RECT 2899.080 88.245 2899.220 89.430 ;
        RECT 2899.010 87.875 2899.290 88.245 ;
      LAYER via2 ;
        RECT 2899.010 87.920 2899.290 88.200 ;
      LAYER met3 ;
        RECT 2898.985 88.210 2899.315 88.225 ;
        RECT 2917.600 88.210 2924.800 88.660 ;
        RECT 2898.985 87.910 2924.800 88.210 ;
        RECT 2898.985 87.895 2899.315 87.910 ;
        RECT 2917.600 87.460 2924.800 87.910 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1234.250 2429.200 1234.570 2429.260 ;
        RECT 2900.830 2429.200 2901.150 2429.260 ;
        RECT 1234.250 2429.060 2901.150 2429.200 ;
        RECT 1234.250 2429.000 1234.570 2429.060 ;
        RECT 2900.830 2429.000 2901.150 2429.060 ;
        RECT 1229.650 2009.300 1229.970 2009.360 ;
        RECT 1234.250 2009.300 1234.570 2009.360 ;
        RECT 1229.650 2009.160 1234.570 2009.300 ;
        RECT 1229.650 2009.100 1229.970 2009.160 ;
        RECT 1234.250 2009.100 1234.570 2009.160 ;
      LAYER via ;
        RECT 1234.280 2429.000 1234.540 2429.260 ;
        RECT 2900.860 2429.000 2901.120 2429.260 ;
        RECT 1229.680 2009.100 1229.940 2009.360 ;
        RECT 1234.280 2009.100 1234.540 2009.360 ;
      LAYER met2 ;
        RECT 2900.850 2433.875 2901.130 2434.245 ;
        RECT 2900.920 2429.290 2901.060 2433.875 ;
        RECT 1234.280 2428.970 1234.540 2429.290 ;
        RECT 2900.860 2428.970 2901.120 2429.290 ;
        RECT 1234.340 2009.390 1234.480 2428.970 ;
        RECT 1229.680 2009.070 1229.940 2009.390 ;
        RECT 1234.280 2009.070 1234.540 2009.390 ;
        RECT 1229.740 2000.000 1229.880 2009.070 ;
        RECT 1229.580 1999.540 1229.880 2000.000 ;
        RECT 1229.580 1996.000 1229.860 1999.540 ;
      LAYER via2 ;
        RECT 2900.850 2433.920 2901.130 2434.200 ;
      LAYER met3 ;
        RECT 2900.825 2434.210 2901.155 2434.225 ;
        RECT 2917.600 2434.210 2924.800 2434.660 ;
        RECT 2900.825 2433.910 2924.800 2434.210 ;
        RECT 2900.825 2433.895 2901.155 2433.910 ;
        RECT 2917.600 2433.460 2924.800 2433.910 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1241.150 2663.800 1241.470 2663.860 ;
        RECT 2900.830 2663.800 2901.150 2663.860 ;
        RECT 1241.150 2663.660 2901.150 2663.800 ;
        RECT 1241.150 2663.600 1241.470 2663.660 ;
        RECT 2900.830 2663.600 2901.150 2663.660 ;
        RECT 1237.470 2009.300 1237.790 2009.360 ;
        RECT 1241.150 2009.300 1241.470 2009.360 ;
        RECT 1237.470 2009.160 1241.470 2009.300 ;
        RECT 1237.470 2009.100 1237.790 2009.160 ;
        RECT 1241.150 2009.100 1241.470 2009.160 ;
      LAYER via ;
        RECT 1241.180 2663.600 1241.440 2663.860 ;
        RECT 2900.860 2663.600 2901.120 2663.860 ;
        RECT 1237.500 2009.100 1237.760 2009.360 ;
        RECT 1241.180 2009.100 1241.440 2009.360 ;
      LAYER met2 ;
        RECT 2900.850 2669.155 2901.130 2669.525 ;
        RECT 2900.920 2663.890 2901.060 2669.155 ;
        RECT 1241.180 2663.570 1241.440 2663.890 ;
        RECT 2900.860 2663.570 2901.120 2663.890 ;
        RECT 1241.240 2009.390 1241.380 2663.570 ;
        RECT 1237.500 2009.070 1237.760 2009.390 ;
        RECT 1241.180 2009.070 1241.440 2009.390 ;
        RECT 1237.560 2000.000 1237.700 2009.070 ;
        RECT 1237.400 1999.540 1237.700 2000.000 ;
        RECT 1237.400 1996.000 1237.680 1999.540 ;
      LAYER via2 ;
        RECT 2900.850 2669.200 2901.130 2669.480 ;
      LAYER met3 ;
        RECT 2900.825 2669.490 2901.155 2669.505 ;
        RECT 2917.600 2669.490 2924.800 2669.940 ;
        RECT 2900.825 2669.190 2924.800 2669.490 ;
        RECT 2900.825 2669.175 2901.155 2669.190 ;
        RECT 2917.600 2668.740 2924.800 2669.190 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1248.050 2898.400 1248.370 2898.460 ;
        RECT 2900.830 2898.400 2901.150 2898.460 ;
        RECT 1248.050 2898.260 2901.150 2898.400 ;
        RECT 1248.050 2898.200 1248.370 2898.260 ;
        RECT 2900.830 2898.200 2901.150 2898.260 ;
      LAYER via ;
        RECT 1248.080 2898.200 1248.340 2898.460 ;
        RECT 2900.860 2898.200 2901.120 2898.460 ;
      LAYER met2 ;
        RECT 2900.850 2903.755 2901.130 2904.125 ;
        RECT 2900.920 2898.490 2901.060 2903.755 ;
        RECT 1248.080 2898.170 1248.340 2898.490 ;
        RECT 2900.860 2898.170 2901.120 2898.490 ;
        RECT 1248.140 2001.650 1248.280 2898.170 ;
        RECT 1247.680 2001.510 1248.280 2001.650 ;
        RECT 1245.220 1999.610 1245.500 2000.000 ;
        RECT 1247.680 1999.610 1247.820 2001.510 ;
        RECT 1245.220 1999.470 1247.820 1999.610 ;
        RECT 1245.220 1996.000 1245.500 1999.470 ;
      LAYER via2 ;
        RECT 2900.850 2903.800 2901.130 2904.080 ;
      LAYER met3 ;
        RECT 2900.825 2904.090 2901.155 2904.105 ;
        RECT 2917.600 2904.090 2924.800 2904.540 ;
        RECT 2900.825 2903.790 2924.800 2904.090 ;
        RECT 2900.825 2903.775 2901.155 2903.790 ;
        RECT 2917.600 2903.340 2924.800 2903.790 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1255.410 3133.000 1255.730 3133.060 ;
        RECT 2900.830 3133.000 2901.150 3133.060 ;
        RECT 1255.410 3132.860 2901.150 3133.000 ;
        RECT 1255.410 3132.800 1255.730 3132.860 ;
        RECT 2900.830 3132.800 2901.150 3132.860 ;
      LAYER via ;
        RECT 1255.440 3132.800 1255.700 3133.060 ;
        RECT 2900.860 3132.800 2901.120 3133.060 ;
      LAYER met2 ;
        RECT 2900.850 3138.355 2901.130 3138.725 ;
        RECT 2900.920 3133.090 2901.060 3138.355 ;
        RECT 1255.440 3132.770 1255.700 3133.090 ;
        RECT 2900.860 3132.770 2901.120 3133.090 ;
        RECT 1253.500 1999.610 1253.780 2000.000 ;
        RECT 1255.500 1999.610 1255.640 3132.770 ;
        RECT 1253.500 1999.470 1255.640 1999.610 ;
        RECT 1253.500 1996.000 1253.780 1999.470 ;
      LAYER via2 ;
        RECT 2900.850 3138.400 2901.130 3138.680 ;
      LAYER met3 ;
        RECT 2900.825 3138.690 2901.155 3138.705 ;
        RECT 2917.600 3138.690 2924.800 3139.140 ;
        RECT 2900.825 3138.390 2924.800 3138.690 ;
        RECT 2900.825 3138.375 2901.155 3138.390 ;
        RECT 2917.600 3137.940 2924.800 3138.390 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1262.310 3367.600 1262.630 3367.660 ;
        RECT 2900.830 3367.600 2901.150 3367.660 ;
        RECT 1262.310 3367.460 2901.150 3367.600 ;
        RECT 1262.310 3367.400 1262.630 3367.460 ;
        RECT 2900.830 3367.400 2901.150 3367.460 ;
      LAYER via ;
        RECT 1262.340 3367.400 1262.600 3367.660 ;
        RECT 2900.860 3367.400 2901.120 3367.660 ;
      LAYER met2 ;
        RECT 2900.850 3372.955 2901.130 3373.325 ;
        RECT 2900.920 3367.690 2901.060 3372.955 ;
        RECT 1262.340 3367.370 1262.600 3367.690 ;
        RECT 2900.860 3367.370 2901.120 3367.690 ;
        RECT 1261.320 1999.610 1261.600 2000.000 ;
        RECT 1262.400 1999.610 1262.540 3367.370 ;
        RECT 1261.320 1999.470 1262.540 1999.610 ;
        RECT 1261.320 1996.000 1261.600 1999.470 ;
      LAYER via2 ;
        RECT 2900.850 3373.000 2901.130 3373.280 ;
      LAYER met3 ;
        RECT 2900.825 3373.290 2901.155 3373.305 ;
        RECT 2917.600 3373.290 2924.800 3373.740 ;
        RECT 2900.825 3372.990 2924.800 3373.290 ;
        RECT 2900.825 3372.975 2901.155 3372.990 ;
        RECT 2917.600 3372.540 2924.800 3372.990 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1269.210 3501.560 1269.530 3501.620 ;
        RECT 2798.250 3501.560 2798.570 3501.620 ;
        RECT 1269.210 3501.420 2798.570 3501.560 ;
        RECT 1269.210 3501.360 1269.530 3501.420 ;
        RECT 2798.250 3501.360 2798.570 3501.420 ;
      LAYER via ;
        RECT 1269.240 3501.360 1269.500 3501.620 ;
        RECT 2798.280 3501.360 2798.540 3501.620 ;
      LAYER met2 ;
        RECT 2798.130 3517.600 2798.690 3524.800 ;
        RECT 2798.340 3501.650 2798.480 3517.600 ;
        RECT 1269.240 3501.330 1269.500 3501.650 ;
        RECT 2798.280 3501.330 2798.540 3501.650 ;
        RECT 1269.300 2000.000 1269.440 3501.330 ;
        RECT 1269.140 1999.540 1269.440 2000.000 ;
        RECT 1269.140 1996.000 1269.420 1999.540 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1282.090 3502.920 1282.410 3502.980 ;
        RECT 2473.950 3502.920 2474.270 3502.980 ;
        RECT 1282.090 3502.780 2474.270 3502.920 ;
        RECT 1282.090 3502.720 1282.410 3502.780 ;
        RECT 2473.950 3502.720 2474.270 3502.780 ;
        RECT 1277.030 2014.400 1277.350 2014.460 ;
        RECT 1282.090 2014.400 1282.410 2014.460 ;
        RECT 1277.030 2014.260 1282.410 2014.400 ;
        RECT 1277.030 2014.200 1277.350 2014.260 ;
        RECT 1282.090 2014.200 1282.410 2014.260 ;
      LAYER via ;
        RECT 1282.120 3502.720 1282.380 3502.980 ;
        RECT 2473.980 3502.720 2474.240 3502.980 ;
        RECT 1277.060 2014.200 1277.320 2014.460 ;
        RECT 1282.120 2014.200 1282.380 2014.460 ;
      LAYER met2 ;
        RECT 2473.830 3517.600 2474.390 3524.800 ;
        RECT 2474.040 3503.010 2474.180 3517.600 ;
        RECT 1282.120 3502.690 1282.380 3503.010 ;
        RECT 2473.980 3502.690 2474.240 3503.010 ;
        RECT 1282.180 2014.490 1282.320 3502.690 ;
        RECT 1277.060 2014.170 1277.320 2014.490 ;
        RECT 1282.120 2014.170 1282.380 2014.490 ;
        RECT 1277.120 2000.000 1277.260 2014.170 ;
        RECT 1276.960 1999.540 1277.260 2000.000 ;
        RECT 1276.960 1996.000 1277.240 1999.540 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1289.910 3504.280 1290.230 3504.340 ;
        RECT 2149.190 3504.280 2149.510 3504.340 ;
        RECT 1289.910 3504.140 2149.510 3504.280 ;
        RECT 1289.910 3504.080 1290.230 3504.140 ;
        RECT 2149.190 3504.080 2149.510 3504.140 ;
        RECT 1284.850 2014.400 1285.170 2014.460 ;
        RECT 1289.910 2014.400 1290.230 2014.460 ;
        RECT 1284.850 2014.260 1290.230 2014.400 ;
        RECT 1284.850 2014.200 1285.170 2014.260 ;
        RECT 1289.910 2014.200 1290.230 2014.260 ;
      LAYER via ;
        RECT 1289.940 3504.080 1290.200 3504.340 ;
        RECT 2149.220 3504.080 2149.480 3504.340 ;
        RECT 1284.880 2014.200 1285.140 2014.460 ;
        RECT 1289.940 2014.200 1290.200 2014.460 ;
      LAYER met2 ;
        RECT 2149.070 3517.600 2149.630 3524.800 ;
        RECT 2149.280 3504.370 2149.420 3517.600 ;
        RECT 1289.940 3504.050 1290.200 3504.370 ;
        RECT 2149.220 3504.050 2149.480 3504.370 ;
        RECT 1290.000 2014.490 1290.140 3504.050 ;
        RECT 1284.880 2014.170 1285.140 2014.490 ;
        RECT 1289.940 2014.170 1290.200 2014.490 ;
        RECT 1284.940 2000.000 1285.080 2014.170 ;
        RECT 1284.780 1999.540 1285.080 2000.000 ;
        RECT 1284.780 1996.000 1285.060 1999.540 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1296.350 3500.880 1296.670 3500.940 ;
        RECT 1824.890 3500.880 1825.210 3500.940 ;
        RECT 1296.350 3500.740 1825.210 3500.880 ;
        RECT 1296.350 3500.680 1296.670 3500.740 ;
        RECT 1824.890 3500.680 1825.210 3500.740 ;
        RECT 1292.670 2014.400 1292.990 2014.460 ;
        RECT 1296.350 2014.400 1296.670 2014.460 ;
        RECT 1292.670 2014.260 1296.670 2014.400 ;
        RECT 1292.670 2014.200 1292.990 2014.260 ;
        RECT 1296.350 2014.200 1296.670 2014.260 ;
      LAYER via ;
        RECT 1296.380 3500.680 1296.640 3500.940 ;
        RECT 1824.920 3500.680 1825.180 3500.940 ;
        RECT 1292.700 2014.200 1292.960 2014.460 ;
        RECT 1296.380 2014.200 1296.640 2014.460 ;
      LAYER met2 ;
        RECT 1824.770 3517.600 1825.330 3524.800 ;
        RECT 1824.980 3500.970 1825.120 3517.600 ;
        RECT 1296.380 3500.650 1296.640 3500.970 ;
        RECT 1824.920 3500.650 1825.180 3500.970 ;
        RECT 1296.440 2014.490 1296.580 3500.650 ;
        RECT 1292.700 2014.170 1292.960 2014.490 ;
        RECT 1296.380 2014.170 1296.640 2014.490 ;
        RECT 1292.760 2000.000 1292.900 2014.170 ;
        RECT 1292.600 1999.540 1292.900 2000.000 ;
        RECT 1292.600 1996.000 1292.880 1999.540 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1499.285 3332.765 1499.455 3422.355 ;
        RECT 1498.365 3008.405 1498.535 3042.915 ;
        RECT 1499.285 2946.525 1499.455 2994.635 ;
        RECT 1498.365 2428.705 1498.535 2463.215 ;
        RECT 1498.365 2331.805 1498.535 2366.655 ;
        RECT 1497.445 2201.245 1497.615 2249.355 ;
        RECT 1497.905 2138.685 1498.075 2184.075 ;
        RECT 1498.365 2028.525 1498.535 2076.975 ;
      LAYER mcon ;
        RECT 1499.285 3422.185 1499.455 3422.355 ;
        RECT 1498.365 3042.745 1498.535 3042.915 ;
        RECT 1499.285 2994.465 1499.455 2994.635 ;
        RECT 1498.365 2463.045 1498.535 2463.215 ;
        RECT 1498.365 2366.485 1498.535 2366.655 ;
        RECT 1497.445 2249.185 1497.615 2249.355 ;
        RECT 1497.905 2183.905 1498.075 2184.075 ;
        RECT 1498.365 2076.805 1498.535 2076.975 ;
      LAYER met1 ;
        RECT 1498.290 3443.080 1498.610 3443.140 ;
        RECT 1500.590 3443.080 1500.910 3443.140 ;
        RECT 1498.290 3442.940 1500.910 3443.080 ;
        RECT 1498.290 3442.880 1498.610 3442.940 ;
        RECT 1500.590 3442.880 1500.910 3442.940 ;
        RECT 1497.830 3422.340 1498.150 3422.400 ;
        RECT 1499.225 3422.340 1499.515 3422.385 ;
        RECT 1497.830 3422.200 1499.515 3422.340 ;
        RECT 1497.830 3422.140 1498.150 3422.200 ;
        RECT 1499.225 3422.155 1499.515 3422.200 ;
        RECT 1499.225 3332.920 1499.515 3332.965 ;
        RECT 1499.670 3332.920 1499.990 3332.980 ;
        RECT 1499.225 3332.780 1499.990 3332.920 ;
        RECT 1499.225 3332.735 1499.515 3332.780 ;
        RECT 1499.670 3332.720 1499.990 3332.780 ;
        RECT 1498.290 3236.360 1498.610 3236.420 ;
        RECT 1498.750 3236.360 1499.070 3236.420 ;
        RECT 1498.290 3236.220 1499.070 3236.360 ;
        RECT 1498.290 3236.160 1498.610 3236.220 ;
        RECT 1498.750 3236.160 1499.070 3236.220 ;
        RECT 1498.290 3202.020 1498.610 3202.080 ;
        RECT 1498.750 3202.020 1499.070 3202.080 ;
        RECT 1498.290 3201.880 1499.070 3202.020 ;
        RECT 1498.290 3201.820 1498.610 3201.880 ;
        RECT 1498.750 3201.820 1499.070 3201.880 ;
        RECT 1497.830 3153.400 1498.150 3153.460 ;
        RECT 1498.750 3153.400 1499.070 3153.460 ;
        RECT 1497.830 3153.260 1499.070 3153.400 ;
        RECT 1497.830 3153.200 1498.150 3153.260 ;
        RECT 1498.750 3153.200 1499.070 3153.260 ;
        RECT 1497.830 3056.840 1498.150 3056.900 ;
        RECT 1498.750 3056.840 1499.070 3056.900 ;
        RECT 1497.830 3056.700 1499.070 3056.840 ;
        RECT 1497.830 3056.640 1498.150 3056.700 ;
        RECT 1498.750 3056.640 1499.070 3056.700 ;
        RECT 1498.290 3042.900 1498.610 3042.960 ;
        RECT 1498.095 3042.760 1498.610 3042.900 ;
        RECT 1498.290 3042.700 1498.610 3042.760 ;
        RECT 1498.305 3008.560 1498.595 3008.605 ;
        RECT 1499.210 3008.560 1499.530 3008.620 ;
        RECT 1498.305 3008.420 1499.530 3008.560 ;
        RECT 1498.305 3008.375 1498.595 3008.420 ;
        RECT 1499.210 3008.360 1499.530 3008.420 ;
        RECT 1499.210 2994.620 1499.530 2994.680 ;
        RECT 1499.015 2994.480 1499.530 2994.620 ;
        RECT 1499.210 2994.420 1499.530 2994.480 ;
        RECT 1499.225 2946.680 1499.515 2946.725 ;
        RECT 1499.670 2946.680 1499.990 2946.740 ;
        RECT 1499.225 2946.540 1499.990 2946.680 ;
        RECT 1499.225 2946.495 1499.515 2946.540 ;
        RECT 1499.670 2946.480 1499.990 2946.540 ;
        RECT 1499.670 2912.340 1499.990 2912.400 ;
        RECT 1499.300 2912.200 1499.990 2912.340 ;
        RECT 1499.300 2911.720 1499.440 2912.200 ;
        RECT 1499.670 2912.140 1499.990 2912.200 ;
        RECT 1499.210 2911.460 1499.530 2911.720 ;
        RECT 1497.830 2815.580 1498.150 2815.840 ;
        RECT 1497.920 2815.160 1498.060 2815.580 ;
        RECT 1497.830 2814.900 1498.150 2815.160 ;
        RECT 1497.830 2767.500 1498.150 2767.560 ;
        RECT 1497.460 2767.360 1498.150 2767.500 ;
        RECT 1497.460 2766.880 1497.600 2767.360 ;
        RECT 1497.830 2767.300 1498.150 2767.360 ;
        RECT 1497.370 2766.620 1497.690 2766.880 ;
        RECT 1496.450 2718.540 1496.770 2718.600 ;
        RECT 1497.370 2718.540 1497.690 2718.600 ;
        RECT 1496.450 2718.400 1497.690 2718.540 ;
        RECT 1496.450 2718.340 1496.770 2718.400 ;
        RECT 1497.370 2718.340 1497.690 2718.400 ;
        RECT 1497.830 2656.660 1498.150 2656.720 ;
        RECT 1498.750 2656.660 1499.070 2656.720 ;
        RECT 1497.830 2656.520 1499.070 2656.660 ;
        RECT 1497.830 2656.460 1498.150 2656.520 ;
        RECT 1498.750 2656.460 1499.070 2656.520 ;
        RECT 1498.750 2622.120 1499.070 2622.380 ;
        RECT 1498.840 2621.980 1498.980 2622.120 ;
        RECT 1499.210 2621.980 1499.530 2622.040 ;
        RECT 1498.840 2621.840 1499.530 2621.980 ;
        RECT 1499.210 2621.780 1499.530 2621.840 ;
        RECT 1498.290 2560.100 1498.610 2560.160 ;
        RECT 1499.670 2560.100 1499.990 2560.160 ;
        RECT 1498.290 2559.960 1499.990 2560.100 ;
        RECT 1498.290 2559.900 1498.610 2559.960 ;
        RECT 1499.670 2559.900 1499.990 2559.960 ;
        RECT 1498.750 2511.820 1499.070 2511.880 ;
        RECT 1499.670 2511.820 1499.990 2511.880 ;
        RECT 1498.750 2511.680 1499.990 2511.820 ;
        RECT 1498.750 2511.620 1499.070 2511.680 ;
        RECT 1499.670 2511.620 1499.990 2511.680 ;
        RECT 1498.290 2463.200 1498.610 2463.260 ;
        RECT 1498.095 2463.060 1498.610 2463.200 ;
        RECT 1498.290 2463.000 1498.610 2463.060 ;
        RECT 1498.290 2428.860 1498.610 2428.920 ;
        RECT 1498.095 2428.720 1498.610 2428.860 ;
        RECT 1498.290 2428.660 1498.610 2428.720 ;
        RECT 1497.830 2380.580 1498.150 2380.640 ;
        RECT 1498.750 2380.580 1499.070 2380.640 ;
        RECT 1497.830 2380.440 1499.070 2380.580 ;
        RECT 1497.830 2380.380 1498.150 2380.440 ;
        RECT 1498.750 2380.380 1499.070 2380.440 ;
        RECT 1498.290 2366.640 1498.610 2366.700 ;
        RECT 1498.095 2366.500 1498.610 2366.640 ;
        RECT 1498.290 2366.440 1498.610 2366.500 ;
        RECT 1498.290 2331.960 1498.610 2332.020 ;
        RECT 1498.095 2331.820 1498.610 2331.960 ;
        RECT 1498.290 2331.760 1498.610 2331.820 ;
        RECT 1496.910 2304.420 1497.230 2304.480 ;
        RECT 1498.750 2304.420 1499.070 2304.480 ;
        RECT 1496.910 2304.280 1499.070 2304.420 ;
        RECT 1496.910 2304.220 1497.230 2304.280 ;
        RECT 1498.750 2304.220 1499.070 2304.280 ;
        RECT 1497.370 2249.340 1497.690 2249.400 ;
        RECT 1497.175 2249.200 1497.690 2249.340 ;
        RECT 1497.370 2249.140 1497.690 2249.200 ;
        RECT 1497.385 2201.400 1497.675 2201.445 ;
        RECT 1497.830 2201.400 1498.150 2201.460 ;
        RECT 1497.385 2201.260 1498.150 2201.400 ;
        RECT 1497.385 2201.215 1497.675 2201.260 ;
        RECT 1497.830 2201.200 1498.150 2201.260 ;
        RECT 1497.830 2184.060 1498.150 2184.120 ;
        RECT 1497.635 2183.920 1498.150 2184.060 ;
        RECT 1497.830 2183.860 1498.150 2183.920 ;
        RECT 1497.830 2138.840 1498.150 2138.900 ;
        RECT 1497.635 2138.700 1498.150 2138.840 ;
        RECT 1497.830 2138.640 1498.150 2138.700 ;
        RECT 1498.305 2076.960 1498.595 2077.005 ;
        RECT 1498.750 2076.960 1499.070 2077.020 ;
        RECT 1498.305 2076.820 1499.070 2076.960 ;
        RECT 1498.305 2076.775 1498.595 2076.820 ;
        RECT 1498.750 2076.760 1499.070 2076.820 ;
        RECT 1498.290 2028.680 1498.610 2028.740 ;
        RECT 1498.095 2028.540 1498.610 2028.680 ;
        RECT 1498.290 2028.480 1498.610 2028.540 ;
        RECT 1300.950 2009.980 1301.270 2010.040 ;
        RECT 1498.290 2009.980 1498.610 2010.040 ;
        RECT 1300.950 2009.840 1498.610 2009.980 ;
        RECT 1300.950 2009.780 1301.270 2009.840 ;
        RECT 1498.290 2009.780 1498.610 2009.840 ;
      LAYER via ;
        RECT 1498.320 3442.880 1498.580 3443.140 ;
        RECT 1500.620 3442.880 1500.880 3443.140 ;
        RECT 1497.860 3422.140 1498.120 3422.400 ;
        RECT 1499.700 3332.720 1499.960 3332.980 ;
        RECT 1498.320 3236.160 1498.580 3236.420 ;
        RECT 1498.780 3236.160 1499.040 3236.420 ;
        RECT 1498.320 3201.820 1498.580 3202.080 ;
        RECT 1498.780 3201.820 1499.040 3202.080 ;
        RECT 1497.860 3153.200 1498.120 3153.460 ;
        RECT 1498.780 3153.200 1499.040 3153.460 ;
        RECT 1497.860 3056.640 1498.120 3056.900 ;
        RECT 1498.780 3056.640 1499.040 3056.900 ;
        RECT 1498.320 3042.700 1498.580 3042.960 ;
        RECT 1499.240 3008.360 1499.500 3008.620 ;
        RECT 1499.240 2994.420 1499.500 2994.680 ;
        RECT 1499.700 2946.480 1499.960 2946.740 ;
        RECT 1499.700 2912.140 1499.960 2912.400 ;
        RECT 1499.240 2911.460 1499.500 2911.720 ;
        RECT 1497.860 2815.580 1498.120 2815.840 ;
        RECT 1497.860 2814.900 1498.120 2815.160 ;
        RECT 1497.860 2767.300 1498.120 2767.560 ;
        RECT 1497.400 2766.620 1497.660 2766.880 ;
        RECT 1496.480 2718.340 1496.740 2718.600 ;
        RECT 1497.400 2718.340 1497.660 2718.600 ;
        RECT 1497.860 2656.460 1498.120 2656.720 ;
        RECT 1498.780 2656.460 1499.040 2656.720 ;
        RECT 1498.780 2622.120 1499.040 2622.380 ;
        RECT 1499.240 2621.780 1499.500 2622.040 ;
        RECT 1498.320 2559.900 1498.580 2560.160 ;
        RECT 1499.700 2559.900 1499.960 2560.160 ;
        RECT 1498.780 2511.620 1499.040 2511.880 ;
        RECT 1499.700 2511.620 1499.960 2511.880 ;
        RECT 1498.320 2463.000 1498.580 2463.260 ;
        RECT 1498.320 2428.660 1498.580 2428.920 ;
        RECT 1497.860 2380.380 1498.120 2380.640 ;
        RECT 1498.780 2380.380 1499.040 2380.640 ;
        RECT 1498.320 2366.440 1498.580 2366.700 ;
        RECT 1498.320 2331.760 1498.580 2332.020 ;
        RECT 1496.940 2304.220 1497.200 2304.480 ;
        RECT 1498.780 2304.220 1499.040 2304.480 ;
        RECT 1497.400 2249.140 1497.660 2249.400 ;
        RECT 1497.860 2201.200 1498.120 2201.460 ;
        RECT 1497.860 2183.860 1498.120 2184.120 ;
        RECT 1497.860 2138.640 1498.120 2138.900 ;
        RECT 1498.780 2076.760 1499.040 2077.020 ;
        RECT 1498.320 2028.480 1498.580 2028.740 ;
        RECT 1300.980 2009.780 1301.240 2010.040 ;
        RECT 1498.320 2009.780 1498.580 2010.040 ;
      LAYER met2 ;
        RECT 1500.470 3517.600 1501.030 3524.800 ;
        RECT 1500.680 3443.170 1500.820 3517.600 ;
        RECT 1498.320 3442.850 1498.580 3443.170 ;
        RECT 1500.620 3442.850 1500.880 3443.170 ;
        RECT 1498.380 3429.650 1498.520 3442.850 ;
        RECT 1497.920 3429.510 1498.520 3429.650 ;
        RECT 1497.920 3422.430 1498.060 3429.510 ;
        RECT 1497.860 3422.110 1498.120 3422.430 ;
        RECT 1499.700 3332.690 1499.960 3333.010 ;
        RECT 1499.760 3298.410 1499.900 3332.690 ;
        RECT 1498.840 3298.270 1499.900 3298.410 ;
        RECT 1498.840 3236.450 1498.980 3298.270 ;
        RECT 1498.320 3236.130 1498.580 3236.450 ;
        RECT 1498.780 3236.130 1499.040 3236.450 ;
        RECT 1498.380 3202.110 1498.520 3236.130 ;
        RECT 1498.320 3201.790 1498.580 3202.110 ;
        RECT 1498.780 3201.790 1499.040 3202.110 ;
        RECT 1498.840 3153.490 1498.980 3201.790 ;
        RECT 1497.860 3153.170 1498.120 3153.490 ;
        RECT 1498.780 3153.170 1499.040 3153.490 ;
        RECT 1497.920 3152.890 1498.060 3153.170 ;
        RECT 1497.920 3152.750 1498.520 3152.890 ;
        RECT 1498.380 3105.290 1498.520 3152.750 ;
        RECT 1498.380 3105.150 1498.980 3105.290 ;
        RECT 1498.840 3056.930 1498.980 3105.150 ;
        RECT 1497.860 3056.610 1498.120 3056.930 ;
        RECT 1498.780 3056.610 1499.040 3056.930 ;
        RECT 1497.920 3056.330 1498.060 3056.610 ;
        RECT 1497.920 3056.190 1498.520 3056.330 ;
        RECT 1498.380 3042.990 1498.520 3056.190 ;
        RECT 1498.320 3042.670 1498.580 3042.990 ;
        RECT 1499.240 3008.330 1499.500 3008.650 ;
        RECT 1499.300 2994.710 1499.440 3008.330 ;
        RECT 1499.240 2994.390 1499.500 2994.710 ;
        RECT 1499.700 2946.450 1499.960 2946.770 ;
        RECT 1499.760 2912.430 1499.900 2946.450 ;
        RECT 1499.700 2912.110 1499.960 2912.430 ;
        RECT 1499.240 2911.430 1499.500 2911.750 ;
        RECT 1499.300 2863.210 1499.440 2911.430 ;
        RECT 1498.380 2863.070 1499.440 2863.210 ;
        RECT 1498.380 2849.610 1498.520 2863.070 ;
        RECT 1497.920 2849.470 1498.520 2849.610 ;
        RECT 1497.920 2815.870 1498.060 2849.470 ;
        RECT 1497.860 2815.550 1498.120 2815.870 ;
        RECT 1497.860 2814.870 1498.120 2815.190 ;
        RECT 1497.920 2802.805 1498.060 2814.870 ;
        RECT 1497.850 2802.435 1498.130 2802.805 ;
        RECT 1497.850 2801.755 1498.130 2802.125 ;
        RECT 1497.920 2767.590 1498.060 2801.755 ;
        RECT 1497.860 2767.270 1498.120 2767.590 ;
        RECT 1497.400 2766.590 1497.660 2766.910 ;
        RECT 1497.460 2746.365 1497.600 2766.590 ;
        RECT 1496.470 2745.995 1496.750 2746.365 ;
        RECT 1497.390 2745.995 1497.670 2746.365 ;
        RECT 1496.540 2718.630 1496.680 2745.995 ;
        RECT 1496.480 2718.310 1496.740 2718.630 ;
        RECT 1497.400 2718.310 1497.660 2718.630 ;
        RECT 1497.460 2697.970 1497.600 2718.310 ;
        RECT 1497.460 2697.830 1498.060 2697.970 ;
        RECT 1497.920 2656.750 1498.060 2697.830 ;
        RECT 1497.860 2656.430 1498.120 2656.750 ;
        RECT 1498.780 2656.430 1499.040 2656.750 ;
        RECT 1498.840 2622.410 1498.980 2656.430 ;
        RECT 1498.780 2622.090 1499.040 2622.410 ;
        RECT 1499.240 2621.750 1499.500 2622.070 ;
        RECT 1499.300 2608.325 1499.440 2621.750 ;
        RECT 1498.310 2607.955 1498.590 2608.325 ;
        RECT 1499.230 2607.955 1499.510 2608.325 ;
        RECT 1498.380 2560.190 1498.520 2607.955 ;
        RECT 1498.320 2559.870 1498.580 2560.190 ;
        RECT 1499.700 2559.870 1499.960 2560.190 ;
        RECT 1499.760 2511.910 1499.900 2559.870 ;
        RECT 1498.780 2511.765 1499.040 2511.910 ;
        RECT 1497.390 2511.395 1497.670 2511.765 ;
        RECT 1498.770 2511.395 1499.050 2511.765 ;
        RECT 1499.700 2511.590 1499.960 2511.910 ;
        RECT 1497.460 2463.485 1497.600 2511.395 ;
        RECT 1497.390 2463.115 1497.670 2463.485 ;
        RECT 1498.310 2463.115 1498.590 2463.485 ;
        RECT 1498.320 2462.970 1498.580 2463.115 ;
        RECT 1498.320 2428.630 1498.580 2428.950 ;
        RECT 1498.380 2415.090 1498.520 2428.630 ;
        RECT 1498.380 2414.950 1498.980 2415.090 ;
        RECT 1498.840 2380.670 1498.980 2414.950 ;
        RECT 1497.860 2380.410 1498.120 2380.670 ;
        RECT 1497.860 2380.350 1498.520 2380.410 ;
        RECT 1498.780 2380.350 1499.040 2380.670 ;
        RECT 1497.920 2380.270 1498.520 2380.350 ;
        RECT 1498.380 2366.730 1498.520 2380.270 ;
        RECT 1498.320 2366.410 1498.580 2366.730 ;
        RECT 1498.320 2331.730 1498.580 2332.050 ;
        RECT 1498.380 2318.530 1498.520 2331.730 ;
        RECT 1498.380 2318.390 1498.980 2318.530 ;
        RECT 1498.840 2304.510 1498.980 2318.390 ;
        RECT 1496.940 2304.190 1497.200 2304.510 ;
        RECT 1498.780 2304.190 1499.040 2304.510 ;
        RECT 1497.000 2256.650 1497.140 2304.190 ;
        RECT 1497.000 2256.510 1497.600 2256.650 ;
        RECT 1497.460 2249.430 1497.600 2256.510 ;
        RECT 1497.400 2249.110 1497.660 2249.430 ;
        RECT 1497.860 2201.170 1498.120 2201.490 ;
        RECT 1497.920 2184.150 1498.060 2201.170 ;
        RECT 1497.860 2183.830 1498.120 2184.150 ;
        RECT 1497.860 2138.610 1498.120 2138.930 ;
        RECT 1497.920 2090.730 1498.060 2138.610 ;
        RECT 1497.920 2090.590 1498.980 2090.730 ;
        RECT 1498.840 2077.050 1498.980 2090.590 ;
        RECT 1498.780 2076.730 1499.040 2077.050 ;
        RECT 1498.320 2028.450 1498.580 2028.770 ;
        RECT 1498.380 2010.070 1498.520 2028.450 ;
        RECT 1300.980 2009.750 1301.240 2010.070 ;
        RECT 1498.320 2009.750 1498.580 2010.070 ;
        RECT 1301.040 2000.000 1301.180 2009.750 ;
        RECT 1300.880 1999.540 1301.180 2000.000 ;
        RECT 1300.880 1996.000 1301.160 1999.540 ;
      LAYER via2 ;
        RECT 1497.850 2802.480 1498.130 2802.760 ;
        RECT 1497.850 2801.800 1498.130 2802.080 ;
        RECT 1496.470 2746.040 1496.750 2746.320 ;
        RECT 1497.390 2746.040 1497.670 2746.320 ;
        RECT 1498.310 2608.000 1498.590 2608.280 ;
        RECT 1499.230 2608.000 1499.510 2608.280 ;
        RECT 1497.390 2511.440 1497.670 2511.720 ;
        RECT 1498.770 2511.440 1499.050 2511.720 ;
        RECT 1497.390 2463.160 1497.670 2463.440 ;
        RECT 1498.310 2463.160 1498.590 2463.440 ;
      LAYER met3 ;
        RECT 1497.825 2802.770 1498.155 2802.785 ;
        RECT 1497.150 2802.470 1498.155 2802.770 ;
        RECT 1497.150 2802.090 1497.450 2802.470 ;
        RECT 1497.825 2802.455 1498.155 2802.470 ;
        RECT 1497.825 2802.090 1498.155 2802.105 ;
        RECT 1497.150 2801.790 1498.155 2802.090 ;
        RECT 1497.825 2801.775 1498.155 2801.790 ;
        RECT 1496.445 2746.330 1496.775 2746.345 ;
        RECT 1497.365 2746.330 1497.695 2746.345 ;
        RECT 1496.445 2746.030 1497.695 2746.330 ;
        RECT 1496.445 2746.015 1496.775 2746.030 ;
        RECT 1497.365 2746.015 1497.695 2746.030 ;
        RECT 1498.285 2608.290 1498.615 2608.305 ;
        RECT 1499.205 2608.290 1499.535 2608.305 ;
        RECT 1498.285 2607.990 1499.535 2608.290 ;
        RECT 1498.285 2607.975 1498.615 2607.990 ;
        RECT 1499.205 2607.975 1499.535 2607.990 ;
        RECT 1497.365 2511.730 1497.695 2511.745 ;
        RECT 1498.745 2511.730 1499.075 2511.745 ;
        RECT 1497.365 2511.430 1499.075 2511.730 ;
        RECT 1497.365 2511.415 1497.695 2511.430 ;
        RECT 1498.745 2511.415 1499.075 2511.430 ;
        RECT 1497.365 2463.450 1497.695 2463.465 ;
        RECT 1498.285 2463.450 1498.615 2463.465 ;
        RECT 1497.365 2463.150 1498.615 2463.450 ;
        RECT 1497.365 2463.135 1497.695 2463.150 ;
        RECT 1498.285 2463.135 1498.615 2463.150 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1158.810 2004.200 1159.130 2004.260 ;
        RECT 1472.990 2004.200 1473.310 2004.260 ;
        RECT 1158.810 2004.060 1473.310 2004.200 ;
        RECT 1158.810 2004.000 1159.130 2004.060 ;
        RECT 1472.990 2004.000 1473.310 2004.060 ;
        RECT 1472.990 324.260 1473.310 324.320 ;
        RECT 2898.990 324.260 2899.310 324.320 ;
        RECT 1472.990 324.120 2899.310 324.260 ;
        RECT 1472.990 324.060 1473.310 324.120 ;
        RECT 2898.990 324.060 2899.310 324.120 ;
      LAYER via ;
        RECT 1158.840 2004.000 1159.100 2004.260 ;
        RECT 1473.020 2004.000 1473.280 2004.260 ;
        RECT 1473.020 324.060 1473.280 324.320 ;
        RECT 2899.020 324.060 2899.280 324.320 ;
      LAYER met2 ;
        RECT 1158.840 2003.970 1159.100 2004.290 ;
        RECT 1473.020 2003.970 1473.280 2004.290 ;
        RECT 1158.900 2000.000 1159.040 2003.970 ;
        RECT 1158.740 1999.540 1159.040 2000.000 ;
        RECT 1158.740 1996.000 1159.020 1999.540 ;
        RECT 1473.080 324.350 1473.220 2003.970 ;
        RECT 1473.020 324.030 1473.280 324.350 ;
        RECT 2899.020 324.030 2899.280 324.350 ;
        RECT 2899.080 322.845 2899.220 324.030 ;
        RECT 2899.010 322.475 2899.290 322.845 ;
      LAYER via2 ;
        RECT 2899.010 322.520 2899.290 322.800 ;
      LAYER met3 ;
        RECT 2898.985 322.810 2899.315 322.825 ;
        RECT 2917.600 322.810 2924.800 323.260 ;
        RECT 2898.985 322.510 2924.800 322.810 ;
        RECT 2898.985 322.495 2899.315 322.510 ;
        RECT 2917.600 322.060 2924.800 322.510 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1175.830 3498.500 1176.150 3498.560 ;
        RECT 1179.510 3498.500 1179.830 3498.560 ;
        RECT 1175.830 3498.360 1179.830 3498.500 ;
        RECT 1175.830 3498.300 1176.150 3498.360 ;
        RECT 1179.510 3498.300 1179.830 3498.360 ;
        RECT 1308.770 2010.660 1309.090 2010.720 ;
        RECT 1297.820 2010.520 1309.090 2010.660 ;
        RECT 1297.820 2009.980 1297.960 2010.520 ;
        RECT 1308.770 2010.460 1309.090 2010.520 ;
        RECT 1269.760 2009.840 1297.960 2009.980 ;
        RECT 1179.510 2009.640 1179.830 2009.700 ;
        RECT 1269.760 2009.640 1269.900 2009.840 ;
        RECT 1179.510 2009.500 1269.900 2009.640 ;
        RECT 1179.510 2009.440 1179.830 2009.500 ;
      LAYER via ;
        RECT 1175.860 3498.300 1176.120 3498.560 ;
        RECT 1179.540 3498.300 1179.800 3498.560 ;
        RECT 1308.800 2010.460 1309.060 2010.720 ;
        RECT 1179.540 2009.440 1179.800 2009.700 ;
      LAYER met2 ;
        RECT 1175.710 3517.600 1176.270 3524.800 ;
        RECT 1175.920 3498.590 1176.060 3517.600 ;
        RECT 1175.860 3498.270 1176.120 3498.590 ;
        RECT 1179.540 3498.270 1179.800 3498.590 ;
        RECT 1179.600 2009.730 1179.740 3498.270 ;
        RECT 1308.800 2010.430 1309.060 2010.750 ;
        RECT 1179.540 2009.410 1179.800 2009.730 ;
        RECT 1308.860 2000.000 1309.000 2010.430 ;
        RECT 1308.700 1999.540 1309.000 2000.000 ;
        RECT 1308.700 1996.000 1308.980 1999.540 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1269.745 2007.785 1269.915 2010.675 ;
      LAYER mcon ;
        RECT 1269.745 2010.505 1269.915 2010.675 ;
      LAYER met1 ;
        RECT 851.530 3498.500 851.850 3498.560 ;
        RECT 855.210 3498.500 855.530 3498.560 ;
        RECT 851.530 3498.360 855.530 3498.500 ;
        RECT 851.530 3498.300 851.850 3498.360 ;
        RECT 855.210 3498.300 855.530 3498.360 ;
        RECT 855.210 2010.660 855.530 2010.720 ;
        RECT 1269.685 2010.660 1269.975 2010.705 ;
        RECT 855.210 2010.520 1269.975 2010.660 ;
        RECT 855.210 2010.460 855.530 2010.520 ;
        RECT 1269.685 2010.475 1269.975 2010.520 ;
        RECT 1269.685 2007.940 1269.975 2007.985 ;
        RECT 1314.750 2007.940 1315.070 2008.000 ;
        RECT 1269.685 2007.800 1315.070 2007.940 ;
        RECT 1269.685 2007.755 1269.975 2007.800 ;
        RECT 1314.750 2007.740 1315.070 2007.800 ;
      LAYER via ;
        RECT 851.560 3498.300 851.820 3498.560 ;
        RECT 855.240 3498.300 855.500 3498.560 ;
        RECT 855.240 2010.460 855.500 2010.720 ;
        RECT 1314.780 2007.740 1315.040 2008.000 ;
      LAYER met2 ;
        RECT 851.410 3517.600 851.970 3524.800 ;
        RECT 851.620 3498.590 851.760 3517.600 ;
        RECT 851.560 3498.270 851.820 3498.590 ;
        RECT 855.240 3498.270 855.500 3498.590 ;
        RECT 855.300 2010.750 855.440 3498.270 ;
        RECT 855.240 2010.430 855.500 2010.750 ;
        RECT 1314.780 2007.710 1315.040 2008.030 ;
        RECT 1314.840 1999.610 1314.980 2007.710 ;
        RECT 1316.520 1999.610 1316.800 2000.000 ;
        RECT 1314.840 1999.470 1316.800 1999.610 ;
        RECT 1316.520 1996.000 1316.800 1999.470 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 772.945 2014.585 773.115 2015.435 ;
        RECT 820.785 2014.585 820.955 2015.435 ;
        RECT 1255.945 2014.585 1256.115 2015.775 ;
        RECT 1303.785 2014.925 1303.955 2015.775 ;
      LAYER mcon ;
        RECT 1255.945 2015.605 1256.115 2015.775 ;
        RECT 772.945 2015.265 773.115 2015.435 ;
        RECT 820.785 2015.265 820.955 2015.435 ;
        RECT 1303.785 2015.605 1303.955 2015.775 ;
      LAYER met1 ;
        RECT 527.230 3498.500 527.550 3498.560 ;
        RECT 530.910 3498.500 531.230 3498.560 ;
        RECT 527.230 3498.360 531.230 3498.500 ;
        RECT 527.230 3498.300 527.550 3498.360 ;
        RECT 530.910 3498.300 531.230 3498.360 ;
        RECT 530.910 2015.760 531.230 2015.820 ;
        RECT 530.540 2015.620 531.230 2015.760 ;
        RECT 530.540 2015.080 530.680 2015.620 ;
        RECT 530.910 2015.560 531.230 2015.620 ;
        RECT 1255.885 2015.760 1256.175 2015.805 ;
        RECT 1303.725 2015.760 1304.015 2015.805 ;
        RECT 1255.885 2015.620 1304.015 2015.760 ;
        RECT 1255.885 2015.575 1256.175 2015.620 ;
        RECT 1303.725 2015.575 1304.015 2015.620 ;
        RECT 772.885 2015.420 773.175 2015.465 ;
        RECT 820.725 2015.420 821.015 2015.465 ;
        RECT 772.885 2015.280 821.015 2015.420 ;
        RECT 772.885 2015.235 773.175 2015.280 ;
        RECT 820.725 2015.235 821.015 2015.280 ;
        RECT 1303.725 2015.080 1304.015 2015.125 ;
        RECT 1324.410 2015.080 1324.730 2015.140 ;
        RECT 530.540 2014.940 531.140 2015.080 ;
        RECT 531.000 2014.740 531.140 2014.940 ;
        RECT 1303.725 2014.940 1324.730 2015.080 ;
        RECT 1303.725 2014.895 1304.015 2014.940 ;
        RECT 1324.410 2014.880 1324.730 2014.940 ;
        RECT 772.885 2014.740 773.175 2014.785 ;
        RECT 531.000 2014.600 773.175 2014.740 ;
        RECT 772.885 2014.555 773.175 2014.600 ;
        RECT 820.725 2014.740 821.015 2014.785 ;
        RECT 1255.885 2014.740 1256.175 2014.785 ;
        RECT 820.725 2014.600 1256.175 2014.740 ;
        RECT 820.725 2014.555 821.015 2014.600 ;
        RECT 1255.885 2014.555 1256.175 2014.600 ;
      LAYER via ;
        RECT 527.260 3498.300 527.520 3498.560 ;
        RECT 530.940 3498.300 531.200 3498.560 ;
        RECT 530.940 2015.560 531.200 2015.820 ;
        RECT 1324.440 2014.880 1324.700 2015.140 ;
      LAYER met2 ;
        RECT 527.110 3517.600 527.670 3524.800 ;
        RECT 527.320 3498.590 527.460 3517.600 ;
        RECT 527.260 3498.270 527.520 3498.590 ;
        RECT 530.940 3498.270 531.200 3498.590 ;
        RECT 531.000 2015.850 531.140 3498.270 ;
        RECT 530.940 2015.530 531.200 2015.850 ;
        RECT 1324.440 2014.850 1324.700 2015.170 ;
        RECT 1324.500 2000.000 1324.640 2014.850 ;
        RECT 1324.340 1999.540 1324.640 2000.000 ;
        RECT 1324.340 1996.000 1324.620 1999.540 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 529.605 2013.905 530.235 2014.075 ;
        RECT 1273.885 2012.885 1274.055 2014.075 ;
      LAYER mcon ;
        RECT 530.065 2013.905 530.235 2014.075 ;
        RECT 1273.885 2013.905 1274.055 2014.075 ;
      LAYER met1 ;
        RECT 202.470 3501.900 202.790 3501.960 ;
        RECT 206.610 3501.900 206.930 3501.960 ;
        RECT 202.470 3501.760 206.930 3501.900 ;
        RECT 202.470 3501.700 202.790 3501.760 ;
        RECT 206.610 3501.700 206.930 3501.760 ;
        RECT 206.610 2014.060 206.930 2014.120 ;
        RECT 529.545 2014.060 529.835 2014.105 ;
        RECT 206.610 2013.920 529.835 2014.060 ;
        RECT 206.610 2013.860 206.930 2013.920 ;
        RECT 529.545 2013.875 529.835 2013.920 ;
        RECT 530.005 2014.060 530.295 2014.105 ;
        RECT 1273.825 2014.060 1274.115 2014.105 ;
        RECT 530.005 2013.920 1274.115 2014.060 ;
        RECT 530.005 2013.875 530.295 2013.920 ;
        RECT 1273.825 2013.875 1274.115 2013.920 ;
        RECT 1273.825 2013.040 1274.115 2013.085 ;
        RECT 1332.230 2013.040 1332.550 2013.100 ;
        RECT 1273.825 2012.900 1332.550 2013.040 ;
        RECT 1273.825 2012.855 1274.115 2012.900 ;
        RECT 1332.230 2012.840 1332.550 2012.900 ;
      LAYER via ;
        RECT 202.500 3501.700 202.760 3501.960 ;
        RECT 206.640 3501.700 206.900 3501.960 ;
        RECT 206.640 2013.860 206.900 2014.120 ;
        RECT 1332.260 2012.840 1332.520 2013.100 ;
      LAYER met2 ;
        RECT 202.350 3517.600 202.910 3524.800 ;
        RECT 202.560 3501.990 202.700 3517.600 ;
        RECT 202.500 3501.670 202.760 3501.990 ;
        RECT 206.640 3501.670 206.900 3501.990 ;
        RECT 206.700 2014.150 206.840 3501.670 ;
        RECT 206.640 2013.830 206.900 2014.150 ;
        RECT 1332.260 2012.810 1332.520 2013.130 ;
        RECT 1332.320 2000.000 1332.460 2012.810 ;
        RECT 1332.160 1999.540 1332.460 2000.000 ;
        RECT 1332.160 1996.000 1332.440 1999.540 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1279.865 2013.225 1280.035 2014.755 ;
        RECT 1306.545 2013.225 1306.715 2014.755 ;
      LAYER mcon ;
        RECT 1279.865 2014.585 1280.035 2014.755 ;
        RECT 1306.545 2014.585 1306.715 2014.755 ;
      LAYER met1 ;
        RECT 1279.805 2014.740 1280.095 2014.785 ;
        RECT 1306.485 2014.740 1306.775 2014.785 ;
        RECT 1279.805 2014.600 1306.775 2014.740 ;
        RECT 1279.805 2014.555 1280.095 2014.600 ;
        RECT 1306.485 2014.555 1306.775 2014.600 ;
        RECT 17.090 2013.380 17.410 2013.440 ;
        RECT 1279.805 2013.380 1280.095 2013.425 ;
        RECT 17.090 2013.240 1280.095 2013.380 ;
        RECT 17.090 2013.180 17.410 2013.240 ;
        RECT 1279.805 2013.195 1280.095 2013.240 ;
        RECT 1306.485 2013.380 1306.775 2013.425 ;
        RECT 1340.050 2013.380 1340.370 2013.440 ;
        RECT 1306.485 2013.240 1340.370 2013.380 ;
        RECT 1306.485 2013.195 1306.775 2013.240 ;
        RECT 1340.050 2013.180 1340.370 2013.240 ;
      LAYER via ;
        RECT 17.120 2013.180 17.380 2013.440 ;
        RECT 1340.080 2013.180 1340.340 2013.440 ;
      LAYER met2 ;
        RECT 17.110 3411.035 17.390 3411.405 ;
        RECT 17.180 2013.470 17.320 3411.035 ;
        RECT 17.120 2013.150 17.380 2013.470 ;
        RECT 1340.080 2013.150 1340.340 2013.470 ;
        RECT 1340.140 2000.000 1340.280 2013.150 ;
        RECT 1339.980 1999.540 1340.280 2000.000 ;
        RECT 1339.980 1996.000 1340.260 1999.540 ;
      LAYER via2 ;
        RECT 17.110 3411.080 17.390 3411.360 ;
      LAYER met3 ;
        RECT -4.800 3411.370 2.400 3411.820 ;
        RECT 17.085 3411.370 17.415 3411.385 ;
        RECT -4.800 3411.070 17.415 3411.370 ;
        RECT -4.800 3410.620 2.400 3411.070 ;
        RECT 17.085 3411.055 17.415 3411.070 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1271.125 2010.505 1271.295 2013.055 ;
      LAYER mcon ;
        RECT 1271.125 2012.885 1271.295 2013.055 ;
      LAYER met1 ;
        RECT 18.010 2013.040 18.330 2013.100 ;
        RECT 1271.065 2013.040 1271.355 2013.085 ;
        RECT 18.010 2012.900 1271.355 2013.040 ;
        RECT 18.010 2012.840 18.330 2012.900 ;
        RECT 1271.065 2012.855 1271.355 2012.900 ;
        RECT 1347.870 2011.000 1348.190 2011.060 ;
        RECT 1297.360 2010.860 1348.190 2011.000 ;
        RECT 1271.065 2010.660 1271.355 2010.705 ;
        RECT 1297.360 2010.660 1297.500 2010.860 ;
        RECT 1347.870 2010.800 1348.190 2010.860 ;
        RECT 1271.065 2010.520 1297.500 2010.660 ;
        RECT 1271.065 2010.475 1271.355 2010.520 ;
      LAYER via ;
        RECT 18.040 2012.840 18.300 2013.100 ;
        RECT 1347.900 2010.800 1348.160 2011.060 ;
      LAYER met2 ;
        RECT 18.030 3124.075 18.310 3124.445 ;
        RECT 18.100 2013.130 18.240 3124.075 ;
        RECT 18.040 2012.810 18.300 2013.130 ;
        RECT 1347.900 2010.770 1348.160 2011.090 ;
        RECT 1347.960 2000.000 1348.100 2010.770 ;
        RECT 1347.800 1999.540 1348.100 2000.000 ;
        RECT 1347.800 1996.000 1348.080 1999.540 ;
      LAYER via2 ;
        RECT 18.030 3124.120 18.310 3124.400 ;
      LAYER met3 ;
        RECT -4.800 3124.410 2.400 3124.860 ;
        RECT 18.005 3124.410 18.335 3124.425 ;
        RECT -4.800 3124.110 18.335 3124.410 ;
        RECT -4.800 3123.660 2.400 3124.110 ;
        RECT 18.005 3124.095 18.335 3124.110 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 19.390 2012.360 19.710 2012.420 ;
        RECT 1356.150 2012.360 1356.470 2012.420 ;
        RECT 19.390 2012.220 1356.470 2012.360 ;
        RECT 19.390 2012.160 19.710 2012.220 ;
        RECT 1356.150 2012.160 1356.470 2012.220 ;
      LAYER via ;
        RECT 19.420 2012.160 19.680 2012.420 ;
        RECT 1356.180 2012.160 1356.440 2012.420 ;
      LAYER met2 ;
        RECT 19.410 2836.435 19.690 2836.805 ;
        RECT 19.480 2012.450 19.620 2836.435 ;
        RECT 19.420 2012.130 19.680 2012.450 ;
        RECT 1356.180 2012.130 1356.440 2012.450 ;
        RECT 1356.240 2000.000 1356.380 2012.130 ;
        RECT 1356.080 1999.540 1356.380 2000.000 ;
        RECT 1356.080 1996.000 1356.360 1999.540 ;
      LAYER via2 ;
        RECT 19.410 2836.480 19.690 2836.760 ;
      LAYER met3 ;
        RECT -4.800 2836.770 2.400 2837.220 ;
        RECT 19.385 2836.770 19.715 2836.785 ;
        RECT -4.800 2836.470 19.715 2836.770 ;
        RECT -4.800 2836.020 2.400 2836.470 ;
        RECT 19.385 2836.455 19.715 2836.470 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 20.310 2011.680 20.630 2011.740 ;
        RECT 1363.970 2011.680 1364.290 2011.740 ;
        RECT 20.310 2011.540 1364.290 2011.680 ;
        RECT 20.310 2011.480 20.630 2011.540 ;
        RECT 1363.970 2011.480 1364.290 2011.540 ;
      LAYER via ;
        RECT 20.340 2011.480 20.600 2011.740 ;
        RECT 1364.000 2011.480 1364.260 2011.740 ;
      LAYER met2 ;
        RECT 20.330 2549.475 20.610 2549.845 ;
        RECT 20.400 2011.770 20.540 2549.475 ;
        RECT 20.340 2011.450 20.600 2011.770 ;
        RECT 1364.000 2011.450 1364.260 2011.770 ;
        RECT 1364.060 2000.000 1364.200 2011.450 ;
        RECT 1363.900 1999.540 1364.200 2000.000 ;
        RECT 1363.900 1996.000 1364.180 1999.540 ;
      LAYER via2 ;
        RECT 20.330 2549.520 20.610 2549.800 ;
      LAYER met3 ;
        RECT -4.800 2549.810 2.400 2550.260 ;
        RECT 20.305 2549.810 20.635 2549.825 ;
        RECT -4.800 2549.510 20.635 2549.810 ;
        RECT -4.800 2549.060 2.400 2549.510 ;
        RECT 20.305 2549.495 20.635 2549.510 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 16.170 2011.340 16.490 2011.400 ;
        RECT 1371.790 2011.340 1372.110 2011.400 ;
        RECT 16.170 2011.200 1372.110 2011.340 ;
        RECT 16.170 2011.140 16.490 2011.200 ;
        RECT 1371.790 2011.140 1372.110 2011.200 ;
      LAYER via ;
        RECT 16.200 2011.140 16.460 2011.400 ;
        RECT 1371.820 2011.140 1372.080 2011.400 ;
      LAYER met2 ;
        RECT 16.190 2261.835 16.470 2262.205 ;
        RECT 16.260 2011.430 16.400 2261.835 ;
        RECT 16.200 2011.110 16.460 2011.430 ;
        RECT 1371.820 2011.110 1372.080 2011.430 ;
        RECT 1371.880 2000.000 1372.020 2011.110 ;
        RECT 1371.720 1999.540 1372.020 2000.000 ;
        RECT 1371.720 1996.000 1372.000 1999.540 ;
      LAYER via2 ;
        RECT 16.190 2261.880 16.470 2262.160 ;
      LAYER met3 ;
        RECT -4.800 2262.170 2.400 2262.620 ;
        RECT 16.165 2262.170 16.495 2262.185 ;
        RECT -4.800 2261.870 16.495 2262.170 ;
        RECT -4.800 2261.420 2.400 2261.870 ;
        RECT 16.165 2261.855 16.495 2261.870 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 54.810 2007.260 55.130 2007.320 ;
        RECT 1379.610 2007.260 1379.930 2007.320 ;
        RECT 54.810 2007.120 1379.930 2007.260 ;
        RECT 54.810 2007.060 55.130 2007.120 ;
        RECT 1379.610 2007.060 1379.930 2007.120 ;
        RECT 15.710 1980.060 16.030 1980.120 ;
        RECT 54.810 1980.060 55.130 1980.120 ;
        RECT 15.710 1979.920 55.130 1980.060 ;
        RECT 15.710 1979.860 16.030 1979.920 ;
        RECT 54.810 1979.860 55.130 1979.920 ;
      LAYER via ;
        RECT 54.840 2007.060 55.100 2007.320 ;
        RECT 1379.640 2007.060 1379.900 2007.320 ;
        RECT 15.740 1979.860 16.000 1980.120 ;
        RECT 54.840 1979.860 55.100 1980.120 ;
      LAYER met2 ;
        RECT 54.840 2007.030 55.100 2007.350 ;
        RECT 1379.640 2007.030 1379.900 2007.350 ;
        RECT 54.900 1980.150 55.040 2007.030 ;
        RECT 1379.700 2000.000 1379.840 2007.030 ;
        RECT 1379.540 1999.540 1379.840 2000.000 ;
        RECT 1379.540 1996.000 1379.820 1999.540 ;
        RECT 15.740 1979.830 16.000 1980.150 ;
        RECT 54.840 1979.830 55.100 1980.150 ;
        RECT 15.800 1975.245 15.940 1979.830 ;
        RECT 15.730 1974.875 16.010 1975.245 ;
      LAYER via2 ;
        RECT 15.730 1974.920 16.010 1975.200 ;
      LAYER met3 ;
        RECT -4.800 1975.210 2.400 1975.660 ;
        RECT 15.705 1975.210 16.035 1975.225 ;
        RECT -4.800 1974.910 16.035 1975.210 ;
        RECT -4.800 1974.460 2.400 1974.910 ;
        RECT 15.705 1974.895 16.035 1974.910 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1166.630 2005.560 1166.950 2005.620 ;
        RECT 1459.650 2005.560 1459.970 2005.620 ;
        RECT 1166.630 2005.420 1459.970 2005.560 ;
        RECT 1166.630 2005.360 1166.950 2005.420 ;
        RECT 1459.650 2005.360 1459.970 2005.420 ;
        RECT 1459.650 558.860 1459.970 558.920 ;
        RECT 2898.990 558.860 2899.310 558.920 ;
        RECT 1459.650 558.720 2899.310 558.860 ;
        RECT 1459.650 558.660 1459.970 558.720 ;
        RECT 2898.990 558.660 2899.310 558.720 ;
      LAYER via ;
        RECT 1166.660 2005.360 1166.920 2005.620 ;
        RECT 1459.680 2005.360 1459.940 2005.620 ;
        RECT 1459.680 558.660 1459.940 558.920 ;
        RECT 2899.020 558.660 2899.280 558.920 ;
      LAYER met2 ;
        RECT 1166.660 2005.330 1166.920 2005.650 ;
        RECT 1459.680 2005.330 1459.940 2005.650 ;
        RECT 1166.720 2000.000 1166.860 2005.330 ;
        RECT 1166.560 1999.540 1166.860 2000.000 ;
        RECT 1166.560 1996.000 1166.840 1999.540 ;
        RECT 1459.740 558.950 1459.880 2005.330 ;
        RECT 1459.680 558.630 1459.940 558.950 ;
        RECT 2899.020 558.630 2899.280 558.950 ;
        RECT 2899.080 557.445 2899.220 558.630 ;
        RECT 2899.010 557.075 2899.290 557.445 ;
      LAYER via2 ;
        RECT 2899.010 557.120 2899.290 557.400 ;
      LAYER met3 ;
        RECT 2898.985 557.410 2899.315 557.425 ;
        RECT 2917.600 557.410 2924.800 557.860 ;
        RECT 2898.985 557.110 2924.800 557.410 ;
        RECT 2898.985 557.095 2899.315 557.110 ;
        RECT 2917.600 556.660 2924.800 557.110 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 72.750 2006.920 73.070 2006.980 ;
        RECT 1387.430 2006.920 1387.750 2006.980 ;
        RECT 72.750 2006.780 1387.750 2006.920 ;
        RECT 72.750 2006.720 73.070 2006.780 ;
        RECT 1387.430 2006.720 1387.750 2006.780 ;
        RECT 17.090 1690.380 17.410 1690.440 ;
        RECT 72.750 1690.380 73.070 1690.440 ;
        RECT 17.090 1690.240 73.070 1690.380 ;
        RECT 17.090 1690.180 17.410 1690.240 ;
        RECT 72.750 1690.180 73.070 1690.240 ;
      LAYER via ;
        RECT 72.780 2006.720 73.040 2006.980 ;
        RECT 1387.460 2006.720 1387.720 2006.980 ;
        RECT 17.120 1690.180 17.380 1690.440 ;
        RECT 72.780 1690.180 73.040 1690.440 ;
      LAYER met2 ;
        RECT 72.780 2006.690 73.040 2007.010 ;
        RECT 1387.460 2006.690 1387.720 2007.010 ;
        RECT 72.840 1690.470 72.980 2006.690 ;
        RECT 1387.520 2000.000 1387.660 2006.690 ;
        RECT 1387.360 1999.540 1387.660 2000.000 ;
        RECT 1387.360 1996.000 1387.640 1999.540 ;
        RECT 17.120 1690.150 17.380 1690.470 ;
        RECT 72.780 1690.150 73.040 1690.470 ;
        RECT 17.180 1687.605 17.320 1690.150 ;
        RECT 17.110 1687.235 17.390 1687.605 ;
      LAYER via2 ;
        RECT 17.110 1687.280 17.390 1687.560 ;
      LAYER met3 ;
        RECT -4.800 1687.570 2.400 1688.020 ;
        RECT 17.085 1687.570 17.415 1687.585 ;
        RECT -4.800 1687.270 17.415 1687.570 ;
        RECT -4.800 1686.820 2.400 1687.270 ;
        RECT 17.085 1687.255 17.415 1687.270 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1135.810 2006.580 1136.130 2006.640 ;
        RECT 1395.250 2006.580 1395.570 2006.640 ;
        RECT 1135.810 2006.440 1395.570 2006.580 ;
        RECT 1135.810 2006.380 1136.130 2006.440 ;
        RECT 1395.250 2006.380 1395.570 2006.440 ;
        RECT 17.550 1476.520 17.870 1476.580 ;
        RECT 1135.810 1476.520 1136.130 1476.580 ;
        RECT 17.550 1476.380 1136.130 1476.520 ;
        RECT 17.550 1476.320 17.870 1476.380 ;
        RECT 1135.810 1476.320 1136.130 1476.380 ;
      LAYER via ;
        RECT 1135.840 2006.380 1136.100 2006.640 ;
        RECT 1395.280 2006.380 1395.540 2006.640 ;
        RECT 17.580 1476.320 17.840 1476.580 ;
        RECT 1135.840 1476.320 1136.100 1476.580 ;
      LAYER met2 ;
        RECT 1135.840 2006.350 1136.100 2006.670 ;
        RECT 1395.280 2006.350 1395.540 2006.670 ;
        RECT 1135.900 1476.610 1136.040 2006.350 ;
        RECT 1395.340 2000.000 1395.480 2006.350 ;
        RECT 1395.180 1999.540 1395.480 2000.000 ;
        RECT 1395.180 1996.000 1395.460 1999.540 ;
        RECT 17.580 1476.290 17.840 1476.610 ;
        RECT 1135.840 1476.290 1136.100 1476.610 ;
        RECT 17.640 1472.045 17.780 1476.290 ;
        RECT 17.570 1471.675 17.850 1472.045 ;
      LAYER via2 ;
        RECT 17.570 1471.720 17.850 1472.000 ;
      LAYER met3 ;
        RECT -4.800 1472.010 2.400 1472.460 ;
        RECT 17.545 1472.010 17.875 1472.025 ;
        RECT -4.800 1471.710 17.875 1472.010 ;
        RECT -4.800 1471.260 2.400 1471.710 ;
        RECT 17.545 1471.695 17.875 1471.710 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1128.910 2006.240 1129.230 2006.300 ;
        RECT 1403.530 2006.240 1403.850 2006.300 ;
        RECT 1128.910 2006.100 1403.850 2006.240 ;
        RECT 1128.910 2006.040 1129.230 2006.100 ;
        RECT 1403.530 2006.040 1403.850 2006.100 ;
        RECT 15.710 1262.660 16.030 1262.720 ;
        RECT 1128.910 1262.660 1129.230 1262.720 ;
        RECT 15.710 1262.520 1129.230 1262.660 ;
        RECT 15.710 1262.460 16.030 1262.520 ;
        RECT 1128.910 1262.460 1129.230 1262.520 ;
      LAYER via ;
        RECT 1128.940 2006.040 1129.200 2006.300 ;
        RECT 1403.560 2006.040 1403.820 2006.300 ;
        RECT 15.740 1262.460 16.000 1262.720 ;
        RECT 1128.940 1262.460 1129.200 1262.720 ;
      LAYER met2 ;
        RECT 1128.940 2006.010 1129.200 2006.330 ;
        RECT 1403.560 2006.010 1403.820 2006.330 ;
        RECT 1129.000 1262.750 1129.140 2006.010 ;
        RECT 1403.620 2000.000 1403.760 2006.010 ;
        RECT 1403.460 1999.540 1403.760 2000.000 ;
        RECT 1403.460 1996.000 1403.740 1999.540 ;
        RECT 15.740 1262.430 16.000 1262.750 ;
        RECT 1128.940 1262.430 1129.200 1262.750 ;
        RECT 15.800 1256.485 15.940 1262.430 ;
        RECT 15.730 1256.115 16.010 1256.485 ;
      LAYER via2 ;
        RECT 15.730 1256.160 16.010 1256.440 ;
      LAYER met3 ;
        RECT -4.800 1256.450 2.400 1256.900 ;
        RECT 15.705 1256.450 16.035 1256.465 ;
        RECT -4.800 1256.150 16.035 1256.450 ;
        RECT -4.800 1255.700 2.400 1256.150 ;
        RECT 15.705 1256.135 16.035 1256.150 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 900.290 1996.720 900.610 1996.780 ;
        RECT 1409.510 1996.720 1409.830 1996.780 ;
        RECT 900.290 1996.580 1409.830 1996.720 ;
        RECT 900.290 1996.520 900.610 1996.580 ;
        RECT 1409.510 1996.520 1409.830 1996.580 ;
        RECT 17.550 1041.660 17.870 1041.720 ;
        RECT 900.290 1041.660 900.610 1041.720 ;
        RECT 17.550 1041.520 900.610 1041.660 ;
        RECT 17.550 1041.460 17.870 1041.520 ;
        RECT 900.290 1041.460 900.610 1041.520 ;
      LAYER via ;
        RECT 900.320 1996.520 900.580 1996.780 ;
        RECT 1409.540 1996.520 1409.800 1996.780 ;
        RECT 17.580 1041.460 17.840 1041.720 ;
        RECT 900.320 1041.460 900.580 1041.720 ;
      LAYER met2 ;
        RECT 1411.280 1996.890 1411.560 2000.000 ;
        RECT 1409.600 1996.810 1411.560 1996.890 ;
        RECT 900.320 1996.490 900.580 1996.810 ;
        RECT 1409.540 1996.750 1411.560 1996.810 ;
        RECT 1409.540 1996.490 1409.800 1996.750 ;
        RECT 900.380 1041.750 900.520 1996.490 ;
        RECT 1411.280 1996.000 1411.560 1996.750 ;
        RECT 17.580 1041.430 17.840 1041.750 ;
        RECT 900.320 1041.430 900.580 1041.750 ;
        RECT 17.640 1040.925 17.780 1041.430 ;
        RECT 17.570 1040.555 17.850 1040.925 ;
      LAYER via2 ;
        RECT 17.570 1040.600 17.850 1040.880 ;
      LAYER met3 ;
        RECT -4.800 1040.890 2.400 1041.340 ;
        RECT 17.545 1040.890 17.875 1040.905 ;
        RECT -4.800 1040.590 17.875 1040.890 ;
        RECT -4.800 1040.140 2.400 1040.590 ;
        RECT 17.545 1040.575 17.875 1040.590 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1114.190 2005.220 1114.510 2005.280 ;
        RECT 1419.170 2005.220 1419.490 2005.280 ;
        RECT 1114.190 2005.080 1419.490 2005.220 ;
        RECT 1114.190 2005.020 1114.510 2005.080 ;
        RECT 1419.170 2005.020 1419.490 2005.080 ;
        RECT 17.550 827.800 17.870 827.860 ;
        RECT 1114.190 827.800 1114.510 827.860 ;
        RECT 17.550 827.660 1114.510 827.800 ;
        RECT 17.550 827.600 17.870 827.660 ;
        RECT 1114.190 827.600 1114.510 827.660 ;
      LAYER via ;
        RECT 1114.220 2005.020 1114.480 2005.280 ;
        RECT 1419.200 2005.020 1419.460 2005.280 ;
        RECT 17.580 827.600 17.840 827.860 ;
        RECT 1114.220 827.600 1114.480 827.860 ;
      LAYER met2 ;
        RECT 1114.220 2004.990 1114.480 2005.310 ;
        RECT 1419.200 2004.990 1419.460 2005.310 ;
        RECT 1114.280 827.890 1114.420 2004.990 ;
        RECT 1419.260 2000.000 1419.400 2004.990 ;
        RECT 1419.100 1999.540 1419.400 2000.000 ;
        RECT 1419.100 1996.000 1419.380 1999.540 ;
        RECT 17.580 827.570 17.840 827.890 ;
        RECT 1114.220 827.570 1114.480 827.890 ;
        RECT 17.640 825.365 17.780 827.570 ;
        RECT 17.570 824.995 17.850 825.365 ;
      LAYER via2 ;
        RECT 17.570 825.040 17.850 825.320 ;
      LAYER met3 ;
        RECT -4.800 825.330 2.400 825.780 ;
        RECT 17.545 825.330 17.875 825.345 ;
        RECT -4.800 825.030 17.875 825.330 ;
        RECT -4.800 824.580 2.400 825.030 ;
        RECT 17.545 825.015 17.875 825.030 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1093.490 1998.760 1093.810 1998.820 ;
        RECT 1425.150 1998.760 1425.470 1998.820 ;
        RECT 1093.490 1998.620 1425.470 1998.760 ;
        RECT 1093.490 1998.560 1093.810 1998.620 ;
        RECT 1425.150 1998.560 1425.470 1998.620 ;
        RECT 14.790 613.940 15.110 614.000 ;
        RECT 1093.490 613.940 1093.810 614.000 ;
        RECT 14.790 613.800 1093.810 613.940 ;
        RECT 14.790 613.740 15.110 613.800 ;
        RECT 1093.490 613.740 1093.810 613.800 ;
      LAYER via ;
        RECT 1093.520 1998.560 1093.780 1998.820 ;
        RECT 1425.180 1998.560 1425.440 1998.820 ;
        RECT 14.820 613.740 15.080 614.000 ;
        RECT 1093.520 613.740 1093.780 614.000 ;
      LAYER met2 ;
        RECT 1426.920 1998.930 1427.200 2000.000 ;
        RECT 1425.240 1998.850 1427.200 1998.930 ;
        RECT 1093.520 1998.530 1093.780 1998.850 ;
        RECT 1425.180 1998.790 1427.200 1998.850 ;
        RECT 1425.180 1998.530 1425.440 1998.790 ;
        RECT 1093.580 614.030 1093.720 1998.530 ;
        RECT 1426.920 1996.000 1427.200 1998.790 ;
        RECT 14.820 613.710 15.080 614.030 ;
        RECT 1093.520 613.710 1093.780 614.030 ;
        RECT 14.880 610.485 15.020 613.710 ;
        RECT 14.810 610.115 15.090 610.485 ;
      LAYER via2 ;
        RECT 14.810 610.160 15.090 610.440 ;
      LAYER met3 ;
        RECT -4.800 610.450 2.400 610.900 ;
        RECT 14.785 610.450 15.115 610.465 ;
        RECT -4.800 610.150 15.115 610.450 ;
        RECT -4.800 609.700 2.400 610.150 ;
        RECT 14.785 610.135 15.115 610.150 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1079.690 2003.180 1080.010 2003.240 ;
        RECT 1434.810 2003.180 1435.130 2003.240 ;
        RECT 1079.690 2003.040 1435.130 2003.180 ;
        RECT 1079.690 2002.980 1080.010 2003.040 ;
        RECT 1434.810 2002.980 1435.130 2003.040 ;
        RECT 16.170 400.080 16.490 400.140 ;
        RECT 1079.690 400.080 1080.010 400.140 ;
        RECT 16.170 399.940 1080.010 400.080 ;
        RECT 16.170 399.880 16.490 399.940 ;
        RECT 1079.690 399.880 1080.010 399.940 ;
      LAYER via ;
        RECT 1079.720 2002.980 1079.980 2003.240 ;
        RECT 1434.840 2002.980 1435.100 2003.240 ;
        RECT 16.200 399.880 16.460 400.140 ;
        RECT 1079.720 399.880 1079.980 400.140 ;
      LAYER met2 ;
        RECT 1079.720 2002.950 1079.980 2003.270 ;
        RECT 1434.840 2002.950 1435.100 2003.270 ;
        RECT 1079.780 400.170 1079.920 2002.950 ;
        RECT 1434.900 2000.000 1435.040 2002.950 ;
        RECT 1434.740 1999.540 1435.040 2000.000 ;
        RECT 1434.740 1996.000 1435.020 1999.540 ;
        RECT 16.200 399.850 16.460 400.170 ;
        RECT 1079.720 399.850 1079.980 400.170 ;
        RECT 16.260 394.925 16.400 399.850 ;
        RECT 16.190 394.555 16.470 394.925 ;
      LAYER via2 ;
        RECT 16.190 394.600 16.470 394.880 ;
      LAYER met3 ;
        RECT -4.800 394.890 2.400 395.340 ;
        RECT 16.165 394.890 16.495 394.905 ;
        RECT -4.800 394.590 16.495 394.890 ;
        RECT -4.800 394.140 2.400 394.590 ;
        RECT 16.165 394.575 16.495 394.590 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1072.790 1998.080 1073.110 1998.140 ;
        RECT 1441.710 1998.080 1442.030 1998.140 ;
        RECT 1072.790 1997.940 1442.030 1998.080 ;
        RECT 1072.790 1997.880 1073.110 1997.940 ;
        RECT 1441.710 1997.880 1442.030 1997.940 ;
        RECT 17.550 179.420 17.870 179.480 ;
        RECT 1072.790 179.420 1073.110 179.480 ;
        RECT 17.550 179.280 1073.110 179.420 ;
        RECT 17.550 179.220 17.870 179.280 ;
        RECT 1072.790 179.220 1073.110 179.280 ;
      LAYER via ;
        RECT 1072.820 1997.880 1073.080 1998.140 ;
        RECT 1441.740 1997.880 1442.000 1998.140 ;
        RECT 17.580 179.220 17.840 179.480 ;
        RECT 1072.820 179.220 1073.080 179.480 ;
      LAYER met2 ;
        RECT 1442.560 1998.250 1442.840 2000.000 ;
        RECT 1441.800 1998.170 1442.840 1998.250 ;
        RECT 1072.820 1997.850 1073.080 1998.170 ;
        RECT 1441.740 1998.110 1442.840 1998.170 ;
        RECT 1441.740 1997.850 1442.000 1998.110 ;
        RECT 1072.880 179.510 1073.020 1997.850 ;
        RECT 1442.560 1996.000 1442.840 1998.110 ;
        RECT 17.580 179.365 17.840 179.510 ;
        RECT 17.570 178.995 17.850 179.365 ;
        RECT 1072.820 179.190 1073.080 179.510 ;
      LAYER via2 ;
        RECT 17.570 179.040 17.850 179.320 ;
      LAYER met3 ;
        RECT -4.800 179.330 2.400 179.780 ;
        RECT 17.545 179.330 17.875 179.345 ;
        RECT -4.800 179.030 17.875 179.330 ;
        RECT -4.800 178.580 2.400 179.030 ;
        RECT 17.545 179.015 17.875 179.030 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1174.450 2004.540 1174.770 2004.600 ;
        RECT 1487.250 2004.540 1487.570 2004.600 ;
        RECT 1174.450 2004.400 1487.570 2004.540 ;
        RECT 1174.450 2004.340 1174.770 2004.400 ;
        RECT 1487.250 2004.340 1487.570 2004.400 ;
        RECT 1487.250 793.460 1487.570 793.520 ;
        RECT 2898.990 793.460 2899.310 793.520 ;
        RECT 1487.250 793.320 2899.310 793.460 ;
        RECT 1487.250 793.260 1487.570 793.320 ;
        RECT 2898.990 793.260 2899.310 793.320 ;
      LAYER via ;
        RECT 1174.480 2004.340 1174.740 2004.600 ;
        RECT 1487.280 2004.340 1487.540 2004.600 ;
        RECT 1487.280 793.260 1487.540 793.520 ;
        RECT 2899.020 793.260 2899.280 793.520 ;
      LAYER met2 ;
        RECT 1174.480 2004.310 1174.740 2004.630 ;
        RECT 1487.280 2004.310 1487.540 2004.630 ;
        RECT 1174.540 2000.000 1174.680 2004.310 ;
        RECT 1174.380 1999.540 1174.680 2000.000 ;
        RECT 1174.380 1996.000 1174.660 1999.540 ;
        RECT 1487.340 793.550 1487.480 2004.310 ;
        RECT 1487.280 793.230 1487.540 793.550 ;
        RECT 2899.020 793.230 2899.280 793.550 ;
        RECT 2899.080 792.045 2899.220 793.230 ;
        RECT 2899.010 791.675 2899.290 792.045 ;
      LAYER via2 ;
        RECT 2899.010 791.720 2899.290 792.000 ;
      LAYER met3 ;
        RECT 2898.985 792.010 2899.315 792.025 ;
        RECT 2917.600 792.010 2924.800 792.460 ;
        RECT 2898.985 791.710 2924.800 792.010 ;
        RECT 2898.985 791.695 2899.315 791.710 ;
        RECT 2917.600 791.260 2924.800 791.710 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1183.650 1999.780 1183.970 1999.840 ;
        RECT 1494.150 1999.780 1494.470 1999.840 ;
        RECT 1183.650 1999.640 1494.470 1999.780 ;
        RECT 1183.650 1999.580 1183.970 1999.640 ;
        RECT 1494.150 1999.580 1494.470 1999.640 ;
        RECT 1494.150 1028.060 1494.470 1028.120 ;
        RECT 2898.990 1028.060 2899.310 1028.120 ;
        RECT 1494.150 1027.920 2899.310 1028.060 ;
        RECT 1494.150 1027.860 1494.470 1027.920 ;
        RECT 2898.990 1027.860 2899.310 1027.920 ;
      LAYER via ;
        RECT 1183.680 1999.580 1183.940 1999.840 ;
        RECT 1494.180 1999.580 1494.440 1999.840 ;
        RECT 1494.180 1027.860 1494.440 1028.120 ;
        RECT 2899.020 1027.860 2899.280 1028.120 ;
      LAYER met2 ;
        RECT 1182.200 1999.610 1182.480 2000.000 ;
        RECT 1183.680 1999.610 1183.940 1999.870 ;
        RECT 1182.200 1999.550 1183.940 1999.610 ;
        RECT 1494.180 1999.550 1494.440 1999.870 ;
        RECT 1182.200 1999.470 1183.880 1999.550 ;
        RECT 1182.200 1996.000 1182.480 1999.470 ;
        RECT 1494.240 1028.150 1494.380 1999.550 ;
        RECT 1494.180 1027.830 1494.440 1028.150 ;
        RECT 2899.020 1027.830 2899.280 1028.150 ;
        RECT 2899.080 1026.645 2899.220 1027.830 ;
        RECT 2899.010 1026.275 2899.290 1026.645 ;
      LAYER via2 ;
        RECT 2899.010 1026.320 2899.290 1026.600 ;
      LAYER met3 ;
        RECT 2898.985 1026.610 2899.315 1026.625 ;
        RECT 2917.600 1026.610 2924.800 1027.060 ;
        RECT 2898.985 1026.310 2924.800 1026.610 ;
        RECT 2898.985 1026.295 2899.315 1026.310 ;
        RECT 2917.600 1025.860 2924.800 1026.310 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1190.090 2003.860 1190.410 2003.920 ;
        RECT 1507.950 2003.860 1508.270 2003.920 ;
        RECT 1190.090 2003.720 1508.270 2003.860 ;
        RECT 1190.090 2003.660 1190.410 2003.720 ;
        RECT 1507.950 2003.660 1508.270 2003.720 ;
        RECT 1507.950 1262.660 1508.270 1262.720 ;
        RECT 2898.990 1262.660 2899.310 1262.720 ;
        RECT 1507.950 1262.520 2899.310 1262.660 ;
        RECT 1507.950 1262.460 1508.270 1262.520 ;
        RECT 2898.990 1262.460 2899.310 1262.520 ;
      LAYER via ;
        RECT 1190.120 2003.660 1190.380 2003.920 ;
        RECT 1507.980 2003.660 1508.240 2003.920 ;
        RECT 1507.980 1262.460 1508.240 1262.720 ;
        RECT 2899.020 1262.460 2899.280 1262.720 ;
      LAYER met2 ;
        RECT 1190.120 2003.630 1190.380 2003.950 ;
        RECT 1507.980 2003.630 1508.240 2003.950 ;
        RECT 1190.180 2000.000 1190.320 2003.630 ;
        RECT 1190.020 1999.540 1190.320 2000.000 ;
        RECT 1190.020 1996.000 1190.300 1999.540 ;
        RECT 1508.040 1262.750 1508.180 2003.630 ;
        RECT 1507.980 1262.430 1508.240 1262.750 ;
        RECT 2899.020 1262.430 2899.280 1262.750 ;
        RECT 2899.080 1261.245 2899.220 1262.430 ;
        RECT 2899.010 1260.875 2899.290 1261.245 ;
      LAYER via2 ;
        RECT 2899.010 1260.920 2899.290 1261.200 ;
      LAYER met3 ;
        RECT 2898.985 1261.210 2899.315 1261.225 ;
        RECT 2917.600 1261.210 2924.800 1261.660 ;
        RECT 2898.985 1260.910 2924.800 1261.210 ;
        RECT 2898.985 1260.895 2899.315 1260.910 ;
        RECT 2917.600 1260.460 2924.800 1260.910 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1199.290 1999.440 1199.610 1999.500 ;
        RECT 1514.850 1999.440 1515.170 1999.500 ;
        RECT 1199.290 1999.300 1515.170 1999.440 ;
        RECT 1199.290 1999.240 1199.610 1999.300 ;
        RECT 1514.850 1999.240 1515.170 1999.300 ;
        RECT 1514.850 1497.260 1515.170 1497.320 ;
        RECT 2898.990 1497.260 2899.310 1497.320 ;
        RECT 1514.850 1497.120 2899.310 1497.260 ;
        RECT 1514.850 1497.060 1515.170 1497.120 ;
        RECT 2898.990 1497.060 2899.310 1497.120 ;
      LAYER via ;
        RECT 1199.320 1999.240 1199.580 1999.500 ;
        RECT 1514.880 1999.240 1515.140 1999.500 ;
        RECT 1514.880 1497.060 1515.140 1497.320 ;
        RECT 2899.020 1497.060 2899.280 1497.320 ;
      LAYER met2 ;
        RECT 1197.840 1999.610 1198.120 2000.000 ;
        RECT 1197.840 1999.530 1199.520 1999.610 ;
        RECT 1197.840 1999.470 1199.580 1999.530 ;
        RECT 1197.840 1996.000 1198.120 1999.470 ;
        RECT 1199.320 1999.210 1199.580 1999.470 ;
        RECT 1514.880 1999.210 1515.140 1999.530 ;
        RECT 1514.940 1497.350 1515.080 1999.210 ;
        RECT 1514.880 1497.030 1515.140 1497.350 ;
        RECT 2899.020 1497.030 2899.280 1497.350 ;
        RECT 2899.080 1495.845 2899.220 1497.030 ;
        RECT 2899.010 1495.475 2899.290 1495.845 ;
      LAYER via2 ;
        RECT 2899.010 1495.520 2899.290 1495.800 ;
      LAYER met3 ;
        RECT 2898.985 1495.810 2899.315 1495.825 ;
        RECT 2917.600 1495.810 2924.800 1496.260 ;
        RECT 2898.985 1495.510 2924.800 1495.810 ;
        RECT 2898.985 1495.495 2899.315 1495.510 ;
        RECT 2917.600 1495.060 2924.800 1495.510 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1206.190 2001.140 1206.510 2001.200 ;
        RECT 1452.290 2001.140 1452.610 2001.200 ;
        RECT 1206.190 2001.000 1452.610 2001.140 ;
        RECT 1206.190 2000.940 1206.510 2001.000 ;
        RECT 1452.290 2000.940 1452.610 2001.000 ;
        RECT 1452.290 1731.860 1452.610 1731.920 ;
        RECT 2898.990 1731.860 2899.310 1731.920 ;
        RECT 1452.290 1731.720 2899.310 1731.860 ;
        RECT 1452.290 1731.660 1452.610 1731.720 ;
        RECT 2898.990 1731.660 2899.310 1731.720 ;
      LAYER via ;
        RECT 1206.220 2000.940 1206.480 2001.200 ;
        RECT 1452.320 2000.940 1452.580 2001.200 ;
        RECT 1452.320 1731.660 1452.580 1731.920 ;
        RECT 2899.020 1731.660 2899.280 1731.920 ;
      LAYER met2 ;
        RECT 1206.220 2000.910 1206.480 2001.230 ;
        RECT 1452.320 2000.910 1452.580 2001.230 ;
        RECT 1206.280 2000.000 1206.420 2000.910 ;
        RECT 1206.120 1999.540 1206.420 2000.000 ;
        RECT 1206.120 1996.000 1206.400 1999.540 ;
        RECT 1452.380 1731.950 1452.520 2000.910 ;
        RECT 1452.320 1731.630 1452.580 1731.950 ;
        RECT 2899.020 1731.630 2899.280 1731.950 ;
        RECT 2899.080 1730.445 2899.220 1731.630 ;
        RECT 2899.010 1730.075 2899.290 1730.445 ;
      LAYER via2 ;
        RECT 2899.010 1730.120 2899.290 1730.400 ;
      LAYER met3 ;
        RECT 2898.985 1730.410 2899.315 1730.425 ;
        RECT 2917.600 1730.410 2924.800 1730.860 ;
        RECT 2898.985 1730.110 2924.800 1730.410 ;
        RECT 2898.985 1730.095 2899.315 1730.110 ;
        RECT 2917.600 1729.660 2924.800 1730.110 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1213.090 2000.120 1213.410 2000.180 ;
        RECT 1453.210 2000.120 1453.530 2000.180 ;
        RECT 1213.090 1999.980 1453.530 2000.120 ;
        RECT 1213.090 1999.920 1213.410 1999.980 ;
        RECT 1453.210 1999.920 1453.530 1999.980 ;
        RECT 1453.210 1966.460 1453.530 1966.520 ;
        RECT 2898.990 1966.460 2899.310 1966.520 ;
        RECT 1453.210 1966.320 2899.310 1966.460 ;
        RECT 1453.210 1966.260 1453.530 1966.320 ;
        RECT 2898.990 1966.260 2899.310 1966.320 ;
      LAYER via ;
        RECT 1213.120 1999.920 1213.380 2000.180 ;
        RECT 1453.240 1999.920 1453.500 2000.180 ;
        RECT 1453.240 1966.260 1453.500 1966.520 ;
        RECT 2899.020 1966.260 2899.280 1966.520 ;
      LAYER met2 ;
        RECT 1213.120 1999.890 1213.380 2000.210 ;
        RECT 1213.180 1999.610 1213.320 1999.890 ;
        RECT 1213.940 1999.610 1214.220 2000.000 ;
        RECT 1453.240 1999.890 1453.500 2000.210 ;
        RECT 1213.180 1999.470 1214.220 1999.610 ;
        RECT 1213.940 1996.000 1214.220 1999.470 ;
        RECT 1453.300 1966.550 1453.440 1999.890 ;
        RECT 1453.240 1966.230 1453.500 1966.550 ;
        RECT 2899.020 1966.230 2899.280 1966.550 ;
        RECT 2899.080 1965.045 2899.220 1966.230 ;
        RECT 2899.010 1964.675 2899.290 1965.045 ;
      LAYER via2 ;
        RECT 2899.010 1964.720 2899.290 1965.000 ;
      LAYER met3 ;
        RECT 2898.985 1965.010 2899.315 1965.025 ;
        RECT 2917.600 1965.010 2924.800 1965.460 ;
        RECT 2898.985 1964.710 2924.800 1965.010 ;
        RECT 2898.985 1964.695 2899.315 1964.710 ;
        RECT 2917.600 1964.260 2924.800 1964.710 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1226.890 2194.600 1227.210 2194.660 ;
        RECT 2900.830 2194.600 2901.150 2194.660 ;
        RECT 1226.890 2194.460 2901.150 2194.600 ;
        RECT 1226.890 2194.400 1227.210 2194.460 ;
        RECT 2900.830 2194.400 2901.150 2194.460 ;
        RECT 1221.830 2009.300 1222.150 2009.360 ;
        RECT 1226.890 2009.300 1227.210 2009.360 ;
        RECT 1221.830 2009.160 1227.210 2009.300 ;
        RECT 1221.830 2009.100 1222.150 2009.160 ;
        RECT 1226.890 2009.100 1227.210 2009.160 ;
      LAYER via ;
        RECT 1226.920 2194.400 1227.180 2194.660 ;
        RECT 2900.860 2194.400 2901.120 2194.660 ;
        RECT 1221.860 2009.100 1222.120 2009.360 ;
        RECT 1226.920 2009.100 1227.180 2009.360 ;
      LAYER met2 ;
        RECT 2900.850 2199.275 2901.130 2199.645 ;
        RECT 2900.920 2194.690 2901.060 2199.275 ;
        RECT 1226.920 2194.370 1227.180 2194.690 ;
        RECT 2900.860 2194.370 2901.120 2194.690 ;
        RECT 1226.980 2009.390 1227.120 2194.370 ;
        RECT 1221.860 2009.070 1222.120 2009.390 ;
        RECT 1226.920 2009.070 1227.180 2009.390 ;
        RECT 1221.920 2000.000 1222.060 2009.070 ;
        RECT 1221.760 1999.540 1222.060 2000.000 ;
        RECT 1221.760 1996.000 1222.040 1999.540 ;
      LAYER via2 ;
        RECT 2900.850 2199.320 2901.130 2199.600 ;
      LAYER met3 ;
        RECT 2900.825 2199.610 2901.155 2199.625 ;
        RECT 2917.600 2199.610 2924.800 2200.060 ;
        RECT 2900.825 2199.310 2924.800 2199.610 ;
        RECT 2900.825 2199.295 2901.155 2199.310 ;
        RECT 2917.600 2198.860 2924.800 2199.310 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1153.290 2002.160 1153.610 2002.220 ;
        RECT 1521.290 2002.160 1521.610 2002.220 ;
        RECT 1153.290 2002.020 1521.610 2002.160 ;
        RECT 1153.290 2001.960 1153.610 2002.020 ;
        RECT 1521.290 2001.960 1521.610 2002.020 ;
        RECT 1521.290 206.960 1521.610 207.020 ;
        RECT 2900.830 206.960 2901.150 207.020 ;
        RECT 1521.290 206.820 2901.150 206.960 ;
        RECT 1521.290 206.760 1521.610 206.820 ;
        RECT 2900.830 206.760 2901.150 206.820 ;
      LAYER via ;
        RECT 1153.320 2001.960 1153.580 2002.220 ;
        RECT 1521.320 2001.960 1521.580 2002.220 ;
        RECT 1521.320 206.760 1521.580 207.020 ;
        RECT 2900.860 206.760 2901.120 207.020 ;
      LAYER met2 ;
        RECT 1153.320 2001.930 1153.580 2002.250 ;
        RECT 1521.320 2001.930 1521.580 2002.250 ;
        RECT 1153.380 2000.000 1153.520 2001.930 ;
        RECT 1153.220 1999.540 1153.520 2000.000 ;
        RECT 1153.220 1996.000 1153.500 1999.540 ;
        RECT 1521.380 207.050 1521.520 2001.930 ;
        RECT 1521.320 206.730 1521.580 207.050 ;
        RECT 2900.860 206.730 2901.120 207.050 ;
        RECT 2900.920 205.205 2901.060 206.730 ;
        RECT 2900.850 204.835 2901.130 205.205 ;
      LAYER via2 ;
        RECT 2900.850 204.880 2901.130 205.160 ;
      LAYER met3 ;
        RECT 2900.825 205.170 2901.155 205.185 ;
        RECT 2917.600 205.170 2924.800 205.620 ;
        RECT 2900.825 204.870 2924.800 205.170 ;
        RECT 2900.825 204.855 2901.155 204.870 ;
        RECT 2917.600 204.420 2924.800 204.870 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1234.710 2546.500 1235.030 2546.560 ;
        RECT 2900.830 2546.500 2901.150 2546.560 ;
        RECT 1234.710 2546.360 2901.150 2546.500 ;
        RECT 1234.710 2546.300 1235.030 2546.360 ;
        RECT 2900.830 2546.300 2901.150 2546.360 ;
      LAYER via ;
        RECT 1234.740 2546.300 1235.000 2546.560 ;
        RECT 2900.860 2546.300 2901.120 2546.560 ;
      LAYER met2 ;
        RECT 2900.850 2551.515 2901.130 2551.885 ;
        RECT 2900.920 2546.590 2901.060 2551.515 ;
        RECT 1234.740 2546.270 1235.000 2546.590 ;
        RECT 2900.860 2546.270 2901.120 2546.590 ;
        RECT 1232.340 1999.610 1232.620 2000.000 ;
        RECT 1234.800 1999.610 1234.940 2546.270 ;
        RECT 1232.340 1999.470 1234.940 1999.610 ;
        RECT 1232.340 1996.000 1232.620 1999.470 ;
      LAYER via2 ;
        RECT 2900.850 2551.560 2901.130 2551.840 ;
      LAYER met3 ;
        RECT 2900.825 2551.850 2901.155 2551.865 ;
        RECT 2917.600 2551.850 2924.800 2552.300 ;
        RECT 2900.825 2551.550 2924.800 2551.850 ;
        RECT 2900.825 2551.535 2901.155 2551.550 ;
        RECT 2917.600 2551.100 2924.800 2551.550 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1241.610 2781.100 1241.930 2781.160 ;
        RECT 2900.830 2781.100 2901.150 2781.160 ;
        RECT 1241.610 2780.960 2901.150 2781.100 ;
        RECT 1241.610 2780.900 1241.930 2780.960 ;
        RECT 2900.830 2780.900 2901.150 2780.960 ;
      LAYER via ;
        RECT 1241.640 2780.900 1241.900 2781.160 ;
        RECT 2900.860 2780.900 2901.120 2781.160 ;
      LAYER met2 ;
        RECT 2900.850 2786.115 2901.130 2786.485 ;
        RECT 2900.920 2781.190 2901.060 2786.115 ;
        RECT 1241.640 2780.870 1241.900 2781.190 ;
        RECT 2900.860 2780.870 2901.120 2781.190 ;
        RECT 1240.160 1999.610 1240.440 2000.000 ;
        RECT 1241.700 1999.610 1241.840 2780.870 ;
        RECT 1240.160 1999.470 1241.840 1999.610 ;
        RECT 1240.160 1996.000 1240.440 1999.470 ;
      LAYER via2 ;
        RECT 2900.850 2786.160 2901.130 2786.440 ;
      LAYER met3 ;
        RECT 2900.825 2786.450 2901.155 2786.465 ;
        RECT 2917.600 2786.450 2924.800 2786.900 ;
        RECT 2900.825 2786.150 2924.800 2786.450 ;
        RECT 2900.825 2786.135 2901.155 2786.150 ;
        RECT 2917.600 2785.700 2924.800 2786.150 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1248.510 3015.700 1248.830 3015.760 ;
        RECT 2900.830 3015.700 2901.150 3015.760 ;
        RECT 1248.510 3015.560 2901.150 3015.700 ;
        RECT 1248.510 3015.500 1248.830 3015.560 ;
        RECT 2900.830 3015.500 2901.150 3015.560 ;
      LAYER via ;
        RECT 1248.540 3015.500 1248.800 3015.760 ;
        RECT 2900.860 3015.500 2901.120 3015.760 ;
      LAYER met2 ;
        RECT 2900.850 3020.715 2901.130 3021.085 ;
        RECT 2900.920 3015.790 2901.060 3020.715 ;
        RECT 1248.540 3015.470 1248.800 3015.790 ;
        RECT 2900.860 3015.470 2901.120 3015.790 ;
        RECT 1247.980 1999.610 1248.260 2000.000 ;
        RECT 1248.600 1999.610 1248.740 3015.470 ;
        RECT 1247.980 1999.470 1248.740 1999.610 ;
        RECT 1247.980 1996.000 1248.260 1999.470 ;
      LAYER via2 ;
        RECT 2900.850 3020.760 2901.130 3021.040 ;
      LAYER met3 ;
        RECT 2900.825 3021.050 2901.155 3021.065 ;
        RECT 2917.600 3021.050 2924.800 3021.500 ;
        RECT 2900.825 3020.750 2924.800 3021.050 ;
        RECT 2900.825 3020.735 2901.155 3020.750 ;
        RECT 2917.600 3020.300 2924.800 3020.750 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1261.850 3250.300 1262.170 3250.360 ;
        RECT 2900.830 3250.300 2901.150 3250.360 ;
        RECT 1261.850 3250.160 2901.150 3250.300 ;
        RECT 1261.850 3250.100 1262.170 3250.160 ;
        RECT 2900.830 3250.100 2901.150 3250.160 ;
        RECT 1255.870 2009.980 1256.190 2010.040 ;
        RECT 1261.850 2009.980 1262.170 2010.040 ;
        RECT 1255.870 2009.840 1262.170 2009.980 ;
        RECT 1255.870 2009.780 1256.190 2009.840 ;
        RECT 1261.850 2009.780 1262.170 2009.840 ;
      LAYER via ;
        RECT 1261.880 3250.100 1262.140 3250.360 ;
        RECT 2900.860 3250.100 2901.120 3250.360 ;
        RECT 1255.900 2009.780 1256.160 2010.040 ;
        RECT 1261.880 2009.780 1262.140 2010.040 ;
      LAYER met2 ;
        RECT 2900.850 3255.315 2901.130 3255.685 ;
        RECT 2900.920 3250.390 2901.060 3255.315 ;
        RECT 1261.880 3250.070 1262.140 3250.390 ;
        RECT 2900.860 3250.070 2901.120 3250.390 ;
        RECT 1261.940 2010.070 1262.080 3250.070 ;
        RECT 1255.900 2009.750 1256.160 2010.070 ;
        RECT 1261.880 2009.750 1262.140 2010.070 ;
        RECT 1255.960 2000.000 1256.100 2009.750 ;
        RECT 1255.800 1999.540 1256.100 2000.000 ;
        RECT 1255.800 1996.000 1256.080 1999.540 ;
      LAYER via2 ;
        RECT 2900.850 3255.360 2901.130 3255.640 ;
      LAYER met3 ;
        RECT 2900.825 3255.650 2901.155 3255.665 ;
        RECT 2917.600 3255.650 2924.800 3256.100 ;
        RECT 2900.825 3255.350 2924.800 3255.650 ;
        RECT 2900.825 3255.335 2901.155 3255.350 ;
        RECT 2917.600 3254.900 2924.800 3255.350 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1268.750 3484.900 1269.070 3484.960 ;
        RECT 2900.830 3484.900 2901.150 3484.960 ;
        RECT 1268.750 3484.760 2901.150 3484.900 ;
        RECT 1268.750 3484.700 1269.070 3484.760 ;
        RECT 2900.830 3484.700 2901.150 3484.760 ;
        RECT 1263.690 2009.980 1264.010 2010.040 ;
        RECT 1268.750 2009.980 1269.070 2010.040 ;
        RECT 1263.690 2009.840 1269.070 2009.980 ;
        RECT 1263.690 2009.780 1264.010 2009.840 ;
        RECT 1268.750 2009.780 1269.070 2009.840 ;
      LAYER via ;
        RECT 1268.780 3484.700 1269.040 3484.960 ;
        RECT 2900.860 3484.700 2901.120 3484.960 ;
        RECT 1263.720 2009.780 1263.980 2010.040 ;
        RECT 1268.780 2009.780 1269.040 2010.040 ;
      LAYER met2 ;
        RECT 2900.850 3489.915 2901.130 3490.285 ;
        RECT 2900.920 3484.990 2901.060 3489.915 ;
        RECT 1268.780 3484.670 1269.040 3484.990 ;
        RECT 2900.860 3484.670 2901.120 3484.990 ;
        RECT 1268.840 2010.070 1268.980 3484.670 ;
        RECT 1263.720 2009.750 1263.980 2010.070 ;
        RECT 1268.780 2009.750 1269.040 2010.070 ;
        RECT 1263.780 2000.000 1263.920 2009.750 ;
        RECT 1263.620 1999.540 1263.920 2000.000 ;
        RECT 1263.620 1996.000 1263.900 1999.540 ;
      LAYER via2 ;
        RECT 2900.850 3489.960 2901.130 3490.240 ;
      LAYER met3 ;
        RECT 2900.825 3490.250 2901.155 3490.265 ;
        RECT 2917.600 3490.250 2924.800 3490.700 ;
        RECT 2900.825 3489.950 2924.800 3490.250 ;
        RECT 2900.825 3489.935 2901.155 3489.950 ;
        RECT 2917.600 3489.500 2924.800 3489.950 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1276.110 3502.240 1276.430 3502.300 ;
        RECT 2635.870 3502.240 2636.190 3502.300 ;
        RECT 1276.110 3502.100 2636.190 3502.240 ;
        RECT 1276.110 3502.040 1276.430 3502.100 ;
        RECT 2635.870 3502.040 2636.190 3502.100 ;
        RECT 1271.970 2013.720 1272.290 2013.780 ;
        RECT 1276.110 2013.720 1276.430 2013.780 ;
        RECT 1271.970 2013.580 1276.430 2013.720 ;
        RECT 1271.970 2013.520 1272.290 2013.580 ;
        RECT 1276.110 2013.520 1276.430 2013.580 ;
      LAYER via ;
        RECT 1276.140 3502.040 1276.400 3502.300 ;
        RECT 2635.900 3502.040 2636.160 3502.300 ;
        RECT 1272.000 2013.520 1272.260 2013.780 ;
        RECT 1276.140 2013.520 1276.400 2013.780 ;
      LAYER met2 ;
        RECT 2635.750 3517.600 2636.310 3524.800 ;
        RECT 2635.960 3502.330 2636.100 3517.600 ;
        RECT 1276.140 3502.010 1276.400 3502.330 ;
        RECT 2635.900 3502.010 2636.160 3502.330 ;
        RECT 1276.200 2013.810 1276.340 3502.010 ;
        RECT 1272.000 2013.490 1272.260 2013.810 ;
        RECT 1276.140 2013.490 1276.400 2013.810 ;
        RECT 1272.060 2000.000 1272.200 2013.490 ;
        RECT 1271.900 1999.540 1272.200 2000.000 ;
        RECT 1271.900 1996.000 1272.180 1999.540 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1282.550 3503.600 1282.870 3503.660 ;
        RECT 2311.570 3503.600 2311.890 3503.660 ;
        RECT 1282.550 3503.460 2311.890 3503.600 ;
        RECT 1282.550 3503.400 1282.870 3503.460 ;
        RECT 2311.570 3503.400 2311.890 3503.460 ;
      LAYER via ;
        RECT 1282.580 3503.400 1282.840 3503.660 ;
        RECT 2311.600 3503.400 2311.860 3503.660 ;
      LAYER met2 ;
        RECT 2311.450 3517.600 2312.010 3524.800 ;
        RECT 2311.660 3503.690 2311.800 3517.600 ;
        RECT 1282.580 3503.370 1282.840 3503.690 ;
        RECT 2311.600 3503.370 2311.860 3503.690 ;
        RECT 1282.640 2000.290 1282.780 3503.370 ;
        RECT 1281.720 2000.150 1282.780 2000.290 ;
        RECT 1279.720 1999.610 1280.000 2000.000 ;
        RECT 1281.720 1999.610 1281.860 2000.150 ;
        RECT 1279.720 1999.470 1281.860 1999.610 ;
        RECT 1279.720 1996.000 1280.000 1999.470 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1289.450 3504.960 1289.770 3505.020 ;
        RECT 1987.270 3504.960 1987.590 3505.020 ;
        RECT 1289.450 3504.820 1987.590 3504.960 ;
        RECT 1289.450 3504.760 1289.770 3504.820 ;
        RECT 1987.270 3504.760 1987.590 3504.820 ;
      LAYER via ;
        RECT 1289.480 3504.760 1289.740 3505.020 ;
        RECT 1987.300 3504.760 1987.560 3505.020 ;
      LAYER met2 ;
        RECT 1987.150 3517.600 1987.710 3524.800 ;
        RECT 1987.360 3505.050 1987.500 3517.600 ;
        RECT 1289.480 3504.730 1289.740 3505.050 ;
        RECT 1987.300 3504.730 1987.560 3505.050 ;
        RECT 1287.540 1999.610 1287.820 2000.000 ;
        RECT 1289.540 1999.610 1289.680 3504.730 ;
        RECT 1287.540 1999.470 1289.680 1999.610 ;
        RECT 1287.540 1996.000 1287.820 1999.470 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1295.890 3500.200 1296.210 3500.260 ;
        RECT 1662.510 3500.200 1662.830 3500.260 ;
        RECT 1295.890 3500.060 1662.830 3500.200 ;
        RECT 1295.890 3500.000 1296.210 3500.060 ;
        RECT 1662.510 3500.000 1662.830 3500.060 ;
      LAYER via ;
        RECT 1295.920 3500.000 1296.180 3500.260 ;
        RECT 1662.540 3500.000 1662.800 3500.260 ;
      LAYER met2 ;
        RECT 1662.390 3517.600 1662.950 3524.800 ;
        RECT 1662.600 3500.290 1662.740 3517.600 ;
        RECT 1295.920 3499.970 1296.180 3500.290 ;
        RECT 1662.540 3499.970 1662.800 3500.290 ;
        RECT 1295.360 1999.610 1295.640 2000.000 ;
        RECT 1295.980 1999.610 1296.120 3499.970 ;
        RECT 1295.360 1999.470 1296.120 1999.610 ;
        RECT 1295.360 1996.000 1295.640 1999.470 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1303.710 3498.500 1304.030 3498.560 ;
        RECT 1338.210 3498.500 1338.530 3498.560 ;
        RECT 1303.710 3498.360 1338.530 3498.500 ;
        RECT 1303.710 3498.300 1304.030 3498.360 ;
        RECT 1338.210 3498.300 1338.530 3498.360 ;
      LAYER via ;
        RECT 1303.740 3498.300 1304.000 3498.560 ;
        RECT 1338.240 3498.300 1338.500 3498.560 ;
      LAYER met2 ;
        RECT 1338.090 3517.600 1338.650 3524.800 ;
        RECT 1338.300 3498.590 1338.440 3517.600 ;
        RECT 1303.740 3498.270 1304.000 3498.590 ;
        RECT 1338.240 3498.270 1338.500 3498.590 ;
        RECT 1303.180 1999.610 1303.460 2000.000 ;
        RECT 1303.800 1999.610 1303.940 3498.270 ;
        RECT 1303.180 1999.470 1303.940 1999.610 ;
        RECT 1303.180 1996.000 1303.460 1999.470 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1162.490 1998.420 1162.810 1998.480 ;
        RECT 1528.190 1998.420 1528.510 1998.480 ;
        RECT 1162.490 1998.280 1528.510 1998.420 ;
        RECT 1162.490 1998.220 1162.810 1998.280 ;
        RECT 1528.190 1998.220 1528.510 1998.280 ;
        RECT 1528.190 441.560 1528.510 441.620 ;
        RECT 2900.830 441.560 2901.150 441.620 ;
        RECT 1528.190 441.420 2901.150 441.560 ;
        RECT 1528.190 441.360 1528.510 441.420 ;
        RECT 2900.830 441.360 2901.150 441.420 ;
      LAYER via ;
        RECT 1162.520 1998.220 1162.780 1998.480 ;
        RECT 1528.220 1998.220 1528.480 1998.480 ;
        RECT 1528.220 441.360 1528.480 441.620 ;
        RECT 2900.860 441.360 2901.120 441.620 ;
      LAYER met2 ;
        RECT 1161.040 1998.250 1161.320 2000.000 ;
        RECT 1162.520 1998.250 1162.780 1998.510 ;
        RECT 1161.040 1998.190 1162.780 1998.250 ;
        RECT 1528.220 1998.190 1528.480 1998.510 ;
        RECT 1161.040 1998.110 1162.720 1998.190 ;
        RECT 1161.040 1996.000 1161.320 1998.110 ;
        RECT 1528.280 441.650 1528.420 1998.190 ;
        RECT 1528.220 441.330 1528.480 441.650 ;
        RECT 2900.860 441.330 2901.120 441.650 ;
        RECT 2900.920 439.805 2901.060 441.330 ;
        RECT 2900.850 439.435 2901.130 439.805 ;
      LAYER via2 ;
        RECT 2900.850 439.480 2901.130 439.760 ;
      LAYER met3 ;
        RECT 2900.825 439.770 2901.155 439.785 ;
        RECT 2917.600 439.770 2924.800 440.220 ;
        RECT 2900.825 439.470 2924.800 439.770 ;
        RECT 2900.825 439.455 2901.155 439.470 ;
        RECT 2917.600 439.020 2924.800 439.470 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1013.910 3499.860 1014.230 3499.920 ;
        RECT 1311.070 3499.860 1311.390 3499.920 ;
        RECT 1013.910 3499.720 1311.390 3499.860 ;
        RECT 1013.910 3499.660 1014.230 3499.720 ;
        RECT 1311.070 3499.660 1311.390 3499.720 ;
      LAYER via ;
        RECT 1013.940 3499.660 1014.200 3499.920 ;
        RECT 1311.100 3499.660 1311.360 3499.920 ;
      LAYER met2 ;
        RECT 1013.790 3517.600 1014.350 3524.800 ;
        RECT 1014.000 3499.950 1014.140 3517.600 ;
        RECT 1013.940 3499.630 1014.200 3499.950 ;
        RECT 1311.100 3499.630 1311.360 3499.950 ;
        RECT 1311.160 2000.000 1311.300 3499.630 ;
        RECT 1311.000 1999.540 1311.300 2000.000 ;
        RECT 1311.000 1996.000 1311.280 1999.540 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 689.150 3501.220 689.470 3501.280 ;
        RECT 1318.890 3501.220 1319.210 3501.280 ;
        RECT 689.150 3501.080 1319.210 3501.220 ;
        RECT 689.150 3501.020 689.470 3501.080 ;
        RECT 1318.890 3501.020 1319.210 3501.080 ;
      LAYER via ;
        RECT 689.180 3501.020 689.440 3501.280 ;
        RECT 1318.920 3501.020 1319.180 3501.280 ;
      LAYER met2 ;
        RECT 689.030 3517.600 689.590 3524.800 ;
        RECT 689.240 3501.310 689.380 3517.600 ;
        RECT 689.180 3500.990 689.440 3501.310 ;
        RECT 1318.920 3500.990 1319.180 3501.310 ;
        RECT 1318.980 1999.610 1319.120 3500.990 ;
        RECT 1319.280 1999.610 1319.560 2000.000 ;
        RECT 1318.980 1999.470 1319.560 1999.610 ;
        RECT 1319.280 1996.000 1319.560 1999.470 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 364.850 3503.940 365.170 3504.000 ;
        RECT 1325.330 3503.940 1325.650 3504.000 ;
        RECT 364.850 3503.800 1325.650 3503.940 ;
        RECT 364.850 3503.740 365.170 3503.800 ;
        RECT 1325.330 3503.740 1325.650 3503.800 ;
      LAYER via ;
        RECT 364.880 3503.740 365.140 3504.000 ;
        RECT 1325.360 3503.740 1325.620 3504.000 ;
      LAYER met2 ;
        RECT 364.730 3517.600 365.290 3524.800 ;
        RECT 364.940 3504.030 365.080 3517.600 ;
        RECT 364.880 3503.710 365.140 3504.030 ;
        RECT 1325.360 3503.710 1325.620 3504.030 ;
        RECT 1325.420 1999.610 1325.560 3503.710 ;
        RECT 1327.100 1999.610 1327.380 2000.000 ;
        RECT 1325.420 1999.470 1327.380 1999.610 ;
        RECT 1327.100 1996.000 1327.380 1999.470 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 40.550 3502.580 40.870 3502.640 ;
        RECT 1332.690 3502.580 1333.010 3502.640 ;
        RECT 40.550 3502.440 1333.010 3502.580 ;
        RECT 40.550 3502.380 40.870 3502.440 ;
        RECT 1332.690 3502.380 1333.010 3502.440 ;
      LAYER via ;
        RECT 40.580 3502.380 40.840 3502.640 ;
        RECT 1332.720 3502.380 1332.980 3502.640 ;
      LAYER met2 ;
        RECT 40.430 3517.600 40.990 3524.800 ;
        RECT 40.640 3502.670 40.780 3517.600 ;
        RECT 40.580 3502.350 40.840 3502.670 ;
        RECT 1332.720 3502.350 1332.980 3502.670 ;
        RECT 1332.780 1999.610 1332.920 3502.350 ;
        RECT 1334.920 1999.610 1335.200 2000.000 ;
        RECT 1332.780 1999.470 1335.200 1999.610 ;
        RECT 1334.920 1996.000 1335.200 1999.470 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.630 3263.900 16.950 3263.960 ;
        RECT 1339.130 3263.900 1339.450 3263.960 ;
        RECT 16.630 3263.760 1339.450 3263.900 ;
        RECT 16.630 3263.700 16.950 3263.760 ;
        RECT 1339.130 3263.700 1339.450 3263.760 ;
      LAYER via ;
        RECT 16.660 3263.700 16.920 3263.960 ;
        RECT 1339.160 3263.700 1339.420 3263.960 ;
      LAYER met2 ;
        RECT 16.650 3267.555 16.930 3267.925 ;
        RECT 16.720 3263.990 16.860 3267.555 ;
        RECT 16.660 3263.670 16.920 3263.990 ;
        RECT 1339.160 3263.670 1339.420 3263.990 ;
        RECT 1339.220 2013.890 1339.360 3263.670 ;
        RECT 1339.220 2013.750 1340.740 2013.890 ;
        RECT 1340.600 1998.930 1340.740 2013.750 ;
        RECT 1342.740 1998.930 1343.020 2000.000 ;
        RECT 1340.600 1998.790 1343.020 1998.930 ;
        RECT 1342.740 1996.000 1343.020 1998.790 ;
      LAYER via2 ;
        RECT 16.650 3267.600 16.930 3267.880 ;
      LAYER met3 ;
        RECT -4.800 3267.890 2.400 3268.340 ;
        RECT 16.625 3267.890 16.955 3267.905 ;
        RECT -4.800 3267.590 16.955 3267.890 ;
        RECT -4.800 3267.140 2.400 3267.590 ;
        RECT 16.625 3267.575 16.955 3267.590 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.250 2974.220 15.570 2974.280 ;
        RECT 1346.490 2974.220 1346.810 2974.280 ;
        RECT 15.250 2974.080 1346.810 2974.220 ;
        RECT 15.250 2974.020 15.570 2974.080 ;
        RECT 1346.490 2974.020 1346.810 2974.080 ;
      LAYER via ;
        RECT 15.280 2974.020 15.540 2974.280 ;
        RECT 1346.520 2974.020 1346.780 2974.280 ;
      LAYER met2 ;
        RECT 15.270 2979.915 15.550 2980.285 ;
        RECT 15.340 2974.310 15.480 2979.915 ;
        RECT 15.280 2973.990 15.540 2974.310 ;
        RECT 1346.520 2973.990 1346.780 2974.310 ;
        RECT 1346.580 2011.850 1346.720 2973.990 ;
        RECT 1346.580 2011.710 1349.480 2011.850 ;
        RECT 1349.340 1999.610 1349.480 2011.710 ;
        RECT 1350.560 1999.610 1350.840 2000.000 ;
        RECT 1349.340 1999.470 1350.840 1999.610 ;
        RECT 1350.560 1996.000 1350.840 1999.470 ;
      LAYER via2 ;
        RECT 15.270 2979.960 15.550 2980.240 ;
      LAYER met3 ;
        RECT -4.800 2980.250 2.400 2980.700 ;
        RECT 15.245 2980.250 15.575 2980.265 ;
        RECT -4.800 2979.950 15.575 2980.250 ;
        RECT -4.800 2979.500 2.400 2979.950 ;
        RECT 15.245 2979.935 15.575 2979.950 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.710 2691.340 16.030 2691.400 ;
        RECT 1353.850 2691.340 1354.170 2691.400 ;
        RECT 15.710 2691.200 1354.170 2691.340 ;
        RECT 15.710 2691.140 16.030 2691.200 ;
        RECT 1353.850 2691.140 1354.170 2691.200 ;
      LAYER via ;
        RECT 15.740 2691.140 16.000 2691.400 ;
        RECT 1353.880 2691.140 1354.140 2691.400 ;
      LAYER met2 ;
        RECT 15.730 2692.955 16.010 2693.325 ;
        RECT 15.800 2691.430 15.940 2692.955 ;
        RECT 15.740 2691.110 16.000 2691.430 ;
        RECT 1353.880 2691.110 1354.140 2691.430 ;
        RECT 1353.940 2013.210 1354.080 2691.110 ;
        RECT 1353.940 2013.070 1357.760 2013.210 ;
        RECT 1357.620 1999.610 1357.760 2013.070 ;
        RECT 1358.380 1999.610 1358.660 2000.000 ;
        RECT 1357.620 1999.470 1358.660 1999.610 ;
        RECT 1358.380 1996.000 1358.660 1999.470 ;
      LAYER via2 ;
        RECT 15.730 2693.000 16.010 2693.280 ;
      LAYER met3 ;
        RECT -4.800 2693.290 2.400 2693.740 ;
        RECT 15.705 2693.290 16.035 2693.305 ;
        RECT -4.800 2692.990 16.035 2693.290 ;
        RECT -4.800 2692.540 2.400 2692.990 ;
        RECT 15.705 2692.975 16.035 2692.990 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 15.710 2401.320 16.030 2401.380 ;
        RECT 1362.590 2401.320 1362.910 2401.380 ;
        RECT 15.710 2401.180 1362.910 2401.320 ;
        RECT 15.710 2401.120 16.030 2401.180 ;
        RECT 1362.590 2401.120 1362.910 2401.180 ;
        RECT 1362.590 2009.640 1362.910 2009.700 ;
        RECT 1366.270 2009.640 1366.590 2009.700 ;
        RECT 1362.590 2009.500 1366.590 2009.640 ;
        RECT 1362.590 2009.440 1362.910 2009.500 ;
        RECT 1366.270 2009.440 1366.590 2009.500 ;
      LAYER via ;
        RECT 15.740 2401.120 16.000 2401.380 ;
        RECT 1362.620 2401.120 1362.880 2401.380 ;
        RECT 1362.620 2009.440 1362.880 2009.700 ;
        RECT 1366.300 2009.440 1366.560 2009.700 ;
      LAYER met2 ;
        RECT 15.730 2405.315 16.010 2405.685 ;
        RECT 15.800 2401.410 15.940 2405.315 ;
        RECT 15.740 2401.090 16.000 2401.410 ;
        RECT 1362.620 2401.090 1362.880 2401.410 ;
        RECT 1362.680 2009.730 1362.820 2401.090 ;
        RECT 1362.620 2009.410 1362.880 2009.730 ;
        RECT 1366.300 2009.410 1366.560 2009.730 ;
        RECT 1366.360 2000.000 1366.500 2009.410 ;
        RECT 1366.200 1999.540 1366.500 2000.000 ;
        RECT 1366.200 1996.000 1366.480 1999.540 ;
      LAYER via2 ;
        RECT 15.730 2405.360 16.010 2405.640 ;
      LAYER met3 ;
        RECT -4.800 2405.650 2.400 2406.100 ;
        RECT 15.705 2405.650 16.035 2405.665 ;
        RECT -4.800 2405.350 16.035 2405.650 ;
        RECT -4.800 2404.900 2.400 2405.350 ;
        RECT 15.705 2405.335 16.035 2405.350 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.630 2118.440 16.950 2118.500 ;
        RECT 1369.490 2118.440 1369.810 2118.500 ;
        RECT 16.630 2118.300 1369.810 2118.440 ;
        RECT 16.630 2118.240 16.950 2118.300 ;
        RECT 1369.490 2118.240 1369.810 2118.300 ;
        RECT 1369.490 2014.740 1369.810 2014.800 ;
        RECT 1374.550 2014.740 1374.870 2014.800 ;
        RECT 1369.490 2014.600 1374.870 2014.740 ;
        RECT 1369.490 2014.540 1369.810 2014.600 ;
        RECT 1374.550 2014.540 1374.870 2014.600 ;
      LAYER via ;
        RECT 16.660 2118.240 16.920 2118.500 ;
        RECT 1369.520 2118.240 1369.780 2118.500 ;
        RECT 1369.520 2014.540 1369.780 2014.800 ;
        RECT 1374.580 2014.540 1374.840 2014.800 ;
      LAYER met2 ;
        RECT 16.650 2118.355 16.930 2118.725 ;
        RECT 16.660 2118.210 16.920 2118.355 ;
        RECT 1369.520 2118.210 1369.780 2118.530 ;
        RECT 1369.580 2014.830 1369.720 2118.210 ;
        RECT 1369.520 2014.510 1369.780 2014.830 ;
        RECT 1374.580 2014.510 1374.840 2014.830 ;
        RECT 1374.640 2000.000 1374.780 2014.510 ;
        RECT 1374.480 1999.540 1374.780 2000.000 ;
        RECT 1374.480 1996.000 1374.760 1999.540 ;
      LAYER via2 ;
        RECT 16.650 2118.400 16.930 2118.680 ;
      LAYER met3 ;
        RECT -4.800 2118.690 2.400 2119.140 ;
        RECT 16.625 2118.690 16.955 2118.705 ;
        RECT -4.800 2118.390 16.955 2118.690 ;
        RECT -4.800 2117.940 2.400 2118.390 ;
        RECT 16.625 2118.375 16.955 2118.390 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1134.890 2000.460 1135.210 2000.520 ;
        RECT 1382.370 2000.460 1382.690 2000.520 ;
        RECT 1134.890 2000.320 1382.690 2000.460 ;
        RECT 1134.890 2000.260 1135.210 2000.320 ;
        RECT 1382.370 2000.260 1382.690 2000.320 ;
        RECT 14.790 1835.220 15.110 1835.280 ;
        RECT 1134.890 1835.220 1135.210 1835.280 ;
        RECT 14.790 1835.080 1135.210 1835.220 ;
        RECT 14.790 1835.020 15.110 1835.080 ;
        RECT 1134.890 1835.020 1135.210 1835.080 ;
      LAYER via ;
        RECT 1134.920 2000.260 1135.180 2000.520 ;
        RECT 1382.400 2000.260 1382.660 2000.520 ;
        RECT 14.820 1835.020 15.080 1835.280 ;
        RECT 1134.920 1835.020 1135.180 1835.280 ;
      LAYER met2 ;
        RECT 1134.920 2000.230 1135.180 2000.550 ;
        RECT 1382.400 2000.230 1382.660 2000.550 ;
        RECT 1134.980 1835.310 1135.120 2000.230 ;
        RECT 1382.460 2000.000 1382.600 2000.230 ;
        RECT 1382.300 1999.540 1382.600 2000.000 ;
        RECT 1382.300 1996.000 1382.580 1999.540 ;
        RECT 14.820 1834.990 15.080 1835.310 ;
        RECT 1134.920 1834.990 1135.180 1835.310 ;
        RECT 14.880 1831.085 15.020 1834.990 ;
        RECT 14.810 1830.715 15.090 1831.085 ;
      LAYER via2 ;
        RECT 14.810 1830.760 15.090 1831.040 ;
      LAYER met3 ;
        RECT -4.800 1831.050 2.400 1831.500 ;
        RECT 14.785 1831.050 15.115 1831.065 ;
        RECT -4.800 1830.750 15.115 1831.050 ;
        RECT -4.800 1830.300 2.400 1830.750 ;
        RECT 14.785 1830.735 15.115 1830.750 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1169.390 2001.820 1169.710 2001.880 ;
        RECT 2480.390 2001.820 2480.710 2001.880 ;
        RECT 1169.390 2001.680 2480.710 2001.820 ;
        RECT 1169.390 2001.620 1169.710 2001.680 ;
        RECT 2480.390 2001.620 2480.710 2001.680 ;
        RECT 2480.390 676.160 2480.710 676.220 ;
        RECT 2900.830 676.160 2901.150 676.220 ;
        RECT 2480.390 676.020 2901.150 676.160 ;
        RECT 2480.390 675.960 2480.710 676.020 ;
        RECT 2900.830 675.960 2901.150 676.020 ;
      LAYER via ;
        RECT 1169.420 2001.620 1169.680 2001.880 ;
        RECT 2480.420 2001.620 2480.680 2001.880 ;
        RECT 2480.420 675.960 2480.680 676.220 ;
        RECT 2900.860 675.960 2901.120 676.220 ;
      LAYER met2 ;
        RECT 1169.420 2001.590 1169.680 2001.910 ;
        RECT 2480.420 2001.590 2480.680 2001.910 ;
        RECT 1169.480 2000.000 1169.620 2001.590 ;
        RECT 1169.320 1999.540 1169.620 2000.000 ;
        RECT 1169.320 1996.000 1169.600 1999.540 ;
        RECT 2480.480 676.250 2480.620 2001.590 ;
        RECT 2480.420 675.930 2480.680 676.250 ;
        RECT 2900.860 675.930 2901.120 676.250 ;
        RECT 2900.920 674.405 2901.060 675.930 ;
        RECT 2900.850 674.035 2901.130 674.405 ;
      LAYER via2 ;
        RECT 2900.850 674.080 2901.130 674.360 ;
      LAYER met3 ;
        RECT 2900.825 674.370 2901.155 674.385 ;
        RECT 2917.600 674.370 2924.800 674.820 ;
        RECT 2900.825 674.070 2924.800 674.370 ;
        RECT 2900.825 674.055 2901.155 674.070 ;
        RECT 2917.600 673.620 2924.800 674.070 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1065.890 1999.100 1066.210 1999.160 ;
        RECT 1388.350 1999.100 1388.670 1999.160 ;
        RECT 1065.890 1998.960 1388.670 1999.100 ;
        RECT 1065.890 1998.900 1066.210 1998.960 ;
        RECT 1388.350 1998.900 1388.670 1998.960 ;
        RECT 16.630 1545.540 16.950 1545.600 ;
        RECT 1065.890 1545.540 1066.210 1545.600 ;
        RECT 16.630 1545.400 1066.210 1545.540 ;
        RECT 16.630 1545.340 16.950 1545.400 ;
        RECT 1065.890 1545.340 1066.210 1545.400 ;
      LAYER via ;
        RECT 1065.920 1998.900 1066.180 1999.160 ;
        RECT 1388.380 1998.900 1388.640 1999.160 ;
        RECT 16.660 1545.340 16.920 1545.600 ;
        RECT 1065.920 1545.340 1066.180 1545.600 ;
      LAYER met2 ;
        RECT 1065.920 1998.870 1066.180 1999.190 ;
        RECT 1388.380 1998.930 1388.640 1999.190 ;
        RECT 1390.120 1998.930 1390.400 2000.000 ;
        RECT 1388.380 1998.870 1390.400 1998.930 ;
        RECT 1065.980 1545.630 1066.120 1998.870 ;
        RECT 1388.440 1998.790 1390.400 1998.870 ;
        RECT 1390.120 1996.000 1390.400 1998.790 ;
        RECT 16.660 1545.310 16.920 1545.630 ;
        RECT 1065.920 1545.310 1066.180 1545.630 ;
        RECT 16.720 1544.125 16.860 1545.310 ;
        RECT 16.650 1543.755 16.930 1544.125 ;
      LAYER via2 ;
        RECT 16.650 1543.800 16.930 1544.080 ;
      LAYER met3 ;
        RECT -4.800 1544.090 2.400 1544.540 ;
        RECT 16.625 1544.090 16.955 1544.105 ;
        RECT -4.800 1543.790 16.955 1544.090 ;
        RECT -4.800 1543.340 2.400 1543.790 ;
        RECT 16.625 1543.775 16.955 1543.790 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1058.990 2003.520 1059.310 2003.580 ;
        RECT 1398.010 2003.520 1398.330 2003.580 ;
        RECT 1058.990 2003.380 1398.330 2003.520 ;
        RECT 1058.990 2003.320 1059.310 2003.380 ;
        RECT 1398.010 2003.320 1398.330 2003.380 ;
        RECT 17.550 1331.680 17.870 1331.740 ;
        RECT 1058.990 1331.680 1059.310 1331.740 ;
        RECT 17.550 1331.540 1059.310 1331.680 ;
        RECT 17.550 1331.480 17.870 1331.540 ;
        RECT 1058.990 1331.480 1059.310 1331.540 ;
      LAYER via ;
        RECT 1059.020 2003.320 1059.280 2003.580 ;
        RECT 1398.040 2003.320 1398.300 2003.580 ;
        RECT 17.580 1331.480 17.840 1331.740 ;
        RECT 1059.020 1331.480 1059.280 1331.740 ;
      LAYER met2 ;
        RECT 1059.020 2003.290 1059.280 2003.610 ;
        RECT 1398.040 2003.290 1398.300 2003.610 ;
        RECT 1059.080 1331.770 1059.220 2003.290 ;
        RECT 1398.100 2000.000 1398.240 2003.290 ;
        RECT 1397.940 1999.540 1398.240 2000.000 ;
        RECT 1397.940 1996.000 1398.220 1999.540 ;
        RECT 17.580 1331.450 17.840 1331.770 ;
        RECT 1059.020 1331.450 1059.280 1331.770 ;
        RECT 17.640 1328.565 17.780 1331.450 ;
        RECT 17.570 1328.195 17.850 1328.565 ;
      LAYER via2 ;
        RECT 17.570 1328.240 17.850 1328.520 ;
      LAYER met3 ;
        RECT -4.800 1328.530 2.400 1328.980 ;
        RECT 17.545 1328.530 17.875 1328.545 ;
        RECT -4.800 1328.230 17.875 1328.530 ;
        RECT -4.800 1327.780 2.400 1328.230 ;
        RECT 17.545 1328.215 17.875 1328.230 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1045.190 2002.840 1045.510 2002.900 ;
        RECT 1405.830 2002.840 1406.150 2002.900 ;
        RECT 1045.190 2002.700 1406.150 2002.840 ;
        RECT 1045.190 2002.640 1045.510 2002.700 ;
        RECT 1405.830 2002.640 1406.150 2002.700 ;
        RECT 15.710 1117.820 16.030 1117.880 ;
        RECT 1045.190 1117.820 1045.510 1117.880 ;
        RECT 15.710 1117.680 1045.510 1117.820 ;
        RECT 15.710 1117.620 16.030 1117.680 ;
        RECT 1045.190 1117.620 1045.510 1117.680 ;
      LAYER via ;
        RECT 1045.220 2002.640 1045.480 2002.900 ;
        RECT 1405.860 2002.640 1406.120 2002.900 ;
        RECT 15.740 1117.620 16.000 1117.880 ;
        RECT 1045.220 1117.620 1045.480 1117.880 ;
      LAYER met2 ;
        RECT 1045.220 2002.610 1045.480 2002.930 ;
        RECT 1405.860 2002.610 1406.120 2002.930 ;
        RECT 1045.280 1117.910 1045.420 2002.610 ;
        RECT 1405.920 2000.000 1406.060 2002.610 ;
        RECT 1405.760 1999.540 1406.060 2000.000 ;
        RECT 1405.760 1996.000 1406.040 1999.540 ;
        RECT 15.740 1117.590 16.000 1117.910 ;
        RECT 1045.220 1117.590 1045.480 1117.910 ;
        RECT 15.800 1113.005 15.940 1117.590 ;
        RECT 15.730 1112.635 16.010 1113.005 ;
      LAYER via2 ;
        RECT 15.730 1112.680 16.010 1112.960 ;
      LAYER met3 ;
        RECT -4.800 1112.970 2.400 1113.420 ;
        RECT 15.705 1112.970 16.035 1112.985 ;
        RECT -4.800 1112.670 16.035 1112.970 ;
        RECT -4.800 1112.220 2.400 1112.670 ;
        RECT 15.705 1112.655 16.035 1112.670 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1038.290 1997.740 1038.610 1997.800 ;
        RECT 1412.270 1997.740 1412.590 1997.800 ;
        RECT 1038.290 1997.600 1412.590 1997.740 ;
        RECT 1038.290 1997.540 1038.610 1997.600 ;
        RECT 1412.270 1997.540 1412.590 1997.600 ;
        RECT 16.170 903.960 16.490 904.020 ;
        RECT 1038.290 903.960 1038.610 904.020 ;
        RECT 16.170 903.820 1038.610 903.960 ;
        RECT 16.170 903.760 16.490 903.820 ;
        RECT 1038.290 903.760 1038.610 903.820 ;
      LAYER via ;
        RECT 1038.320 1997.540 1038.580 1997.800 ;
        RECT 1412.300 1997.540 1412.560 1997.800 ;
        RECT 16.200 903.760 16.460 904.020 ;
        RECT 1038.320 903.760 1038.580 904.020 ;
      LAYER met2 ;
        RECT 1038.320 1997.510 1038.580 1997.830 ;
        RECT 1412.300 1997.570 1412.560 1997.830 ;
        RECT 1413.580 1997.570 1413.860 2000.000 ;
        RECT 1412.300 1997.510 1413.860 1997.570 ;
        RECT 1038.380 904.050 1038.520 1997.510 ;
        RECT 1412.360 1997.430 1413.860 1997.510 ;
        RECT 1413.580 1996.000 1413.860 1997.430 ;
        RECT 16.200 903.730 16.460 904.050 ;
        RECT 1038.320 903.730 1038.580 904.050 ;
        RECT 16.260 897.445 16.400 903.730 ;
        RECT 16.190 897.075 16.470 897.445 ;
      LAYER via2 ;
        RECT 16.190 897.120 16.470 897.400 ;
      LAYER met3 ;
        RECT -4.800 897.410 2.400 897.860 ;
        RECT 16.165 897.410 16.495 897.425 ;
        RECT -4.800 897.110 16.495 897.410 ;
        RECT -4.800 896.660 2.400 897.110 ;
        RECT 16.165 897.095 16.495 897.110 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1135.350 2005.900 1135.670 2005.960 ;
        RECT 1421.930 2005.900 1422.250 2005.960 ;
        RECT 1135.350 2005.760 1422.250 2005.900 ;
        RECT 1135.350 2005.700 1135.670 2005.760 ;
        RECT 1421.930 2005.700 1422.250 2005.760 ;
        RECT 17.550 682.960 17.870 683.020 ;
        RECT 1135.350 682.960 1135.670 683.020 ;
        RECT 17.550 682.820 1135.670 682.960 ;
        RECT 17.550 682.760 17.870 682.820 ;
        RECT 1135.350 682.760 1135.670 682.820 ;
      LAYER via ;
        RECT 1135.380 2005.700 1135.640 2005.960 ;
        RECT 1421.960 2005.700 1422.220 2005.960 ;
        RECT 17.580 682.760 17.840 683.020 ;
        RECT 1135.380 682.760 1135.640 683.020 ;
      LAYER met2 ;
        RECT 1135.380 2005.670 1135.640 2005.990 ;
        RECT 1421.960 2005.670 1422.220 2005.990 ;
        RECT 1135.440 683.050 1135.580 2005.670 ;
        RECT 1422.020 2000.000 1422.160 2005.670 ;
        RECT 1421.860 1999.540 1422.160 2000.000 ;
        RECT 1421.860 1996.000 1422.140 1999.540 ;
        RECT 17.580 682.730 17.840 683.050 ;
        RECT 1135.380 682.730 1135.640 683.050 ;
        RECT 17.640 681.885 17.780 682.730 ;
        RECT 17.570 681.515 17.850 681.885 ;
      LAYER via2 ;
        RECT 17.570 681.560 17.850 681.840 ;
      LAYER met3 ;
        RECT -4.800 681.850 2.400 682.300 ;
        RECT 17.545 681.850 17.875 681.865 ;
        RECT -4.800 681.550 17.875 681.850 ;
        RECT -4.800 681.100 2.400 681.550 ;
        RECT 17.545 681.535 17.875 681.550 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1399.465 1996.905 1400.095 1997.075 ;
        RECT 1414.185 1996.905 1414.355 1997.755 ;
      LAYER mcon ;
        RECT 1414.185 1997.585 1414.355 1997.755 ;
        RECT 1399.925 1996.905 1400.095 1997.075 ;
      LAYER met1 ;
        RECT 1414.125 1997.740 1414.415 1997.785 ;
        RECT 1427.910 1997.740 1428.230 1997.800 ;
        RECT 1414.125 1997.600 1428.230 1997.740 ;
        RECT 1414.125 1997.555 1414.415 1997.600 ;
        RECT 1427.910 1997.540 1428.230 1997.600 ;
        RECT 1024.490 1997.060 1024.810 1997.120 ;
        RECT 1399.405 1997.060 1399.695 1997.105 ;
        RECT 1024.490 1996.920 1399.695 1997.060 ;
        RECT 1024.490 1996.860 1024.810 1996.920 ;
        RECT 1399.405 1996.875 1399.695 1996.920 ;
        RECT 1399.865 1997.060 1400.155 1997.105 ;
        RECT 1414.125 1997.060 1414.415 1997.105 ;
        RECT 1399.865 1996.920 1414.415 1997.060 ;
        RECT 1399.865 1996.875 1400.155 1996.920 ;
        RECT 1414.125 1996.875 1414.415 1996.920 ;
        RECT 17.550 469.100 17.870 469.160 ;
        RECT 1024.490 469.100 1024.810 469.160 ;
        RECT 17.550 468.960 1024.810 469.100 ;
        RECT 17.550 468.900 17.870 468.960 ;
        RECT 1024.490 468.900 1024.810 468.960 ;
      LAYER via ;
        RECT 1427.940 1997.540 1428.200 1997.800 ;
        RECT 1024.520 1996.860 1024.780 1997.120 ;
        RECT 17.580 468.900 17.840 469.160 ;
        RECT 1024.520 468.900 1024.780 469.160 ;
      LAYER met2 ;
        RECT 1427.940 1997.570 1428.200 1997.830 ;
        RECT 1429.680 1997.570 1429.960 2000.000 ;
        RECT 1427.940 1997.510 1429.960 1997.570 ;
        RECT 1428.000 1997.430 1429.960 1997.510 ;
        RECT 1024.520 1996.830 1024.780 1997.150 ;
        RECT 1024.580 469.190 1024.720 1996.830 ;
        RECT 1429.680 1996.000 1429.960 1997.430 ;
        RECT 17.580 468.870 17.840 469.190 ;
        RECT 1024.520 468.870 1024.780 469.190 ;
        RECT 17.640 466.325 17.780 468.870 ;
        RECT 17.570 465.955 17.850 466.325 ;
      LAYER via2 ;
        RECT 17.570 466.000 17.850 466.280 ;
      LAYER met3 ;
        RECT -4.800 466.290 2.400 466.740 ;
        RECT 17.545 466.290 17.875 466.305 ;
        RECT -4.800 465.990 17.875 466.290 ;
        RECT -4.800 465.540 2.400 465.990 ;
        RECT 17.545 465.975 17.875 465.990 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1127.990 2004.880 1128.310 2004.940 ;
        RECT 1437.570 2004.880 1437.890 2004.940 ;
        RECT 1127.990 2004.740 1437.890 2004.880 ;
        RECT 1127.990 2004.680 1128.310 2004.740 ;
        RECT 1437.570 2004.680 1437.890 2004.740 ;
        RECT 15.250 255.240 15.570 255.300 ;
        RECT 1127.990 255.240 1128.310 255.300 ;
        RECT 15.250 255.100 1128.310 255.240 ;
        RECT 15.250 255.040 15.570 255.100 ;
        RECT 1127.990 255.040 1128.310 255.100 ;
      LAYER via ;
        RECT 1128.020 2004.680 1128.280 2004.940 ;
        RECT 1437.600 2004.680 1437.860 2004.940 ;
        RECT 15.280 255.040 15.540 255.300 ;
        RECT 1128.020 255.040 1128.280 255.300 ;
      LAYER met2 ;
        RECT 1128.020 2004.650 1128.280 2004.970 ;
        RECT 1437.600 2004.650 1437.860 2004.970 ;
        RECT 1128.080 255.330 1128.220 2004.650 ;
        RECT 1437.660 2000.000 1437.800 2004.650 ;
        RECT 1437.500 1999.540 1437.800 2000.000 ;
        RECT 1437.500 1996.000 1437.780 1999.540 ;
        RECT 15.280 255.010 15.540 255.330 ;
        RECT 1128.020 255.010 1128.280 255.330 ;
        RECT 15.340 250.765 15.480 255.010 ;
        RECT 15.270 250.395 15.550 250.765 ;
      LAYER via2 ;
        RECT 15.270 250.440 15.550 250.720 ;
      LAYER met3 ;
        RECT -4.800 250.730 2.400 251.180 ;
        RECT 15.245 250.730 15.575 250.745 ;
        RECT -4.800 250.430 15.575 250.730 ;
        RECT -4.800 249.980 2.400 250.430 ;
        RECT 15.245 250.415 15.575 250.430 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1443.550 1996.520 1443.870 1996.780 ;
        RECT 65.390 1996.040 65.710 1996.100 ;
        RECT 1443.640 1996.040 1443.780 1996.520 ;
        RECT 65.390 1995.900 1443.780 1996.040 ;
        RECT 65.390 1995.840 65.710 1995.900 ;
        RECT 17.090 41.380 17.410 41.440 ;
        RECT 65.390 41.380 65.710 41.440 ;
        RECT 17.090 41.240 65.710 41.380 ;
        RECT 17.090 41.180 17.410 41.240 ;
        RECT 65.390 41.180 65.710 41.240 ;
      LAYER via ;
        RECT 1443.580 1996.520 1443.840 1996.780 ;
        RECT 65.420 1995.840 65.680 1996.100 ;
        RECT 17.120 41.180 17.380 41.440 ;
        RECT 65.420 41.180 65.680 41.440 ;
      LAYER met2 ;
        RECT 1445.320 1996.890 1445.600 2000.000 ;
        RECT 1443.640 1996.810 1445.600 1996.890 ;
        RECT 1443.580 1996.750 1445.600 1996.810 ;
        RECT 1443.580 1996.490 1443.840 1996.750 ;
        RECT 65.420 1995.810 65.680 1996.130 ;
        RECT 1445.320 1996.000 1445.600 1996.750 ;
        RECT 65.480 41.470 65.620 1995.810 ;
        RECT 17.120 41.150 17.380 41.470 ;
        RECT 65.420 41.150 65.680 41.470 ;
        RECT 17.180 35.885 17.320 41.150 ;
        RECT 17.110 35.515 17.390 35.885 ;
      LAYER via2 ;
        RECT 17.110 35.560 17.390 35.840 ;
      LAYER met3 ;
        RECT -4.800 35.850 2.400 36.300 ;
        RECT 17.085 35.850 17.415 35.865 ;
        RECT -4.800 35.550 17.415 35.850 ;
        RECT -4.800 35.100 2.400 35.550 ;
        RECT 17.085 35.535 17.415 35.550 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1177.210 2002.500 1177.530 2002.560 ;
        RECT 1541.990 2002.500 1542.310 2002.560 ;
        RECT 1177.210 2002.360 1542.310 2002.500 ;
        RECT 1177.210 2002.300 1177.530 2002.360 ;
        RECT 1541.990 2002.300 1542.310 2002.360 ;
        RECT 1541.990 910.760 1542.310 910.820 ;
        RECT 2900.830 910.760 2901.150 910.820 ;
        RECT 1541.990 910.620 2901.150 910.760 ;
        RECT 1541.990 910.560 1542.310 910.620 ;
        RECT 2900.830 910.560 2901.150 910.620 ;
      LAYER via ;
        RECT 1177.240 2002.300 1177.500 2002.560 ;
        RECT 1542.020 2002.300 1542.280 2002.560 ;
        RECT 1542.020 910.560 1542.280 910.820 ;
        RECT 2900.860 910.560 2901.120 910.820 ;
      LAYER met2 ;
        RECT 1177.240 2002.270 1177.500 2002.590 ;
        RECT 1542.020 2002.270 1542.280 2002.590 ;
        RECT 1177.300 2000.000 1177.440 2002.270 ;
        RECT 1177.140 1999.540 1177.440 2000.000 ;
        RECT 1177.140 1996.000 1177.420 1999.540 ;
        RECT 1542.080 910.850 1542.220 2002.270 ;
        RECT 1542.020 910.530 1542.280 910.850 ;
        RECT 2900.860 910.530 2901.120 910.850 ;
        RECT 2900.920 909.685 2901.060 910.530 ;
        RECT 2900.850 909.315 2901.130 909.685 ;
      LAYER via2 ;
        RECT 2900.850 909.360 2901.130 909.640 ;
      LAYER met3 ;
        RECT 2900.825 909.650 2901.155 909.665 ;
        RECT 2917.600 909.650 2924.800 910.100 ;
        RECT 2900.825 909.350 2924.800 909.650 ;
        RECT 2900.825 909.335 2901.155 909.350 ;
        RECT 2917.600 908.900 2924.800 909.350 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1297.270 1139.920 1297.590 1139.980 ;
        RECT 1352.010 1139.920 1352.330 1139.980 ;
        RECT 1297.270 1139.780 1352.330 1139.920 ;
        RECT 1297.270 1139.720 1297.590 1139.780 ;
        RECT 1352.010 1139.720 1352.330 1139.780 ;
        RECT 1607.310 1139.580 1607.630 1139.640 ;
        RECT 1615.130 1139.580 1615.450 1139.640 ;
        RECT 1607.310 1139.440 1615.450 1139.580 ;
        RECT 1607.310 1139.380 1607.630 1139.440 ;
        RECT 1615.130 1139.380 1615.450 1139.440 ;
        RECT 1510.710 1139.240 1511.030 1139.300 ;
        RECT 1545.210 1139.240 1545.530 1139.300 ;
        RECT 1510.710 1139.100 1545.530 1139.240 ;
        RECT 1510.710 1139.040 1511.030 1139.100 ;
        RECT 1545.210 1139.040 1545.530 1139.100 ;
        RECT 2186.910 1139.240 2187.230 1139.300 ;
        RECT 2221.410 1139.240 2221.730 1139.300 ;
        RECT 2186.910 1139.100 2221.730 1139.240 ;
        RECT 2186.910 1139.040 2187.230 1139.100 ;
        RECT 2221.410 1139.040 2221.730 1139.100 ;
        RECT 2380.110 1139.240 2380.430 1139.300 ;
        RECT 2414.610 1139.240 2414.930 1139.300 ;
        RECT 2380.110 1139.100 2414.930 1139.240 ;
        RECT 2380.110 1139.040 2380.430 1139.100 ;
        RECT 2414.610 1139.040 2414.930 1139.100 ;
        RECT 2669.910 1139.240 2670.230 1139.300 ;
        RECT 2704.410 1139.240 2704.730 1139.300 ;
        RECT 2669.910 1139.100 2704.730 1139.240 ;
        RECT 2669.910 1139.040 2670.230 1139.100 ;
        RECT 2704.410 1139.040 2704.730 1139.100 ;
        RECT 2766.510 1139.240 2766.830 1139.300 ;
        RECT 2801.010 1139.240 2801.330 1139.300 ;
        RECT 2766.510 1139.100 2801.330 1139.240 ;
        RECT 2766.510 1139.040 2766.830 1139.100 ;
        RECT 2801.010 1139.040 2801.330 1139.100 ;
        RECT 2863.110 1139.240 2863.430 1139.300 ;
        RECT 2897.610 1139.240 2897.930 1139.300 ;
        RECT 2863.110 1139.100 2897.930 1139.240 ;
        RECT 2863.110 1139.040 2863.430 1139.100 ;
        RECT 2897.610 1139.040 2897.930 1139.100 ;
      LAYER via ;
        RECT 1297.300 1139.720 1297.560 1139.980 ;
        RECT 1352.040 1139.720 1352.300 1139.980 ;
        RECT 1607.340 1139.380 1607.600 1139.640 ;
        RECT 1615.160 1139.380 1615.420 1139.640 ;
        RECT 1510.740 1139.040 1511.000 1139.300 ;
        RECT 1545.240 1139.040 1545.500 1139.300 ;
        RECT 2186.940 1139.040 2187.200 1139.300 ;
        RECT 2221.440 1139.040 2221.700 1139.300 ;
        RECT 2380.140 1139.040 2380.400 1139.300 ;
        RECT 2414.640 1139.040 2414.900 1139.300 ;
        RECT 2669.940 1139.040 2670.200 1139.300 ;
        RECT 2704.440 1139.040 2704.700 1139.300 ;
        RECT 2766.540 1139.040 2766.800 1139.300 ;
        RECT 2801.040 1139.040 2801.300 1139.300 ;
        RECT 2863.140 1139.040 2863.400 1139.300 ;
        RECT 2897.640 1139.040 2897.900 1139.300 ;
      LAYER met2 ;
        RECT 1184.960 1996.890 1185.240 2000.000 ;
        RECT 1185.970 1996.890 1186.250 1997.005 ;
        RECT 1184.960 1996.750 1186.250 1996.890 ;
        RECT 1184.960 1996.000 1185.240 1996.750 ;
        RECT 1185.970 1996.635 1186.250 1996.750 ;
        RECT 1220.930 1140.515 1221.210 1140.885 ;
        RECT 1221.000 1140.090 1221.140 1140.515 ;
        RECT 1221.850 1140.090 1222.130 1140.205 ;
        RECT 1221.000 1139.950 1222.130 1140.090 ;
        RECT 1221.850 1139.835 1222.130 1139.950 ;
        RECT 1242.090 1139.835 1242.370 1140.205 ;
        RECT 1297.290 1139.835 1297.570 1140.205 ;
        RECT 1242.160 1138.165 1242.300 1139.835 ;
        RECT 1297.300 1139.690 1297.560 1139.835 ;
        RECT 1352.040 1139.690 1352.300 1140.010 ;
        RECT 1352.100 1139.525 1352.240 1139.690 ;
        RECT 1607.340 1139.525 1607.600 1139.670 ;
        RECT 1615.160 1139.525 1615.420 1139.670 ;
        RECT 1352.030 1139.155 1352.310 1139.525 ;
        RECT 1510.730 1139.155 1511.010 1139.525 ;
        RECT 1510.740 1139.010 1511.000 1139.155 ;
        RECT 1545.240 1139.010 1545.500 1139.330 ;
        RECT 1607.330 1139.155 1607.610 1139.525 ;
        RECT 1615.150 1139.155 1615.430 1139.525 ;
        RECT 2076.530 1139.155 2076.810 1139.525 ;
        RECT 2186.930 1139.155 2187.210 1139.525 ;
        RECT 2283.530 1139.410 2283.810 1139.525 ;
        RECT 2284.450 1139.410 2284.730 1139.525 ;
        RECT 1545.300 1138.845 1545.440 1139.010 ;
        RECT 2076.600 1138.845 2076.740 1139.155 ;
        RECT 2186.940 1139.010 2187.200 1139.155 ;
        RECT 2221.440 1139.010 2221.700 1139.330 ;
        RECT 2283.530 1139.270 2284.730 1139.410 ;
        RECT 2283.530 1139.155 2283.810 1139.270 ;
        RECT 2284.450 1139.155 2284.730 1139.270 ;
        RECT 2380.130 1139.155 2380.410 1139.525 ;
        RECT 2380.140 1139.010 2380.400 1139.155 ;
        RECT 2414.640 1139.010 2414.900 1139.330 ;
        RECT 2669.930 1139.155 2670.210 1139.525 ;
        RECT 2669.940 1139.010 2670.200 1139.155 ;
        RECT 2704.440 1139.010 2704.700 1139.330 ;
        RECT 2766.530 1139.155 2766.810 1139.525 ;
        RECT 2766.540 1139.010 2766.800 1139.155 ;
        RECT 2801.040 1139.010 2801.300 1139.330 ;
        RECT 2863.130 1139.155 2863.410 1139.525 ;
        RECT 2863.140 1139.010 2863.400 1139.155 ;
        RECT 2897.640 1139.010 2897.900 1139.330 ;
        RECT 2221.500 1138.845 2221.640 1139.010 ;
        RECT 2414.700 1138.845 2414.840 1139.010 ;
        RECT 2704.500 1138.845 2704.640 1139.010 ;
        RECT 2801.100 1138.845 2801.240 1139.010 ;
        RECT 2897.700 1138.845 2897.840 1139.010 ;
        RECT 1545.230 1138.475 1545.510 1138.845 ;
        RECT 2076.530 1138.475 2076.810 1138.845 ;
        RECT 2221.430 1138.475 2221.710 1138.845 ;
        RECT 2414.630 1138.475 2414.910 1138.845 ;
        RECT 2704.430 1138.475 2704.710 1138.845 ;
        RECT 2801.030 1138.475 2801.310 1138.845 ;
        RECT 2897.630 1138.475 2897.910 1138.845 ;
        RECT 1242.090 1137.795 1242.370 1138.165 ;
      LAYER via2 ;
        RECT 1185.970 1996.680 1186.250 1996.960 ;
        RECT 1220.930 1140.560 1221.210 1140.840 ;
        RECT 1221.850 1139.880 1222.130 1140.160 ;
        RECT 1242.090 1139.880 1242.370 1140.160 ;
        RECT 1297.290 1139.880 1297.570 1140.160 ;
        RECT 1352.030 1139.200 1352.310 1139.480 ;
        RECT 1510.730 1139.200 1511.010 1139.480 ;
        RECT 1607.330 1139.200 1607.610 1139.480 ;
        RECT 1615.150 1139.200 1615.430 1139.480 ;
        RECT 2076.530 1139.200 2076.810 1139.480 ;
        RECT 2186.930 1139.200 2187.210 1139.480 ;
        RECT 2283.530 1139.200 2283.810 1139.480 ;
        RECT 2284.450 1139.200 2284.730 1139.480 ;
        RECT 2380.130 1139.200 2380.410 1139.480 ;
        RECT 2669.930 1139.200 2670.210 1139.480 ;
        RECT 2766.530 1139.200 2766.810 1139.480 ;
        RECT 2863.130 1139.200 2863.410 1139.480 ;
        RECT 1545.230 1138.520 1545.510 1138.800 ;
        RECT 2076.530 1138.520 2076.810 1138.800 ;
        RECT 2221.430 1138.520 2221.710 1138.800 ;
        RECT 2414.630 1138.520 2414.910 1138.800 ;
        RECT 2704.430 1138.520 2704.710 1138.800 ;
        RECT 2801.030 1138.520 2801.310 1138.800 ;
        RECT 2897.630 1138.520 2897.910 1138.800 ;
        RECT 1242.090 1137.840 1242.370 1138.120 ;
      LAYER met3 ;
        RECT 1185.945 1996.980 1186.275 1996.985 ;
        RECT 1185.945 1996.970 1186.530 1996.980 ;
        RECT 1185.945 1996.670 1186.730 1996.970 ;
        RECT 1185.945 1996.660 1186.530 1996.670 ;
        RECT 1185.945 1996.655 1186.275 1996.660 ;
        RECT 2917.600 1144.250 2924.800 1144.700 ;
        RECT 2916.710 1143.950 2924.800 1144.250 ;
        RECT 1186.150 1140.850 1186.530 1140.860 ;
        RECT 1220.905 1140.850 1221.235 1140.865 ;
        RECT 1186.150 1140.550 1221.235 1140.850 ;
        RECT 1186.150 1140.540 1186.530 1140.550 ;
        RECT 1220.905 1140.535 1221.235 1140.550 ;
        RECT 1221.825 1140.170 1222.155 1140.185 ;
        RECT 1242.065 1140.170 1242.395 1140.185 ;
        RECT 1221.825 1139.870 1242.395 1140.170 ;
        RECT 1221.825 1139.855 1222.155 1139.870 ;
        RECT 1242.065 1139.855 1242.395 1139.870 ;
        RECT 1289.190 1140.170 1289.570 1140.180 ;
        RECT 1297.265 1140.170 1297.595 1140.185 ;
        RECT 1289.190 1139.870 1297.595 1140.170 ;
        RECT 1289.190 1139.860 1289.570 1139.870 ;
        RECT 1297.265 1139.855 1297.595 1139.870 ;
        RECT 1366.510 1139.870 1414.650 1140.170 ;
        RECT 1352.005 1139.490 1352.335 1139.505 ;
        RECT 1366.510 1139.490 1366.810 1139.870 ;
        RECT 1352.005 1139.190 1366.810 1139.490 ;
        RECT 1352.005 1139.175 1352.335 1139.190 ;
        RECT 1414.350 1138.810 1414.650 1139.870 ;
        RECT 1676.550 1139.870 1724.690 1140.170 ;
        RECT 1510.705 1139.490 1511.035 1139.505 ;
        RECT 1607.305 1139.490 1607.635 1139.505 ;
        RECT 1463.110 1139.190 1511.035 1139.490 ;
        RECT 1463.110 1138.810 1463.410 1139.190 ;
        RECT 1510.705 1139.175 1511.035 1139.190 ;
        RECT 1559.710 1139.190 1607.635 1139.490 ;
        RECT 1414.350 1138.510 1463.410 1138.810 ;
        RECT 1545.205 1138.810 1545.535 1138.825 ;
        RECT 1559.710 1138.810 1560.010 1139.190 ;
        RECT 1607.305 1139.175 1607.635 1139.190 ;
        RECT 1615.125 1139.490 1615.455 1139.505 ;
        RECT 1615.125 1139.190 1655.690 1139.490 ;
        RECT 1615.125 1139.175 1615.455 1139.190 ;
        RECT 1545.205 1138.510 1560.010 1138.810 ;
        RECT 1655.390 1138.810 1655.690 1139.190 ;
        RECT 1676.550 1138.810 1676.850 1139.870 ;
        RECT 1655.390 1138.510 1676.850 1138.810 ;
        RECT 1724.390 1138.810 1724.690 1139.870 ;
        RECT 1725.310 1139.870 1773.450 1140.170 ;
        RECT 1725.310 1138.810 1725.610 1139.870 ;
        RECT 1773.150 1139.490 1773.450 1139.870 ;
        RECT 1821.910 1139.870 1870.050 1140.170 ;
        RECT 1773.150 1139.190 1821.290 1139.490 ;
        RECT 1724.390 1138.510 1725.610 1138.810 ;
        RECT 1820.990 1138.810 1821.290 1139.190 ;
        RECT 1821.910 1138.810 1822.210 1139.870 ;
        RECT 1869.750 1139.490 1870.050 1139.870 ;
        RECT 1918.510 1139.870 2029.210 1140.170 ;
        RECT 1869.750 1139.190 1917.890 1139.490 ;
        RECT 1820.990 1138.510 1822.210 1138.810 ;
        RECT 1917.590 1138.810 1917.890 1139.190 ;
        RECT 1918.510 1138.810 1918.810 1139.870 ;
        RECT 2028.910 1139.490 2029.210 1139.870 ;
        RECT 2476.950 1139.870 2573.850 1140.170 ;
        RECT 2076.505 1139.490 2076.835 1139.505 ;
        RECT 2186.905 1139.490 2187.235 1139.505 ;
        RECT 2283.505 1139.490 2283.835 1139.505 ;
        RECT 2028.910 1139.190 2076.835 1139.490 ;
        RECT 2076.505 1139.175 2076.835 1139.190 ;
        RECT 2139.310 1139.190 2187.235 1139.490 ;
        RECT 1917.590 1138.510 1918.810 1138.810 ;
        RECT 2076.505 1138.810 2076.835 1138.825 ;
        RECT 2139.310 1138.810 2139.610 1139.190 ;
        RECT 2186.905 1139.175 2187.235 1139.190 ;
        RECT 2235.910 1139.190 2283.835 1139.490 ;
        RECT 2076.505 1138.510 2139.610 1138.810 ;
        RECT 2221.405 1138.810 2221.735 1138.825 ;
        RECT 2235.910 1138.810 2236.210 1139.190 ;
        RECT 2283.505 1139.175 2283.835 1139.190 ;
        RECT 2284.425 1139.490 2284.755 1139.505 ;
        RECT 2380.105 1139.490 2380.435 1139.505 ;
        RECT 2284.425 1139.190 2331.890 1139.490 ;
        RECT 2284.425 1139.175 2284.755 1139.190 ;
        RECT 2221.405 1138.510 2236.210 1138.810 ;
        RECT 2331.590 1138.810 2331.890 1139.190 ;
        RECT 2332.510 1139.190 2380.435 1139.490 ;
        RECT 2332.510 1138.810 2332.810 1139.190 ;
        RECT 2380.105 1139.175 2380.435 1139.190 ;
        RECT 2331.590 1138.510 2332.810 1138.810 ;
        RECT 2414.605 1138.810 2414.935 1138.825 ;
        RECT 2476.950 1138.810 2477.250 1139.870 ;
        RECT 2414.605 1138.510 2477.250 1138.810 ;
        RECT 2573.550 1138.810 2573.850 1139.870 ;
        RECT 2669.905 1139.490 2670.235 1139.505 ;
        RECT 2766.505 1139.490 2766.835 1139.505 ;
        RECT 2863.105 1139.490 2863.435 1139.505 ;
        RECT 2622.310 1139.190 2670.235 1139.490 ;
        RECT 2622.310 1138.810 2622.610 1139.190 ;
        RECT 2669.905 1139.175 2670.235 1139.190 ;
        RECT 2718.910 1139.190 2766.835 1139.490 ;
        RECT 2573.550 1138.510 2622.610 1138.810 ;
        RECT 2704.405 1138.810 2704.735 1138.825 ;
        RECT 2718.910 1138.810 2719.210 1139.190 ;
        RECT 2766.505 1139.175 2766.835 1139.190 ;
        RECT 2815.510 1139.190 2863.435 1139.490 ;
        RECT 2704.405 1138.510 2719.210 1138.810 ;
        RECT 2801.005 1138.810 2801.335 1138.825 ;
        RECT 2815.510 1138.810 2815.810 1139.190 ;
        RECT 2863.105 1139.175 2863.435 1139.190 ;
        RECT 2801.005 1138.510 2815.810 1138.810 ;
        RECT 2897.605 1138.810 2897.935 1138.825 ;
        RECT 2916.710 1138.810 2917.010 1143.950 ;
        RECT 2917.600 1143.500 2924.800 1143.950 ;
        RECT 2897.605 1138.510 2917.010 1138.810 ;
        RECT 1545.205 1138.495 1545.535 1138.510 ;
        RECT 2076.505 1138.495 2076.835 1138.510 ;
        RECT 2221.405 1138.495 2221.735 1138.510 ;
        RECT 2414.605 1138.495 2414.935 1138.510 ;
        RECT 2704.405 1138.495 2704.735 1138.510 ;
        RECT 2801.005 1138.495 2801.335 1138.510 ;
        RECT 2897.605 1138.495 2897.935 1138.510 ;
        RECT 1242.065 1138.130 1242.395 1138.145 ;
        RECT 1289.190 1138.130 1289.570 1138.140 ;
        RECT 1242.065 1137.830 1289.570 1138.130 ;
        RECT 1242.065 1137.815 1242.395 1137.830 ;
        RECT 1289.190 1137.820 1289.570 1137.830 ;
      LAYER via3 ;
        RECT 1186.180 1996.660 1186.500 1996.980 ;
        RECT 1186.180 1140.540 1186.500 1140.860 ;
        RECT 1289.220 1139.860 1289.540 1140.180 ;
        RECT 1289.220 1137.820 1289.540 1138.140 ;
      LAYER met4 ;
        RECT 1186.175 1996.655 1186.505 1996.985 ;
        RECT 1186.190 1140.865 1186.490 1996.655 ;
        RECT 1186.175 1140.535 1186.505 1140.865 ;
        RECT 1289.215 1139.855 1289.545 1140.185 ;
        RECT 1289.230 1138.145 1289.530 1139.855 ;
        RECT 1289.215 1137.815 1289.545 1138.145 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1220.985 1996.225 1221.155 2000.815 ;
        RECT 1269.745 1996.225 1269.915 2000.815 ;
        RECT 1317.585 1996.225 1317.755 2000.815 ;
        RECT 1399.005 1997.245 1400.555 1997.415 ;
        RECT 1399.005 1996.225 1399.175 1997.245 ;
        RECT 1400.845 1996.225 1401.015 1997.415 ;
        RECT 1449.145 1996.905 1449.315 1997.755 ;
        RECT 1496.985 1995.885 1497.155 1997.755 ;
        RECT 1690.645 1997.245 1690.815 1998.095 ;
        RECT 1655.685 1996.905 1656.315 1997.075 ;
        RECT 1738.485 1996.905 1738.655 1998.095 ;
        RECT 1787.245 1997.245 1787.415 1998.095 ;
        RECT 1752.285 1996.905 1752.915 1997.075 ;
        RECT 1835.085 1996.905 1835.255 1998.095 ;
        RECT 1883.845 1997.245 1884.015 1998.095 ;
        RECT 1848.885 1996.905 1849.515 1997.075 ;
        RECT 1931.685 1996.905 1931.855 1998.095 ;
        RECT 1545.745 1995.205 1545.915 1996.055 ;
        RECT 1593.585 1995.205 1593.755 1996.395 ;
        RECT 1934.905 1990.785 1935.075 1997.075 ;
      LAYER mcon ;
        RECT 1220.985 2000.645 1221.155 2000.815 ;
        RECT 1269.745 2000.645 1269.915 2000.815 ;
        RECT 1317.585 2000.645 1317.755 2000.815 ;
        RECT 1690.645 1997.925 1690.815 1998.095 ;
        RECT 1449.145 1997.585 1449.315 1997.755 ;
        RECT 1400.385 1997.245 1400.555 1997.415 ;
        RECT 1400.845 1997.245 1401.015 1997.415 ;
        RECT 1496.985 1997.585 1497.155 1997.755 ;
        RECT 1738.485 1997.925 1738.655 1998.095 ;
        RECT 1787.245 1997.925 1787.415 1998.095 ;
        RECT 1835.085 1997.925 1835.255 1998.095 ;
        RECT 1883.845 1997.925 1884.015 1998.095 ;
        RECT 1931.685 1997.925 1931.855 1998.095 ;
        RECT 1656.145 1996.905 1656.315 1997.075 ;
        RECT 1752.745 1996.905 1752.915 1997.075 ;
        RECT 1849.345 1996.905 1849.515 1997.075 ;
        RECT 1934.905 1996.905 1935.075 1997.075 ;
        RECT 1593.585 1996.225 1593.755 1996.395 ;
        RECT 1545.745 1995.885 1545.915 1996.055 ;
      LAYER met1 ;
        RECT 1192.850 2000.800 1193.170 2000.860 ;
        RECT 1220.925 2000.800 1221.215 2000.845 ;
        RECT 1192.850 2000.660 1221.215 2000.800 ;
        RECT 1192.850 2000.600 1193.170 2000.660 ;
        RECT 1220.925 2000.615 1221.215 2000.660 ;
        RECT 1269.685 2000.800 1269.975 2000.845 ;
        RECT 1317.525 2000.800 1317.815 2000.845 ;
        RECT 1269.685 2000.660 1317.815 2000.800 ;
        RECT 1269.685 2000.615 1269.975 2000.660 ;
        RECT 1317.525 2000.615 1317.815 2000.660 ;
        RECT 1690.585 1998.080 1690.875 1998.125 ;
        RECT 1738.425 1998.080 1738.715 1998.125 ;
        RECT 1690.585 1997.940 1738.715 1998.080 ;
        RECT 1690.585 1997.895 1690.875 1997.940 ;
        RECT 1738.425 1997.895 1738.715 1997.940 ;
        RECT 1787.185 1998.080 1787.475 1998.125 ;
        RECT 1835.025 1998.080 1835.315 1998.125 ;
        RECT 1787.185 1997.940 1835.315 1998.080 ;
        RECT 1787.185 1997.895 1787.475 1997.940 ;
        RECT 1835.025 1997.895 1835.315 1997.940 ;
        RECT 1883.785 1998.080 1884.075 1998.125 ;
        RECT 1931.625 1998.080 1931.915 1998.125 ;
        RECT 1883.785 1997.940 1931.915 1998.080 ;
        RECT 1883.785 1997.895 1884.075 1997.940 ;
        RECT 1931.625 1997.895 1931.915 1997.940 ;
        RECT 1449.085 1997.740 1449.375 1997.785 ;
        RECT 1496.925 1997.740 1497.215 1997.785 ;
        RECT 1449.085 1997.600 1497.215 1997.740 ;
        RECT 1449.085 1997.555 1449.375 1997.600 ;
        RECT 1496.925 1997.555 1497.215 1997.600 ;
        RECT 1400.325 1997.400 1400.615 1997.445 ;
        RECT 1400.785 1997.400 1401.075 1997.445 ;
        RECT 1690.585 1997.400 1690.875 1997.445 ;
        RECT 1787.185 1997.400 1787.475 1997.445 ;
        RECT 1883.785 1997.400 1884.075 1997.445 ;
        RECT 1400.325 1997.260 1401.075 1997.400 ;
        RECT 1400.325 1997.215 1400.615 1997.260 ;
        RECT 1400.785 1997.215 1401.075 1997.260 ;
        RECT 1662.140 1997.260 1690.875 1997.400 ;
        RECT 1449.085 1997.060 1449.375 1997.105 ;
        RECT 1655.625 1997.060 1655.915 1997.105 ;
        RECT 1429.380 1996.920 1449.375 1997.060 ;
        RECT 1220.925 1996.380 1221.215 1996.425 ;
        RECT 1269.685 1996.380 1269.975 1996.425 ;
        RECT 1220.925 1996.240 1269.975 1996.380 ;
        RECT 1220.925 1996.195 1221.215 1996.240 ;
        RECT 1269.685 1996.195 1269.975 1996.240 ;
        RECT 1317.525 1996.380 1317.815 1996.425 ;
        RECT 1398.945 1996.380 1399.235 1996.425 ;
        RECT 1317.525 1996.240 1399.235 1996.380 ;
        RECT 1317.525 1996.195 1317.815 1996.240 ;
        RECT 1398.945 1996.195 1399.235 1996.240 ;
        RECT 1400.785 1996.380 1401.075 1996.425 ;
        RECT 1429.380 1996.380 1429.520 1996.920 ;
        RECT 1449.085 1996.875 1449.375 1996.920 ;
        RECT 1607.400 1996.920 1655.915 1997.060 ;
        RECT 1400.785 1996.240 1429.520 1996.380 ;
        RECT 1593.525 1996.380 1593.815 1996.425 ;
        RECT 1607.400 1996.380 1607.540 1996.920 ;
        RECT 1655.625 1996.875 1655.915 1996.920 ;
        RECT 1656.085 1997.060 1656.375 1997.105 ;
        RECT 1662.140 1997.060 1662.280 1997.260 ;
        RECT 1690.585 1997.215 1690.875 1997.260 ;
        RECT 1758.740 1997.260 1787.475 1997.400 ;
        RECT 1656.085 1996.920 1662.280 1997.060 ;
        RECT 1738.425 1997.060 1738.715 1997.105 ;
        RECT 1752.225 1997.060 1752.515 1997.105 ;
        RECT 1738.425 1996.920 1752.515 1997.060 ;
        RECT 1656.085 1996.875 1656.375 1996.920 ;
        RECT 1738.425 1996.875 1738.715 1996.920 ;
        RECT 1752.225 1996.875 1752.515 1996.920 ;
        RECT 1752.685 1997.060 1752.975 1997.105 ;
        RECT 1758.740 1997.060 1758.880 1997.260 ;
        RECT 1787.185 1997.215 1787.475 1997.260 ;
        RECT 1855.340 1997.260 1884.075 1997.400 ;
        RECT 1752.685 1996.920 1758.880 1997.060 ;
        RECT 1835.025 1997.060 1835.315 1997.105 ;
        RECT 1848.825 1997.060 1849.115 1997.105 ;
        RECT 1835.025 1996.920 1849.115 1997.060 ;
        RECT 1752.685 1996.875 1752.975 1996.920 ;
        RECT 1835.025 1996.875 1835.315 1996.920 ;
        RECT 1848.825 1996.875 1849.115 1996.920 ;
        RECT 1849.285 1997.060 1849.575 1997.105 ;
        RECT 1855.340 1997.060 1855.480 1997.260 ;
        RECT 1883.785 1997.215 1884.075 1997.260 ;
        RECT 1849.285 1996.920 1855.480 1997.060 ;
        RECT 1931.625 1997.060 1931.915 1997.105 ;
        RECT 1934.845 1997.060 1935.135 1997.105 ;
        RECT 1931.625 1996.920 1935.135 1997.060 ;
        RECT 1849.285 1996.875 1849.575 1996.920 ;
        RECT 1931.625 1996.875 1931.915 1996.920 ;
        RECT 1934.845 1996.875 1935.135 1996.920 ;
        RECT 1593.525 1996.240 1607.540 1996.380 ;
        RECT 1400.785 1996.195 1401.075 1996.240 ;
        RECT 1593.525 1996.195 1593.815 1996.240 ;
        RECT 1496.925 1996.040 1497.215 1996.085 ;
        RECT 1545.685 1996.040 1545.975 1996.085 ;
        RECT 1496.925 1995.900 1545.975 1996.040 ;
        RECT 1496.925 1995.855 1497.215 1995.900 ;
        RECT 1545.685 1995.855 1545.975 1995.900 ;
        RECT 1545.685 1995.360 1545.975 1995.405 ;
        RECT 1593.525 1995.360 1593.815 1995.405 ;
        RECT 1545.685 1995.220 1593.815 1995.360 ;
        RECT 1545.685 1995.175 1545.975 1995.220 ;
        RECT 1593.525 1995.175 1593.815 1995.220 ;
        RECT 1934.845 1990.940 1935.135 1990.985 ;
        RECT 1969.790 1990.940 1970.110 1991.000 ;
        RECT 1934.845 1990.800 1970.110 1990.940 ;
        RECT 1934.845 1990.755 1935.135 1990.800 ;
        RECT 1969.790 1990.740 1970.110 1990.800 ;
        RECT 1969.790 1379.960 1970.110 1380.020 ;
        RECT 2900.830 1379.960 2901.150 1380.020 ;
        RECT 1969.790 1379.820 2901.150 1379.960 ;
        RECT 1969.790 1379.760 1970.110 1379.820 ;
        RECT 2900.830 1379.760 2901.150 1379.820 ;
      LAYER via ;
        RECT 1192.880 2000.600 1193.140 2000.860 ;
        RECT 1969.820 1990.740 1970.080 1991.000 ;
        RECT 1969.820 1379.760 1970.080 1380.020 ;
        RECT 2900.860 1379.760 2901.120 1380.020 ;
      LAYER met2 ;
        RECT 1192.880 2000.570 1193.140 2000.890 ;
        RECT 1192.940 2000.000 1193.080 2000.570 ;
        RECT 1192.780 1999.540 1193.080 2000.000 ;
        RECT 1192.780 1996.000 1193.060 1999.540 ;
        RECT 1969.820 1990.710 1970.080 1991.030 ;
        RECT 1969.880 1380.050 1970.020 1990.710 ;
        RECT 1969.820 1379.730 1970.080 1380.050 ;
        RECT 2900.860 1379.730 2901.120 1380.050 ;
        RECT 2900.920 1378.885 2901.060 1379.730 ;
        RECT 2900.850 1378.515 2901.130 1378.885 ;
      LAYER via2 ;
        RECT 2900.850 1378.560 2901.130 1378.840 ;
      LAYER met3 ;
        RECT 2900.825 1378.850 2901.155 1378.865 ;
        RECT 2917.600 1378.850 2924.800 1379.300 ;
        RECT 2900.825 1378.550 2924.800 1378.850 ;
        RECT 2900.825 1378.535 2901.155 1378.550 ;
        RECT 2917.600 1378.100 2924.800 1378.550 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1448.150 1608.780 1448.470 1608.840 ;
        RECT 1490.010 1608.780 1490.330 1608.840 ;
        RECT 1448.150 1608.640 1490.330 1608.780 ;
        RECT 1448.150 1608.580 1448.470 1608.640 ;
        RECT 1490.010 1608.580 1490.330 1608.640 ;
        RECT 1897.110 1608.780 1897.430 1608.840 ;
        RECT 1931.610 1608.780 1931.930 1608.840 ;
        RECT 1897.110 1608.640 1931.930 1608.780 ;
        RECT 1897.110 1608.580 1897.430 1608.640 ;
        RECT 1931.610 1608.580 1931.930 1608.640 ;
      LAYER via ;
        RECT 1448.180 1608.580 1448.440 1608.840 ;
        RECT 1490.040 1608.580 1490.300 1608.840 ;
        RECT 1897.140 1608.580 1897.400 1608.840 ;
        RECT 1931.640 1608.580 1931.900 1608.840 ;
      LAYER met2 ;
        RECT 1200.600 1997.570 1200.880 2000.000 ;
        RECT 1201.610 1997.570 1201.890 1997.685 ;
        RECT 1200.600 1997.430 1201.890 1997.570 ;
        RECT 1200.600 1996.000 1200.880 1997.430 ;
        RECT 1201.610 1997.315 1201.890 1997.430 ;
        RECT 1545.230 1610.395 1545.510 1610.765 ;
        RECT 1811.110 1610.395 1811.390 1610.765 ;
        RECT 2004.310 1610.395 2004.590 1610.765 ;
        RECT 1545.300 1609.405 1545.440 1610.395 ;
        RECT 1811.180 1609.405 1811.320 1610.395 ;
        RECT 2004.380 1609.405 2004.520 1610.395 ;
        RECT 1545.230 1609.035 1545.510 1609.405 ;
        RECT 1608.250 1609.035 1608.530 1609.405 ;
        RECT 1704.850 1609.035 1705.130 1609.405 ;
        RECT 1811.110 1609.035 1811.390 1609.405 ;
        RECT 1931.630 1609.035 1931.910 1609.405 ;
        RECT 2004.310 1609.035 2004.590 1609.405 ;
        RECT 2091.250 1609.035 2091.530 1609.405 ;
        RECT 2187.850 1609.035 2188.130 1609.405 ;
        RECT 2284.450 1609.035 2284.730 1609.405 ;
        RECT 2381.050 1609.035 2381.330 1609.405 ;
        RECT 2476.730 1609.290 2477.010 1609.405 ;
        RECT 2477.650 1609.290 2477.930 1609.405 ;
        RECT 2476.730 1609.150 2477.930 1609.290 ;
        RECT 2476.730 1609.035 2477.010 1609.150 ;
        RECT 2477.650 1609.035 2477.930 1609.150 ;
        RECT 2573.330 1609.290 2573.610 1609.405 ;
        RECT 2574.250 1609.290 2574.530 1609.405 ;
        RECT 2573.330 1609.150 2574.530 1609.290 ;
        RECT 2573.330 1609.035 2573.610 1609.150 ;
        RECT 2574.250 1609.035 2574.530 1609.150 ;
        RECT 2669.930 1609.290 2670.210 1609.405 ;
        RECT 2670.850 1609.290 2671.130 1609.405 ;
        RECT 2669.930 1609.150 2671.130 1609.290 ;
        RECT 2669.930 1609.035 2670.210 1609.150 ;
        RECT 2670.850 1609.035 2671.130 1609.150 ;
        RECT 2863.130 1609.035 2863.410 1609.405 ;
        RECT 1425.170 1608.355 1425.450 1608.725 ;
        RECT 1448.180 1608.550 1448.440 1608.870 ;
        RECT 1490.040 1608.725 1490.300 1608.870 ;
        RECT 1425.240 1607.365 1425.380 1608.355 ;
        RECT 1448.240 1607.365 1448.380 1608.550 ;
        RECT 1490.030 1608.355 1490.310 1608.725 ;
        RECT 1607.330 1608.610 1607.610 1608.725 ;
        RECT 1608.320 1608.610 1608.460 1609.035 ;
        RECT 1607.330 1608.470 1608.460 1608.610 ;
        RECT 1703.930 1608.610 1704.210 1608.725 ;
        RECT 1704.920 1608.610 1705.060 1609.035 ;
        RECT 1931.700 1608.870 1931.840 1609.035 ;
        RECT 1897.140 1608.725 1897.400 1608.870 ;
        RECT 1703.930 1608.470 1705.060 1608.610 ;
        RECT 1607.330 1608.355 1607.610 1608.470 ;
        RECT 1703.930 1608.355 1704.210 1608.470 ;
        RECT 1897.130 1608.355 1897.410 1608.725 ;
        RECT 1931.640 1608.550 1931.900 1608.870 ;
        RECT 2090.330 1608.610 2090.610 1608.725 ;
        RECT 2091.320 1608.610 2091.460 1609.035 ;
        RECT 2090.330 1608.470 2091.460 1608.610 ;
        RECT 2186.930 1608.610 2187.210 1608.725 ;
        RECT 2187.920 1608.610 2188.060 1609.035 ;
        RECT 2186.930 1608.470 2188.060 1608.610 ;
        RECT 2283.530 1608.610 2283.810 1608.725 ;
        RECT 2284.520 1608.610 2284.660 1609.035 ;
        RECT 2283.530 1608.470 2284.660 1608.610 ;
        RECT 2380.130 1608.610 2380.410 1608.725 ;
        RECT 2381.120 1608.610 2381.260 1609.035 ;
        RECT 2380.130 1608.470 2381.260 1608.610 ;
        RECT 2814.370 1608.610 2814.650 1608.725 ;
        RECT 2815.750 1608.610 2816.030 1608.725 ;
        RECT 2814.370 1608.470 2816.030 1608.610 ;
        RECT 2863.200 1608.610 2863.340 1609.035 ;
        RECT 2863.590 1608.610 2863.870 1608.725 ;
        RECT 2863.200 1608.470 2863.870 1608.610 ;
        RECT 2090.330 1608.355 2090.610 1608.470 ;
        RECT 2186.930 1608.355 2187.210 1608.470 ;
        RECT 2283.530 1608.355 2283.810 1608.470 ;
        RECT 2380.130 1608.355 2380.410 1608.470 ;
        RECT 2814.370 1608.355 2814.650 1608.470 ;
        RECT 2815.750 1608.355 2816.030 1608.470 ;
        RECT 2863.590 1608.355 2863.870 1608.470 ;
        RECT 1425.170 1606.995 1425.450 1607.365 ;
        RECT 1448.170 1606.995 1448.450 1607.365 ;
      LAYER via2 ;
        RECT 1201.610 1997.360 1201.890 1997.640 ;
        RECT 1545.230 1610.440 1545.510 1610.720 ;
        RECT 1811.110 1610.440 1811.390 1610.720 ;
        RECT 2004.310 1610.440 2004.590 1610.720 ;
        RECT 1545.230 1609.080 1545.510 1609.360 ;
        RECT 1608.250 1609.080 1608.530 1609.360 ;
        RECT 1704.850 1609.080 1705.130 1609.360 ;
        RECT 1811.110 1609.080 1811.390 1609.360 ;
        RECT 1931.630 1609.080 1931.910 1609.360 ;
        RECT 2004.310 1609.080 2004.590 1609.360 ;
        RECT 2091.250 1609.080 2091.530 1609.360 ;
        RECT 2187.850 1609.080 2188.130 1609.360 ;
        RECT 2284.450 1609.080 2284.730 1609.360 ;
        RECT 2381.050 1609.080 2381.330 1609.360 ;
        RECT 2476.730 1609.080 2477.010 1609.360 ;
        RECT 2477.650 1609.080 2477.930 1609.360 ;
        RECT 2573.330 1609.080 2573.610 1609.360 ;
        RECT 2574.250 1609.080 2574.530 1609.360 ;
        RECT 2669.930 1609.080 2670.210 1609.360 ;
        RECT 2670.850 1609.080 2671.130 1609.360 ;
        RECT 2863.130 1609.080 2863.410 1609.360 ;
        RECT 1425.170 1608.400 1425.450 1608.680 ;
        RECT 1490.030 1608.400 1490.310 1608.680 ;
        RECT 1607.330 1608.400 1607.610 1608.680 ;
        RECT 1703.930 1608.400 1704.210 1608.680 ;
        RECT 1897.130 1608.400 1897.410 1608.680 ;
        RECT 2090.330 1608.400 2090.610 1608.680 ;
        RECT 2186.930 1608.400 2187.210 1608.680 ;
        RECT 2283.530 1608.400 2283.810 1608.680 ;
        RECT 2380.130 1608.400 2380.410 1608.680 ;
        RECT 2814.370 1608.400 2814.650 1608.680 ;
        RECT 2815.750 1608.400 2816.030 1608.680 ;
        RECT 2863.590 1608.400 2863.870 1608.680 ;
        RECT 1425.170 1607.040 1425.450 1607.320 ;
        RECT 1448.170 1607.040 1448.450 1607.320 ;
      LAYER met3 ;
        RECT 1201.585 1997.650 1201.915 1997.665 ;
        RECT 1217.430 1997.650 1217.810 1997.660 ;
        RECT 1201.585 1997.350 1217.810 1997.650 ;
        RECT 1201.585 1997.335 1201.915 1997.350 ;
        RECT 1217.430 1997.340 1217.810 1997.350 ;
        RECT 2917.600 1613.450 2924.800 1613.900 ;
        RECT 2916.710 1613.150 2924.800 1613.450 ;
        RECT 1497.110 1610.730 1497.490 1610.740 ;
        RECT 1545.205 1610.730 1545.535 1610.745 ;
        RECT 1497.110 1610.430 1545.535 1610.730 ;
        RECT 1497.110 1610.420 1497.490 1610.430 ;
        RECT 1545.205 1610.415 1545.535 1610.430 ;
        RECT 1786.910 1610.730 1787.290 1610.740 ;
        RECT 1811.085 1610.730 1811.415 1610.745 ;
        RECT 1786.910 1610.430 1811.415 1610.730 ;
        RECT 1786.910 1610.420 1787.290 1610.430 ;
        RECT 1811.085 1610.415 1811.415 1610.430 ;
        RECT 1980.110 1610.730 1980.490 1610.740 ;
        RECT 2004.285 1610.730 2004.615 1610.745 ;
        RECT 1980.110 1610.430 2004.615 1610.730 ;
        RECT 1980.110 1610.420 1980.490 1610.430 ;
        RECT 2004.285 1610.415 2004.615 1610.430 ;
        RECT 1545.205 1609.370 1545.535 1609.385 ;
        RECT 1608.225 1609.370 1608.555 1609.385 ;
        RECT 1704.825 1609.370 1705.155 1609.385 ;
        RECT 1811.085 1609.370 1811.415 1609.385 ;
        RECT 1931.605 1609.370 1931.935 1609.385 ;
        RECT 2004.285 1609.370 2004.615 1609.385 ;
        RECT 2091.225 1609.370 2091.555 1609.385 ;
        RECT 2187.825 1609.370 2188.155 1609.385 ;
        RECT 2284.425 1609.370 2284.755 1609.385 ;
        RECT 2381.025 1609.370 2381.355 1609.385 ;
        RECT 2476.705 1609.370 2477.035 1609.385 ;
        RECT 1255.190 1609.070 1400.850 1609.370 ;
        RECT 1217.430 1608.010 1217.810 1608.020 ;
        RECT 1255.190 1608.010 1255.490 1609.070 ;
        RECT 1400.550 1608.690 1400.850 1609.070 ;
        RECT 1545.205 1609.070 1560.010 1609.370 ;
        RECT 1545.205 1609.055 1545.535 1609.070 ;
        RECT 1425.145 1608.690 1425.475 1608.705 ;
        RECT 1400.550 1608.390 1425.475 1608.690 ;
        RECT 1425.145 1608.375 1425.475 1608.390 ;
        RECT 1490.005 1608.690 1490.335 1608.705 ;
        RECT 1497.110 1608.690 1497.490 1608.700 ;
        RECT 1490.005 1608.390 1497.490 1608.690 ;
        RECT 1559.710 1608.690 1560.010 1609.070 ;
        RECT 1608.225 1609.070 1656.610 1609.370 ;
        RECT 1608.225 1609.055 1608.555 1609.070 ;
        RECT 1607.305 1608.690 1607.635 1608.705 ;
        RECT 1559.710 1608.390 1607.635 1608.690 ;
        RECT 1656.310 1608.690 1656.610 1609.070 ;
        RECT 1704.825 1609.070 1753.210 1609.370 ;
        RECT 1704.825 1609.055 1705.155 1609.070 ;
        RECT 1703.905 1608.690 1704.235 1608.705 ;
        RECT 1656.310 1608.390 1704.235 1608.690 ;
        RECT 1752.910 1608.690 1753.210 1609.070 ;
        RECT 1811.085 1609.070 1849.810 1609.370 ;
        RECT 1811.085 1609.055 1811.415 1609.070 ;
        RECT 1786.910 1608.690 1787.290 1608.700 ;
        RECT 1752.910 1608.390 1787.290 1608.690 ;
        RECT 1849.510 1608.690 1849.810 1609.070 ;
        RECT 1931.605 1609.070 1946.410 1609.370 ;
        RECT 1931.605 1609.055 1931.935 1609.070 ;
        RECT 1897.105 1608.690 1897.435 1608.705 ;
        RECT 1849.510 1608.390 1897.435 1608.690 ;
        RECT 1946.110 1608.690 1946.410 1609.070 ;
        RECT 2004.285 1609.070 2043.010 1609.370 ;
        RECT 2004.285 1609.055 2004.615 1609.070 ;
        RECT 1980.110 1608.690 1980.490 1608.700 ;
        RECT 1946.110 1608.390 1980.490 1608.690 ;
        RECT 2042.710 1608.690 2043.010 1609.070 ;
        RECT 2091.225 1609.070 2139.610 1609.370 ;
        RECT 2091.225 1609.055 2091.555 1609.070 ;
        RECT 2090.305 1608.690 2090.635 1608.705 ;
        RECT 2042.710 1608.390 2090.635 1608.690 ;
        RECT 2139.310 1608.690 2139.610 1609.070 ;
        RECT 2187.825 1609.070 2236.210 1609.370 ;
        RECT 2187.825 1609.055 2188.155 1609.070 ;
        RECT 2186.905 1608.690 2187.235 1608.705 ;
        RECT 2139.310 1608.390 2187.235 1608.690 ;
        RECT 2235.910 1608.690 2236.210 1609.070 ;
        RECT 2284.425 1609.070 2332.810 1609.370 ;
        RECT 2284.425 1609.055 2284.755 1609.070 ;
        RECT 2283.505 1608.690 2283.835 1608.705 ;
        RECT 2235.910 1608.390 2283.835 1608.690 ;
        RECT 2332.510 1608.690 2332.810 1609.070 ;
        RECT 2381.025 1609.070 2429.410 1609.370 ;
        RECT 2381.025 1609.055 2381.355 1609.070 ;
        RECT 2380.105 1608.690 2380.435 1608.705 ;
        RECT 2332.510 1608.390 2380.435 1608.690 ;
        RECT 2429.110 1608.690 2429.410 1609.070 ;
        RECT 2475.110 1609.070 2477.035 1609.370 ;
        RECT 2475.110 1608.690 2475.410 1609.070 ;
        RECT 2476.705 1609.055 2477.035 1609.070 ;
        RECT 2477.625 1609.370 2477.955 1609.385 ;
        RECT 2573.305 1609.370 2573.635 1609.385 ;
        RECT 2477.625 1609.070 2526.010 1609.370 ;
        RECT 2477.625 1609.055 2477.955 1609.070 ;
        RECT 2429.110 1608.390 2475.410 1608.690 ;
        RECT 2525.710 1608.690 2526.010 1609.070 ;
        RECT 2571.710 1609.070 2573.635 1609.370 ;
        RECT 2571.710 1608.690 2572.010 1609.070 ;
        RECT 2573.305 1609.055 2573.635 1609.070 ;
        RECT 2574.225 1609.370 2574.555 1609.385 ;
        RECT 2669.905 1609.370 2670.235 1609.385 ;
        RECT 2574.225 1609.070 2622.610 1609.370 ;
        RECT 2574.225 1609.055 2574.555 1609.070 ;
        RECT 2525.710 1608.390 2572.010 1608.690 ;
        RECT 2622.310 1608.690 2622.610 1609.070 ;
        RECT 2668.310 1609.070 2670.235 1609.370 ;
        RECT 2668.310 1608.690 2668.610 1609.070 ;
        RECT 2669.905 1609.055 2670.235 1609.070 ;
        RECT 2670.825 1609.370 2671.155 1609.385 ;
        RECT 2863.105 1609.370 2863.435 1609.385 ;
        RECT 2670.825 1609.070 2767.050 1609.370 ;
        RECT 2670.825 1609.055 2671.155 1609.070 ;
        RECT 2622.310 1608.390 2668.610 1608.690 ;
        RECT 2766.750 1608.690 2767.050 1609.070 ;
        RECT 2849.550 1609.070 2863.435 1609.370 ;
        RECT 2814.345 1608.690 2814.675 1608.705 ;
        RECT 2766.750 1608.390 2814.675 1608.690 ;
        RECT 1490.005 1608.375 1490.335 1608.390 ;
        RECT 1497.110 1608.380 1497.490 1608.390 ;
        RECT 1607.305 1608.375 1607.635 1608.390 ;
        RECT 1703.905 1608.375 1704.235 1608.390 ;
        RECT 1786.910 1608.380 1787.290 1608.390 ;
        RECT 1897.105 1608.375 1897.435 1608.390 ;
        RECT 1980.110 1608.380 1980.490 1608.390 ;
        RECT 2090.305 1608.375 2090.635 1608.390 ;
        RECT 2186.905 1608.375 2187.235 1608.390 ;
        RECT 2283.505 1608.375 2283.835 1608.390 ;
        RECT 2380.105 1608.375 2380.435 1608.390 ;
        RECT 2814.345 1608.375 2814.675 1608.390 ;
        RECT 2815.725 1608.690 2816.055 1608.705 ;
        RECT 2849.550 1608.690 2849.850 1609.070 ;
        RECT 2863.105 1609.055 2863.435 1609.070 ;
        RECT 2815.725 1608.390 2849.850 1608.690 ;
        RECT 2863.565 1608.690 2863.895 1608.705 ;
        RECT 2916.710 1608.690 2917.010 1613.150 ;
        RECT 2917.600 1612.700 2924.800 1613.150 ;
        RECT 2863.565 1608.390 2917.010 1608.690 ;
        RECT 2815.725 1608.375 2816.055 1608.390 ;
        RECT 2863.565 1608.375 2863.895 1608.390 ;
        RECT 1217.430 1607.710 1255.490 1608.010 ;
        RECT 1217.430 1607.700 1217.810 1607.710 ;
        RECT 1425.145 1607.330 1425.475 1607.345 ;
        RECT 1448.145 1607.330 1448.475 1607.345 ;
        RECT 1425.145 1607.030 1448.475 1607.330 ;
        RECT 1425.145 1607.015 1425.475 1607.030 ;
        RECT 1448.145 1607.015 1448.475 1607.030 ;
      LAYER via3 ;
        RECT 1217.460 1997.340 1217.780 1997.660 ;
        RECT 1497.140 1610.420 1497.460 1610.740 ;
        RECT 1786.940 1610.420 1787.260 1610.740 ;
        RECT 1980.140 1610.420 1980.460 1610.740 ;
        RECT 1217.460 1607.700 1217.780 1608.020 ;
        RECT 1497.140 1608.380 1497.460 1608.700 ;
        RECT 1786.940 1608.380 1787.260 1608.700 ;
        RECT 1980.140 1608.380 1980.460 1608.700 ;
      LAYER met4 ;
        RECT 1217.455 1997.335 1217.785 1997.665 ;
        RECT 1217.470 1608.025 1217.770 1997.335 ;
        RECT 1497.135 1610.415 1497.465 1610.745 ;
        RECT 1786.935 1610.415 1787.265 1610.745 ;
        RECT 1980.135 1610.415 1980.465 1610.745 ;
        RECT 1497.150 1608.705 1497.450 1610.415 ;
        RECT 1786.950 1608.705 1787.250 1610.415 ;
        RECT 1980.150 1608.705 1980.450 1610.415 ;
        RECT 1497.135 1608.375 1497.465 1608.705 ;
        RECT 1786.935 1608.375 1787.265 1608.705 ;
        RECT 1980.135 1608.375 1980.465 1608.705 ;
        RECT 1217.455 1607.695 1217.785 1608.025 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1208.490 2001.480 1208.810 2001.540 ;
        RECT 1452.750 2001.480 1453.070 2001.540 ;
        RECT 1208.490 2001.340 1453.070 2001.480 ;
        RECT 1208.490 2001.280 1208.810 2001.340 ;
        RECT 1452.750 2001.280 1453.070 2001.340 ;
        RECT 1452.750 1849.160 1453.070 1849.220 ;
        RECT 2900.830 1849.160 2901.150 1849.220 ;
        RECT 1452.750 1849.020 2901.150 1849.160 ;
        RECT 1452.750 1848.960 1453.070 1849.020 ;
        RECT 2900.830 1848.960 2901.150 1849.020 ;
      LAYER via ;
        RECT 1208.520 2001.280 1208.780 2001.540 ;
        RECT 1452.780 2001.280 1453.040 2001.540 ;
        RECT 1452.780 1848.960 1453.040 1849.220 ;
        RECT 2900.860 1848.960 2901.120 1849.220 ;
      LAYER met2 ;
        RECT 1208.520 2001.250 1208.780 2001.570 ;
        RECT 1452.780 2001.250 1453.040 2001.570 ;
        RECT 1208.580 2000.000 1208.720 2001.250 ;
        RECT 1208.420 1999.540 1208.720 2000.000 ;
        RECT 1208.420 1996.000 1208.700 1999.540 ;
        RECT 1452.840 1849.250 1452.980 2001.250 ;
        RECT 1452.780 1848.930 1453.040 1849.250 ;
        RECT 2900.860 1848.930 2901.120 1849.250 ;
        RECT 2900.920 1848.085 2901.060 1848.930 ;
        RECT 2900.850 1847.715 2901.130 1848.085 ;
      LAYER via2 ;
        RECT 2900.850 1847.760 2901.130 1848.040 ;
      LAYER met3 ;
        RECT 2900.825 1848.050 2901.155 1848.065 ;
        RECT 2917.600 1848.050 2924.800 1848.500 ;
        RECT 2900.825 1847.750 2924.800 1848.050 ;
        RECT 2900.825 1847.735 2901.155 1847.750 ;
        RECT 2917.600 1847.300 2924.800 1847.750 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1220.910 2077.300 1221.230 2077.360 ;
        RECT 2900.830 2077.300 2901.150 2077.360 ;
        RECT 1220.910 2077.160 2901.150 2077.300 ;
        RECT 1220.910 2077.100 1221.230 2077.160 ;
        RECT 2900.830 2077.100 2901.150 2077.160 ;
        RECT 1216.310 2009.300 1216.630 2009.360 ;
        RECT 1220.910 2009.300 1221.230 2009.360 ;
        RECT 1216.310 2009.160 1221.230 2009.300 ;
        RECT 1216.310 2009.100 1216.630 2009.160 ;
        RECT 1220.910 2009.100 1221.230 2009.160 ;
      LAYER via ;
        RECT 1220.940 2077.100 1221.200 2077.360 ;
        RECT 2900.860 2077.100 2901.120 2077.360 ;
        RECT 1216.340 2009.100 1216.600 2009.360 ;
        RECT 1220.940 2009.100 1221.200 2009.360 ;
      LAYER met2 ;
        RECT 2900.850 2082.315 2901.130 2082.685 ;
        RECT 2900.920 2077.390 2901.060 2082.315 ;
        RECT 1220.940 2077.070 1221.200 2077.390 ;
        RECT 2900.860 2077.070 2901.120 2077.390 ;
        RECT 1221.000 2009.390 1221.140 2077.070 ;
        RECT 1216.340 2009.070 1216.600 2009.390 ;
        RECT 1220.940 2009.070 1221.200 2009.390 ;
        RECT 1216.400 2000.000 1216.540 2009.070 ;
        RECT 1216.240 1999.540 1216.540 2000.000 ;
        RECT 1216.240 1996.000 1216.520 1999.540 ;
      LAYER via2 ;
        RECT 2900.850 2082.360 2901.130 2082.640 ;
      LAYER met3 ;
        RECT 2900.825 2082.650 2901.155 2082.665 ;
        RECT 2917.600 2082.650 2924.800 2083.100 ;
        RECT 2900.825 2082.350 2924.800 2082.650 ;
        RECT 2900.825 2082.335 2901.155 2082.350 ;
        RECT 2917.600 2081.900 2924.800 2082.350 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1227.810 2311.900 1228.130 2311.960 ;
        RECT 2900.830 2311.900 2901.150 2311.960 ;
        RECT 1227.810 2311.760 2901.150 2311.900 ;
        RECT 1227.810 2311.700 1228.130 2311.760 ;
        RECT 2900.830 2311.700 2901.150 2311.760 ;
        RECT 1224.590 2009.980 1224.910 2010.040 ;
        RECT 1227.810 2009.980 1228.130 2010.040 ;
        RECT 1224.590 2009.840 1228.130 2009.980 ;
        RECT 1224.590 2009.780 1224.910 2009.840 ;
        RECT 1227.810 2009.780 1228.130 2009.840 ;
      LAYER via ;
        RECT 1227.840 2311.700 1228.100 2311.960 ;
        RECT 2900.860 2311.700 2901.120 2311.960 ;
        RECT 1224.620 2009.780 1224.880 2010.040 ;
        RECT 1227.840 2009.780 1228.100 2010.040 ;
      LAYER met2 ;
        RECT 2900.850 2316.915 2901.130 2317.285 ;
        RECT 2900.920 2311.990 2901.060 2316.915 ;
        RECT 1227.840 2311.670 1228.100 2311.990 ;
        RECT 2900.860 2311.670 2901.120 2311.990 ;
        RECT 1227.900 2010.070 1228.040 2311.670 ;
        RECT 1224.620 2009.750 1224.880 2010.070 ;
        RECT 1227.840 2009.750 1228.100 2010.070 ;
        RECT 1224.680 2000.000 1224.820 2009.750 ;
        RECT 1224.520 1999.540 1224.820 2000.000 ;
        RECT 1224.520 1996.000 1224.800 1999.540 ;
      LAYER via2 ;
        RECT 2900.850 2316.960 2901.130 2317.240 ;
      LAYER met3 ;
        RECT 2900.825 2317.250 2901.155 2317.265 ;
        RECT 2917.600 2317.250 2924.800 2317.700 ;
        RECT 2900.825 2316.950 2924.800 2317.250 ;
        RECT 2900.825 2316.935 2901.155 2316.950 ;
        RECT 2917.600 2316.500 2924.800 2316.950 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1607.310 146.100 1607.630 146.160 ;
        RECT 1608.230 146.100 1608.550 146.160 ;
        RECT 1607.310 145.960 1608.550 146.100 ;
        RECT 1607.310 145.900 1607.630 145.960 ;
        RECT 1608.230 145.900 1608.550 145.960 ;
        RECT 1510.710 145.760 1511.030 145.820 ;
        RECT 1544.750 145.760 1545.070 145.820 ;
        RECT 1510.710 145.620 1545.070 145.760 ;
        RECT 1510.710 145.560 1511.030 145.620 ;
        RECT 1544.750 145.560 1545.070 145.620 ;
        RECT 2186.910 145.760 2187.230 145.820 ;
        RECT 2220.950 145.760 2221.270 145.820 ;
        RECT 2186.910 145.620 2221.270 145.760 ;
        RECT 2186.910 145.560 2187.230 145.620 ;
        RECT 2220.950 145.560 2221.270 145.620 ;
        RECT 2573.310 145.760 2573.630 145.820 ;
        RECT 2607.350 145.760 2607.670 145.820 ;
        RECT 2573.310 145.620 2607.670 145.760 ;
        RECT 2573.310 145.560 2573.630 145.620 ;
        RECT 2607.350 145.560 2607.670 145.620 ;
        RECT 2669.910 145.760 2670.230 145.820 ;
        RECT 2703.950 145.760 2704.270 145.820 ;
        RECT 2669.910 145.620 2704.270 145.760 ;
        RECT 2669.910 145.560 2670.230 145.620 ;
        RECT 2703.950 145.560 2704.270 145.620 ;
        RECT 2766.510 145.760 2766.830 145.820 ;
        RECT 2800.550 145.760 2800.870 145.820 ;
        RECT 2766.510 145.620 2800.870 145.760 ;
        RECT 2766.510 145.560 2766.830 145.620 ;
        RECT 2800.550 145.560 2800.870 145.620 ;
        RECT 2863.110 145.760 2863.430 145.820 ;
        RECT 2897.150 145.760 2897.470 145.820 ;
        RECT 2863.110 145.620 2897.470 145.760 ;
        RECT 2863.110 145.560 2863.430 145.620 ;
        RECT 2897.150 145.560 2897.470 145.620 ;
      LAYER via ;
        RECT 1607.340 145.900 1607.600 146.160 ;
        RECT 1608.260 145.900 1608.520 146.160 ;
        RECT 1510.740 145.560 1511.000 145.820 ;
        RECT 1544.780 145.560 1545.040 145.820 ;
        RECT 2186.940 145.560 2187.200 145.820 ;
        RECT 2220.980 145.560 2221.240 145.820 ;
        RECT 2573.340 145.560 2573.600 145.820 ;
        RECT 2607.380 145.560 2607.640 145.820 ;
        RECT 2669.940 145.560 2670.200 145.820 ;
        RECT 2703.980 145.560 2704.240 145.820 ;
        RECT 2766.540 145.560 2766.800 145.820 ;
        RECT 2800.580 145.560 2800.840 145.820 ;
        RECT 2863.140 145.560 2863.400 145.820 ;
        RECT 2897.180 145.560 2897.440 145.820 ;
      LAYER met2 ;
        RECT 1155.980 1996.890 1156.260 2000.000 ;
        RECT 1157.910 1996.890 1158.190 1997.005 ;
        RECT 1155.980 1996.750 1158.190 1996.890 ;
        RECT 1155.980 1996.000 1156.260 1996.750 ;
        RECT 1157.910 1996.635 1158.190 1996.750 ;
        RECT 2487.310 147.035 2487.590 147.405 ;
        RECT 1607.340 146.045 1607.600 146.190 ;
        RECT 1608.260 146.045 1608.520 146.190 ;
        RECT 1510.730 145.675 1511.010 146.045 ;
        RECT 1510.740 145.530 1511.000 145.675 ;
        RECT 1544.780 145.530 1545.040 145.850 ;
        RECT 1607.330 145.675 1607.610 146.045 ;
        RECT 1608.250 145.675 1608.530 146.045 ;
        RECT 2075.610 145.675 2075.890 146.045 ;
        RECT 2186.930 145.675 2187.210 146.045 ;
        RECT 2283.530 145.930 2283.810 146.045 ;
        RECT 2284.450 145.930 2284.730 146.045 ;
        RECT 1544.840 145.250 1544.980 145.530 ;
        RECT 1545.230 145.250 1545.510 145.365 ;
        RECT 1544.840 145.110 1545.510 145.250 ;
        RECT 2075.680 145.250 2075.820 145.675 ;
        RECT 2186.940 145.530 2187.200 145.675 ;
        RECT 2220.980 145.530 2221.240 145.850 ;
        RECT 2283.530 145.790 2284.730 145.930 ;
        RECT 2283.530 145.675 2283.810 145.790 ;
        RECT 2284.450 145.675 2284.730 145.790 ;
        RECT 2456.030 145.675 2456.310 146.045 ;
        RECT 2076.530 145.250 2076.810 145.365 ;
        RECT 2075.680 145.110 2076.810 145.250 ;
        RECT 2221.040 145.250 2221.180 145.530 ;
        RECT 2221.430 145.250 2221.710 145.365 ;
        RECT 2221.040 145.110 2221.710 145.250 ;
        RECT 1545.230 144.995 1545.510 145.110 ;
        RECT 2076.530 144.995 2076.810 145.110 ;
        RECT 2221.430 144.995 2221.710 145.110 ;
        RECT 2456.100 144.005 2456.240 145.675 ;
        RECT 2487.380 145.365 2487.520 147.035 ;
        RECT 2573.330 145.675 2573.610 146.045 ;
        RECT 2573.340 145.530 2573.600 145.675 ;
        RECT 2607.380 145.530 2607.640 145.850 ;
        RECT 2669.930 145.675 2670.210 146.045 ;
        RECT 2669.940 145.530 2670.200 145.675 ;
        RECT 2703.980 145.530 2704.240 145.850 ;
        RECT 2766.530 145.675 2766.810 146.045 ;
        RECT 2766.540 145.530 2766.800 145.675 ;
        RECT 2800.580 145.530 2800.840 145.850 ;
        RECT 2863.130 145.675 2863.410 146.045 ;
        RECT 2863.140 145.530 2863.400 145.675 ;
        RECT 2897.180 145.530 2897.440 145.850 ;
        RECT 2487.310 144.995 2487.590 145.365 ;
        RECT 2607.440 145.250 2607.580 145.530 ;
        RECT 2607.830 145.250 2608.110 145.365 ;
        RECT 2607.440 145.110 2608.110 145.250 ;
        RECT 2704.040 145.250 2704.180 145.530 ;
        RECT 2704.430 145.250 2704.710 145.365 ;
        RECT 2704.040 145.110 2704.710 145.250 ;
        RECT 2800.640 145.250 2800.780 145.530 ;
        RECT 2801.030 145.250 2801.310 145.365 ;
        RECT 2800.640 145.110 2801.310 145.250 ;
        RECT 2897.240 145.250 2897.380 145.530 ;
        RECT 2897.630 145.250 2897.910 145.365 ;
        RECT 2897.240 145.110 2897.910 145.250 ;
        RECT 2607.830 144.995 2608.110 145.110 ;
        RECT 2704.430 144.995 2704.710 145.110 ;
        RECT 2801.030 144.995 2801.310 145.110 ;
        RECT 2897.630 144.995 2897.910 145.110 ;
        RECT 2456.030 143.635 2456.310 144.005 ;
      LAYER via2 ;
        RECT 1157.910 1996.680 1158.190 1996.960 ;
        RECT 2487.310 147.080 2487.590 147.360 ;
        RECT 1510.730 145.720 1511.010 146.000 ;
        RECT 1607.330 145.720 1607.610 146.000 ;
        RECT 1608.250 145.720 1608.530 146.000 ;
        RECT 2075.610 145.720 2075.890 146.000 ;
        RECT 2186.930 145.720 2187.210 146.000 ;
        RECT 1545.230 145.040 1545.510 145.320 ;
        RECT 2283.530 145.720 2283.810 146.000 ;
        RECT 2284.450 145.720 2284.730 146.000 ;
        RECT 2456.030 145.720 2456.310 146.000 ;
        RECT 2076.530 145.040 2076.810 145.320 ;
        RECT 2221.430 145.040 2221.710 145.320 ;
        RECT 2573.330 145.720 2573.610 146.000 ;
        RECT 2669.930 145.720 2670.210 146.000 ;
        RECT 2766.530 145.720 2766.810 146.000 ;
        RECT 2863.130 145.720 2863.410 146.000 ;
        RECT 2487.310 145.040 2487.590 145.320 ;
        RECT 2607.830 145.040 2608.110 145.320 ;
        RECT 2704.430 145.040 2704.710 145.320 ;
        RECT 2801.030 145.040 2801.310 145.320 ;
        RECT 2897.630 145.040 2897.910 145.320 ;
        RECT 2456.030 143.680 2456.310 143.960 ;
      LAYER met3 ;
        RECT 1157.885 1996.970 1158.215 1996.985 ;
        RECT 1158.550 1996.970 1158.930 1996.980 ;
        RECT 1157.885 1996.670 1158.930 1996.970 ;
        RECT 1157.885 1996.655 1158.215 1996.670 ;
        RECT 1158.550 1996.660 1158.930 1996.670 ;
        RECT 2487.285 147.370 2487.615 147.385 ;
        RECT 2463.150 147.070 2487.615 147.370 ;
        RECT 1345.310 146.690 1345.690 146.700 ;
        RECT 1345.310 146.390 1414.650 146.690 ;
        RECT 1345.310 146.380 1345.690 146.390 ;
        RECT 1158.550 146.010 1158.930 146.020 ;
        RECT 1248.710 146.010 1249.090 146.020 ;
        RECT 1158.550 145.710 1249.090 146.010 ;
        RECT 1158.550 145.700 1158.930 145.710 ;
        RECT 1248.710 145.700 1249.090 145.710 ;
        RECT 1249.630 145.330 1250.010 145.340 ;
        RECT 1345.310 145.330 1345.690 145.340 ;
        RECT 1249.630 145.030 1345.690 145.330 ;
        RECT 1414.350 145.330 1414.650 146.390 ;
        RECT 1676.550 146.390 1724.690 146.690 ;
        RECT 1510.705 146.010 1511.035 146.025 ;
        RECT 1607.305 146.010 1607.635 146.025 ;
        RECT 1463.110 145.710 1511.035 146.010 ;
        RECT 1463.110 145.330 1463.410 145.710 ;
        RECT 1510.705 145.695 1511.035 145.710 ;
        RECT 1559.710 145.710 1607.635 146.010 ;
        RECT 1414.350 145.030 1463.410 145.330 ;
        RECT 1545.205 145.330 1545.535 145.345 ;
        RECT 1559.710 145.330 1560.010 145.710 ;
        RECT 1607.305 145.695 1607.635 145.710 ;
        RECT 1608.225 146.010 1608.555 146.025 ;
        RECT 1608.225 145.710 1655.690 146.010 ;
        RECT 1608.225 145.695 1608.555 145.710 ;
        RECT 1545.205 145.030 1560.010 145.330 ;
        RECT 1655.390 145.330 1655.690 145.710 ;
        RECT 1676.550 145.330 1676.850 146.390 ;
        RECT 1655.390 145.030 1676.850 145.330 ;
        RECT 1724.390 145.330 1724.690 146.390 ;
        RECT 1725.310 146.390 1773.450 146.690 ;
        RECT 1725.310 145.330 1725.610 146.390 ;
        RECT 1773.150 146.010 1773.450 146.390 ;
        RECT 1821.910 146.390 1870.050 146.690 ;
        RECT 1773.150 145.710 1821.290 146.010 ;
        RECT 1724.390 145.030 1725.610 145.330 ;
        RECT 1820.990 145.330 1821.290 145.710 ;
        RECT 1821.910 145.330 1822.210 146.390 ;
        RECT 1869.750 146.010 1870.050 146.390 ;
        RECT 1918.510 146.390 2029.210 146.690 ;
        RECT 1869.750 145.710 1917.890 146.010 ;
        RECT 1820.990 145.030 1822.210 145.330 ;
        RECT 1917.590 145.330 1917.890 145.710 ;
        RECT 1918.510 145.330 1918.810 146.390 ;
        RECT 2028.910 146.010 2029.210 146.390 ;
        RECT 2075.585 146.010 2075.915 146.025 ;
        RECT 2186.905 146.010 2187.235 146.025 ;
        RECT 2283.505 146.010 2283.835 146.025 ;
        RECT 2028.910 145.710 2075.915 146.010 ;
        RECT 2075.585 145.695 2075.915 145.710 ;
        RECT 2139.310 145.710 2187.235 146.010 ;
        RECT 1917.590 145.030 1918.810 145.330 ;
        RECT 2076.505 145.330 2076.835 145.345 ;
        RECT 2139.310 145.330 2139.610 145.710 ;
        RECT 2186.905 145.695 2187.235 145.710 ;
        RECT 2235.910 145.710 2283.835 146.010 ;
        RECT 2076.505 145.030 2139.610 145.330 ;
        RECT 2221.405 145.330 2221.735 145.345 ;
        RECT 2235.910 145.330 2236.210 145.710 ;
        RECT 2283.505 145.695 2283.835 145.710 ;
        RECT 2284.425 146.010 2284.755 146.025 ;
        RECT 2456.005 146.010 2456.335 146.025 ;
        RECT 2463.150 146.010 2463.450 147.070 ;
        RECT 2487.285 147.055 2487.615 147.070 ;
        RECT 2917.600 146.690 2924.800 147.140 ;
        RECT 2916.710 146.390 2924.800 146.690 ;
        RECT 2573.305 146.010 2573.635 146.025 ;
        RECT 2669.905 146.010 2670.235 146.025 ;
        RECT 2766.505 146.010 2766.835 146.025 ;
        RECT 2863.105 146.010 2863.435 146.025 ;
        RECT 2284.425 145.710 2331.890 146.010 ;
        RECT 2284.425 145.695 2284.755 145.710 ;
        RECT 2221.405 145.030 2236.210 145.330 ;
        RECT 2331.590 145.330 2331.890 145.710 ;
        RECT 2332.510 145.710 2390.770 146.010 ;
        RECT 2332.510 145.330 2332.810 145.710 ;
        RECT 2331.590 145.030 2332.810 145.330 ;
        RECT 2390.470 145.330 2390.770 145.710 ;
        RECT 2456.005 145.710 2463.450 146.010 ;
        RECT 2525.710 145.710 2573.635 146.010 ;
        RECT 2456.005 145.695 2456.335 145.710 ;
        RECT 2407.910 145.330 2408.290 145.340 ;
        RECT 2390.470 145.030 2408.290 145.330 ;
        RECT 1249.630 145.020 1250.010 145.030 ;
        RECT 1345.310 145.020 1345.690 145.030 ;
        RECT 1545.205 145.015 1545.535 145.030 ;
        RECT 2076.505 145.015 2076.835 145.030 ;
        RECT 2221.405 145.015 2221.735 145.030 ;
        RECT 2407.910 145.020 2408.290 145.030 ;
        RECT 2487.285 145.330 2487.615 145.345 ;
        RECT 2525.710 145.330 2526.010 145.710 ;
        RECT 2573.305 145.695 2573.635 145.710 ;
        RECT 2622.310 145.710 2670.235 146.010 ;
        RECT 2487.285 145.030 2526.010 145.330 ;
        RECT 2607.805 145.330 2608.135 145.345 ;
        RECT 2622.310 145.330 2622.610 145.710 ;
        RECT 2669.905 145.695 2670.235 145.710 ;
        RECT 2718.910 145.710 2766.835 146.010 ;
        RECT 2607.805 145.030 2622.610 145.330 ;
        RECT 2704.405 145.330 2704.735 145.345 ;
        RECT 2718.910 145.330 2719.210 145.710 ;
        RECT 2766.505 145.695 2766.835 145.710 ;
        RECT 2815.510 145.710 2863.435 146.010 ;
        RECT 2704.405 145.030 2719.210 145.330 ;
        RECT 2801.005 145.330 2801.335 145.345 ;
        RECT 2815.510 145.330 2815.810 145.710 ;
        RECT 2863.105 145.695 2863.435 145.710 ;
        RECT 2801.005 145.030 2815.810 145.330 ;
        RECT 2897.605 145.330 2897.935 145.345 ;
        RECT 2916.710 145.330 2917.010 146.390 ;
        RECT 2917.600 145.940 2924.800 146.390 ;
        RECT 2897.605 145.030 2917.010 145.330 ;
        RECT 2487.285 145.015 2487.615 145.030 ;
        RECT 2607.805 145.015 2608.135 145.030 ;
        RECT 2704.405 145.015 2704.735 145.030 ;
        RECT 2801.005 145.015 2801.335 145.030 ;
        RECT 2897.605 145.015 2897.935 145.030 ;
        RECT 2407.910 143.970 2408.290 143.980 ;
        RECT 2456.005 143.970 2456.335 143.985 ;
        RECT 2407.910 143.670 2456.335 143.970 ;
        RECT 2407.910 143.660 2408.290 143.670 ;
        RECT 2456.005 143.655 2456.335 143.670 ;
      LAYER via3 ;
        RECT 1158.580 1996.660 1158.900 1996.980 ;
        RECT 1345.340 146.380 1345.660 146.700 ;
        RECT 1158.580 145.700 1158.900 146.020 ;
        RECT 1248.740 145.700 1249.060 146.020 ;
        RECT 1249.660 145.020 1249.980 145.340 ;
        RECT 1345.340 145.020 1345.660 145.340 ;
        RECT 2407.940 145.020 2408.260 145.340 ;
        RECT 2407.940 143.660 2408.260 143.980 ;
      LAYER met4 ;
        RECT 1158.575 1996.655 1158.905 1996.985 ;
        RECT 1158.590 146.025 1158.890 1996.655 ;
        RECT 1345.335 146.375 1345.665 146.705 ;
        RECT 1158.575 145.695 1158.905 146.025 ;
        RECT 1248.735 146.010 1249.065 146.025 ;
        RECT 1248.735 145.710 1249.970 146.010 ;
        RECT 1248.735 145.695 1249.065 145.710 ;
        RECT 1249.670 145.345 1249.970 145.710 ;
        RECT 1345.350 145.345 1345.650 146.375 ;
        RECT 1249.655 145.015 1249.985 145.345 ;
        RECT 1345.335 145.015 1345.665 145.345 ;
        RECT 2407.935 145.015 2408.265 145.345 ;
        RECT 2407.950 143.985 2408.250 145.015 ;
        RECT 2407.935 143.655 2408.265 143.985 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1240.690 2491.080 1241.010 2491.140 ;
        RECT 2900.830 2491.080 2901.150 2491.140 ;
        RECT 1240.690 2490.940 2901.150 2491.080 ;
        RECT 1240.690 2490.880 1241.010 2490.940 ;
        RECT 2900.830 2490.880 2901.150 2490.940 ;
        RECT 1235.170 2009.980 1235.490 2010.040 ;
        RECT 1240.690 2009.980 1241.010 2010.040 ;
        RECT 1235.170 2009.840 1241.010 2009.980 ;
        RECT 1235.170 2009.780 1235.490 2009.840 ;
        RECT 1240.690 2009.780 1241.010 2009.840 ;
      LAYER via ;
        RECT 1240.720 2490.880 1240.980 2491.140 ;
        RECT 2900.860 2490.880 2901.120 2491.140 ;
        RECT 1235.200 2009.780 1235.460 2010.040 ;
        RECT 1240.720 2009.780 1240.980 2010.040 ;
      LAYER met2 ;
        RECT 2900.850 2493.035 2901.130 2493.405 ;
        RECT 2900.920 2491.170 2901.060 2493.035 ;
        RECT 1240.720 2490.850 1240.980 2491.170 ;
        RECT 2900.860 2490.850 2901.120 2491.170 ;
        RECT 1240.780 2010.070 1240.920 2490.850 ;
        RECT 1235.200 2009.750 1235.460 2010.070 ;
        RECT 1240.720 2009.750 1240.980 2010.070 ;
        RECT 1235.260 2000.000 1235.400 2009.750 ;
        RECT 1235.100 1999.540 1235.400 2000.000 ;
        RECT 1235.100 1996.000 1235.380 1999.540 ;
      LAYER via2 ;
        RECT 2900.850 2493.080 2901.130 2493.360 ;
      LAYER met3 ;
        RECT 2900.825 2493.370 2901.155 2493.385 ;
        RECT 2917.600 2493.370 2924.800 2493.820 ;
        RECT 2900.825 2493.070 2924.800 2493.370 ;
        RECT 2900.825 2493.055 2901.155 2493.070 ;
        RECT 2917.600 2492.620 2924.800 2493.070 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1247.590 2725.680 1247.910 2725.740 ;
        RECT 2900.830 2725.680 2901.150 2725.740 ;
        RECT 1247.590 2725.540 2901.150 2725.680 ;
        RECT 1247.590 2725.480 1247.910 2725.540 ;
        RECT 2900.830 2725.480 2901.150 2725.540 ;
        RECT 1242.990 2009.980 1243.310 2010.040 ;
        RECT 1247.590 2009.980 1247.910 2010.040 ;
        RECT 1242.990 2009.840 1247.910 2009.980 ;
        RECT 1242.990 2009.780 1243.310 2009.840 ;
        RECT 1247.590 2009.780 1247.910 2009.840 ;
      LAYER via ;
        RECT 1247.620 2725.480 1247.880 2725.740 ;
        RECT 2900.860 2725.480 2901.120 2725.740 ;
        RECT 1243.020 2009.780 1243.280 2010.040 ;
        RECT 1247.620 2009.780 1247.880 2010.040 ;
      LAYER met2 ;
        RECT 2900.850 2727.635 2901.130 2728.005 ;
        RECT 2900.920 2725.770 2901.060 2727.635 ;
        RECT 1247.620 2725.450 1247.880 2725.770 ;
        RECT 2900.860 2725.450 2901.120 2725.770 ;
        RECT 1247.680 2010.070 1247.820 2725.450 ;
        RECT 1243.020 2009.750 1243.280 2010.070 ;
        RECT 1247.620 2009.750 1247.880 2010.070 ;
        RECT 1243.080 2000.000 1243.220 2009.750 ;
        RECT 1242.920 1999.540 1243.220 2000.000 ;
        RECT 1242.920 1996.000 1243.200 1999.540 ;
      LAYER via2 ;
        RECT 2900.850 2727.680 2901.130 2727.960 ;
      LAYER met3 ;
        RECT 2900.825 2727.970 2901.155 2727.985 ;
        RECT 2917.600 2727.970 2924.800 2728.420 ;
        RECT 2900.825 2727.670 2924.800 2727.970 ;
        RECT 2900.825 2727.655 2901.155 2727.670 ;
        RECT 2917.600 2727.220 2924.800 2727.670 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1254.950 2960.280 1255.270 2960.340 ;
        RECT 2900.830 2960.280 2901.150 2960.340 ;
        RECT 1254.950 2960.140 2901.150 2960.280 ;
        RECT 1254.950 2960.080 1255.270 2960.140 ;
        RECT 2900.830 2960.080 2901.150 2960.140 ;
        RECT 1250.810 2009.980 1251.130 2010.040 ;
        RECT 1254.950 2009.980 1255.270 2010.040 ;
        RECT 1250.810 2009.840 1255.270 2009.980 ;
        RECT 1250.810 2009.780 1251.130 2009.840 ;
        RECT 1254.950 2009.780 1255.270 2009.840 ;
      LAYER via ;
        RECT 1254.980 2960.080 1255.240 2960.340 ;
        RECT 2900.860 2960.080 2901.120 2960.340 ;
        RECT 1250.840 2009.780 1251.100 2010.040 ;
        RECT 1254.980 2009.780 1255.240 2010.040 ;
      LAYER met2 ;
        RECT 2900.850 2962.235 2901.130 2962.605 ;
        RECT 2900.920 2960.370 2901.060 2962.235 ;
        RECT 1254.980 2960.050 1255.240 2960.370 ;
        RECT 2900.860 2960.050 2901.120 2960.370 ;
        RECT 1255.040 2010.070 1255.180 2960.050 ;
        RECT 1250.840 2009.750 1251.100 2010.070 ;
        RECT 1254.980 2009.750 1255.240 2010.070 ;
        RECT 1250.900 2000.000 1251.040 2009.750 ;
        RECT 1250.740 1999.540 1251.040 2000.000 ;
        RECT 1250.740 1996.000 1251.020 1999.540 ;
      LAYER via2 ;
        RECT 2900.850 2962.280 2901.130 2962.560 ;
      LAYER met3 ;
        RECT 2900.825 2962.570 2901.155 2962.585 ;
        RECT 2917.600 2962.570 2924.800 2963.020 ;
        RECT 2900.825 2962.270 2924.800 2962.570 ;
        RECT 2900.825 2962.255 2901.155 2962.270 ;
        RECT 2917.600 2961.820 2924.800 2962.270 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1261.390 3194.880 1261.710 3194.940 ;
        RECT 2900.830 3194.880 2901.150 3194.940 ;
        RECT 1261.390 3194.740 2901.150 3194.880 ;
        RECT 1261.390 3194.680 1261.710 3194.740 ;
        RECT 2900.830 3194.680 2901.150 3194.740 ;
      LAYER via ;
        RECT 1261.420 3194.680 1261.680 3194.940 ;
        RECT 2900.860 3194.680 2901.120 3194.940 ;
      LAYER met2 ;
        RECT 2900.850 3196.835 2901.130 3197.205 ;
        RECT 2900.920 3194.970 2901.060 3196.835 ;
        RECT 1261.420 3194.650 1261.680 3194.970 ;
        RECT 2900.860 3194.650 2901.120 3194.970 ;
        RECT 1261.480 2001.650 1261.620 3194.650 ;
        RECT 1261.020 2001.510 1261.620 2001.650 ;
        RECT 1258.560 1998.930 1258.840 2000.000 ;
        RECT 1261.020 1998.930 1261.160 2001.510 ;
        RECT 1258.560 1998.790 1261.160 1998.930 ;
        RECT 1258.560 1996.000 1258.840 1998.790 ;
      LAYER via2 ;
        RECT 2900.850 3196.880 2901.130 3197.160 ;
      LAYER met3 ;
        RECT 2900.825 3197.170 2901.155 3197.185 ;
        RECT 2917.600 3197.170 2924.800 3197.620 ;
        RECT 2900.825 3196.870 2924.800 3197.170 ;
        RECT 2900.825 3196.855 2901.155 3196.870 ;
        RECT 2917.600 3196.420 2924.800 3196.870 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1497.460 3429.680 1506.340 3429.820 ;
        RECT 1268.290 3429.480 1268.610 3429.540 ;
        RECT 1497.460 3429.480 1497.600 3429.680 ;
        RECT 1268.290 3429.340 1497.600 3429.480 ;
        RECT 1506.200 3429.480 1506.340 3429.680 ;
        RECT 2900.830 3429.480 2901.150 3429.540 ;
        RECT 1506.200 3429.340 2901.150 3429.480 ;
        RECT 1268.290 3429.280 1268.610 3429.340 ;
        RECT 2900.830 3429.280 2901.150 3429.340 ;
      LAYER via ;
        RECT 1268.320 3429.280 1268.580 3429.540 ;
        RECT 2900.860 3429.280 2901.120 3429.540 ;
      LAYER met2 ;
        RECT 2900.850 3431.435 2901.130 3431.805 ;
        RECT 2900.920 3429.570 2901.060 3431.435 ;
        RECT 1268.320 3429.250 1268.580 3429.570 ;
        RECT 2900.860 3429.250 2901.120 3429.570 ;
        RECT 1266.380 1999.610 1266.660 2000.000 ;
        RECT 1268.380 1999.610 1268.520 3429.250 ;
        RECT 1266.380 1999.470 1268.520 1999.610 ;
        RECT 1266.380 1996.000 1266.660 1999.470 ;
      LAYER via2 ;
        RECT 2900.850 3431.480 2901.130 3431.760 ;
      LAYER met3 ;
        RECT 2900.825 3431.770 2901.155 3431.785 ;
        RECT 2917.600 3431.770 2924.800 3432.220 ;
        RECT 2900.825 3431.470 2924.800 3431.770 ;
        RECT 2900.825 3431.455 2901.155 3431.470 ;
        RECT 2917.600 3431.020 2924.800 3431.470 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1275.650 3501.900 1275.970 3501.960 ;
        RECT 2717.290 3501.900 2717.610 3501.960 ;
        RECT 1275.650 3501.760 2717.610 3501.900 ;
        RECT 1275.650 3501.700 1275.970 3501.760 ;
        RECT 2717.290 3501.700 2717.610 3501.760 ;
      LAYER via ;
        RECT 1275.680 3501.700 1275.940 3501.960 ;
        RECT 2717.320 3501.700 2717.580 3501.960 ;
      LAYER met2 ;
        RECT 2717.170 3517.600 2717.730 3524.800 ;
        RECT 2717.380 3501.990 2717.520 3517.600 ;
        RECT 1275.680 3501.670 1275.940 3501.990 ;
        RECT 2717.320 3501.670 2717.580 3501.990 ;
        RECT 1274.200 1999.610 1274.480 2000.000 ;
        RECT 1275.740 1999.610 1275.880 3501.670 ;
        RECT 1274.200 1999.470 1275.880 1999.610 ;
        RECT 1274.200 1996.000 1274.480 1999.470 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1283.010 3503.260 1283.330 3503.320 ;
        RECT 2392.530 3503.260 2392.850 3503.320 ;
        RECT 1283.010 3503.120 2392.850 3503.260 ;
        RECT 1283.010 3503.060 1283.330 3503.120 ;
        RECT 2392.530 3503.060 2392.850 3503.120 ;
      LAYER via ;
        RECT 1283.040 3503.060 1283.300 3503.320 ;
        RECT 2392.560 3503.060 2392.820 3503.320 ;
      LAYER met2 ;
        RECT 2392.410 3517.600 2392.970 3524.800 ;
        RECT 2392.620 3503.350 2392.760 3517.600 ;
        RECT 1283.040 3503.030 1283.300 3503.350 ;
        RECT 2392.560 3503.030 2392.820 3503.350 ;
        RECT 1282.020 1999.610 1282.300 2000.000 ;
        RECT 1283.100 1999.610 1283.240 3503.030 ;
        RECT 1282.020 1999.470 1283.240 1999.610 ;
        RECT 1282.020 1996.000 1282.300 1999.470 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1296.810 3504.620 1297.130 3504.680 ;
        RECT 2068.230 3504.620 2068.550 3504.680 ;
        RECT 1296.810 3504.480 2068.550 3504.620 ;
        RECT 1296.810 3504.420 1297.130 3504.480 ;
        RECT 2068.230 3504.420 2068.550 3504.480 ;
        RECT 1290.370 2011.000 1290.690 2011.060 ;
        RECT 1296.810 2011.000 1297.130 2011.060 ;
        RECT 1290.370 2010.860 1297.130 2011.000 ;
        RECT 1290.370 2010.800 1290.690 2010.860 ;
        RECT 1296.810 2010.800 1297.130 2010.860 ;
      LAYER via ;
        RECT 1296.840 3504.420 1297.100 3504.680 ;
        RECT 2068.260 3504.420 2068.520 3504.680 ;
        RECT 1290.400 2010.800 1290.660 2011.060 ;
        RECT 1296.840 2010.800 1297.100 2011.060 ;
      LAYER met2 ;
        RECT 2068.110 3517.600 2068.670 3524.800 ;
        RECT 2068.320 3504.710 2068.460 3517.600 ;
        RECT 1296.840 3504.390 1297.100 3504.710 ;
        RECT 2068.260 3504.390 2068.520 3504.710 ;
        RECT 1296.900 2011.090 1297.040 3504.390 ;
        RECT 1290.400 2010.770 1290.660 2011.090 ;
        RECT 1296.840 2010.770 1297.100 2011.090 ;
        RECT 1290.460 2000.000 1290.600 2010.770 ;
        RECT 1290.300 1999.540 1290.600 2000.000 ;
        RECT 1290.300 1996.000 1290.580 1999.540 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1303.250 3500.540 1303.570 3500.600 ;
        RECT 1743.930 3500.540 1744.250 3500.600 ;
        RECT 1303.250 3500.400 1744.250 3500.540 ;
        RECT 1303.250 3500.340 1303.570 3500.400 ;
        RECT 1743.930 3500.340 1744.250 3500.400 ;
        RECT 1298.190 2014.400 1298.510 2014.460 ;
        RECT 1303.250 2014.400 1303.570 2014.460 ;
        RECT 1298.190 2014.260 1303.570 2014.400 ;
        RECT 1298.190 2014.200 1298.510 2014.260 ;
        RECT 1303.250 2014.200 1303.570 2014.260 ;
      LAYER via ;
        RECT 1303.280 3500.340 1303.540 3500.600 ;
        RECT 1743.960 3500.340 1744.220 3500.600 ;
        RECT 1298.220 2014.200 1298.480 2014.460 ;
        RECT 1303.280 2014.200 1303.540 2014.460 ;
      LAYER met2 ;
        RECT 1743.810 3517.600 1744.370 3524.800 ;
        RECT 1744.020 3500.630 1744.160 3517.600 ;
        RECT 1303.280 3500.310 1303.540 3500.630 ;
        RECT 1743.960 3500.310 1744.220 3500.630 ;
        RECT 1303.340 2014.490 1303.480 3500.310 ;
        RECT 1298.220 2014.170 1298.480 2014.490 ;
        RECT 1303.280 2014.170 1303.540 2014.490 ;
        RECT 1298.280 2000.000 1298.420 2014.170 ;
        RECT 1298.120 1999.540 1298.420 2000.000 ;
        RECT 1298.120 1996.000 1298.400 1999.540 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1310.610 3499.520 1310.930 3499.580 ;
        RECT 1419.170 3499.520 1419.490 3499.580 ;
        RECT 1310.610 3499.380 1419.490 3499.520 ;
        RECT 1310.610 3499.320 1310.930 3499.380 ;
        RECT 1419.170 3499.320 1419.490 3499.380 ;
        RECT 1306.010 2014.400 1306.330 2014.460 ;
        RECT 1310.610 2014.400 1310.930 2014.460 ;
        RECT 1306.010 2014.260 1310.930 2014.400 ;
        RECT 1306.010 2014.200 1306.330 2014.260 ;
        RECT 1310.610 2014.200 1310.930 2014.260 ;
      LAYER via ;
        RECT 1310.640 3499.320 1310.900 3499.580 ;
        RECT 1419.200 3499.320 1419.460 3499.580 ;
        RECT 1306.040 2014.200 1306.300 2014.460 ;
        RECT 1310.640 2014.200 1310.900 2014.460 ;
      LAYER met2 ;
        RECT 1419.050 3517.600 1419.610 3524.800 ;
        RECT 1419.260 3499.610 1419.400 3517.600 ;
        RECT 1310.640 3499.290 1310.900 3499.610 ;
        RECT 1419.200 3499.290 1419.460 3499.610 ;
        RECT 1310.700 2014.490 1310.840 3499.290 ;
        RECT 1306.040 2014.170 1306.300 2014.490 ;
        RECT 1310.640 2014.170 1310.900 2014.490 ;
        RECT 1306.100 2000.000 1306.240 2014.170 ;
        RECT 1305.940 1999.540 1306.240 2000.000 ;
        RECT 1305.940 1996.000 1306.220 1999.540 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1607.310 380.700 1607.630 380.760 ;
        RECT 1615.130 380.700 1615.450 380.760 ;
        RECT 1607.310 380.560 1615.450 380.700 ;
        RECT 1607.310 380.500 1607.630 380.560 ;
        RECT 1615.130 380.500 1615.450 380.560 ;
        RECT 1401.230 380.360 1401.550 380.420 ;
        RECT 1448.610 380.360 1448.930 380.420 ;
        RECT 1401.230 380.220 1448.930 380.360 ;
        RECT 1401.230 380.160 1401.550 380.220 ;
        RECT 1448.610 380.160 1448.930 380.220 ;
        RECT 1510.710 380.360 1511.030 380.420 ;
        RECT 1545.210 380.360 1545.530 380.420 ;
        RECT 1510.710 380.220 1545.530 380.360 ;
        RECT 1510.710 380.160 1511.030 380.220 ;
        RECT 1545.210 380.160 1545.530 380.220 ;
        RECT 2186.910 380.360 2187.230 380.420 ;
        RECT 2221.410 380.360 2221.730 380.420 ;
        RECT 2186.910 380.220 2221.730 380.360 ;
        RECT 2186.910 380.160 2187.230 380.220 ;
        RECT 2221.410 380.160 2221.730 380.220 ;
        RECT 2511.210 380.360 2511.530 380.420 ;
        RECT 2552.610 380.360 2552.930 380.420 ;
        RECT 2511.210 380.220 2552.930 380.360 ;
        RECT 2511.210 380.160 2511.530 380.220 ;
        RECT 2552.610 380.160 2552.930 380.220 ;
        RECT 2669.910 380.360 2670.230 380.420 ;
        RECT 2704.410 380.360 2704.730 380.420 ;
        RECT 2669.910 380.220 2704.730 380.360 ;
        RECT 2669.910 380.160 2670.230 380.220 ;
        RECT 2704.410 380.160 2704.730 380.220 ;
        RECT 2766.510 380.360 2766.830 380.420 ;
        RECT 2801.010 380.360 2801.330 380.420 ;
        RECT 2766.510 380.220 2801.330 380.360 ;
        RECT 2766.510 380.160 2766.830 380.220 ;
        RECT 2801.010 380.160 2801.330 380.220 ;
        RECT 2863.110 380.360 2863.430 380.420 ;
        RECT 2897.610 380.360 2897.930 380.420 ;
        RECT 2863.110 380.220 2897.930 380.360 ;
        RECT 2863.110 380.160 2863.430 380.220 ;
        RECT 2897.610 380.160 2897.930 380.220 ;
      LAYER via ;
        RECT 1607.340 380.500 1607.600 380.760 ;
        RECT 1615.160 380.500 1615.420 380.760 ;
        RECT 1401.260 380.160 1401.520 380.420 ;
        RECT 1448.640 380.160 1448.900 380.420 ;
        RECT 1510.740 380.160 1511.000 380.420 ;
        RECT 1545.240 380.160 1545.500 380.420 ;
        RECT 2186.940 380.160 2187.200 380.420 ;
        RECT 2221.440 380.160 2221.700 380.420 ;
        RECT 2511.240 380.160 2511.500 380.420 ;
        RECT 2552.640 380.160 2552.900 380.420 ;
        RECT 2669.940 380.160 2670.200 380.420 ;
        RECT 2704.440 380.160 2704.700 380.420 ;
        RECT 2766.540 380.160 2766.800 380.420 ;
        RECT 2801.040 380.160 2801.300 380.420 ;
        RECT 2863.140 380.160 2863.400 380.420 ;
        RECT 2897.640 380.160 2897.900 380.420 ;
      LAYER met2 ;
        RECT 1163.800 1996.890 1164.080 2000.000 ;
        RECT 1164.810 1996.890 1165.090 1997.005 ;
        RECT 1163.800 1996.750 1165.090 1996.890 ;
        RECT 1163.800 1996.000 1164.080 1996.750 ;
        RECT 1164.810 1996.635 1165.090 1996.750 ;
        RECT 2607.830 382.315 2608.110 382.685 ;
        RECT 2552.630 380.955 2552.910 381.325 ;
        RECT 1607.340 380.645 1607.600 380.790 ;
        RECT 1615.160 380.645 1615.420 380.790 ;
        RECT 1401.250 380.275 1401.530 380.645 ;
        RECT 1401.260 380.130 1401.520 380.275 ;
        RECT 1448.640 380.130 1448.900 380.450 ;
        RECT 1510.730 380.275 1511.010 380.645 ;
        RECT 1510.740 380.130 1511.000 380.275 ;
        RECT 1545.240 380.130 1545.500 380.450 ;
        RECT 1607.330 380.275 1607.610 380.645 ;
        RECT 1615.150 380.275 1615.430 380.645 ;
        RECT 2076.530 380.275 2076.810 380.645 ;
        RECT 2186.930 380.275 2187.210 380.645 ;
        RECT 2283.530 380.530 2283.810 380.645 ;
        RECT 2284.450 380.530 2284.730 380.645 ;
        RECT 1448.700 379.965 1448.840 380.130 ;
        RECT 1545.300 379.965 1545.440 380.130 ;
        RECT 2076.600 379.965 2076.740 380.275 ;
        RECT 2186.940 380.130 2187.200 380.275 ;
        RECT 2221.440 380.130 2221.700 380.450 ;
        RECT 2283.530 380.390 2284.730 380.530 ;
        RECT 2283.530 380.275 2283.810 380.390 ;
        RECT 2284.450 380.275 2284.730 380.390 ;
        RECT 2414.630 380.275 2414.910 380.645 ;
        RECT 2552.700 380.450 2552.840 380.955 ;
        RECT 2221.500 379.965 2221.640 380.130 ;
        RECT 2414.700 379.965 2414.840 380.275 ;
        RECT 2511.240 380.130 2511.500 380.450 ;
        RECT 2552.640 380.130 2552.900 380.450 ;
        RECT 1221.390 379.850 1221.670 379.965 ;
        RECT 1222.310 379.850 1222.590 379.965 ;
        RECT 1221.390 379.710 1222.590 379.850 ;
        RECT 1221.390 379.595 1221.670 379.710 ;
        RECT 1222.310 379.595 1222.590 379.710 ;
        RECT 1448.630 379.595 1448.910 379.965 ;
        RECT 1545.230 379.595 1545.510 379.965 ;
        RECT 2076.530 379.595 2076.810 379.965 ;
        RECT 2221.430 379.595 2221.710 379.965 ;
        RECT 2414.630 379.595 2414.910 379.965 ;
        RECT 2511.300 379.285 2511.440 380.130 ;
        RECT 2607.900 379.965 2608.040 382.315 ;
        RECT 2669.930 380.275 2670.210 380.645 ;
        RECT 2669.940 380.130 2670.200 380.275 ;
        RECT 2704.440 380.130 2704.700 380.450 ;
        RECT 2766.530 380.275 2766.810 380.645 ;
        RECT 2766.540 380.130 2766.800 380.275 ;
        RECT 2801.040 380.130 2801.300 380.450 ;
        RECT 2863.130 380.275 2863.410 380.645 ;
        RECT 2863.140 380.130 2863.400 380.275 ;
        RECT 2897.640 380.130 2897.900 380.450 ;
        RECT 2704.500 379.965 2704.640 380.130 ;
        RECT 2801.100 379.965 2801.240 380.130 ;
        RECT 2897.700 379.965 2897.840 380.130 ;
        RECT 2607.830 379.595 2608.110 379.965 ;
        RECT 2704.430 379.595 2704.710 379.965 ;
        RECT 2801.030 379.595 2801.310 379.965 ;
        RECT 2897.630 379.595 2897.910 379.965 ;
        RECT 2511.230 378.915 2511.510 379.285 ;
      LAYER via2 ;
        RECT 1164.810 1996.680 1165.090 1996.960 ;
        RECT 2607.830 382.360 2608.110 382.640 ;
        RECT 2552.630 381.000 2552.910 381.280 ;
        RECT 1401.250 380.320 1401.530 380.600 ;
        RECT 1510.730 380.320 1511.010 380.600 ;
        RECT 1607.330 380.320 1607.610 380.600 ;
        RECT 1615.150 380.320 1615.430 380.600 ;
        RECT 2076.530 380.320 2076.810 380.600 ;
        RECT 2186.930 380.320 2187.210 380.600 ;
        RECT 2283.530 380.320 2283.810 380.600 ;
        RECT 2284.450 380.320 2284.730 380.600 ;
        RECT 2414.630 380.320 2414.910 380.600 ;
        RECT 1221.390 379.640 1221.670 379.920 ;
        RECT 1222.310 379.640 1222.590 379.920 ;
        RECT 1448.630 379.640 1448.910 379.920 ;
        RECT 1545.230 379.640 1545.510 379.920 ;
        RECT 2076.530 379.640 2076.810 379.920 ;
        RECT 2221.430 379.640 2221.710 379.920 ;
        RECT 2414.630 379.640 2414.910 379.920 ;
        RECT 2669.930 380.320 2670.210 380.600 ;
        RECT 2766.530 380.320 2766.810 380.600 ;
        RECT 2863.130 380.320 2863.410 380.600 ;
        RECT 2607.830 379.640 2608.110 379.920 ;
        RECT 2704.430 379.640 2704.710 379.920 ;
        RECT 2801.030 379.640 2801.310 379.920 ;
        RECT 2897.630 379.640 2897.910 379.920 ;
        RECT 2511.230 378.960 2511.510 379.240 ;
      LAYER met3 ;
        RECT 1164.785 1996.980 1165.115 1996.985 ;
        RECT 1164.785 1996.970 1165.370 1996.980 ;
        RECT 1164.785 1996.670 1165.570 1996.970 ;
        RECT 1164.785 1996.660 1165.370 1996.670 ;
        RECT 1164.785 1996.655 1165.115 1996.660 ;
        RECT 2607.805 382.650 2608.135 382.665 ;
        RECT 2559.750 382.350 2608.135 382.650 ;
        RECT 1164.990 381.290 1165.370 381.300 ;
        RECT 1207.310 381.290 1207.690 381.300 ;
        RECT 2552.605 381.290 2552.935 381.305 ;
        RECT 2559.750 381.290 2560.050 382.350 ;
        RECT 2607.805 382.335 2608.135 382.350 ;
        RECT 2917.600 381.290 2924.800 381.740 ;
        RECT 1164.990 380.990 1207.690 381.290 ;
        RECT 1164.990 380.980 1165.370 380.990 ;
        RECT 1207.310 380.980 1207.690 380.990 ;
        RECT 1676.550 380.990 1724.690 381.290 ;
        RECT 1304.830 380.610 1305.210 380.620 ;
        RECT 1401.225 380.610 1401.555 380.625 ;
        RECT 1510.705 380.610 1511.035 380.625 ;
        RECT 1607.305 380.610 1607.635 380.625 ;
        RECT 1304.830 380.310 1401.555 380.610 ;
        RECT 1304.830 380.300 1305.210 380.310 ;
        RECT 1401.225 380.295 1401.555 380.310 ;
        RECT 1463.110 380.310 1511.035 380.610 ;
        RECT 1207.310 379.930 1207.690 379.940 ;
        RECT 1221.365 379.930 1221.695 379.945 ;
        RECT 1207.310 379.630 1221.695 379.930 ;
        RECT 1207.310 379.620 1207.690 379.630 ;
        RECT 1221.365 379.615 1221.695 379.630 ;
        RECT 1222.285 379.930 1222.615 379.945 ;
        RECT 1303.910 379.930 1304.290 379.940 ;
        RECT 1222.285 379.630 1304.290 379.930 ;
        RECT 1222.285 379.615 1222.615 379.630 ;
        RECT 1303.910 379.620 1304.290 379.630 ;
        RECT 1448.605 379.930 1448.935 379.945 ;
        RECT 1463.110 379.930 1463.410 380.310 ;
        RECT 1510.705 380.295 1511.035 380.310 ;
        RECT 1559.710 380.310 1607.635 380.610 ;
        RECT 1448.605 379.630 1463.410 379.930 ;
        RECT 1545.205 379.930 1545.535 379.945 ;
        RECT 1559.710 379.930 1560.010 380.310 ;
        RECT 1607.305 380.295 1607.635 380.310 ;
        RECT 1615.125 380.610 1615.455 380.625 ;
        RECT 1615.125 380.310 1655.690 380.610 ;
        RECT 1615.125 380.295 1615.455 380.310 ;
        RECT 1545.205 379.630 1560.010 379.930 ;
        RECT 1655.390 379.930 1655.690 380.310 ;
        RECT 1676.550 379.930 1676.850 380.990 ;
        RECT 1655.390 379.630 1676.850 379.930 ;
        RECT 1724.390 379.930 1724.690 380.990 ;
        RECT 1725.310 380.990 1773.450 381.290 ;
        RECT 1725.310 379.930 1725.610 380.990 ;
        RECT 1773.150 380.610 1773.450 380.990 ;
        RECT 1821.910 380.990 1870.050 381.290 ;
        RECT 1773.150 380.310 1821.290 380.610 ;
        RECT 1724.390 379.630 1725.610 379.930 ;
        RECT 1820.990 379.930 1821.290 380.310 ;
        RECT 1821.910 379.930 1822.210 380.990 ;
        RECT 1869.750 380.610 1870.050 380.990 ;
        RECT 1918.510 380.990 2029.210 381.290 ;
        RECT 1869.750 380.310 1917.890 380.610 ;
        RECT 1820.990 379.630 1822.210 379.930 ;
        RECT 1917.590 379.930 1917.890 380.310 ;
        RECT 1918.510 379.930 1918.810 380.990 ;
        RECT 2028.910 380.610 2029.210 380.990 ;
        RECT 2552.605 380.990 2560.050 381.290 ;
        RECT 2916.710 380.990 2924.800 381.290 ;
        RECT 2552.605 380.975 2552.935 380.990 ;
        RECT 2076.505 380.610 2076.835 380.625 ;
        RECT 2186.905 380.610 2187.235 380.625 ;
        RECT 2283.505 380.610 2283.835 380.625 ;
        RECT 2028.910 380.310 2076.835 380.610 ;
        RECT 2076.505 380.295 2076.835 380.310 ;
        RECT 2139.310 380.310 2187.235 380.610 ;
        RECT 1917.590 379.630 1918.810 379.930 ;
        RECT 2076.505 379.930 2076.835 379.945 ;
        RECT 2139.310 379.930 2139.610 380.310 ;
        RECT 2186.905 380.295 2187.235 380.310 ;
        RECT 2235.910 380.310 2283.835 380.610 ;
        RECT 2076.505 379.630 2139.610 379.930 ;
        RECT 2221.405 379.930 2221.735 379.945 ;
        RECT 2235.910 379.930 2236.210 380.310 ;
        RECT 2283.505 380.295 2283.835 380.310 ;
        RECT 2284.425 380.610 2284.755 380.625 ;
        RECT 2414.605 380.610 2414.935 380.625 ;
        RECT 2463.110 380.610 2463.490 380.620 ;
        RECT 2669.905 380.610 2670.235 380.625 ;
        RECT 2766.505 380.610 2766.835 380.625 ;
        RECT 2863.105 380.610 2863.435 380.625 ;
        RECT 2284.425 380.310 2331.890 380.610 ;
        RECT 2284.425 380.295 2284.755 380.310 ;
        RECT 2221.405 379.630 2236.210 379.930 ;
        RECT 2331.590 379.930 2331.890 380.310 ;
        RECT 2332.510 380.310 2414.935 380.610 ;
        RECT 2332.510 379.930 2332.810 380.310 ;
        RECT 2414.605 380.295 2414.935 380.310 ;
        RECT 2415.310 380.310 2463.490 380.610 ;
        RECT 2331.590 379.630 2332.810 379.930 ;
        RECT 2414.605 379.930 2414.935 379.945 ;
        RECT 2415.310 379.930 2415.610 380.310 ;
        RECT 2463.110 380.300 2463.490 380.310 ;
        RECT 2622.310 380.310 2670.235 380.610 ;
        RECT 2414.605 379.630 2415.610 379.930 ;
        RECT 2607.805 379.930 2608.135 379.945 ;
        RECT 2622.310 379.930 2622.610 380.310 ;
        RECT 2669.905 380.295 2670.235 380.310 ;
        RECT 2718.910 380.310 2766.835 380.610 ;
        RECT 2607.805 379.630 2622.610 379.930 ;
        RECT 2704.405 379.930 2704.735 379.945 ;
        RECT 2718.910 379.930 2719.210 380.310 ;
        RECT 2766.505 380.295 2766.835 380.310 ;
        RECT 2815.510 380.310 2863.435 380.610 ;
        RECT 2704.405 379.630 2719.210 379.930 ;
        RECT 2801.005 379.930 2801.335 379.945 ;
        RECT 2815.510 379.930 2815.810 380.310 ;
        RECT 2863.105 380.295 2863.435 380.310 ;
        RECT 2801.005 379.630 2815.810 379.930 ;
        RECT 2897.605 379.930 2897.935 379.945 ;
        RECT 2916.710 379.930 2917.010 380.990 ;
        RECT 2917.600 380.540 2924.800 380.990 ;
        RECT 2897.605 379.630 2917.010 379.930 ;
        RECT 1448.605 379.615 1448.935 379.630 ;
        RECT 1545.205 379.615 1545.535 379.630 ;
        RECT 2076.505 379.615 2076.835 379.630 ;
        RECT 2221.405 379.615 2221.735 379.630 ;
        RECT 2414.605 379.615 2414.935 379.630 ;
        RECT 2607.805 379.615 2608.135 379.630 ;
        RECT 2704.405 379.615 2704.735 379.630 ;
        RECT 2801.005 379.615 2801.335 379.630 ;
        RECT 2897.605 379.615 2897.935 379.630 ;
        RECT 2463.110 379.250 2463.490 379.260 ;
        RECT 2511.205 379.250 2511.535 379.265 ;
        RECT 2463.110 378.950 2511.535 379.250 ;
        RECT 2463.110 378.940 2463.490 378.950 ;
        RECT 2511.205 378.935 2511.535 378.950 ;
      LAYER via3 ;
        RECT 1165.020 1996.660 1165.340 1996.980 ;
        RECT 1165.020 380.980 1165.340 381.300 ;
        RECT 1207.340 380.980 1207.660 381.300 ;
        RECT 1304.860 380.300 1305.180 380.620 ;
        RECT 1207.340 379.620 1207.660 379.940 ;
        RECT 1303.940 379.620 1304.260 379.940 ;
        RECT 2463.140 380.300 2463.460 380.620 ;
        RECT 2463.140 378.940 2463.460 379.260 ;
      LAYER met4 ;
        RECT 1165.015 1996.655 1165.345 1996.985 ;
        RECT 1165.030 381.305 1165.330 1996.655 ;
        RECT 1165.015 380.975 1165.345 381.305 ;
        RECT 1207.335 380.975 1207.665 381.305 ;
        RECT 1207.350 379.945 1207.650 380.975 ;
        RECT 1304.855 380.295 1305.185 380.625 ;
        RECT 2463.135 380.295 2463.465 380.625 ;
        RECT 1207.335 379.615 1207.665 379.945 ;
        RECT 1303.935 379.615 1304.265 379.945 ;
        RECT 1303.950 379.250 1304.250 379.615 ;
        RECT 1304.870 379.250 1305.170 380.295 ;
        RECT 2463.150 379.265 2463.450 380.295 ;
        RECT 1303.950 378.950 1305.170 379.250 ;
        RECT 2463.135 378.935 2463.465 379.265 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1095.405 3429.325 1095.575 3477.435 ;
        RECT 1094.945 3332.765 1095.115 3380.875 ;
        RECT 1096.325 3236.205 1096.495 3284.315 ;
        RECT 1096.785 3084.225 1096.955 3132.675 ;
        RECT 1095.405 3043.425 1095.575 3057.195 ;
        RECT 1096.325 3007.725 1096.495 3042.915 ;
        RECT 1095.865 2946.525 1096.035 2994.635 ;
        RECT 1094.485 2849.625 1094.655 2898.075 ;
        RECT 1094.485 2753.065 1094.655 2767.175 ;
        RECT 1095.405 2525.265 1095.575 2552.975 ;
        RECT 1094.945 2221.985 1095.115 2270.095 ;
        RECT 1270.205 2009.485 1270.375 2010.335 ;
        RECT 1289.525 2009.485 1289.695 2013.735 ;
      LAYER mcon ;
        RECT 1095.405 3477.265 1095.575 3477.435 ;
        RECT 1094.945 3380.705 1095.115 3380.875 ;
        RECT 1096.325 3284.145 1096.495 3284.315 ;
        RECT 1096.785 3132.505 1096.955 3132.675 ;
        RECT 1095.405 3057.025 1095.575 3057.195 ;
        RECT 1096.325 3042.745 1096.495 3042.915 ;
        RECT 1095.865 2994.465 1096.035 2994.635 ;
        RECT 1094.485 2897.905 1094.655 2898.075 ;
        RECT 1094.485 2767.005 1094.655 2767.175 ;
        RECT 1095.405 2552.805 1095.575 2552.975 ;
        RECT 1094.945 2269.925 1095.115 2270.095 ;
        RECT 1289.525 2013.565 1289.695 2013.735 ;
        RECT 1270.205 2010.165 1270.375 2010.335 ;
      LAYER met1 ;
        RECT 1095.345 3477.420 1095.635 3477.465 ;
        RECT 1095.790 3477.420 1096.110 3477.480 ;
        RECT 1095.345 3477.280 1096.110 3477.420 ;
        RECT 1095.345 3477.235 1095.635 3477.280 ;
        RECT 1095.790 3477.220 1096.110 3477.280 ;
        RECT 1095.330 3429.480 1095.650 3429.540 ;
        RECT 1095.135 3429.340 1095.650 3429.480 ;
        RECT 1095.330 3429.280 1095.650 3429.340 ;
        RECT 1094.870 3380.860 1095.190 3380.920 ;
        RECT 1094.675 3380.720 1095.190 3380.860 ;
        RECT 1094.870 3380.660 1095.190 3380.720 ;
        RECT 1094.885 3332.920 1095.175 3332.965 ;
        RECT 1095.330 3332.920 1095.650 3332.980 ;
        RECT 1094.885 3332.780 1095.650 3332.920 ;
        RECT 1094.885 3332.735 1095.175 3332.780 ;
        RECT 1095.330 3332.720 1095.650 3332.780 ;
        RECT 1095.790 3298.240 1096.110 3298.300 ;
        RECT 1096.710 3298.240 1097.030 3298.300 ;
        RECT 1095.790 3298.100 1097.030 3298.240 ;
        RECT 1095.790 3298.040 1096.110 3298.100 ;
        RECT 1096.710 3298.040 1097.030 3298.100 ;
        RECT 1096.265 3284.300 1096.555 3284.345 ;
        RECT 1096.710 3284.300 1097.030 3284.360 ;
        RECT 1096.265 3284.160 1097.030 3284.300 ;
        RECT 1096.265 3284.115 1096.555 3284.160 ;
        RECT 1096.710 3284.100 1097.030 3284.160 ;
        RECT 1096.250 3236.360 1096.570 3236.420 ;
        RECT 1096.055 3236.220 1096.570 3236.360 ;
        RECT 1096.250 3236.160 1096.570 3236.220 ;
        RECT 1096.250 3202.020 1096.570 3202.080 ;
        RECT 1095.420 3201.880 1096.570 3202.020 ;
        RECT 1095.420 3201.400 1095.560 3201.880 ;
        RECT 1096.250 3201.820 1096.570 3201.880 ;
        RECT 1095.330 3201.140 1095.650 3201.400 ;
        RECT 1095.330 3187.740 1095.650 3187.800 ;
        RECT 1095.790 3187.740 1096.110 3187.800 ;
        RECT 1095.330 3187.600 1096.110 3187.740 ;
        RECT 1095.330 3187.540 1095.650 3187.600 ;
        RECT 1095.790 3187.540 1096.110 3187.600 ;
        RECT 1096.710 3132.660 1097.030 3132.720 ;
        RECT 1096.515 3132.520 1097.030 3132.660 ;
        RECT 1096.710 3132.460 1097.030 3132.520 ;
        RECT 1096.710 3084.380 1097.030 3084.440 ;
        RECT 1096.515 3084.240 1097.030 3084.380 ;
        RECT 1096.710 3084.180 1097.030 3084.240 ;
        RECT 1095.345 3057.180 1095.635 3057.225 ;
        RECT 1096.710 3057.180 1097.030 3057.240 ;
        RECT 1095.345 3057.040 1097.030 3057.180 ;
        RECT 1095.345 3056.995 1095.635 3057.040 ;
        RECT 1096.710 3056.980 1097.030 3057.040 ;
        RECT 1095.330 3043.580 1095.650 3043.640 ;
        RECT 1095.135 3043.440 1095.650 3043.580 ;
        RECT 1095.330 3043.380 1095.650 3043.440 ;
        RECT 1095.330 3042.900 1095.650 3042.960 ;
        RECT 1096.265 3042.900 1096.555 3042.945 ;
        RECT 1095.330 3042.760 1096.555 3042.900 ;
        RECT 1095.330 3042.700 1095.650 3042.760 ;
        RECT 1096.265 3042.715 1096.555 3042.760 ;
        RECT 1096.250 3007.880 1096.570 3007.940 ;
        RECT 1096.055 3007.740 1096.570 3007.880 ;
        RECT 1096.250 3007.680 1096.570 3007.740 ;
        RECT 1095.805 2994.620 1096.095 2994.665 ;
        RECT 1096.250 2994.620 1096.570 2994.680 ;
        RECT 1095.805 2994.480 1096.570 2994.620 ;
        RECT 1095.805 2994.435 1096.095 2994.480 ;
        RECT 1096.250 2994.420 1096.570 2994.480 ;
        RECT 1095.790 2946.680 1096.110 2946.740 ;
        RECT 1095.595 2946.540 1096.110 2946.680 ;
        RECT 1095.790 2946.480 1096.110 2946.540 ;
        RECT 1094.870 2912.000 1095.190 2912.060 ;
        RECT 1095.790 2912.000 1096.110 2912.060 ;
        RECT 1094.870 2911.860 1096.110 2912.000 ;
        RECT 1094.870 2911.800 1095.190 2911.860 ;
        RECT 1095.790 2911.800 1096.110 2911.860 ;
        RECT 1094.425 2898.060 1094.715 2898.105 ;
        RECT 1094.870 2898.060 1095.190 2898.120 ;
        RECT 1094.425 2897.920 1095.190 2898.060 ;
        RECT 1094.425 2897.875 1094.715 2897.920 ;
        RECT 1094.870 2897.860 1095.190 2897.920 ;
        RECT 1094.410 2849.780 1094.730 2849.840 ;
        RECT 1094.215 2849.640 1094.730 2849.780 ;
        RECT 1094.410 2849.580 1094.730 2849.640 ;
        RECT 1094.410 2815.240 1094.730 2815.500 ;
        RECT 1094.500 2814.760 1094.640 2815.240 ;
        RECT 1094.870 2814.760 1095.190 2814.820 ;
        RECT 1094.500 2814.620 1095.190 2814.760 ;
        RECT 1094.870 2814.560 1095.190 2814.620 ;
        RECT 1094.410 2767.160 1094.730 2767.220 ;
        RECT 1094.215 2767.020 1094.730 2767.160 ;
        RECT 1094.410 2766.960 1094.730 2767.020 ;
        RECT 1094.410 2753.220 1094.730 2753.280 ;
        RECT 1094.215 2753.080 1094.730 2753.220 ;
        RECT 1094.410 2753.020 1094.730 2753.080 ;
        RECT 1094.410 2718.680 1094.730 2718.940 ;
        RECT 1094.500 2718.200 1094.640 2718.680 ;
        RECT 1094.870 2718.200 1095.190 2718.260 ;
        RECT 1094.500 2718.060 1095.190 2718.200 ;
        RECT 1094.870 2718.000 1095.190 2718.060 ;
        RECT 1094.870 2621.640 1095.190 2621.700 ;
        RECT 1095.790 2621.640 1096.110 2621.700 ;
        RECT 1094.870 2621.500 1096.110 2621.640 ;
        RECT 1094.870 2621.440 1095.190 2621.500 ;
        RECT 1095.790 2621.440 1096.110 2621.500 ;
        RECT 1093.950 2573.360 1094.270 2573.420 ;
        RECT 1095.330 2573.360 1095.650 2573.420 ;
        RECT 1093.950 2573.220 1095.650 2573.360 ;
        RECT 1093.950 2573.160 1094.270 2573.220 ;
        RECT 1095.330 2573.160 1095.650 2573.220 ;
        RECT 1095.330 2552.960 1095.650 2553.020 ;
        RECT 1095.135 2552.820 1095.650 2552.960 ;
        RECT 1095.330 2552.760 1095.650 2552.820 ;
        RECT 1095.330 2525.420 1095.650 2525.480 ;
        RECT 1095.135 2525.280 1095.650 2525.420 ;
        RECT 1095.330 2525.220 1095.650 2525.280 ;
        RECT 1095.330 2463.540 1095.650 2463.600 ;
        RECT 1095.790 2463.540 1096.110 2463.600 ;
        RECT 1095.330 2463.400 1096.110 2463.540 ;
        RECT 1095.330 2463.340 1095.650 2463.400 ;
        RECT 1095.790 2463.340 1096.110 2463.400 ;
        RECT 1095.790 2429.000 1096.110 2429.260 ;
        RECT 1095.880 2428.520 1096.020 2429.000 ;
        RECT 1096.250 2428.520 1096.570 2428.580 ;
        RECT 1095.880 2428.380 1096.570 2428.520 ;
        RECT 1096.250 2428.320 1096.570 2428.380 ;
        RECT 1094.870 2332.100 1095.190 2332.360 ;
        RECT 1094.960 2331.620 1095.100 2332.100 ;
        RECT 1096.710 2331.620 1097.030 2331.680 ;
        RECT 1094.960 2331.480 1097.030 2331.620 ;
        RECT 1096.710 2331.420 1097.030 2331.480 ;
        RECT 1094.885 2270.080 1095.175 2270.125 ;
        RECT 1095.330 2270.080 1095.650 2270.140 ;
        RECT 1094.885 2269.940 1095.650 2270.080 ;
        RECT 1094.885 2269.895 1095.175 2269.940 ;
        RECT 1095.330 2269.880 1095.650 2269.940 ;
        RECT 1094.870 2222.140 1095.190 2222.200 ;
        RECT 1094.675 2222.000 1095.190 2222.140 ;
        RECT 1094.870 2221.940 1095.190 2222.000 ;
        RECT 1094.870 2173.520 1095.190 2173.580 ;
        RECT 1095.330 2173.520 1095.650 2173.580 ;
        RECT 1094.870 2173.380 1095.650 2173.520 ;
        RECT 1094.870 2173.320 1095.190 2173.380 ;
        RECT 1095.330 2173.320 1095.650 2173.380 ;
        RECT 1289.465 2013.720 1289.755 2013.765 ;
        RECT 1313.830 2013.720 1314.150 2013.780 ;
        RECT 1289.465 2013.580 1314.150 2013.720 ;
        RECT 1289.465 2013.535 1289.755 2013.580 ;
        RECT 1313.830 2013.520 1314.150 2013.580 ;
        RECT 1096.710 2010.320 1097.030 2010.380 ;
        RECT 1270.145 2010.320 1270.435 2010.365 ;
        RECT 1096.710 2010.180 1270.435 2010.320 ;
        RECT 1096.710 2010.120 1097.030 2010.180 ;
        RECT 1270.145 2010.135 1270.435 2010.180 ;
        RECT 1270.145 2009.640 1270.435 2009.685 ;
        RECT 1289.465 2009.640 1289.755 2009.685 ;
        RECT 1270.145 2009.500 1289.755 2009.640 ;
        RECT 1270.145 2009.455 1270.435 2009.500 ;
        RECT 1289.465 2009.455 1289.755 2009.500 ;
      LAYER via ;
        RECT 1095.820 3477.220 1096.080 3477.480 ;
        RECT 1095.360 3429.280 1095.620 3429.540 ;
        RECT 1094.900 3380.660 1095.160 3380.920 ;
        RECT 1095.360 3332.720 1095.620 3332.980 ;
        RECT 1095.820 3298.040 1096.080 3298.300 ;
        RECT 1096.740 3298.040 1097.000 3298.300 ;
        RECT 1096.740 3284.100 1097.000 3284.360 ;
        RECT 1096.280 3236.160 1096.540 3236.420 ;
        RECT 1096.280 3201.820 1096.540 3202.080 ;
        RECT 1095.360 3201.140 1095.620 3201.400 ;
        RECT 1095.360 3187.540 1095.620 3187.800 ;
        RECT 1095.820 3187.540 1096.080 3187.800 ;
        RECT 1096.740 3132.460 1097.000 3132.720 ;
        RECT 1096.740 3084.180 1097.000 3084.440 ;
        RECT 1096.740 3056.980 1097.000 3057.240 ;
        RECT 1095.360 3043.380 1095.620 3043.640 ;
        RECT 1095.360 3042.700 1095.620 3042.960 ;
        RECT 1096.280 3007.680 1096.540 3007.940 ;
        RECT 1096.280 2994.420 1096.540 2994.680 ;
        RECT 1095.820 2946.480 1096.080 2946.740 ;
        RECT 1094.900 2911.800 1095.160 2912.060 ;
        RECT 1095.820 2911.800 1096.080 2912.060 ;
        RECT 1094.900 2897.860 1095.160 2898.120 ;
        RECT 1094.440 2849.580 1094.700 2849.840 ;
        RECT 1094.440 2815.240 1094.700 2815.500 ;
        RECT 1094.900 2814.560 1095.160 2814.820 ;
        RECT 1094.440 2766.960 1094.700 2767.220 ;
        RECT 1094.440 2753.020 1094.700 2753.280 ;
        RECT 1094.440 2718.680 1094.700 2718.940 ;
        RECT 1094.900 2718.000 1095.160 2718.260 ;
        RECT 1094.900 2621.440 1095.160 2621.700 ;
        RECT 1095.820 2621.440 1096.080 2621.700 ;
        RECT 1093.980 2573.160 1094.240 2573.420 ;
        RECT 1095.360 2573.160 1095.620 2573.420 ;
        RECT 1095.360 2552.760 1095.620 2553.020 ;
        RECT 1095.360 2525.220 1095.620 2525.480 ;
        RECT 1095.360 2463.340 1095.620 2463.600 ;
        RECT 1095.820 2463.340 1096.080 2463.600 ;
        RECT 1095.820 2429.000 1096.080 2429.260 ;
        RECT 1096.280 2428.320 1096.540 2428.580 ;
        RECT 1094.900 2332.100 1095.160 2332.360 ;
        RECT 1096.740 2331.420 1097.000 2331.680 ;
        RECT 1095.360 2269.880 1095.620 2270.140 ;
        RECT 1094.900 2221.940 1095.160 2222.200 ;
        RECT 1094.900 2173.320 1095.160 2173.580 ;
        RECT 1095.360 2173.320 1095.620 2173.580 ;
        RECT 1313.860 2013.520 1314.120 2013.780 ;
        RECT 1096.740 2010.120 1097.000 2010.380 ;
      LAYER met2 ;
        RECT 1094.750 3517.600 1095.310 3524.800 ;
        RECT 1094.960 3517.370 1095.100 3517.600 ;
        RECT 1094.500 3517.230 1095.100 3517.370 ;
        RECT 1094.500 3478.725 1094.640 3517.230 ;
        RECT 1094.430 3478.355 1094.710 3478.725 ;
        RECT 1096.270 3477.930 1096.550 3478.045 ;
        RECT 1095.880 3477.790 1096.550 3477.930 ;
        RECT 1095.880 3477.510 1096.020 3477.790 ;
        RECT 1096.270 3477.675 1096.550 3477.790 ;
        RECT 1095.820 3477.190 1096.080 3477.510 ;
        RECT 1095.360 3429.250 1095.620 3429.570 ;
        RECT 1095.420 3394.970 1095.560 3429.250 ;
        RECT 1094.960 3394.830 1095.560 3394.970 ;
        RECT 1094.960 3380.950 1095.100 3394.830 ;
        RECT 1094.900 3380.630 1095.160 3380.950 ;
        RECT 1095.360 3332.690 1095.620 3333.010 ;
        RECT 1095.420 3298.410 1095.560 3332.690 ;
        RECT 1095.420 3298.330 1096.020 3298.410 ;
        RECT 1095.420 3298.270 1096.080 3298.330 ;
        RECT 1095.820 3298.010 1096.080 3298.270 ;
        RECT 1096.740 3298.010 1097.000 3298.330 ;
        RECT 1096.800 3284.390 1096.940 3298.010 ;
        RECT 1096.740 3284.070 1097.000 3284.390 ;
        RECT 1096.280 3236.130 1096.540 3236.450 ;
        RECT 1096.340 3202.110 1096.480 3236.130 ;
        RECT 1096.280 3201.790 1096.540 3202.110 ;
        RECT 1095.360 3201.110 1095.620 3201.430 ;
        RECT 1095.420 3187.830 1095.560 3201.110 ;
        RECT 1095.360 3187.510 1095.620 3187.830 ;
        RECT 1095.820 3187.510 1096.080 3187.830 ;
        RECT 1095.880 3152.890 1096.020 3187.510 ;
        RECT 1095.880 3152.750 1096.940 3152.890 ;
        RECT 1096.800 3132.750 1096.940 3152.750 ;
        RECT 1096.740 3132.430 1097.000 3132.750 ;
        RECT 1096.740 3084.150 1097.000 3084.470 ;
        RECT 1096.800 3057.270 1096.940 3084.150 ;
        RECT 1096.740 3056.950 1097.000 3057.270 ;
        RECT 1095.360 3043.350 1095.620 3043.670 ;
        RECT 1095.420 3042.990 1095.560 3043.350 ;
        RECT 1095.360 3042.670 1095.620 3042.990 ;
        RECT 1096.280 3007.650 1096.540 3007.970 ;
        RECT 1096.340 2994.710 1096.480 3007.650 ;
        RECT 1096.280 2994.390 1096.540 2994.710 ;
        RECT 1095.820 2946.450 1096.080 2946.770 ;
        RECT 1095.880 2912.090 1096.020 2946.450 ;
        RECT 1094.900 2911.770 1095.160 2912.090 ;
        RECT 1095.820 2911.770 1096.080 2912.090 ;
        RECT 1094.960 2898.150 1095.100 2911.770 ;
        RECT 1094.900 2897.830 1095.160 2898.150 ;
        RECT 1094.440 2849.550 1094.700 2849.870 ;
        RECT 1094.500 2815.530 1094.640 2849.550 ;
        RECT 1094.440 2815.210 1094.700 2815.530 ;
        RECT 1094.900 2814.530 1095.160 2814.850 ;
        RECT 1094.960 2801.330 1095.100 2814.530 ;
        RECT 1094.500 2801.190 1095.100 2801.330 ;
        RECT 1094.500 2767.250 1094.640 2801.190 ;
        RECT 1094.440 2766.930 1094.700 2767.250 ;
        RECT 1094.440 2752.990 1094.700 2753.310 ;
        RECT 1094.500 2718.970 1094.640 2752.990 ;
        RECT 1094.440 2718.650 1094.700 2718.970 ;
        RECT 1094.900 2717.970 1095.160 2718.290 ;
        RECT 1094.960 2704.885 1095.100 2717.970 ;
        RECT 1094.890 2704.515 1095.170 2704.885 ;
        RECT 1095.810 2704.515 1096.090 2704.885 ;
        RECT 1095.880 2669.410 1096.020 2704.515 ;
        RECT 1094.960 2669.270 1096.020 2669.410 ;
        RECT 1094.960 2656.605 1095.100 2669.270 ;
        RECT 1094.890 2656.235 1095.170 2656.605 ;
        RECT 1095.810 2656.235 1096.090 2656.605 ;
        RECT 1095.880 2621.730 1096.020 2656.235 ;
        RECT 1094.900 2621.410 1095.160 2621.730 ;
        RECT 1095.820 2621.410 1096.080 2621.730 ;
        RECT 1094.960 2608.325 1095.100 2621.410 ;
        RECT 1093.970 2607.955 1094.250 2608.325 ;
        RECT 1094.890 2607.955 1095.170 2608.325 ;
        RECT 1094.040 2573.450 1094.180 2607.955 ;
        RECT 1093.980 2573.130 1094.240 2573.450 ;
        RECT 1095.360 2573.130 1095.620 2573.450 ;
        RECT 1095.420 2553.050 1095.560 2573.130 ;
        RECT 1095.360 2552.730 1095.620 2553.050 ;
        RECT 1095.360 2525.190 1095.620 2525.510 ;
        RECT 1095.420 2463.630 1095.560 2525.190 ;
        RECT 1095.360 2463.310 1095.620 2463.630 ;
        RECT 1095.820 2463.310 1096.080 2463.630 ;
        RECT 1095.880 2429.290 1096.020 2463.310 ;
        RECT 1095.820 2428.970 1096.080 2429.290 ;
        RECT 1096.280 2428.290 1096.540 2428.610 ;
        RECT 1096.340 2366.925 1096.480 2428.290 ;
        RECT 1094.890 2366.555 1095.170 2366.925 ;
        RECT 1096.270 2366.555 1096.550 2366.925 ;
        RECT 1094.960 2332.390 1095.100 2366.555 ;
        RECT 1094.900 2332.070 1095.160 2332.390 ;
        RECT 1096.740 2331.390 1097.000 2331.710 ;
        RECT 1096.800 2283.850 1096.940 2331.390 ;
        RECT 1095.420 2283.710 1096.940 2283.850 ;
        RECT 1095.420 2270.170 1095.560 2283.710 ;
        RECT 1095.360 2269.850 1095.620 2270.170 ;
        RECT 1094.900 2221.910 1095.160 2222.230 ;
        RECT 1094.960 2187.290 1095.100 2221.910 ;
        RECT 1094.960 2187.150 1095.560 2187.290 ;
        RECT 1095.420 2173.610 1095.560 2187.150 ;
        RECT 1094.900 2173.290 1095.160 2173.610 ;
        RECT 1095.360 2173.290 1095.620 2173.610 ;
        RECT 1094.960 2125.525 1095.100 2173.290 ;
        RECT 1094.890 2125.155 1095.170 2125.525 ;
        RECT 1096.730 2125.155 1097.010 2125.525 ;
        RECT 1096.800 2010.410 1096.940 2125.155 ;
        RECT 1313.860 2013.490 1314.120 2013.810 ;
        RECT 1096.740 2010.090 1097.000 2010.410 ;
        RECT 1313.920 2000.000 1314.060 2013.490 ;
        RECT 1313.760 1999.540 1314.060 2000.000 ;
        RECT 1313.760 1996.000 1314.040 1999.540 ;
      LAYER via2 ;
        RECT 1094.430 3478.400 1094.710 3478.680 ;
        RECT 1096.270 3477.720 1096.550 3478.000 ;
        RECT 1094.890 2704.560 1095.170 2704.840 ;
        RECT 1095.810 2704.560 1096.090 2704.840 ;
        RECT 1094.890 2656.280 1095.170 2656.560 ;
        RECT 1095.810 2656.280 1096.090 2656.560 ;
        RECT 1093.970 2608.000 1094.250 2608.280 ;
        RECT 1094.890 2608.000 1095.170 2608.280 ;
        RECT 1094.890 2366.600 1095.170 2366.880 ;
        RECT 1096.270 2366.600 1096.550 2366.880 ;
        RECT 1094.890 2125.200 1095.170 2125.480 ;
        RECT 1096.730 2125.200 1097.010 2125.480 ;
      LAYER met3 ;
        RECT 1094.405 3478.690 1094.735 3478.705 ;
        RECT 1094.405 3478.390 1097.250 3478.690 ;
        RECT 1094.405 3478.375 1094.735 3478.390 ;
        RECT 1096.245 3478.010 1096.575 3478.025 ;
        RECT 1096.950 3478.010 1097.250 3478.390 ;
        RECT 1096.245 3477.710 1097.250 3478.010 ;
        RECT 1096.245 3477.695 1096.575 3477.710 ;
        RECT 1094.865 2704.850 1095.195 2704.865 ;
        RECT 1095.785 2704.850 1096.115 2704.865 ;
        RECT 1094.865 2704.550 1096.115 2704.850 ;
        RECT 1094.865 2704.535 1095.195 2704.550 ;
        RECT 1095.785 2704.535 1096.115 2704.550 ;
        RECT 1094.865 2656.570 1095.195 2656.585 ;
        RECT 1095.785 2656.570 1096.115 2656.585 ;
        RECT 1094.865 2656.270 1096.115 2656.570 ;
        RECT 1094.865 2656.255 1095.195 2656.270 ;
        RECT 1095.785 2656.255 1096.115 2656.270 ;
        RECT 1093.945 2608.290 1094.275 2608.305 ;
        RECT 1094.865 2608.290 1095.195 2608.305 ;
        RECT 1093.945 2607.990 1095.195 2608.290 ;
        RECT 1093.945 2607.975 1094.275 2607.990 ;
        RECT 1094.865 2607.975 1095.195 2607.990 ;
        RECT 1094.865 2366.890 1095.195 2366.905 ;
        RECT 1096.245 2366.890 1096.575 2366.905 ;
        RECT 1094.865 2366.590 1096.575 2366.890 ;
        RECT 1094.865 2366.575 1095.195 2366.590 ;
        RECT 1096.245 2366.575 1096.575 2366.590 ;
        RECT 1094.865 2125.490 1095.195 2125.505 ;
        RECT 1096.705 2125.490 1097.035 2125.505 ;
        RECT 1094.865 2125.190 1097.035 2125.490 ;
        RECT 1094.865 2125.175 1095.195 2125.190 ;
        RECT 1096.705 2125.175 1097.035 2125.190 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 771.565 3381.045 771.735 3429.155 ;
        RECT 771.565 2898.585 771.735 2946.355 ;
        RECT 772.025 2608.225 772.195 2656.335 ;
        RECT 772.025 2511.665 772.195 2559.775 ;
        RECT 771.105 2221.985 771.275 2270.095 ;
        RECT 1289.985 2009.485 1290.155 2011.015 ;
      LAYER mcon ;
        RECT 771.565 3428.985 771.735 3429.155 ;
        RECT 771.565 2946.185 771.735 2946.355 ;
        RECT 772.025 2656.165 772.195 2656.335 ;
        RECT 772.025 2559.605 772.195 2559.775 ;
        RECT 771.105 2269.925 771.275 2270.095 ;
        RECT 1289.985 2010.845 1290.155 2011.015 ;
      LAYER met1 ;
        RECT 770.570 3477.760 770.890 3477.820 ;
        RECT 771.030 3477.760 771.350 3477.820 ;
        RECT 770.570 3477.620 771.350 3477.760 ;
        RECT 770.570 3477.560 770.890 3477.620 ;
        RECT 771.030 3477.560 771.350 3477.620 ;
        RECT 771.030 3443.080 771.350 3443.140 ;
        RECT 771.950 3443.080 772.270 3443.140 ;
        RECT 771.030 3442.940 772.270 3443.080 ;
        RECT 771.030 3442.880 771.350 3442.940 ;
        RECT 771.950 3442.880 772.270 3442.940 ;
        RECT 771.505 3429.140 771.795 3429.185 ;
        RECT 771.950 3429.140 772.270 3429.200 ;
        RECT 771.505 3429.000 772.270 3429.140 ;
        RECT 771.505 3428.955 771.795 3429.000 ;
        RECT 771.950 3428.940 772.270 3429.000 ;
        RECT 771.490 3381.200 771.810 3381.260 ;
        RECT 771.295 3381.060 771.810 3381.200 ;
        RECT 771.490 3381.000 771.810 3381.060 ;
        RECT 771.490 3367.600 771.810 3367.660 ;
        RECT 772.410 3367.600 772.730 3367.660 ;
        RECT 771.490 3367.460 772.730 3367.600 ;
        RECT 771.490 3367.400 771.810 3367.460 ;
        RECT 772.410 3367.400 772.730 3367.460 ;
        RECT 771.490 3270.700 771.810 3270.760 ;
        RECT 772.410 3270.700 772.730 3270.760 ;
        RECT 771.490 3270.560 772.730 3270.700 ;
        RECT 771.490 3270.500 771.810 3270.560 ;
        RECT 772.410 3270.500 772.730 3270.560 ;
        RECT 771.490 3174.140 771.810 3174.200 ;
        RECT 772.410 3174.140 772.730 3174.200 ;
        RECT 771.490 3174.000 772.730 3174.140 ;
        RECT 771.490 3173.940 771.810 3174.000 ;
        RECT 772.410 3173.940 772.730 3174.000 ;
        RECT 771.490 3077.580 771.810 3077.640 ;
        RECT 772.410 3077.580 772.730 3077.640 ;
        RECT 771.490 3077.440 772.730 3077.580 ;
        RECT 771.490 3077.380 771.810 3077.440 ;
        RECT 772.410 3077.380 772.730 3077.440 ;
        RECT 771.490 2981.020 771.810 2981.080 ;
        RECT 772.410 2981.020 772.730 2981.080 ;
        RECT 771.490 2980.880 772.730 2981.020 ;
        RECT 771.490 2980.820 771.810 2980.880 ;
        RECT 772.410 2980.820 772.730 2980.880 ;
        RECT 771.490 2946.340 771.810 2946.400 ;
        RECT 771.295 2946.200 771.810 2946.340 ;
        RECT 771.490 2946.140 771.810 2946.200 ;
        RECT 771.490 2898.740 771.810 2898.800 ;
        RECT 771.295 2898.600 771.810 2898.740 ;
        RECT 771.490 2898.540 771.810 2898.600 ;
        RECT 771.030 2898.060 771.350 2898.120 ;
        RECT 771.950 2898.060 772.270 2898.120 ;
        RECT 771.030 2897.920 772.270 2898.060 ;
        RECT 771.030 2897.860 771.350 2897.920 ;
        RECT 771.950 2897.860 772.270 2897.920 ;
        RECT 771.030 2814.760 771.350 2814.820 ;
        RECT 771.950 2814.760 772.270 2814.820 ;
        RECT 771.030 2814.620 772.270 2814.760 ;
        RECT 771.030 2814.560 771.350 2814.620 ;
        RECT 771.950 2814.560 772.270 2814.620 ;
        RECT 771.950 2656.320 772.270 2656.380 ;
        RECT 771.755 2656.180 772.270 2656.320 ;
        RECT 771.950 2656.120 772.270 2656.180 ;
        RECT 771.965 2608.380 772.255 2608.425 ;
        RECT 772.410 2608.380 772.730 2608.440 ;
        RECT 771.965 2608.240 772.730 2608.380 ;
        RECT 771.965 2608.195 772.255 2608.240 ;
        RECT 772.410 2608.180 772.730 2608.240 ;
        RECT 771.950 2559.760 772.270 2559.820 ;
        RECT 771.755 2559.620 772.270 2559.760 ;
        RECT 771.950 2559.560 772.270 2559.620 ;
        RECT 771.965 2511.820 772.255 2511.865 ;
        RECT 772.410 2511.820 772.730 2511.880 ;
        RECT 771.965 2511.680 772.730 2511.820 ;
        RECT 771.965 2511.635 772.255 2511.680 ;
        RECT 772.410 2511.620 772.730 2511.680 ;
        RECT 771.030 2463.200 771.350 2463.260 ;
        RECT 771.950 2463.200 772.270 2463.260 ;
        RECT 771.030 2463.060 772.270 2463.200 ;
        RECT 771.030 2463.000 771.350 2463.060 ;
        RECT 771.950 2463.000 772.270 2463.060 ;
        RECT 771.490 2332.300 771.810 2332.360 ;
        RECT 772.410 2332.300 772.730 2332.360 ;
        RECT 771.490 2332.160 772.730 2332.300 ;
        RECT 771.490 2332.100 771.810 2332.160 ;
        RECT 772.410 2332.100 772.730 2332.160 ;
        RECT 771.045 2270.080 771.335 2270.125 ;
        RECT 771.490 2270.080 771.810 2270.140 ;
        RECT 771.045 2269.940 771.810 2270.080 ;
        RECT 771.045 2269.895 771.335 2269.940 ;
        RECT 771.490 2269.880 771.810 2269.940 ;
        RECT 771.030 2222.140 771.350 2222.200 ;
        RECT 770.835 2222.000 771.350 2222.140 ;
        RECT 771.030 2221.940 771.350 2222.000 ;
        RECT 771.490 2138.980 771.810 2139.240 ;
        RECT 771.580 2138.840 771.720 2138.980 ;
        RECT 771.950 2138.840 772.270 2138.900 ;
        RECT 771.580 2138.700 772.270 2138.840 ;
        RECT 771.950 2138.640 772.270 2138.700 ;
        RECT 770.570 2125.240 770.890 2125.300 ;
        RECT 771.950 2125.240 772.270 2125.300 ;
        RECT 770.570 2125.100 772.270 2125.240 ;
        RECT 770.570 2125.040 770.890 2125.100 ;
        RECT 771.950 2125.040 772.270 2125.100 ;
        RECT 772.410 2042.420 772.730 2042.680 ;
        RECT 772.500 2042.000 772.640 2042.420 ;
        RECT 772.410 2041.740 772.730 2042.000 ;
        RECT 772.410 2011.000 772.730 2011.060 ;
        RECT 1289.925 2011.000 1290.215 2011.045 ;
        RECT 772.410 2010.860 1290.215 2011.000 ;
        RECT 772.410 2010.800 772.730 2010.860 ;
        RECT 1289.925 2010.815 1290.215 2010.860 ;
        RECT 1289.925 2009.640 1290.215 2009.685 ;
        RECT 1321.650 2009.640 1321.970 2009.700 ;
        RECT 1289.925 2009.500 1321.970 2009.640 ;
        RECT 1289.925 2009.455 1290.215 2009.500 ;
        RECT 1321.650 2009.440 1321.970 2009.500 ;
      LAYER via ;
        RECT 770.600 3477.560 770.860 3477.820 ;
        RECT 771.060 3477.560 771.320 3477.820 ;
        RECT 771.060 3442.880 771.320 3443.140 ;
        RECT 771.980 3442.880 772.240 3443.140 ;
        RECT 771.980 3428.940 772.240 3429.200 ;
        RECT 771.520 3381.000 771.780 3381.260 ;
        RECT 771.520 3367.400 771.780 3367.660 ;
        RECT 772.440 3367.400 772.700 3367.660 ;
        RECT 771.520 3270.500 771.780 3270.760 ;
        RECT 772.440 3270.500 772.700 3270.760 ;
        RECT 771.520 3173.940 771.780 3174.200 ;
        RECT 772.440 3173.940 772.700 3174.200 ;
        RECT 771.520 3077.380 771.780 3077.640 ;
        RECT 772.440 3077.380 772.700 3077.640 ;
        RECT 771.520 2980.820 771.780 2981.080 ;
        RECT 772.440 2980.820 772.700 2981.080 ;
        RECT 771.520 2946.140 771.780 2946.400 ;
        RECT 771.520 2898.540 771.780 2898.800 ;
        RECT 771.060 2897.860 771.320 2898.120 ;
        RECT 771.980 2897.860 772.240 2898.120 ;
        RECT 771.060 2814.560 771.320 2814.820 ;
        RECT 771.980 2814.560 772.240 2814.820 ;
        RECT 771.980 2656.120 772.240 2656.380 ;
        RECT 772.440 2608.180 772.700 2608.440 ;
        RECT 771.980 2559.560 772.240 2559.820 ;
        RECT 772.440 2511.620 772.700 2511.880 ;
        RECT 771.060 2463.000 771.320 2463.260 ;
        RECT 771.980 2463.000 772.240 2463.260 ;
        RECT 771.520 2332.100 771.780 2332.360 ;
        RECT 772.440 2332.100 772.700 2332.360 ;
        RECT 771.520 2269.880 771.780 2270.140 ;
        RECT 771.060 2221.940 771.320 2222.200 ;
        RECT 771.520 2138.980 771.780 2139.240 ;
        RECT 771.980 2138.640 772.240 2138.900 ;
        RECT 770.600 2125.040 770.860 2125.300 ;
        RECT 771.980 2125.040 772.240 2125.300 ;
        RECT 772.440 2042.420 772.700 2042.680 ;
        RECT 772.440 2041.740 772.700 2042.000 ;
        RECT 772.440 2010.800 772.700 2011.060 ;
        RECT 1321.680 2009.440 1321.940 2009.700 ;
      LAYER met2 ;
        RECT 770.450 3517.600 771.010 3524.800 ;
        RECT 770.660 3477.850 770.800 3517.600 ;
        RECT 770.600 3477.530 770.860 3477.850 ;
        RECT 771.060 3477.530 771.320 3477.850 ;
        RECT 771.120 3443.170 771.260 3477.530 ;
        RECT 771.060 3442.850 771.320 3443.170 ;
        RECT 771.980 3442.850 772.240 3443.170 ;
        RECT 772.040 3429.230 772.180 3442.850 ;
        RECT 771.980 3428.910 772.240 3429.230 ;
        RECT 771.520 3380.970 771.780 3381.290 ;
        RECT 771.580 3367.690 771.720 3380.970 ;
        RECT 771.520 3367.370 771.780 3367.690 ;
        RECT 772.440 3367.370 772.700 3367.690 ;
        RECT 772.500 3318.810 772.640 3367.370 ;
        RECT 771.580 3318.670 772.640 3318.810 ;
        RECT 771.580 3270.790 771.720 3318.670 ;
        RECT 771.520 3270.470 771.780 3270.790 ;
        RECT 772.440 3270.470 772.700 3270.790 ;
        RECT 772.500 3222.250 772.640 3270.470 ;
        RECT 771.580 3222.110 772.640 3222.250 ;
        RECT 771.580 3174.230 771.720 3222.110 ;
        RECT 771.520 3173.910 771.780 3174.230 ;
        RECT 772.440 3173.910 772.700 3174.230 ;
        RECT 772.500 3125.690 772.640 3173.910 ;
        RECT 771.580 3125.550 772.640 3125.690 ;
        RECT 771.580 3077.670 771.720 3125.550 ;
        RECT 771.520 3077.350 771.780 3077.670 ;
        RECT 772.440 3077.350 772.700 3077.670 ;
        RECT 772.500 3029.130 772.640 3077.350 ;
        RECT 771.580 3028.990 772.640 3029.130 ;
        RECT 771.580 2981.110 771.720 3028.990 ;
        RECT 771.520 2980.790 771.780 2981.110 ;
        RECT 772.440 2980.850 772.700 2981.110 ;
        RECT 772.040 2980.790 772.700 2980.850 ;
        RECT 772.040 2980.710 772.640 2980.790 ;
        RECT 772.040 2959.770 772.180 2980.710 ;
        RECT 771.580 2959.630 772.180 2959.770 ;
        RECT 771.580 2946.430 771.720 2959.630 ;
        RECT 771.520 2946.110 771.780 2946.430 ;
        RECT 771.520 2898.570 771.780 2898.830 ;
        RECT 771.120 2898.510 771.780 2898.570 ;
        RECT 771.120 2898.430 771.720 2898.510 ;
        RECT 771.120 2898.150 771.260 2898.430 ;
        RECT 771.060 2897.830 771.320 2898.150 ;
        RECT 771.980 2897.830 772.240 2898.150 ;
        RECT 772.040 2814.850 772.180 2897.830 ;
        RECT 771.060 2814.530 771.320 2814.850 ;
        RECT 771.980 2814.530 772.240 2814.850 ;
        RECT 771.120 2766.650 771.260 2814.530 ;
        RECT 771.120 2766.510 771.720 2766.650 ;
        RECT 771.580 2719.050 771.720 2766.510 ;
        RECT 771.580 2718.910 772.640 2719.050 ;
        RECT 772.500 2670.090 772.640 2718.910 ;
        RECT 772.040 2669.950 772.640 2670.090 ;
        RECT 772.040 2656.410 772.180 2669.950 ;
        RECT 771.980 2656.090 772.240 2656.410 ;
        RECT 772.440 2608.150 772.700 2608.470 ;
        RECT 772.500 2573.530 772.640 2608.150 ;
        RECT 772.040 2573.390 772.640 2573.530 ;
        RECT 772.040 2559.850 772.180 2573.390 ;
        RECT 771.980 2559.530 772.240 2559.850 ;
        RECT 772.440 2511.590 772.700 2511.910 ;
        RECT 772.500 2476.970 772.640 2511.590 ;
        RECT 772.040 2476.830 772.640 2476.970 ;
        RECT 772.040 2463.290 772.180 2476.830 ;
        RECT 771.060 2462.970 771.320 2463.290 ;
        RECT 771.980 2462.970 772.240 2463.290 ;
        RECT 771.120 2415.205 771.260 2462.970 ;
        RECT 771.050 2414.835 771.330 2415.205 ;
        RECT 772.430 2414.835 772.710 2415.205 ;
        RECT 772.500 2380.410 772.640 2414.835 ;
        RECT 771.580 2380.270 772.640 2380.410 ;
        RECT 771.580 2332.390 771.720 2380.270 ;
        RECT 771.520 2332.070 771.780 2332.390 ;
        RECT 772.440 2332.070 772.700 2332.390 ;
        RECT 772.500 2283.850 772.640 2332.070 ;
        RECT 771.580 2283.710 772.640 2283.850 ;
        RECT 771.580 2270.170 771.720 2283.710 ;
        RECT 771.520 2269.850 771.780 2270.170 ;
        RECT 771.060 2221.910 771.320 2222.230 ;
        RECT 771.120 2187.290 771.260 2221.910 ;
        RECT 771.120 2187.150 771.720 2187.290 ;
        RECT 771.580 2139.270 771.720 2187.150 ;
        RECT 771.520 2138.950 771.780 2139.270 ;
        RECT 771.980 2138.610 772.240 2138.930 ;
        RECT 772.040 2125.330 772.180 2138.610 ;
        RECT 770.600 2125.010 770.860 2125.330 ;
        RECT 771.980 2125.010 772.240 2125.330 ;
        RECT 770.660 2077.245 770.800 2125.010 ;
        RECT 770.590 2076.875 770.870 2077.245 ;
        RECT 771.510 2076.875 771.790 2077.245 ;
        RECT 771.580 2076.565 771.720 2076.875 ;
        RECT 771.510 2076.195 771.790 2076.565 ;
        RECT 772.430 2076.195 772.710 2076.565 ;
        RECT 772.500 2042.710 772.640 2076.195 ;
        RECT 772.440 2042.390 772.700 2042.710 ;
        RECT 772.440 2041.710 772.700 2042.030 ;
        RECT 772.500 2011.090 772.640 2041.710 ;
        RECT 772.440 2010.770 772.700 2011.090 ;
        RECT 1321.680 2009.410 1321.940 2009.730 ;
        RECT 1321.740 2000.000 1321.880 2009.410 ;
        RECT 1321.580 1999.540 1321.880 2000.000 ;
        RECT 1321.580 1996.000 1321.860 1999.540 ;
      LAYER via2 ;
        RECT 771.050 2414.880 771.330 2415.160 ;
        RECT 772.430 2414.880 772.710 2415.160 ;
        RECT 770.590 2076.920 770.870 2077.200 ;
        RECT 771.510 2076.920 771.790 2077.200 ;
        RECT 771.510 2076.240 771.790 2076.520 ;
        RECT 772.430 2076.240 772.710 2076.520 ;
      LAYER met3 ;
        RECT 771.025 2415.170 771.355 2415.185 ;
        RECT 772.405 2415.170 772.735 2415.185 ;
        RECT 771.025 2414.870 772.735 2415.170 ;
        RECT 771.025 2414.855 771.355 2414.870 ;
        RECT 772.405 2414.855 772.735 2414.870 ;
        RECT 770.565 2077.210 770.895 2077.225 ;
        RECT 771.485 2077.210 771.815 2077.225 ;
        RECT 770.565 2076.910 771.815 2077.210 ;
        RECT 770.565 2076.895 770.895 2076.910 ;
        RECT 771.485 2076.895 771.815 2076.910 ;
        RECT 771.485 2076.530 771.815 2076.545 ;
        RECT 772.405 2076.530 772.735 2076.545 ;
        RECT 771.485 2076.230 772.735 2076.530 ;
        RECT 771.485 2076.215 771.815 2076.230 ;
        RECT 772.405 2076.215 772.735 2076.230 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 445.810 3498.500 446.130 3498.560 ;
        RECT 448.110 3498.500 448.430 3498.560 ;
        RECT 445.810 3498.360 448.430 3498.500 ;
        RECT 445.810 3498.300 446.130 3498.360 ;
        RECT 448.110 3498.300 448.430 3498.360 ;
        RECT 448.110 2014.400 448.430 2014.460 ;
        RECT 448.110 2014.260 1274.500 2014.400 ;
        RECT 448.110 2014.200 448.430 2014.260 ;
        RECT 1274.360 2014.060 1274.500 2014.260 ;
        RECT 1329.470 2014.060 1329.790 2014.120 ;
        RECT 1274.360 2013.920 1329.790 2014.060 ;
        RECT 1329.470 2013.860 1329.790 2013.920 ;
      LAYER via ;
        RECT 445.840 3498.300 446.100 3498.560 ;
        RECT 448.140 3498.300 448.400 3498.560 ;
        RECT 448.140 2014.200 448.400 2014.460 ;
        RECT 1329.500 2013.860 1329.760 2014.120 ;
      LAYER met2 ;
        RECT 445.690 3517.600 446.250 3524.800 ;
        RECT 445.900 3498.590 446.040 3517.600 ;
        RECT 445.840 3498.270 446.100 3498.590 ;
        RECT 448.140 3498.270 448.400 3498.590 ;
        RECT 448.200 2014.490 448.340 3498.270 ;
        RECT 448.140 2014.170 448.400 2014.490 ;
        RECT 1329.500 2013.830 1329.760 2014.150 ;
        RECT 1329.560 2000.000 1329.700 2013.830 ;
        RECT 1329.400 1999.540 1329.700 2000.000 ;
        RECT 1329.400 1996.000 1329.680 1999.540 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 528.685 2013.565 530.695 2013.735 ;
        RECT 1270.665 2010.165 1270.835 2013.735 ;
        RECT 1297.345 2010.165 1298.435 2010.335 ;
      LAYER mcon ;
        RECT 530.525 2013.565 530.695 2013.735 ;
        RECT 1270.665 2013.565 1270.835 2013.735 ;
        RECT 1298.265 2010.165 1298.435 2010.335 ;
      LAYER met1 ;
        RECT 121.510 3498.500 121.830 3498.560 ;
        RECT 123.810 3498.500 124.130 3498.560 ;
        RECT 121.510 3498.360 124.130 3498.500 ;
        RECT 121.510 3498.300 121.830 3498.360 ;
        RECT 123.810 3498.300 124.130 3498.360 ;
        RECT 123.810 2013.720 124.130 2013.780 ;
        RECT 528.625 2013.720 528.915 2013.765 ;
        RECT 123.810 2013.580 528.915 2013.720 ;
        RECT 123.810 2013.520 124.130 2013.580 ;
        RECT 528.625 2013.535 528.915 2013.580 ;
        RECT 530.465 2013.720 530.755 2013.765 ;
        RECT 1270.605 2013.720 1270.895 2013.765 ;
        RECT 530.465 2013.580 1270.895 2013.720 ;
        RECT 530.465 2013.535 530.755 2013.580 ;
        RECT 1270.605 2013.535 1270.895 2013.580 ;
        RECT 1270.605 2010.320 1270.895 2010.365 ;
        RECT 1297.285 2010.320 1297.575 2010.365 ;
        RECT 1270.605 2010.180 1297.575 2010.320 ;
        RECT 1270.605 2010.135 1270.895 2010.180 ;
        RECT 1297.285 2010.135 1297.575 2010.180 ;
        RECT 1298.205 2010.320 1298.495 2010.365 ;
        RECT 1337.750 2010.320 1338.070 2010.380 ;
        RECT 1298.205 2010.180 1338.070 2010.320 ;
        RECT 1298.205 2010.135 1298.495 2010.180 ;
        RECT 1337.750 2010.120 1338.070 2010.180 ;
      LAYER via ;
        RECT 121.540 3498.300 121.800 3498.560 ;
        RECT 123.840 3498.300 124.100 3498.560 ;
        RECT 123.840 2013.520 124.100 2013.780 ;
        RECT 1337.780 2010.120 1338.040 2010.380 ;
      LAYER met2 ;
        RECT 121.390 3517.600 121.950 3524.800 ;
        RECT 121.600 3498.590 121.740 3517.600 ;
        RECT 121.540 3498.270 121.800 3498.590 ;
        RECT 123.840 3498.270 124.100 3498.590 ;
        RECT 123.900 2013.810 124.040 3498.270 ;
        RECT 123.840 2013.490 124.100 2013.810 ;
        RECT 1337.780 2010.090 1338.040 2010.410 ;
        RECT 1337.840 2000.000 1337.980 2010.090 ;
        RECT 1337.680 1999.540 1337.980 2000.000 ;
        RECT 1337.680 1996.000 1337.960 1999.540 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 17.550 2012.700 17.870 2012.760 ;
        RECT 1345.570 2012.700 1345.890 2012.760 ;
        RECT 17.550 2012.560 1345.890 2012.700 ;
        RECT 17.550 2012.500 17.870 2012.560 ;
        RECT 1345.570 2012.500 1345.890 2012.560 ;
      LAYER via ;
        RECT 17.580 2012.500 17.840 2012.760 ;
        RECT 1345.600 2012.500 1345.860 2012.760 ;
      LAYER met2 ;
        RECT 17.570 3339.635 17.850 3340.005 ;
        RECT 17.640 2012.790 17.780 3339.635 ;
        RECT 17.580 2012.470 17.840 2012.790 ;
        RECT 1345.600 2012.470 1345.860 2012.790 ;
        RECT 1345.660 2000.000 1345.800 2012.470 ;
        RECT 1345.500 1999.540 1345.800 2000.000 ;
        RECT 1345.500 1996.000 1345.780 1999.540 ;
      LAYER via2 ;
        RECT 17.570 3339.680 17.850 3339.960 ;
      LAYER met3 ;
        RECT -4.800 3339.970 2.400 3340.420 ;
        RECT 17.545 3339.970 17.875 3339.985 ;
        RECT -4.800 3339.670 17.875 3339.970 ;
        RECT -4.800 3339.220 2.400 3339.670 ;
        RECT 17.545 3339.655 17.875 3339.670 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 18.470 2012.020 18.790 2012.080 ;
        RECT 1353.390 2012.020 1353.710 2012.080 ;
        RECT 18.470 2011.880 1353.710 2012.020 ;
        RECT 18.470 2011.820 18.790 2011.880 ;
        RECT 1353.390 2011.820 1353.710 2011.880 ;
      LAYER via ;
        RECT 18.500 2011.820 18.760 2012.080 ;
        RECT 1353.420 2011.820 1353.680 2012.080 ;
      LAYER met2 ;
        RECT 18.490 3051.995 18.770 3052.365 ;
        RECT 18.560 2012.110 18.700 3051.995 ;
        RECT 18.500 2011.790 18.760 2012.110 ;
        RECT 1353.420 2011.790 1353.680 2012.110 ;
        RECT 1353.480 2000.000 1353.620 2011.790 ;
        RECT 1353.320 1999.540 1353.620 2000.000 ;
        RECT 1353.320 1996.000 1353.600 1999.540 ;
      LAYER via2 ;
        RECT 18.490 3052.040 18.770 3052.320 ;
      LAYER met3 ;
        RECT -4.800 3052.330 2.400 3052.780 ;
        RECT 18.465 3052.330 18.795 3052.345 ;
        RECT -4.800 3052.030 18.795 3052.330 ;
        RECT -4.800 3051.580 2.400 3052.030 ;
        RECT 18.465 3052.015 18.795 3052.030 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 14.790 2760.360 15.110 2760.420 ;
        RECT 1314.290 2760.360 1314.610 2760.420 ;
        RECT 14.790 2760.220 1314.610 2760.360 ;
        RECT 14.790 2760.160 15.110 2760.220 ;
        RECT 1314.290 2760.160 1314.610 2760.220 ;
        RECT 1314.290 2010.660 1314.610 2010.720 ;
        RECT 1361.210 2010.660 1361.530 2010.720 ;
        RECT 1314.290 2010.520 1361.530 2010.660 ;
        RECT 1314.290 2010.460 1314.610 2010.520 ;
        RECT 1361.210 2010.460 1361.530 2010.520 ;
      LAYER via ;
        RECT 14.820 2760.160 15.080 2760.420 ;
        RECT 1314.320 2760.160 1314.580 2760.420 ;
        RECT 1314.320 2010.460 1314.580 2010.720 ;
        RECT 1361.240 2010.460 1361.500 2010.720 ;
      LAYER met2 ;
        RECT 14.810 2765.035 15.090 2765.405 ;
        RECT 14.880 2760.450 15.020 2765.035 ;
        RECT 14.820 2760.130 15.080 2760.450 ;
        RECT 1314.320 2760.130 1314.580 2760.450 ;
        RECT 1314.380 2010.750 1314.520 2760.130 ;
        RECT 1314.320 2010.430 1314.580 2010.750 ;
        RECT 1361.240 2010.430 1361.500 2010.750 ;
        RECT 1361.300 2000.000 1361.440 2010.430 ;
        RECT 1361.140 1999.540 1361.440 2000.000 ;
        RECT 1361.140 1996.000 1361.420 1999.540 ;
      LAYER via2 ;
        RECT 14.810 2765.080 15.090 2765.360 ;
      LAYER met3 ;
        RECT -4.800 2765.370 2.400 2765.820 ;
        RECT 14.785 2765.370 15.115 2765.385 ;
        RECT -4.800 2765.070 15.115 2765.370 ;
        RECT -4.800 2764.620 2.400 2765.070 ;
        RECT 14.785 2765.055 15.115 2765.070 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.630 2477.480 16.950 2477.540 ;
        RECT 1321.190 2477.480 1321.510 2477.540 ;
        RECT 16.630 2477.340 1321.510 2477.480 ;
        RECT 16.630 2477.280 16.950 2477.340 ;
        RECT 1321.190 2477.280 1321.510 2477.340 ;
        RECT 1321.190 2014.740 1321.510 2014.800 ;
        RECT 1369.030 2014.740 1369.350 2014.800 ;
        RECT 1321.190 2014.600 1369.350 2014.740 ;
        RECT 1321.190 2014.540 1321.510 2014.600 ;
        RECT 1369.030 2014.540 1369.350 2014.600 ;
      LAYER via ;
        RECT 16.660 2477.280 16.920 2477.540 ;
        RECT 1321.220 2477.280 1321.480 2477.540 ;
        RECT 1321.220 2014.540 1321.480 2014.800 ;
        RECT 1369.060 2014.540 1369.320 2014.800 ;
      LAYER met2 ;
        RECT 16.650 2477.395 16.930 2477.765 ;
        RECT 16.660 2477.250 16.920 2477.395 ;
        RECT 1321.220 2477.250 1321.480 2477.570 ;
        RECT 1321.280 2014.830 1321.420 2477.250 ;
        RECT 1321.220 2014.510 1321.480 2014.830 ;
        RECT 1369.060 2014.510 1369.320 2014.830 ;
        RECT 1369.120 2000.000 1369.260 2014.510 ;
        RECT 1368.960 1999.540 1369.260 2000.000 ;
        RECT 1368.960 1996.000 1369.240 1999.540 ;
      LAYER via2 ;
        RECT 16.650 2477.440 16.930 2477.720 ;
      LAYER met3 ;
        RECT -4.800 2477.730 2.400 2478.180 ;
        RECT 16.625 2477.730 16.955 2477.745 ;
        RECT -4.800 2477.430 16.955 2477.730 ;
        RECT -4.800 2476.980 2.400 2477.430 ;
        RECT 16.625 2477.415 16.955 2477.430 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 14.790 2187.460 15.110 2187.520 ;
        RECT 1328.090 2187.460 1328.410 2187.520 ;
        RECT 14.790 2187.320 1328.410 2187.460 ;
        RECT 14.790 2187.260 15.110 2187.320 ;
        RECT 1328.090 2187.260 1328.410 2187.320 ;
        RECT 1328.090 2014.400 1328.410 2014.460 ;
        RECT 1376.850 2014.400 1377.170 2014.460 ;
        RECT 1328.090 2014.260 1377.170 2014.400 ;
        RECT 1328.090 2014.200 1328.410 2014.260 ;
        RECT 1376.850 2014.200 1377.170 2014.260 ;
      LAYER via ;
        RECT 14.820 2187.260 15.080 2187.520 ;
        RECT 1328.120 2187.260 1328.380 2187.520 ;
        RECT 1328.120 2014.200 1328.380 2014.460 ;
        RECT 1376.880 2014.200 1377.140 2014.460 ;
      LAYER met2 ;
        RECT 14.810 2189.755 15.090 2190.125 ;
        RECT 14.880 2187.550 15.020 2189.755 ;
        RECT 14.820 2187.230 15.080 2187.550 ;
        RECT 1328.120 2187.230 1328.380 2187.550 ;
        RECT 1328.180 2014.490 1328.320 2187.230 ;
        RECT 1328.120 2014.170 1328.380 2014.490 ;
        RECT 1376.880 2014.170 1377.140 2014.490 ;
        RECT 1376.940 2000.000 1377.080 2014.170 ;
        RECT 1376.780 1999.540 1377.080 2000.000 ;
        RECT 1376.780 1996.000 1377.060 1999.540 ;
      LAYER via2 ;
        RECT 14.810 2189.800 15.090 2190.080 ;
      LAYER met3 ;
        RECT -4.800 2190.090 2.400 2190.540 ;
        RECT 14.785 2190.090 15.115 2190.105 ;
        RECT -4.800 2189.790 15.115 2190.090 ;
        RECT -4.800 2189.340 2.400 2189.790 ;
        RECT 14.785 2189.775 15.115 2189.790 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1361.745 2009.485 1361.915 2010.335 ;
      LAYER mcon ;
        RECT 1361.745 2010.165 1361.915 2010.335 ;
      LAYER met1 ;
        RECT 1361.685 2010.320 1361.975 2010.365 ;
        RECT 1385.130 2010.320 1385.450 2010.380 ;
        RECT 1361.685 2010.180 1385.450 2010.320 ;
        RECT 1361.685 2010.135 1361.975 2010.180 ;
        RECT 1385.130 2010.120 1385.450 2010.180 ;
        RECT 1324.870 2009.640 1325.190 2009.700 ;
        RECT 1361.685 2009.640 1361.975 2009.685 ;
        RECT 1324.870 2009.500 1361.975 2009.640 ;
        RECT 1324.870 2009.440 1325.190 2009.500 ;
        RECT 1361.685 2009.455 1361.975 2009.500 ;
        RECT 17.090 1997.400 17.410 1997.460 ;
        RECT 1324.870 1997.400 1325.190 1997.460 ;
        RECT 17.090 1997.260 1325.190 1997.400 ;
        RECT 17.090 1997.200 17.410 1997.260 ;
        RECT 1324.870 1997.200 1325.190 1997.260 ;
      LAYER via ;
        RECT 1385.160 2010.120 1385.420 2010.380 ;
        RECT 1324.900 2009.440 1325.160 2009.700 ;
        RECT 17.120 1997.200 17.380 1997.460 ;
        RECT 1324.900 1997.200 1325.160 1997.460 ;
      LAYER met2 ;
        RECT 1385.160 2010.090 1385.420 2010.410 ;
        RECT 1324.900 2009.410 1325.160 2009.730 ;
        RECT 1324.960 1997.490 1325.100 2009.410 ;
        RECT 1385.220 2000.000 1385.360 2010.090 ;
        RECT 1385.060 1999.540 1385.360 2000.000 ;
        RECT 17.120 1997.170 17.380 1997.490 ;
        RECT 1324.900 1997.170 1325.160 1997.490 ;
        RECT 17.180 1903.165 17.320 1997.170 ;
        RECT 1385.060 1996.000 1385.340 1999.540 ;
        RECT 17.110 1902.795 17.390 1903.165 ;
      LAYER via2 ;
        RECT 17.110 1902.840 17.390 1903.120 ;
      LAYER met3 ;
        RECT -4.800 1903.130 2.400 1903.580 ;
        RECT 17.085 1903.130 17.415 1903.145 ;
        RECT -4.800 1902.830 17.415 1903.130 ;
        RECT -4.800 1902.380 2.400 1902.830 ;
        RECT 17.085 1902.815 17.415 1902.830 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1548.890 620.740 1549.210 620.800 ;
        RECT 2900.830 620.740 2901.150 620.800 ;
        RECT 1548.890 620.600 2901.150 620.740 ;
        RECT 1548.890 620.540 1549.210 620.600 ;
        RECT 2900.830 620.540 2901.150 620.600 ;
      LAYER via ;
        RECT 1548.920 620.540 1549.180 620.800 ;
        RECT 2900.860 620.540 2901.120 620.800 ;
      LAYER met2 ;
        RECT 1170.330 1996.890 1170.610 1997.005 ;
        RECT 1171.620 1996.890 1171.900 2000.000 ;
        RECT 1170.330 1996.750 1171.900 1996.890 ;
        RECT 1170.330 1996.635 1170.610 1996.750 ;
        RECT 1171.620 1996.000 1171.900 1996.750 ;
        RECT 1548.910 1693.355 1549.190 1693.725 ;
        RECT 1548.980 620.830 1549.120 1693.355 ;
        RECT 1548.920 620.510 1549.180 620.830 ;
        RECT 2900.860 620.510 2901.120 620.830 ;
        RECT 2900.920 615.925 2901.060 620.510 ;
        RECT 2900.850 615.555 2901.130 615.925 ;
      LAYER via2 ;
        RECT 1170.330 1996.680 1170.610 1996.960 ;
        RECT 1548.910 1693.400 1549.190 1693.680 ;
        RECT 2900.850 615.600 2901.130 615.880 ;
      LAYER met3 ;
        RECT 1169.590 1996.970 1169.970 1996.980 ;
        RECT 1170.305 1996.970 1170.635 1996.985 ;
        RECT 1169.590 1996.670 1170.635 1996.970 ;
        RECT 1169.590 1996.660 1169.970 1996.670 ;
        RECT 1170.305 1996.655 1170.635 1996.670 ;
        RECT 1169.590 1693.690 1169.970 1693.700 ;
        RECT 1548.885 1693.690 1549.215 1693.705 ;
        RECT 1169.590 1693.390 1549.215 1693.690 ;
        RECT 1169.590 1693.380 1169.970 1693.390 ;
        RECT 1548.885 1693.375 1549.215 1693.390 ;
        RECT 2900.825 615.890 2901.155 615.905 ;
        RECT 2917.600 615.890 2924.800 616.340 ;
        RECT 2900.825 615.590 2924.800 615.890 ;
        RECT 2900.825 615.575 2901.155 615.590 ;
        RECT 2917.600 615.140 2924.800 615.590 ;
      LAYER via3 ;
        RECT 1169.620 1996.660 1169.940 1996.980 ;
        RECT 1169.620 1693.380 1169.940 1693.700 ;
      LAYER met4 ;
        RECT 1169.615 1996.655 1169.945 1996.985 ;
        RECT 1169.630 1693.705 1169.930 1996.655 ;
        RECT 1169.615 1693.375 1169.945 1693.705 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 16.630 2008.960 16.950 2009.020 ;
        RECT 1392.950 2008.960 1393.270 2009.020 ;
        RECT 16.630 2008.820 1393.270 2008.960 ;
        RECT 16.630 2008.760 16.950 2008.820 ;
        RECT 1392.950 2008.760 1393.270 2008.820 ;
      LAYER via ;
        RECT 16.660 2008.760 16.920 2009.020 ;
        RECT 1392.980 2008.760 1393.240 2009.020 ;
      LAYER met2 ;
        RECT 16.660 2008.730 16.920 2009.050 ;
        RECT 1392.980 2008.730 1393.240 2009.050 ;
        RECT 16.720 1615.525 16.860 2008.730 ;
        RECT 1393.040 2000.000 1393.180 2008.730 ;
        RECT 1392.880 1999.540 1393.180 2000.000 ;
        RECT 1392.880 1996.000 1393.160 1999.540 ;
        RECT 16.650 1615.155 16.930 1615.525 ;
      LAYER via2 ;
        RECT 16.650 1615.200 16.930 1615.480 ;
      LAYER met3 ;
        RECT -4.800 1615.490 2.400 1615.940 ;
        RECT 16.625 1615.490 16.955 1615.505 ;
        RECT -4.800 1615.190 16.955 1615.490 ;
        RECT -4.800 1614.740 2.400 1615.190 ;
        RECT 16.625 1615.175 16.955 1615.190 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 19.850 2008.620 20.170 2008.680 ;
        RECT 1400.770 2008.620 1401.090 2008.680 ;
        RECT 19.850 2008.480 1401.090 2008.620 ;
        RECT 19.850 2008.420 20.170 2008.480 ;
        RECT 1400.770 2008.420 1401.090 2008.480 ;
      LAYER via ;
        RECT 19.880 2008.420 20.140 2008.680 ;
        RECT 1400.800 2008.420 1401.060 2008.680 ;
      LAYER met2 ;
        RECT 19.880 2008.390 20.140 2008.710 ;
        RECT 1400.800 2008.390 1401.060 2008.710 ;
        RECT 19.940 1400.645 20.080 2008.390 ;
        RECT 1400.860 2000.000 1401.000 2008.390 ;
        RECT 1400.700 1999.540 1401.000 2000.000 ;
        RECT 1400.700 1996.000 1400.980 1999.540 ;
        RECT 19.870 1400.275 20.150 1400.645 ;
      LAYER via2 ;
        RECT 19.870 1400.320 20.150 1400.600 ;
      LAYER met3 ;
        RECT -4.800 1400.610 2.400 1401.060 ;
        RECT 19.845 1400.610 20.175 1400.625 ;
        RECT -4.800 1400.310 20.175 1400.610 ;
        RECT -4.800 1399.860 2.400 1400.310 ;
        RECT 19.845 1400.295 20.175 1400.310 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 18.930 2008.280 19.250 2008.340 ;
        RECT 1408.590 2008.280 1408.910 2008.340 ;
        RECT 18.930 2008.140 1408.910 2008.280 ;
        RECT 18.930 2008.080 19.250 2008.140 ;
        RECT 1408.590 2008.080 1408.910 2008.140 ;
      LAYER via ;
        RECT 18.960 2008.080 19.220 2008.340 ;
        RECT 1408.620 2008.080 1408.880 2008.340 ;
      LAYER met2 ;
        RECT 18.960 2008.050 19.220 2008.370 ;
        RECT 1408.620 2008.050 1408.880 2008.370 ;
        RECT 19.020 1185.085 19.160 2008.050 ;
        RECT 1408.680 2000.000 1408.820 2008.050 ;
        RECT 1408.520 1999.540 1408.820 2000.000 ;
        RECT 1408.520 1996.000 1408.800 1999.540 ;
        RECT 18.950 1184.715 19.230 1185.085 ;
      LAYER via2 ;
        RECT 18.950 1184.760 19.230 1185.040 ;
      LAYER met3 ;
        RECT -4.800 1185.050 2.400 1185.500 ;
        RECT 18.925 1185.050 19.255 1185.065 ;
        RECT -4.800 1184.750 19.255 1185.050 ;
        RECT -4.800 1184.300 2.400 1184.750 ;
        RECT 18.925 1184.735 19.255 1184.750 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1415.050 1996.890 1415.330 1997.005 ;
        RECT 1416.340 1996.890 1416.620 2000.000 ;
        RECT 1415.050 1996.750 1416.620 1996.890 ;
        RECT 1415.050 1996.635 1415.330 1996.750 ;
        RECT 1416.340 1996.000 1416.620 1996.750 ;
        RECT 17.570 972.555 17.850 972.925 ;
        RECT 17.640 969.525 17.780 972.555 ;
        RECT 17.570 969.155 17.850 969.525 ;
      LAYER via2 ;
        RECT 1415.050 1996.680 1415.330 1996.960 ;
        RECT 17.570 972.600 17.850 972.880 ;
        RECT 17.570 969.200 17.850 969.480 ;
      LAYER met3 ;
        RECT 1414.310 1996.970 1414.690 1996.980 ;
        RECT 1415.025 1996.970 1415.355 1996.985 ;
        RECT 1414.310 1996.670 1415.355 1996.970 ;
        RECT 1414.310 1996.660 1414.690 1996.670 ;
        RECT 1415.025 1996.655 1415.355 1996.670 ;
        RECT 17.545 972.890 17.875 972.905 ;
        RECT 1414.310 972.890 1414.690 972.900 ;
        RECT 17.545 972.590 1414.690 972.890 ;
        RECT 17.545 972.575 17.875 972.590 ;
        RECT 1414.310 972.580 1414.690 972.590 ;
        RECT -4.800 969.490 2.400 969.940 ;
        RECT 17.545 969.490 17.875 969.505 ;
        RECT -4.800 969.190 17.875 969.490 ;
        RECT -4.800 968.740 2.400 969.190 ;
        RECT 17.545 969.175 17.875 969.190 ;
      LAYER via3 ;
        RECT 1414.340 1996.660 1414.660 1996.980 ;
        RECT 1414.340 972.580 1414.660 972.900 ;
      LAYER met4 ;
        RECT 1414.335 1996.655 1414.665 1996.985 ;
        RECT 1414.350 972.905 1414.650 1996.655 ;
        RECT 1414.335 972.575 1414.665 972.905 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1422.410 1996.890 1422.690 1997.005 ;
        RECT 1424.160 1996.890 1424.440 2000.000 ;
        RECT 1422.410 1996.750 1424.440 1996.890 ;
        RECT 1422.410 1996.635 1422.690 1996.750 ;
        RECT 1424.160 1996.000 1424.440 1996.750 ;
        RECT 17.570 758.355 17.850 758.725 ;
        RECT 17.640 753.965 17.780 758.355 ;
        RECT 17.570 753.595 17.850 753.965 ;
      LAYER via2 ;
        RECT 1422.410 1996.680 1422.690 1996.960 ;
        RECT 17.570 758.400 17.850 758.680 ;
        RECT 17.570 753.640 17.850 753.920 ;
      LAYER met3 ;
        RECT 1421.670 1996.970 1422.050 1996.980 ;
        RECT 1422.385 1996.970 1422.715 1996.985 ;
        RECT 1421.670 1996.670 1422.715 1996.970 ;
        RECT 1421.670 1996.660 1422.050 1996.670 ;
        RECT 1422.385 1996.655 1422.715 1996.670 ;
        RECT 17.545 758.690 17.875 758.705 ;
        RECT 1421.670 758.690 1422.050 758.700 ;
        RECT 17.545 758.390 1422.050 758.690 ;
        RECT 17.545 758.375 17.875 758.390 ;
        RECT 1421.670 758.380 1422.050 758.390 ;
        RECT -4.800 753.930 2.400 754.380 ;
        RECT 17.545 753.930 17.875 753.945 ;
        RECT -4.800 753.630 17.875 753.930 ;
        RECT -4.800 753.180 2.400 753.630 ;
        RECT 17.545 753.615 17.875 753.630 ;
      LAYER via3 ;
        RECT 1421.700 1996.660 1422.020 1996.980 ;
        RECT 1421.700 758.380 1422.020 758.700 ;
      LAYER met4 ;
        RECT 1421.695 1996.655 1422.025 1996.985 ;
        RECT 1421.710 758.705 1422.010 1996.655 ;
        RECT 1421.695 758.375 1422.025 758.705 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1430.690 1996.890 1430.970 1997.005 ;
        RECT 1431.980 1996.890 1432.260 2000.000 ;
        RECT 1430.690 1996.750 1432.260 1996.890 ;
        RECT 1430.690 1996.635 1430.970 1996.750 ;
        RECT 1431.980 1996.000 1432.260 1996.750 ;
        RECT 17.570 544.835 17.850 545.205 ;
        RECT 17.640 538.405 17.780 544.835 ;
        RECT 17.570 538.035 17.850 538.405 ;
      LAYER via2 ;
        RECT 1430.690 1996.680 1430.970 1996.960 ;
        RECT 17.570 544.880 17.850 545.160 ;
        RECT 17.570 538.080 17.850 538.360 ;
      LAYER met3 ;
        RECT 1428.110 1996.970 1428.490 1996.980 ;
        RECT 1430.665 1996.970 1430.995 1996.985 ;
        RECT 1428.110 1996.670 1430.995 1996.970 ;
        RECT 1428.110 1996.660 1428.490 1996.670 ;
        RECT 1430.665 1996.655 1430.995 1996.670 ;
        RECT 17.545 545.170 17.875 545.185 ;
        RECT 1428.110 545.170 1428.490 545.180 ;
        RECT 17.545 544.870 1428.490 545.170 ;
        RECT 17.545 544.855 17.875 544.870 ;
        RECT 1428.110 544.860 1428.490 544.870 ;
        RECT -4.800 538.370 2.400 538.820 ;
        RECT 17.545 538.370 17.875 538.385 ;
        RECT -4.800 538.070 17.875 538.370 ;
        RECT -4.800 537.620 2.400 538.070 ;
        RECT 17.545 538.055 17.875 538.070 ;
      LAYER via3 ;
        RECT 1428.140 1996.660 1428.460 1996.980 ;
        RECT 1428.140 544.860 1428.460 545.180 ;
      LAYER met4 ;
        RECT 1428.135 1996.655 1428.465 1996.985 ;
        RECT 1428.150 545.185 1428.450 1996.655 ;
        RECT 1428.135 544.855 1428.465 545.185 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1438.970 1996.890 1439.250 1997.005 ;
        RECT 1440.260 1996.890 1440.540 2000.000 ;
        RECT 1438.970 1996.750 1440.540 1996.890 ;
        RECT 1438.970 1996.635 1439.250 1996.750 ;
        RECT 1440.260 1996.000 1440.540 1996.750 ;
      LAYER via2 ;
        RECT 1438.970 1996.680 1439.250 1996.960 ;
      LAYER met3 ;
        RECT 1435.470 1996.970 1435.850 1996.980 ;
        RECT 1438.945 1996.970 1439.275 1996.985 ;
        RECT 1435.470 1996.670 1439.275 1996.970 ;
        RECT 1435.470 1996.660 1435.850 1996.670 ;
        RECT 1438.945 1996.655 1439.275 1996.670 ;
        RECT 1435.470 324.170 1435.850 324.180 ;
        RECT 3.070 323.870 1435.850 324.170 ;
        RECT -4.800 322.810 2.400 323.260 ;
        RECT 3.070 322.810 3.370 323.870 ;
        RECT 1435.470 323.860 1435.850 323.870 ;
        RECT -4.800 322.510 3.370 322.810 ;
        RECT -4.800 322.060 2.400 322.510 ;
      LAYER via3 ;
        RECT 1435.500 1996.660 1435.820 1996.980 ;
        RECT 1435.500 323.860 1435.820 324.180 ;
      LAYER met4 ;
        RECT 1435.495 1996.655 1435.825 1996.985 ;
        RECT 1435.510 324.185 1435.810 1996.655 ;
        RECT 1435.495 323.855 1435.825 324.185 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1448.170 2008.875 1448.450 2009.245 ;
        RECT 1448.240 2000.000 1448.380 2008.875 ;
        RECT 1448.080 1999.540 1448.380 2000.000 ;
        RECT 1448.080 1996.000 1448.360 1999.540 ;
        RECT 17.110 1679.755 17.390 1680.125 ;
        RECT 17.180 107.285 17.320 1679.755 ;
        RECT 17.110 106.915 17.390 107.285 ;
      LAYER via2 ;
        RECT 1448.170 2008.920 1448.450 2009.200 ;
        RECT 17.110 1679.800 17.390 1680.080 ;
        RECT 17.110 106.960 17.390 107.240 ;
      LAYER met3 ;
        RECT 1314.030 2009.210 1314.410 2009.220 ;
        RECT 1448.145 2009.210 1448.475 2009.225 ;
        RECT 1314.030 2008.910 1448.475 2009.210 ;
        RECT 1314.030 2008.900 1314.410 2008.910 ;
        RECT 1448.145 2008.895 1448.475 2008.910 ;
        RECT 17.085 1680.090 17.415 1680.105 ;
        RECT 1314.030 1680.090 1314.410 1680.100 ;
        RECT 17.085 1679.790 1314.410 1680.090 ;
        RECT 17.085 1679.775 17.415 1679.790 ;
        RECT 1314.030 1679.780 1314.410 1679.790 ;
        RECT -4.800 107.250 2.400 107.700 ;
        RECT 17.085 107.250 17.415 107.265 ;
        RECT -4.800 106.950 17.415 107.250 ;
        RECT -4.800 106.500 2.400 106.950 ;
        RECT 17.085 106.935 17.415 106.950 ;
      LAYER via3 ;
        RECT 1314.060 2008.900 1314.380 2009.220 ;
        RECT 1314.060 1679.780 1314.380 1680.100 ;
      LAYER met4 ;
        RECT 1314.055 2008.895 1314.385 2009.225 ;
        RECT 1314.070 1680.105 1314.370 2008.895 ;
        RECT 1314.055 1679.775 1314.385 1680.105 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 2425.190 855.340 2425.510 855.400 ;
        RECT 2900.830 855.340 2901.150 855.400 ;
        RECT 2425.190 855.200 2901.150 855.340 ;
        RECT 2425.190 855.140 2425.510 855.200 ;
        RECT 2900.830 855.140 2901.150 855.200 ;
      LAYER via ;
        RECT 2425.220 855.140 2425.480 855.400 ;
        RECT 2900.860 855.140 2901.120 855.400 ;
      LAYER met2 ;
        RECT 1179.070 2009.555 1179.350 2009.925 ;
        RECT 2425.210 2009.555 2425.490 2009.925 ;
        RECT 1179.140 1999.610 1179.280 2009.555 ;
        RECT 1179.440 1999.610 1179.720 2000.000 ;
        RECT 1179.140 1999.470 1179.720 1999.610 ;
        RECT 1179.440 1996.000 1179.720 1999.470 ;
        RECT 2425.280 855.430 2425.420 2009.555 ;
        RECT 2425.220 855.110 2425.480 855.430 ;
        RECT 2900.860 855.110 2901.120 855.430 ;
        RECT 2900.920 850.525 2901.060 855.110 ;
        RECT 2900.850 850.155 2901.130 850.525 ;
      LAYER via2 ;
        RECT 1179.070 2009.600 1179.350 2009.880 ;
        RECT 2425.210 2009.600 2425.490 2009.880 ;
        RECT 2900.850 850.200 2901.130 850.480 ;
      LAYER met3 ;
        RECT 1179.045 2009.890 1179.375 2009.905 ;
        RECT 2425.185 2009.890 2425.515 2009.905 ;
        RECT 1179.045 2009.590 2425.515 2009.890 ;
        RECT 1179.045 2009.575 1179.375 2009.590 ;
        RECT 2425.185 2009.575 2425.515 2009.590 ;
        RECT 2900.825 850.490 2901.155 850.505 ;
        RECT 2917.600 850.490 2924.800 850.940 ;
        RECT 2900.825 850.190 2924.800 850.490 ;
        RECT 2900.825 850.175 2901.155 850.190 ;
        RECT 2917.600 849.740 2924.800 850.190 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1562.690 1089.940 1563.010 1090.000 ;
        RECT 2900.830 1089.940 2901.150 1090.000 ;
        RECT 1562.690 1089.800 2901.150 1089.940 ;
        RECT 1562.690 1089.740 1563.010 1089.800 ;
        RECT 2900.830 1089.740 2901.150 1089.800 ;
      LAYER via ;
        RECT 1562.720 1089.740 1562.980 1090.000 ;
        RECT 2900.860 1089.740 2901.120 1090.000 ;
      LAYER met2 ;
        RECT 1187.720 1996.890 1188.000 2000.000 ;
        RECT 1189.190 1996.890 1189.470 1997.005 ;
        RECT 1187.720 1996.750 1189.470 1996.890 ;
        RECT 1187.720 1996.000 1188.000 1996.750 ;
        RECT 1189.190 1996.635 1189.470 1996.750 ;
        RECT 1562.710 1700.155 1562.990 1700.525 ;
        RECT 1562.780 1090.030 1562.920 1700.155 ;
        RECT 1562.720 1089.710 1562.980 1090.030 ;
        RECT 2900.860 1089.710 2901.120 1090.030 ;
        RECT 2900.920 1085.125 2901.060 1089.710 ;
        RECT 2900.850 1084.755 2901.130 1085.125 ;
      LAYER via2 ;
        RECT 1189.190 1996.680 1189.470 1996.960 ;
        RECT 1562.710 1700.200 1562.990 1700.480 ;
        RECT 2900.850 1084.800 2901.130 1085.080 ;
      LAYER met3 ;
        RECT 1189.165 1996.970 1189.495 1996.985 ;
        RECT 1190.750 1996.970 1191.130 1996.980 ;
        RECT 1189.165 1996.670 1191.130 1996.970 ;
        RECT 1189.165 1996.655 1189.495 1996.670 ;
        RECT 1190.750 1996.660 1191.130 1996.670 ;
        RECT 1190.750 1700.490 1191.130 1700.500 ;
        RECT 1562.685 1700.490 1563.015 1700.505 ;
        RECT 1190.750 1700.190 1563.015 1700.490 ;
        RECT 1190.750 1700.180 1191.130 1700.190 ;
        RECT 1562.685 1700.175 1563.015 1700.190 ;
        RECT 2900.825 1085.090 2901.155 1085.105 ;
        RECT 2917.600 1085.090 2924.800 1085.540 ;
        RECT 2900.825 1084.790 2924.800 1085.090 ;
        RECT 2900.825 1084.775 2901.155 1084.790 ;
        RECT 2917.600 1084.340 2924.800 1084.790 ;
      LAYER via3 ;
        RECT 1190.780 1996.660 1191.100 1996.980 ;
        RECT 1190.780 1700.180 1191.100 1700.500 ;
      LAYER met4 ;
        RECT 1190.775 1996.655 1191.105 1996.985 ;
        RECT 1190.790 1700.505 1191.090 1996.655 ;
        RECT 1190.775 1700.175 1191.105 1700.505 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1576.490 1324.540 1576.810 1324.600 ;
        RECT 2900.830 1324.540 2901.150 1324.600 ;
        RECT 1576.490 1324.400 2901.150 1324.540 ;
        RECT 1576.490 1324.340 1576.810 1324.400 ;
        RECT 2900.830 1324.340 2901.150 1324.400 ;
      LAYER via ;
        RECT 1576.520 1324.340 1576.780 1324.600 ;
        RECT 2900.860 1324.340 2901.120 1324.600 ;
      LAYER met2 ;
        RECT 1195.540 1996.890 1195.820 2000.000 ;
        RECT 1197.010 1996.890 1197.290 1997.005 ;
        RECT 1195.540 1996.750 1197.290 1996.890 ;
        RECT 1195.540 1996.000 1195.820 1996.750 ;
        RECT 1197.010 1996.635 1197.290 1996.750 ;
        RECT 1576.510 1694.035 1576.790 1694.405 ;
        RECT 1576.580 1324.630 1576.720 1694.035 ;
        RECT 1576.520 1324.310 1576.780 1324.630 ;
        RECT 2900.860 1324.310 2901.120 1324.630 ;
        RECT 2900.920 1319.725 2901.060 1324.310 ;
        RECT 2900.850 1319.355 2901.130 1319.725 ;
      LAYER via2 ;
        RECT 1197.010 1996.680 1197.290 1996.960 ;
        RECT 1576.510 1694.080 1576.790 1694.360 ;
        RECT 2900.850 1319.400 2901.130 1319.680 ;
      LAYER met3 ;
        RECT 1196.985 1996.970 1197.315 1996.985 ;
        RECT 1199.950 1996.970 1200.330 1996.980 ;
        RECT 1196.985 1996.670 1200.330 1996.970 ;
        RECT 1196.985 1996.655 1197.315 1996.670 ;
        RECT 1199.950 1996.660 1200.330 1996.670 ;
        RECT 1199.950 1694.370 1200.330 1694.380 ;
        RECT 1576.485 1694.370 1576.815 1694.385 ;
        RECT 1199.950 1694.070 1576.815 1694.370 ;
        RECT 1199.950 1694.060 1200.330 1694.070 ;
        RECT 1576.485 1694.055 1576.815 1694.070 ;
        RECT 2900.825 1319.690 2901.155 1319.705 ;
        RECT 2917.600 1319.690 2924.800 1320.140 ;
        RECT 2900.825 1319.390 2924.800 1319.690 ;
        RECT 2900.825 1319.375 2901.155 1319.390 ;
        RECT 2917.600 1318.940 2924.800 1319.390 ;
      LAYER via3 ;
        RECT 1199.980 1996.660 1200.300 1996.980 ;
        RECT 1199.980 1694.060 1200.300 1694.380 ;
      LAYER met4 ;
        RECT 1199.975 1996.655 1200.305 1996.985 ;
        RECT 1199.990 1694.385 1200.290 1996.655 ;
        RECT 1199.975 1694.055 1200.305 1694.385 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1497.830 1554.040 1498.150 1554.100 ;
        RECT 1521.750 1554.040 1522.070 1554.100 ;
        RECT 1497.830 1553.900 1522.070 1554.040 ;
        RECT 1497.830 1553.840 1498.150 1553.900 ;
        RECT 1521.750 1553.840 1522.070 1553.900 ;
        RECT 1603.630 1554.040 1603.950 1554.100 ;
        RECT 1641.810 1554.040 1642.130 1554.100 ;
        RECT 1603.630 1553.900 1642.130 1554.040 ;
        RECT 1603.630 1553.840 1603.950 1553.900 ;
        RECT 1641.810 1553.840 1642.130 1553.900 ;
        RECT 1798.210 1554.040 1798.530 1554.100 ;
        RECT 1835.010 1554.040 1835.330 1554.100 ;
        RECT 1798.210 1553.900 1835.330 1554.040 ;
        RECT 1798.210 1553.840 1798.530 1553.900 ;
        RECT 1835.010 1553.840 1835.330 1553.900 ;
        RECT 2377.810 1554.040 2378.130 1554.100 ;
        RECT 2414.610 1554.040 2414.930 1554.100 ;
        RECT 2377.810 1553.900 2414.930 1554.040 ;
        RECT 2377.810 1553.840 2378.130 1553.900 ;
        RECT 2414.610 1553.840 2414.930 1553.900 ;
        RECT 2705.330 1554.040 2705.650 1554.100 ;
        RECT 2719.130 1554.040 2719.450 1554.100 ;
        RECT 2705.330 1553.900 2719.450 1554.040 ;
        RECT 2705.330 1553.840 2705.650 1553.900 ;
        RECT 2719.130 1553.840 2719.450 1553.900 ;
        RECT 1441.710 1553.700 1442.030 1553.760 ;
        RECT 1483.110 1553.700 1483.430 1553.760 ;
        RECT 1441.710 1553.560 1483.430 1553.700 ;
        RECT 1441.710 1553.500 1442.030 1553.560 ;
        RECT 1483.110 1553.500 1483.430 1553.560 ;
        RECT 1703.910 1553.700 1704.230 1553.760 ;
        RECT 1738.410 1553.700 1738.730 1553.760 ;
        RECT 1703.910 1553.560 1738.730 1553.700 ;
        RECT 1703.910 1553.500 1704.230 1553.560 ;
        RECT 1738.410 1553.500 1738.730 1553.560 ;
        RECT 1897.110 1553.700 1897.430 1553.760 ;
        RECT 1931.610 1553.700 1931.930 1553.760 ;
        RECT 1897.110 1553.560 1931.930 1553.700 ;
        RECT 1897.110 1553.500 1897.430 1553.560 ;
        RECT 1931.610 1553.500 1931.930 1553.560 ;
        RECT 1993.710 1553.700 1994.030 1553.760 ;
        RECT 2028.210 1553.700 2028.530 1553.760 ;
        RECT 1993.710 1553.560 2028.530 1553.700 ;
        RECT 1993.710 1553.500 1994.030 1553.560 ;
        RECT 2028.210 1553.500 2028.530 1553.560 ;
        RECT 2090.310 1553.700 2090.630 1553.760 ;
        RECT 2124.810 1553.700 2125.130 1553.760 ;
        RECT 2090.310 1553.560 2125.130 1553.700 ;
        RECT 2090.310 1553.500 2090.630 1553.560 ;
        RECT 2124.810 1553.500 2125.130 1553.560 ;
        RECT 2186.910 1553.700 2187.230 1553.760 ;
        RECT 2221.410 1553.700 2221.730 1553.760 ;
        RECT 2186.910 1553.560 2221.730 1553.700 ;
        RECT 2186.910 1553.500 2187.230 1553.560 ;
        RECT 2221.410 1553.500 2221.730 1553.560 ;
        RECT 2283.510 1553.700 2283.830 1553.760 ;
        RECT 2318.010 1553.700 2318.330 1553.760 ;
        RECT 2283.510 1553.560 2318.330 1553.700 ;
        RECT 2283.510 1553.500 2283.830 1553.560 ;
        RECT 2318.010 1553.500 2318.330 1553.560 ;
        RECT 2476.710 1553.700 2477.030 1553.760 ;
        RECT 2511.210 1553.700 2511.530 1553.760 ;
        RECT 2476.710 1553.560 2511.530 1553.700 ;
        RECT 2476.710 1553.500 2477.030 1553.560 ;
        RECT 2511.210 1553.500 2511.530 1553.560 ;
        RECT 2573.310 1553.700 2573.630 1553.760 ;
        RECT 2607.810 1553.700 2608.130 1553.760 ;
        RECT 2573.310 1553.560 2608.130 1553.700 ;
        RECT 2573.310 1553.500 2573.630 1553.560 ;
        RECT 2607.810 1553.500 2608.130 1553.560 ;
        RECT 2669.910 1553.700 2670.230 1553.760 ;
        RECT 2704.410 1553.700 2704.730 1553.760 ;
        RECT 2669.910 1553.560 2704.730 1553.700 ;
        RECT 2669.910 1553.500 2670.230 1553.560 ;
        RECT 2704.410 1553.500 2704.730 1553.560 ;
      LAYER via ;
        RECT 1497.860 1553.840 1498.120 1554.100 ;
        RECT 1521.780 1553.840 1522.040 1554.100 ;
        RECT 1603.660 1553.840 1603.920 1554.100 ;
        RECT 1641.840 1553.840 1642.100 1554.100 ;
        RECT 1798.240 1553.840 1798.500 1554.100 ;
        RECT 1835.040 1553.840 1835.300 1554.100 ;
        RECT 2377.840 1553.840 2378.100 1554.100 ;
        RECT 2414.640 1553.840 2414.900 1554.100 ;
        RECT 2705.360 1553.840 2705.620 1554.100 ;
        RECT 2719.160 1553.840 2719.420 1554.100 ;
        RECT 1441.740 1553.500 1442.000 1553.760 ;
        RECT 1483.140 1553.500 1483.400 1553.760 ;
        RECT 1703.940 1553.500 1704.200 1553.760 ;
        RECT 1738.440 1553.500 1738.700 1553.760 ;
        RECT 1897.140 1553.500 1897.400 1553.760 ;
        RECT 1931.640 1553.500 1931.900 1553.760 ;
        RECT 1993.740 1553.500 1994.000 1553.760 ;
        RECT 2028.240 1553.500 2028.500 1553.760 ;
        RECT 2090.340 1553.500 2090.600 1553.760 ;
        RECT 2124.840 1553.500 2125.100 1553.760 ;
        RECT 2186.940 1553.500 2187.200 1553.760 ;
        RECT 2221.440 1553.500 2221.700 1553.760 ;
        RECT 2283.540 1553.500 2283.800 1553.760 ;
        RECT 2318.040 1553.500 2318.300 1553.760 ;
        RECT 2476.740 1553.500 2477.000 1553.760 ;
        RECT 2511.240 1553.500 2511.500 1553.760 ;
        RECT 2573.340 1553.500 2573.600 1553.760 ;
        RECT 2607.840 1553.500 2608.100 1553.760 ;
        RECT 2669.940 1553.500 2670.200 1553.760 ;
        RECT 2704.440 1553.500 2704.700 1553.760 ;
      LAYER met2 ;
        RECT 1203.360 1996.890 1203.640 2000.000 ;
        RECT 1204.830 1996.890 1205.110 1997.005 ;
        RECT 1203.360 1996.750 1205.110 1996.890 ;
        RECT 1203.360 1996.000 1203.640 1996.750 ;
        RECT 1204.830 1996.635 1205.110 1996.750 ;
        RECT 1338.230 1554.635 1338.510 1555.005 ;
        RECT 1338.300 1552.965 1338.440 1554.635 ;
        RECT 1483.130 1553.955 1483.410 1554.325 ;
        RECT 1497.850 1553.955 1498.130 1554.325 ;
        RECT 1521.770 1553.955 1522.050 1554.325 ;
        RECT 1483.200 1553.790 1483.340 1553.955 ;
        RECT 1497.860 1553.810 1498.120 1553.955 ;
        RECT 1521.780 1553.810 1522.040 1553.955 ;
        RECT 1603.660 1553.810 1603.920 1554.130 ;
        RECT 1641.830 1553.955 1642.110 1554.325 ;
        RECT 1738.430 1553.955 1738.710 1554.325 ;
        RECT 1641.840 1553.810 1642.100 1553.955 ;
        RECT 1441.740 1553.645 1442.000 1553.790 ;
        RECT 1441.730 1553.275 1442.010 1553.645 ;
        RECT 1483.140 1553.470 1483.400 1553.790 ;
        RECT 1603.720 1553.645 1603.860 1553.810 ;
        RECT 1738.500 1553.790 1738.640 1553.955 ;
        RECT 1798.240 1553.810 1798.500 1554.130 ;
        RECT 1835.030 1553.955 1835.310 1554.325 ;
        RECT 1931.630 1553.955 1931.910 1554.325 ;
        RECT 2028.230 1553.955 2028.510 1554.325 ;
        RECT 2124.830 1553.955 2125.110 1554.325 ;
        RECT 2221.430 1553.955 2221.710 1554.325 ;
        RECT 2318.030 1553.955 2318.310 1554.325 ;
        RECT 1835.040 1553.810 1835.300 1553.955 ;
        RECT 1703.940 1553.645 1704.200 1553.790 ;
        RECT 1603.650 1553.275 1603.930 1553.645 ;
        RECT 1703.930 1553.275 1704.210 1553.645 ;
        RECT 1738.440 1553.470 1738.700 1553.790 ;
        RECT 1798.300 1553.645 1798.440 1553.810 ;
        RECT 1931.700 1553.790 1931.840 1553.955 ;
        RECT 2028.300 1553.790 2028.440 1553.955 ;
        RECT 2124.900 1553.790 2125.040 1553.955 ;
        RECT 2221.500 1553.790 2221.640 1553.955 ;
        RECT 2318.100 1553.790 2318.240 1553.955 ;
        RECT 2377.840 1553.810 2378.100 1554.130 ;
        RECT 2414.630 1553.955 2414.910 1554.325 ;
        RECT 2511.230 1553.955 2511.510 1554.325 ;
        RECT 2607.830 1553.955 2608.110 1554.325 ;
        RECT 2704.430 1553.955 2704.710 1554.325 ;
        RECT 2705.350 1553.955 2705.630 1554.325 ;
        RECT 2414.640 1553.810 2414.900 1553.955 ;
        RECT 1897.140 1553.645 1897.400 1553.790 ;
        RECT 1798.230 1553.275 1798.510 1553.645 ;
        RECT 1897.130 1553.275 1897.410 1553.645 ;
        RECT 1931.640 1553.470 1931.900 1553.790 ;
        RECT 1993.740 1553.645 1994.000 1553.790 ;
        RECT 1993.730 1553.275 1994.010 1553.645 ;
        RECT 2028.240 1553.470 2028.500 1553.790 ;
        RECT 2090.340 1553.645 2090.600 1553.790 ;
        RECT 2090.330 1553.275 2090.610 1553.645 ;
        RECT 2124.840 1553.470 2125.100 1553.790 ;
        RECT 2186.940 1553.645 2187.200 1553.790 ;
        RECT 2186.930 1553.275 2187.210 1553.645 ;
        RECT 2221.440 1553.470 2221.700 1553.790 ;
        RECT 2283.540 1553.645 2283.800 1553.790 ;
        RECT 2283.530 1553.275 2283.810 1553.645 ;
        RECT 2318.040 1553.470 2318.300 1553.790 ;
        RECT 2377.900 1553.645 2378.040 1553.810 ;
        RECT 2511.300 1553.790 2511.440 1553.955 ;
        RECT 2607.900 1553.790 2608.040 1553.955 ;
        RECT 2704.500 1553.790 2704.640 1553.955 ;
        RECT 2705.360 1553.810 2705.620 1553.955 ;
        RECT 2719.160 1553.810 2719.420 1554.130 ;
        RECT 2476.740 1553.645 2477.000 1553.790 ;
        RECT 2377.830 1553.275 2378.110 1553.645 ;
        RECT 2476.730 1553.275 2477.010 1553.645 ;
        RECT 2511.240 1553.470 2511.500 1553.790 ;
        RECT 2573.340 1553.645 2573.600 1553.790 ;
        RECT 2573.330 1553.275 2573.610 1553.645 ;
        RECT 2607.840 1553.470 2608.100 1553.790 ;
        RECT 2669.940 1553.645 2670.200 1553.790 ;
        RECT 2669.930 1553.275 2670.210 1553.645 ;
        RECT 2704.440 1553.470 2704.700 1553.790 ;
        RECT 2719.220 1552.965 2719.360 1553.810 ;
        RECT 1338.230 1552.595 1338.510 1552.965 ;
        RECT 2719.150 1552.595 2719.430 1552.965 ;
        RECT 2777.110 1552.595 2777.390 1552.965 ;
        RECT 2777.180 1551.605 2777.320 1552.595 ;
        RECT 2777.110 1551.235 2777.390 1551.605 ;
      LAYER via2 ;
        RECT 1204.830 1996.680 1205.110 1996.960 ;
        RECT 1338.230 1554.680 1338.510 1554.960 ;
        RECT 1483.130 1554.000 1483.410 1554.280 ;
        RECT 1497.850 1554.000 1498.130 1554.280 ;
        RECT 1521.770 1554.000 1522.050 1554.280 ;
        RECT 1641.830 1554.000 1642.110 1554.280 ;
        RECT 1738.430 1554.000 1738.710 1554.280 ;
        RECT 1441.730 1553.320 1442.010 1553.600 ;
        RECT 1835.030 1554.000 1835.310 1554.280 ;
        RECT 1931.630 1554.000 1931.910 1554.280 ;
        RECT 2028.230 1554.000 2028.510 1554.280 ;
        RECT 2124.830 1554.000 2125.110 1554.280 ;
        RECT 2221.430 1554.000 2221.710 1554.280 ;
        RECT 2318.030 1554.000 2318.310 1554.280 ;
        RECT 1603.650 1553.320 1603.930 1553.600 ;
        RECT 1703.930 1553.320 1704.210 1553.600 ;
        RECT 2414.630 1554.000 2414.910 1554.280 ;
        RECT 2511.230 1554.000 2511.510 1554.280 ;
        RECT 2607.830 1554.000 2608.110 1554.280 ;
        RECT 2704.430 1554.000 2704.710 1554.280 ;
        RECT 2705.350 1554.000 2705.630 1554.280 ;
        RECT 1798.230 1553.320 1798.510 1553.600 ;
        RECT 1897.130 1553.320 1897.410 1553.600 ;
        RECT 1993.730 1553.320 1994.010 1553.600 ;
        RECT 2090.330 1553.320 2090.610 1553.600 ;
        RECT 2186.930 1553.320 2187.210 1553.600 ;
        RECT 2283.530 1553.320 2283.810 1553.600 ;
        RECT 2377.830 1553.320 2378.110 1553.600 ;
        RECT 2476.730 1553.320 2477.010 1553.600 ;
        RECT 2573.330 1553.320 2573.610 1553.600 ;
        RECT 2669.930 1553.320 2670.210 1553.600 ;
        RECT 1338.230 1552.640 1338.510 1552.920 ;
        RECT 2719.150 1552.640 2719.430 1552.920 ;
        RECT 2777.110 1552.640 2777.390 1552.920 ;
        RECT 2777.110 1551.280 2777.390 1551.560 ;
      LAYER met3 ;
        RECT 1204.805 1996.970 1205.135 1996.985 ;
        RECT 1206.390 1996.970 1206.770 1996.980 ;
        RECT 1204.805 1996.670 1206.770 1996.970 ;
        RECT 1204.805 1996.655 1205.135 1996.670 ;
        RECT 1206.390 1996.660 1206.770 1996.670 ;
        RECT 1206.390 1554.970 1206.770 1554.980 ;
        RECT 1289.190 1554.970 1289.570 1554.980 ;
        RECT 1206.390 1554.670 1289.570 1554.970 ;
        RECT 1206.390 1554.660 1206.770 1554.670 ;
        RECT 1289.190 1554.660 1289.570 1554.670 ;
        RECT 1290.110 1554.970 1290.490 1554.980 ;
        RECT 1338.205 1554.970 1338.535 1554.985 ;
        RECT 1290.110 1554.670 1338.535 1554.970 ;
        RECT 1290.110 1554.660 1290.490 1554.670 ;
        RECT 1338.205 1554.655 1338.535 1554.670 ;
        RECT 1483.105 1554.290 1483.435 1554.305 ;
        RECT 1497.825 1554.290 1498.155 1554.305 ;
        RECT 1483.105 1553.990 1498.155 1554.290 ;
        RECT 1483.105 1553.975 1483.435 1553.990 ;
        RECT 1497.825 1553.975 1498.155 1553.990 ;
        RECT 1521.745 1554.290 1522.075 1554.305 ;
        RECT 1641.805 1554.290 1642.135 1554.305 ;
        RECT 1738.405 1554.290 1738.735 1554.305 ;
        RECT 1835.005 1554.290 1835.335 1554.305 ;
        RECT 1931.605 1554.290 1931.935 1554.305 ;
        RECT 2028.205 1554.290 2028.535 1554.305 ;
        RECT 2124.805 1554.290 2125.135 1554.305 ;
        RECT 2221.405 1554.290 2221.735 1554.305 ;
        RECT 2318.005 1554.290 2318.335 1554.305 ;
        RECT 2414.605 1554.290 2414.935 1554.305 ;
        RECT 2511.205 1554.290 2511.535 1554.305 ;
        RECT 2607.805 1554.290 2608.135 1554.305 ;
        RECT 2704.405 1554.290 2704.735 1554.305 ;
        RECT 2705.325 1554.290 2705.655 1554.305 ;
        RECT 1521.745 1553.990 1560.010 1554.290 ;
        RECT 1521.745 1553.975 1522.075 1553.990 ;
        RECT 1289.190 1553.610 1289.570 1553.620 ;
        RECT 1290.110 1553.610 1290.490 1553.620 ;
        RECT 1441.705 1553.610 1442.035 1553.625 ;
        RECT 1289.190 1553.310 1290.490 1553.610 ;
        RECT 1289.190 1553.300 1289.570 1553.310 ;
        RECT 1290.110 1553.300 1290.490 1553.310 ;
        RECT 1394.110 1553.310 1442.035 1553.610 ;
        RECT 1559.710 1553.610 1560.010 1553.990 ;
        RECT 1641.805 1553.990 1656.610 1554.290 ;
        RECT 1641.805 1553.975 1642.135 1553.990 ;
        RECT 1603.625 1553.610 1603.955 1553.625 ;
        RECT 1559.710 1553.310 1603.955 1553.610 ;
        RECT 1656.310 1553.610 1656.610 1553.990 ;
        RECT 1738.405 1553.990 1753.210 1554.290 ;
        RECT 1738.405 1553.975 1738.735 1553.990 ;
        RECT 1703.905 1553.610 1704.235 1553.625 ;
        RECT 1656.310 1553.310 1704.235 1553.610 ;
        RECT 1752.910 1553.610 1753.210 1553.990 ;
        RECT 1835.005 1553.990 1849.810 1554.290 ;
        RECT 1835.005 1553.975 1835.335 1553.990 ;
        RECT 1798.205 1553.610 1798.535 1553.625 ;
        RECT 1752.910 1553.310 1798.535 1553.610 ;
        RECT 1849.510 1553.610 1849.810 1553.990 ;
        RECT 1931.605 1553.990 1946.410 1554.290 ;
        RECT 1931.605 1553.975 1931.935 1553.990 ;
        RECT 1897.105 1553.610 1897.435 1553.625 ;
        RECT 1849.510 1553.310 1897.435 1553.610 ;
        RECT 1946.110 1553.610 1946.410 1553.990 ;
        RECT 2028.205 1553.990 2043.010 1554.290 ;
        RECT 2028.205 1553.975 2028.535 1553.990 ;
        RECT 1993.705 1553.610 1994.035 1553.625 ;
        RECT 1946.110 1553.310 1994.035 1553.610 ;
        RECT 2042.710 1553.610 2043.010 1553.990 ;
        RECT 2124.805 1553.990 2139.610 1554.290 ;
        RECT 2124.805 1553.975 2125.135 1553.990 ;
        RECT 2090.305 1553.610 2090.635 1553.625 ;
        RECT 2042.710 1553.310 2090.635 1553.610 ;
        RECT 2139.310 1553.610 2139.610 1553.990 ;
        RECT 2221.405 1553.990 2236.210 1554.290 ;
        RECT 2221.405 1553.975 2221.735 1553.990 ;
        RECT 2186.905 1553.610 2187.235 1553.625 ;
        RECT 2139.310 1553.310 2187.235 1553.610 ;
        RECT 2235.910 1553.610 2236.210 1553.990 ;
        RECT 2318.005 1553.990 2332.810 1554.290 ;
        RECT 2318.005 1553.975 2318.335 1553.990 ;
        RECT 2283.505 1553.610 2283.835 1553.625 ;
        RECT 2235.910 1553.310 2283.835 1553.610 ;
        RECT 2332.510 1553.610 2332.810 1553.990 ;
        RECT 2414.605 1553.990 2429.410 1554.290 ;
        RECT 2414.605 1553.975 2414.935 1553.990 ;
        RECT 2377.805 1553.610 2378.135 1553.625 ;
        RECT 2332.510 1553.310 2378.135 1553.610 ;
        RECT 2429.110 1553.610 2429.410 1553.990 ;
        RECT 2511.205 1553.990 2526.010 1554.290 ;
        RECT 2511.205 1553.975 2511.535 1553.990 ;
        RECT 2476.705 1553.610 2477.035 1553.625 ;
        RECT 2429.110 1553.310 2477.035 1553.610 ;
        RECT 2525.710 1553.610 2526.010 1553.990 ;
        RECT 2607.805 1553.990 2622.610 1554.290 ;
        RECT 2607.805 1553.975 2608.135 1553.990 ;
        RECT 2573.305 1553.610 2573.635 1553.625 ;
        RECT 2525.710 1553.310 2573.635 1553.610 ;
        RECT 2622.310 1553.610 2622.610 1553.990 ;
        RECT 2704.405 1553.990 2705.655 1554.290 ;
        RECT 2704.405 1553.975 2704.735 1553.990 ;
        RECT 2705.325 1553.975 2705.655 1553.990 ;
        RECT 2801.670 1553.980 2802.050 1554.300 ;
        RECT 2917.600 1554.290 2924.800 1554.740 ;
        RECT 2916.710 1553.990 2924.800 1554.290 ;
        RECT 2669.905 1553.610 2670.235 1553.625 ;
        RECT 2801.710 1553.610 2802.010 1553.980 ;
        RECT 2622.310 1553.310 2670.235 1553.610 ;
        RECT 1338.205 1552.930 1338.535 1552.945 ;
        RECT 1394.110 1552.930 1394.410 1553.310 ;
        RECT 1441.705 1553.295 1442.035 1553.310 ;
        RECT 1603.625 1553.295 1603.955 1553.310 ;
        RECT 1703.905 1553.295 1704.235 1553.310 ;
        RECT 1798.205 1553.295 1798.535 1553.310 ;
        RECT 1897.105 1553.295 1897.435 1553.310 ;
        RECT 1993.705 1553.295 1994.035 1553.310 ;
        RECT 2090.305 1553.295 2090.635 1553.310 ;
        RECT 2186.905 1553.295 2187.235 1553.310 ;
        RECT 2283.505 1553.295 2283.835 1553.310 ;
        RECT 2377.805 1553.295 2378.135 1553.310 ;
        RECT 2476.705 1553.295 2477.035 1553.310 ;
        RECT 2573.305 1553.295 2573.635 1553.310 ;
        RECT 2669.905 1553.295 2670.235 1553.310 ;
        RECT 2800.790 1553.310 2802.010 1553.610 ;
        RECT 2802.590 1553.610 2802.970 1553.620 ;
        RECT 2916.710 1553.610 2917.010 1553.990 ;
        RECT 2802.590 1553.310 2883.890 1553.610 ;
        RECT 1338.205 1552.630 1394.410 1552.930 ;
        RECT 2719.125 1552.930 2719.455 1552.945 ;
        RECT 2752.910 1552.930 2753.290 1552.940 ;
        RECT 2719.125 1552.630 2753.290 1552.930 ;
        RECT 1338.205 1552.615 1338.535 1552.630 ;
        RECT 2719.125 1552.615 2719.455 1552.630 ;
        RECT 2752.910 1552.620 2753.290 1552.630 ;
        RECT 2777.085 1552.930 2777.415 1552.945 ;
        RECT 2800.790 1552.930 2801.090 1553.310 ;
        RECT 2802.590 1553.300 2802.970 1553.310 ;
        RECT 2777.085 1552.630 2801.090 1552.930 ;
        RECT 2883.590 1552.930 2883.890 1553.310 ;
        RECT 2884.510 1553.310 2917.010 1553.610 ;
        RECT 2917.600 1553.540 2924.800 1553.990 ;
        RECT 2884.510 1552.930 2884.810 1553.310 ;
        RECT 2883.590 1552.630 2884.810 1552.930 ;
        RECT 2777.085 1552.615 2777.415 1552.630 ;
        RECT 2752.910 1551.570 2753.290 1551.580 ;
        RECT 2777.085 1551.570 2777.415 1551.585 ;
        RECT 2752.910 1551.270 2777.415 1551.570 ;
        RECT 2752.910 1551.260 2753.290 1551.270 ;
        RECT 2777.085 1551.255 2777.415 1551.270 ;
      LAYER via3 ;
        RECT 1206.420 1996.660 1206.740 1996.980 ;
        RECT 1206.420 1554.660 1206.740 1554.980 ;
        RECT 1289.220 1554.660 1289.540 1554.980 ;
        RECT 1290.140 1554.660 1290.460 1554.980 ;
        RECT 1289.220 1553.300 1289.540 1553.620 ;
        RECT 1290.140 1553.300 1290.460 1553.620 ;
        RECT 2801.700 1553.980 2802.020 1554.300 ;
        RECT 2752.940 1552.620 2753.260 1552.940 ;
        RECT 2802.620 1553.300 2802.940 1553.620 ;
        RECT 2752.940 1551.260 2753.260 1551.580 ;
      LAYER met4 ;
        RECT 1206.415 1996.655 1206.745 1996.985 ;
        RECT 1206.430 1554.985 1206.730 1996.655 ;
        RECT 2801.710 1555.350 2802.930 1555.650 ;
        RECT 1206.415 1554.655 1206.745 1554.985 ;
        RECT 1289.215 1554.655 1289.545 1554.985 ;
        RECT 1290.135 1554.655 1290.465 1554.985 ;
        RECT 1289.230 1553.625 1289.530 1554.655 ;
        RECT 1290.150 1553.625 1290.450 1554.655 ;
        RECT 2801.710 1554.305 2802.010 1555.350 ;
        RECT 2801.695 1553.975 2802.025 1554.305 ;
        RECT 2802.630 1553.625 2802.930 1555.350 ;
        RECT 1289.215 1553.295 1289.545 1553.625 ;
        RECT 1290.135 1553.295 1290.465 1553.625 ;
        RECT 2802.615 1553.295 2802.945 1553.625 ;
        RECT 2752.935 1552.615 2753.265 1552.945 ;
        RECT 2752.950 1551.585 2753.250 1552.615 ;
        RECT 2752.935 1551.255 2753.265 1551.585 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1224.205 2007.785 1224.375 2009.995 ;
        RECT 1241.685 2007.785 1241.855 2009.315 ;
      LAYER mcon ;
        RECT 1224.205 2009.825 1224.375 2009.995 ;
        RECT 1241.685 2009.145 1241.855 2009.315 ;
      LAYER met1 ;
        RECT 1211.250 2009.980 1211.570 2010.040 ;
        RECT 1224.145 2009.980 1224.435 2010.025 ;
        RECT 1211.250 2009.840 1224.435 2009.980 ;
        RECT 1211.250 2009.780 1211.570 2009.840 ;
        RECT 1224.145 2009.795 1224.435 2009.840 ;
        RECT 1241.625 2009.300 1241.915 2009.345 ;
        RECT 2445.890 2009.300 2446.210 2009.360 ;
        RECT 1241.625 2009.160 2446.210 2009.300 ;
        RECT 1241.625 2009.115 1241.915 2009.160 ;
        RECT 2445.890 2009.100 2446.210 2009.160 ;
        RECT 1224.145 2007.940 1224.435 2007.985 ;
        RECT 1241.625 2007.940 1241.915 2007.985 ;
        RECT 1224.145 2007.800 1241.915 2007.940 ;
        RECT 1224.145 2007.755 1224.435 2007.800 ;
        RECT 1241.625 2007.755 1241.915 2007.800 ;
        RECT 2445.890 1793.740 2446.210 1793.800 ;
        RECT 2900.370 1793.740 2900.690 1793.800 ;
        RECT 2445.890 1793.600 2900.690 1793.740 ;
        RECT 2445.890 1793.540 2446.210 1793.600 ;
        RECT 2900.370 1793.540 2900.690 1793.600 ;
      LAYER via ;
        RECT 1211.280 2009.780 1211.540 2010.040 ;
        RECT 2445.920 2009.100 2446.180 2009.360 ;
        RECT 2445.920 1793.540 2446.180 1793.800 ;
        RECT 2900.400 1793.540 2900.660 1793.800 ;
      LAYER met2 ;
        RECT 1211.280 2009.750 1211.540 2010.070 ;
        RECT 1211.340 2000.000 1211.480 2009.750 ;
        RECT 2445.920 2009.070 2446.180 2009.390 ;
        RECT 1211.180 1999.540 1211.480 2000.000 ;
        RECT 1211.180 1996.000 1211.460 1999.540 ;
        RECT 2445.980 1793.830 2446.120 2009.070 ;
        RECT 2445.920 1793.510 2446.180 1793.830 ;
        RECT 2900.400 1793.510 2900.660 1793.830 ;
        RECT 2900.460 1789.605 2900.600 1793.510 ;
        RECT 2900.390 1789.235 2900.670 1789.605 ;
      LAYER via2 ;
        RECT 2900.390 1789.280 2900.670 1789.560 ;
      LAYER met3 ;
        RECT 2900.365 1789.570 2900.695 1789.585 ;
        RECT 2917.600 1789.570 2924.800 1790.020 ;
        RECT 2900.365 1789.270 2924.800 1789.570 ;
        RECT 2900.365 1789.255 2900.695 1789.270 ;
        RECT 2917.600 1788.820 2924.800 1789.270 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1219.070 2021.880 1219.390 2021.940 ;
        RECT 2900.830 2021.880 2901.150 2021.940 ;
        RECT 1219.070 2021.740 2901.150 2021.880 ;
        RECT 1219.070 2021.680 1219.390 2021.740 ;
        RECT 2900.830 2021.680 2901.150 2021.740 ;
      LAYER via ;
        RECT 1219.100 2021.680 1219.360 2021.940 ;
        RECT 2900.860 2021.680 2901.120 2021.940 ;
      LAYER met2 ;
        RECT 2900.850 2023.835 2901.130 2024.205 ;
        RECT 2900.920 2021.970 2901.060 2023.835 ;
        RECT 1219.100 2021.650 1219.360 2021.970 ;
        RECT 2900.860 2021.650 2901.120 2021.970 ;
        RECT 1219.160 2000.000 1219.300 2021.650 ;
        RECT 1219.000 1999.540 1219.300 2000.000 ;
        RECT 1219.000 1996.000 1219.280 1999.540 ;
      LAYER via2 ;
        RECT 2900.850 2023.880 2901.130 2024.160 ;
      LAYER met3 ;
        RECT 2900.825 2024.170 2901.155 2024.185 ;
        RECT 2917.600 2024.170 2924.800 2024.620 ;
        RECT 2900.825 2023.870 2924.800 2024.170 ;
        RECT 2900.825 2023.855 2901.155 2023.870 ;
        RECT 2917.600 2023.420 2924.800 2023.870 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1497.000 2256.680 1499.440 2256.820 ;
        RECT 1227.350 2256.480 1227.670 2256.540 ;
        RECT 1497.000 2256.480 1497.140 2256.680 ;
        RECT 1227.350 2256.340 1497.140 2256.480 ;
        RECT 1499.300 2256.480 1499.440 2256.680 ;
        RECT 2900.830 2256.480 2901.150 2256.540 ;
        RECT 1499.300 2256.340 2901.150 2256.480 ;
        RECT 1227.350 2256.280 1227.670 2256.340 ;
        RECT 2900.830 2256.280 2901.150 2256.340 ;
      LAYER via ;
        RECT 1227.380 2256.280 1227.640 2256.540 ;
        RECT 2900.860 2256.280 2901.120 2256.540 ;
      LAYER met2 ;
        RECT 2900.850 2258.435 2901.130 2258.805 ;
        RECT 2900.920 2256.570 2901.060 2258.435 ;
        RECT 1227.380 2256.250 1227.640 2256.570 ;
        RECT 2900.860 2256.250 2901.120 2256.570 ;
        RECT 1226.820 1999.610 1227.100 2000.000 ;
        RECT 1227.440 1999.610 1227.580 2256.250 ;
        RECT 1226.820 1999.470 1227.580 1999.610 ;
        RECT 1226.820 1996.000 1227.100 1999.470 ;
      LAYER via2 ;
        RECT 2900.850 2258.480 2901.130 2258.760 ;
      LAYER met3 ;
        RECT 2900.825 2258.770 2901.155 2258.785 ;
        RECT 2917.600 2258.770 2924.800 2259.220 ;
        RECT 2900.825 2258.470 2924.800 2258.770 ;
        RECT 2900.825 2258.455 2901.155 2258.470 ;
        RECT 2917.600 2258.020 2924.800 2258.470 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1205.730 1687.660 1206.050 1687.720 ;
        RECT 1214.930 1687.660 1215.250 1687.720 ;
        RECT 1205.730 1687.520 1215.250 1687.660 ;
        RECT 1205.730 1687.460 1206.050 1687.520 ;
        RECT 1214.930 1687.460 1215.250 1687.520 ;
        RECT 634.410 1673.720 634.730 1673.780 ;
        RECT 1205.730 1673.720 1206.050 1673.780 ;
        RECT 634.410 1673.580 1206.050 1673.720 ;
        RECT 634.410 1673.520 634.730 1673.580 ;
        RECT 1205.730 1673.520 1206.050 1673.580 ;
      LAYER via ;
        RECT 1205.760 1687.460 1206.020 1687.720 ;
        RECT 1214.960 1687.460 1215.220 1687.720 ;
        RECT 634.440 1673.520 634.700 1673.780 ;
        RECT 1205.760 1673.520 1206.020 1673.780 ;
      LAYER met2 ;
        RECT 1214.860 1700.340 1215.140 1704.000 ;
        RECT 1214.860 1700.000 1215.160 1700.340 ;
        RECT 1215.020 1687.750 1215.160 1700.000 ;
        RECT 1205.760 1687.430 1206.020 1687.750 ;
        RECT 1214.960 1687.430 1215.220 1687.750 ;
        RECT 1205.820 1673.810 1205.960 1687.430 ;
        RECT 634.440 1673.490 634.700 1673.810 ;
        RECT 1205.760 1673.490 1206.020 1673.810 ;
        RECT 634.500 17.410 634.640 1673.490 ;
        RECT 633.120 17.270 634.640 17.410 ;
        RECT 633.120 2.400 633.260 17.270 ;
        RECT 632.910 -4.800 633.470 2.400 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1398.470 1690.380 1398.790 1690.440 ;
        RECT 1449.990 1690.380 1450.310 1690.440 ;
        RECT 1398.470 1690.240 1450.310 1690.380 ;
        RECT 1398.470 1690.180 1398.790 1690.240 ;
        RECT 1449.990 1690.180 1450.310 1690.240 ;
        RECT 1449.990 1680.860 1450.310 1680.920 ;
        RECT 2415.070 1680.860 2415.390 1680.920 ;
        RECT 1449.990 1680.720 2415.390 1680.860 ;
        RECT 1449.990 1680.660 1450.310 1680.720 ;
        RECT 2415.070 1680.660 2415.390 1680.720 ;
      LAYER via ;
        RECT 1398.500 1690.180 1398.760 1690.440 ;
        RECT 1450.020 1690.180 1450.280 1690.440 ;
        RECT 1450.020 1680.660 1450.280 1680.920 ;
        RECT 2415.100 1680.660 2415.360 1680.920 ;
      LAYER met2 ;
        RECT 1398.400 1700.340 1398.680 1704.000 ;
        RECT 1398.400 1700.000 1398.700 1700.340 ;
        RECT 1398.560 1690.470 1398.700 1700.000 ;
        RECT 1398.500 1690.150 1398.760 1690.470 ;
        RECT 1450.020 1690.150 1450.280 1690.470 ;
        RECT 1450.080 1680.950 1450.220 1690.150 ;
        RECT 1450.020 1680.630 1450.280 1680.950 ;
        RECT 2415.100 1680.630 2415.360 1680.950 ;
        RECT 2415.160 17.410 2415.300 1680.630 ;
        RECT 2415.160 17.270 2417.600 17.410 ;
        RECT 2417.460 2.400 2417.600 17.270 ;
        RECT 2417.250 -4.800 2417.810 2.400 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1407.285 1684.445 1407.455 1686.315 ;
        RECT 1420.165 1684.445 1420.335 1687.675 ;
      LAYER mcon ;
        RECT 1420.165 1687.505 1420.335 1687.675 ;
        RECT 1407.285 1686.145 1407.455 1686.315 ;
      LAYER met1 ;
        RECT 1583.390 1688.000 1583.710 1688.060 ;
        RECT 1438.120 1687.860 1583.710 1688.000 ;
        RECT 1420.105 1687.660 1420.395 1687.705 ;
        RECT 1438.120 1687.660 1438.260 1687.860 ;
        RECT 1583.390 1687.800 1583.710 1687.860 ;
        RECT 1420.105 1687.520 1438.260 1687.660 ;
        RECT 1420.105 1687.475 1420.395 1687.520 ;
        RECT 1400.310 1686.300 1400.630 1686.360 ;
        RECT 1407.225 1686.300 1407.515 1686.345 ;
        RECT 1400.310 1686.160 1407.515 1686.300 ;
        RECT 1400.310 1686.100 1400.630 1686.160 ;
        RECT 1407.225 1686.115 1407.515 1686.160 ;
        RECT 1407.225 1684.600 1407.515 1684.645 ;
        RECT 1420.105 1684.600 1420.395 1684.645 ;
        RECT 1407.225 1684.460 1420.395 1684.600 ;
        RECT 1407.225 1684.415 1407.515 1684.460 ;
        RECT 1420.105 1684.415 1420.395 1684.460 ;
        RECT 1583.390 24.040 1583.710 24.100 ;
        RECT 2434.850 24.040 2435.170 24.100 ;
        RECT 1583.390 23.900 2435.170 24.040 ;
        RECT 1583.390 23.840 1583.710 23.900 ;
        RECT 2434.850 23.840 2435.170 23.900 ;
      LAYER via ;
        RECT 1583.420 1687.800 1583.680 1688.060 ;
        RECT 1400.340 1686.100 1400.600 1686.360 ;
        RECT 1583.420 23.840 1583.680 24.100 ;
        RECT 2434.880 23.840 2435.140 24.100 ;
      LAYER met2 ;
        RECT 1400.240 1700.340 1400.520 1704.000 ;
        RECT 1400.240 1700.000 1400.540 1700.340 ;
        RECT 1400.400 1686.390 1400.540 1700.000 ;
        RECT 1583.420 1687.770 1583.680 1688.090 ;
        RECT 1400.340 1686.070 1400.600 1686.390 ;
        RECT 1583.480 24.130 1583.620 1687.770 ;
        RECT 1583.420 23.810 1583.680 24.130 ;
        RECT 2434.880 23.810 2435.140 24.130 ;
        RECT 2434.940 2.400 2435.080 23.810 ;
        RECT 2434.730 -4.800 2435.290 2.400 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1413.725 1683.765 1413.895 1685.295 ;
        RECT 1439.025 1685.125 1439.195 1687.675 ;
      LAYER mcon ;
        RECT 1439.025 1687.505 1439.195 1687.675 ;
        RECT 1413.725 1685.125 1413.895 1685.295 ;
      LAYER met1 ;
        RECT 1438.965 1687.660 1439.255 1687.705 ;
        RECT 1597.190 1687.660 1597.510 1687.720 ;
        RECT 1438.965 1687.520 1597.510 1687.660 ;
        RECT 1438.965 1687.475 1439.255 1687.520 ;
        RECT 1597.190 1687.460 1597.510 1687.520 ;
        RECT 1402.150 1685.280 1402.470 1685.340 ;
        RECT 1413.665 1685.280 1413.955 1685.325 ;
        RECT 1438.965 1685.280 1439.255 1685.325 ;
        RECT 1402.150 1685.140 1413.955 1685.280 ;
        RECT 1402.150 1685.080 1402.470 1685.140 ;
        RECT 1413.665 1685.095 1413.955 1685.140 ;
        RECT 1421.100 1685.140 1439.255 1685.280 ;
        RECT 1413.665 1683.920 1413.955 1683.965 ;
        RECT 1421.100 1683.920 1421.240 1685.140 ;
        RECT 1438.965 1685.095 1439.255 1685.140 ;
        RECT 1413.665 1683.780 1421.240 1683.920 ;
        RECT 1413.665 1683.735 1413.955 1683.780 ;
        RECT 1597.190 37.980 1597.510 38.040 ;
        RECT 2452.790 37.980 2453.110 38.040 ;
        RECT 1597.190 37.840 2453.110 37.980 ;
        RECT 1597.190 37.780 1597.510 37.840 ;
        RECT 2452.790 37.780 2453.110 37.840 ;
      LAYER via ;
        RECT 1597.220 1687.460 1597.480 1687.720 ;
        RECT 1402.180 1685.080 1402.440 1685.340 ;
        RECT 1597.220 37.780 1597.480 38.040 ;
        RECT 2452.820 37.780 2453.080 38.040 ;
      LAYER met2 ;
        RECT 1402.080 1700.340 1402.360 1704.000 ;
        RECT 1402.080 1700.000 1402.380 1700.340 ;
        RECT 1402.240 1685.370 1402.380 1700.000 ;
        RECT 1597.220 1687.430 1597.480 1687.750 ;
        RECT 1402.180 1685.050 1402.440 1685.370 ;
        RECT 1597.280 38.070 1597.420 1687.430 ;
        RECT 1597.220 37.750 1597.480 38.070 ;
        RECT 2452.820 37.750 2453.080 38.070 ;
        RECT 2452.880 2.400 2453.020 37.750 ;
        RECT 2452.670 -4.800 2453.230 2.400 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1438.565 1685.465 1438.735 1688.695 ;
      LAYER mcon ;
        RECT 1438.565 1688.525 1438.735 1688.695 ;
      LAYER met1 ;
        RECT 1438.505 1688.680 1438.795 1688.725 ;
        RECT 1514.390 1688.680 1514.710 1688.740 ;
        RECT 1438.505 1688.540 1514.710 1688.680 ;
        RECT 1438.505 1688.495 1438.795 1688.540 ;
        RECT 1514.390 1688.480 1514.710 1688.540 ;
        RECT 1403.990 1685.620 1404.310 1685.680 ;
        RECT 1438.505 1685.620 1438.795 1685.665 ;
        RECT 1403.990 1685.480 1438.795 1685.620 ;
        RECT 1403.990 1685.420 1404.310 1685.480 ;
        RECT 1438.505 1685.435 1438.795 1685.480 ;
        RECT 1514.390 44.780 1514.710 44.840 ;
        RECT 2470.730 44.780 2471.050 44.840 ;
        RECT 1514.390 44.640 2471.050 44.780 ;
        RECT 1514.390 44.580 1514.710 44.640 ;
        RECT 2470.730 44.580 2471.050 44.640 ;
      LAYER via ;
        RECT 1514.420 1688.480 1514.680 1688.740 ;
        RECT 1404.020 1685.420 1404.280 1685.680 ;
        RECT 1514.420 44.580 1514.680 44.840 ;
        RECT 2470.760 44.580 2471.020 44.840 ;
      LAYER met2 ;
        RECT 1403.920 1700.340 1404.200 1704.000 ;
        RECT 1403.920 1700.000 1404.220 1700.340 ;
        RECT 1404.080 1685.710 1404.220 1700.000 ;
        RECT 1514.420 1688.450 1514.680 1688.770 ;
        RECT 1404.020 1685.390 1404.280 1685.710 ;
        RECT 1514.480 44.870 1514.620 1688.450 ;
        RECT 1514.420 44.550 1514.680 44.870 ;
        RECT 2470.760 44.550 2471.020 44.870 ;
        RECT 2470.820 2.400 2470.960 44.550 ;
        RECT 2470.610 -4.800 2471.170 2.400 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1437.645 1686.825 1437.815 1688.015 ;
      LAYER mcon ;
        RECT 1437.645 1687.845 1437.815 1688.015 ;
      LAYER met1 ;
        RECT 1405.830 1688.000 1406.150 1688.060 ;
        RECT 1437.585 1688.000 1437.875 1688.045 ;
        RECT 1405.830 1687.860 1437.875 1688.000 ;
        RECT 1405.830 1687.800 1406.150 1687.860 ;
        RECT 1437.585 1687.815 1437.875 1687.860 ;
        RECT 1437.585 1686.980 1437.875 1687.025 ;
        RECT 2445.890 1686.980 2446.210 1687.040 ;
        RECT 1437.585 1686.840 2446.210 1686.980 ;
        RECT 1437.585 1686.795 1437.875 1686.840 ;
        RECT 2445.890 1686.780 2446.210 1686.840 ;
        RECT 2445.890 24.040 2446.210 24.100 ;
        RECT 2488.670 24.040 2488.990 24.100 ;
        RECT 2445.890 23.900 2488.990 24.040 ;
        RECT 2445.890 23.840 2446.210 23.900 ;
        RECT 2488.670 23.840 2488.990 23.900 ;
      LAYER via ;
        RECT 1405.860 1687.800 1406.120 1688.060 ;
        RECT 2445.920 1686.780 2446.180 1687.040 ;
        RECT 2445.920 23.840 2446.180 24.100 ;
        RECT 2488.700 23.840 2488.960 24.100 ;
      LAYER met2 ;
        RECT 1405.760 1700.340 1406.040 1704.000 ;
        RECT 1405.760 1700.000 1406.060 1700.340 ;
        RECT 1405.920 1688.090 1406.060 1700.000 ;
        RECT 1405.860 1687.770 1406.120 1688.090 ;
        RECT 2445.920 1686.750 2446.180 1687.070 ;
        RECT 2445.980 24.130 2446.120 1686.750 ;
        RECT 2445.920 23.810 2446.180 24.130 ;
        RECT 2488.700 23.810 2488.960 24.130 ;
        RECT 2488.760 2.400 2488.900 23.810 ;
        RECT 2488.550 -4.800 2489.110 2.400 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1415.565 1684.955 1415.735 1686.655 ;
        RECT 1415.105 1684.785 1415.735 1684.955 ;
      LAYER mcon ;
        RECT 1415.565 1686.485 1415.735 1686.655 ;
      LAYER met1 ;
        RECT 1415.505 1686.640 1415.795 1686.685 ;
        RECT 1449.530 1686.640 1449.850 1686.700 ;
        RECT 1415.505 1686.500 1449.850 1686.640 ;
        RECT 1415.505 1686.455 1415.795 1686.500 ;
        RECT 1449.530 1686.440 1449.850 1686.500 ;
        RECT 1407.670 1684.940 1407.990 1685.000 ;
        RECT 1415.045 1684.940 1415.335 1684.985 ;
        RECT 1407.670 1684.800 1415.335 1684.940 ;
        RECT 1407.670 1684.740 1407.990 1684.800 ;
        RECT 1415.045 1684.755 1415.335 1684.800 ;
        RECT 1449.530 1673.720 1449.850 1673.780 ;
        RECT 2504.770 1673.720 2505.090 1673.780 ;
        RECT 1449.530 1673.580 2505.090 1673.720 ;
        RECT 1449.530 1673.520 1449.850 1673.580 ;
        RECT 2504.770 1673.520 2505.090 1673.580 ;
      LAYER via ;
        RECT 1449.560 1686.440 1449.820 1686.700 ;
        RECT 1407.700 1684.740 1407.960 1685.000 ;
        RECT 1449.560 1673.520 1449.820 1673.780 ;
        RECT 2504.800 1673.520 2505.060 1673.780 ;
      LAYER met2 ;
        RECT 1407.600 1700.340 1407.880 1704.000 ;
        RECT 1407.600 1700.000 1407.900 1700.340 ;
        RECT 1407.760 1685.030 1407.900 1700.000 ;
        RECT 1449.560 1686.410 1449.820 1686.730 ;
        RECT 1407.700 1684.710 1407.960 1685.030 ;
        RECT 1449.620 1673.810 1449.760 1686.410 ;
        RECT 1449.560 1673.490 1449.820 1673.810 ;
        RECT 2504.800 1673.490 2505.060 1673.810 ;
        RECT 2504.860 17.410 2505.000 1673.490 ;
        RECT 2504.860 17.270 2506.380 17.410 ;
        RECT 2506.240 2.400 2506.380 17.270 ;
        RECT 2506.030 -4.800 2506.590 2.400 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1437.185 1686.825 1437.355 1689.035 ;
      LAYER mcon ;
        RECT 1437.185 1688.865 1437.355 1689.035 ;
      LAYER met1 ;
        RECT 1437.125 1689.020 1437.415 1689.065 ;
        RECT 1507.490 1689.020 1507.810 1689.080 ;
        RECT 1437.125 1688.880 1507.810 1689.020 ;
        RECT 1437.125 1688.835 1437.415 1688.880 ;
        RECT 1507.490 1688.820 1507.810 1688.880 ;
        RECT 1409.510 1686.980 1409.830 1687.040 ;
        RECT 1437.125 1686.980 1437.415 1687.025 ;
        RECT 1409.510 1686.840 1437.415 1686.980 ;
        RECT 1409.510 1686.780 1409.830 1686.840 ;
        RECT 1437.125 1686.795 1437.415 1686.840 ;
        RECT 1507.490 58.720 1507.810 58.780 ;
        RECT 2518.570 58.720 2518.890 58.780 ;
        RECT 1507.490 58.580 2518.890 58.720 ;
        RECT 1507.490 58.520 1507.810 58.580 ;
        RECT 2518.570 58.520 2518.890 58.580 ;
      LAYER via ;
        RECT 1507.520 1688.820 1507.780 1689.080 ;
        RECT 1409.540 1686.780 1409.800 1687.040 ;
        RECT 1507.520 58.520 1507.780 58.780 ;
        RECT 2518.600 58.520 2518.860 58.780 ;
      LAYER met2 ;
        RECT 1409.440 1700.340 1409.720 1704.000 ;
        RECT 1409.440 1700.000 1409.740 1700.340 ;
        RECT 1409.600 1687.070 1409.740 1700.000 ;
        RECT 1507.520 1688.790 1507.780 1689.110 ;
        RECT 1409.540 1686.750 1409.800 1687.070 ;
        RECT 1507.580 58.810 1507.720 1688.790 ;
        RECT 1507.520 58.490 1507.780 58.810 ;
        RECT 2518.600 58.490 2518.860 58.810 ;
        RECT 2518.660 17.410 2518.800 58.490 ;
        RECT 2518.660 17.270 2524.320 17.410 ;
        RECT 2524.180 2.400 2524.320 17.270 ;
        RECT 2523.970 -4.800 2524.530 2.400 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1438.105 1688.865 1439.655 1689.035 ;
        RECT 1414.645 1686.485 1414.815 1688.695 ;
        RECT 1438.105 1688.525 1438.275 1688.865 ;
        RECT 1439.485 1685.465 1439.655 1688.865 ;
      LAYER mcon ;
        RECT 1414.645 1688.525 1414.815 1688.695 ;
      LAYER met1 ;
        RECT 1414.585 1688.680 1414.875 1688.725 ;
        RECT 1438.045 1688.680 1438.335 1688.725 ;
        RECT 1414.585 1688.540 1438.335 1688.680 ;
        RECT 1414.585 1688.495 1414.875 1688.540 ;
        RECT 1438.045 1688.495 1438.335 1688.540 ;
        RECT 1414.585 1686.455 1414.875 1686.685 ;
        RECT 1411.350 1686.300 1411.670 1686.360 ;
        RECT 1414.660 1686.300 1414.800 1686.455 ;
        RECT 1411.350 1686.160 1414.800 1686.300 ;
        RECT 1411.350 1686.100 1411.670 1686.160 ;
        RECT 1439.425 1685.620 1439.715 1685.665 ;
        RECT 1459.190 1685.620 1459.510 1685.680 ;
        RECT 1439.425 1685.480 1459.510 1685.620 ;
        RECT 1439.425 1685.435 1439.715 1685.480 ;
        RECT 1459.190 1685.420 1459.510 1685.480 ;
        RECT 1459.190 65.520 1459.510 65.580 ;
        RECT 2539.270 65.520 2539.590 65.580 ;
        RECT 1459.190 65.380 2539.590 65.520 ;
        RECT 1459.190 65.320 1459.510 65.380 ;
        RECT 2539.270 65.320 2539.590 65.380 ;
      LAYER via ;
        RECT 1411.380 1686.100 1411.640 1686.360 ;
        RECT 1459.220 1685.420 1459.480 1685.680 ;
        RECT 1459.220 65.320 1459.480 65.580 ;
        RECT 2539.300 65.320 2539.560 65.580 ;
      LAYER met2 ;
        RECT 1411.280 1700.340 1411.560 1704.000 ;
        RECT 1411.280 1700.000 1411.580 1700.340 ;
        RECT 1411.440 1686.390 1411.580 1700.000 ;
        RECT 1411.380 1686.070 1411.640 1686.390 ;
        RECT 1459.220 1685.390 1459.480 1685.710 ;
        RECT 1459.280 65.610 1459.420 1685.390 ;
        RECT 1459.220 65.290 1459.480 65.610 ;
        RECT 2539.300 65.290 2539.560 65.610 ;
        RECT 2539.360 17.410 2539.500 65.290 ;
        RECT 2539.360 17.270 2542.260 17.410 ;
        RECT 2542.120 2.400 2542.260 17.270 ;
        RECT 2541.910 -4.800 2542.470 2.400 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1413.190 1689.360 1413.510 1689.420 ;
        RECT 1493.690 1689.360 1494.010 1689.420 ;
        RECT 1413.190 1689.220 1494.010 1689.360 ;
        RECT 1413.190 1689.160 1413.510 1689.220 ;
        RECT 1493.690 1689.160 1494.010 1689.220 ;
        RECT 1493.690 72.320 1494.010 72.380 ;
        RECT 2560.430 72.320 2560.750 72.380 ;
        RECT 1493.690 72.180 2560.750 72.320 ;
        RECT 1493.690 72.120 1494.010 72.180 ;
        RECT 2560.430 72.120 2560.750 72.180 ;
      LAYER via ;
        RECT 1413.220 1689.160 1413.480 1689.420 ;
        RECT 1493.720 1689.160 1493.980 1689.420 ;
        RECT 1493.720 72.120 1493.980 72.380 ;
        RECT 2560.460 72.120 2560.720 72.380 ;
      LAYER met2 ;
        RECT 1413.120 1700.340 1413.400 1704.000 ;
        RECT 1413.120 1700.000 1413.420 1700.340 ;
        RECT 1413.280 1689.450 1413.420 1700.000 ;
        RECT 1413.220 1689.130 1413.480 1689.450 ;
        RECT 1493.720 1689.130 1493.980 1689.450 ;
        RECT 1493.780 72.410 1493.920 1689.130 ;
        RECT 1493.720 72.090 1493.980 72.410 ;
        RECT 2560.460 72.090 2560.720 72.410 ;
        RECT 2560.520 7.210 2560.660 72.090 ;
        RECT 2560.060 7.070 2560.660 7.210 ;
        RECT 2560.060 2.400 2560.200 7.070 ;
        RECT 2559.850 -4.800 2560.410 2.400 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1436.725 1689.205 1440.115 1689.375 ;
        RECT 1436.725 1688.865 1436.895 1689.205 ;
        RECT 1439.945 1685.125 1440.115 1689.205 ;
      LAYER met1 ;
        RECT 1415.030 1689.020 1415.350 1689.080 ;
        RECT 1436.665 1689.020 1436.955 1689.065 ;
        RECT 1415.030 1688.880 1436.955 1689.020 ;
        RECT 1415.030 1688.820 1415.350 1688.880 ;
        RECT 1436.665 1688.835 1436.955 1688.880 ;
        RECT 1439.885 1685.280 1440.175 1685.325 ;
        RECT 1452.290 1685.280 1452.610 1685.340 ;
        RECT 1439.885 1685.140 1452.610 1685.280 ;
        RECT 1439.885 1685.095 1440.175 1685.140 ;
        RECT 1452.290 1685.080 1452.610 1685.140 ;
        RECT 1452.290 79.460 1452.610 79.520 ;
        RECT 2573.770 79.460 2574.090 79.520 ;
        RECT 1452.290 79.320 2574.090 79.460 ;
        RECT 1452.290 79.260 1452.610 79.320 ;
        RECT 2573.770 79.260 2574.090 79.320 ;
      LAYER via ;
        RECT 1415.060 1688.820 1415.320 1689.080 ;
        RECT 1452.320 1685.080 1452.580 1685.340 ;
        RECT 1452.320 79.260 1452.580 79.520 ;
        RECT 2573.800 79.260 2574.060 79.520 ;
      LAYER met2 ;
        RECT 1414.960 1700.340 1415.240 1704.000 ;
        RECT 1414.960 1700.000 1415.260 1700.340 ;
        RECT 1415.120 1689.110 1415.260 1700.000 ;
        RECT 1415.060 1688.790 1415.320 1689.110 ;
        RECT 1452.320 1685.050 1452.580 1685.370 ;
        RECT 1452.380 79.550 1452.520 1685.050 ;
        RECT 1452.320 79.230 1452.580 79.550 ;
        RECT 2573.800 79.230 2574.060 79.550 ;
        RECT 2573.860 17.410 2574.000 79.230 ;
        RECT 2573.860 17.270 2578.140 17.410 ;
        RECT 2578.000 2.400 2578.140 17.270 ;
        RECT 2577.790 -4.800 2578.350 2.400 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1174.985 1681.045 1175.155 1686.995 ;
        RECT 1207.645 1686.825 1207.815 1688.355 ;
      LAYER mcon ;
        RECT 1207.645 1688.185 1207.815 1688.355 ;
        RECT 1174.985 1686.825 1175.155 1686.995 ;
      LAYER met1 ;
        RECT 1207.585 1688.340 1207.875 1688.385 ;
        RECT 1232.870 1688.340 1233.190 1688.400 ;
        RECT 1207.585 1688.200 1233.190 1688.340 ;
        RECT 1207.585 1688.155 1207.875 1688.200 ;
        RECT 1232.870 1688.140 1233.190 1688.200 ;
        RECT 1174.925 1686.980 1175.215 1687.025 ;
        RECT 1207.585 1686.980 1207.875 1687.025 ;
        RECT 1174.925 1686.840 1207.875 1686.980 ;
        RECT 1174.925 1686.795 1175.215 1686.840 ;
        RECT 1207.585 1686.795 1207.875 1686.840 ;
        RECT 813.810 1681.200 814.130 1681.260 ;
        RECT 1174.925 1681.200 1175.215 1681.245 ;
        RECT 813.810 1681.060 1175.215 1681.200 ;
        RECT 813.810 1681.000 814.130 1681.060 ;
        RECT 1174.925 1681.015 1175.215 1681.060 ;
      LAYER via ;
        RECT 1232.900 1688.140 1233.160 1688.400 ;
        RECT 813.840 1681.000 814.100 1681.260 ;
      LAYER met2 ;
        RECT 1232.800 1700.340 1233.080 1704.000 ;
        RECT 1232.800 1700.000 1233.100 1700.340 ;
        RECT 1232.960 1688.430 1233.100 1700.000 ;
        RECT 1232.900 1688.110 1233.160 1688.430 ;
        RECT 813.840 1680.970 814.100 1681.290 ;
        RECT 813.900 17.410 814.040 1680.970 ;
        RECT 811.600 17.270 814.040 17.410 ;
        RECT 811.600 2.400 811.740 17.270 ;
        RECT 811.390 -4.800 811.950 2.400 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1416.870 1666.580 1417.190 1666.640 ;
        RECT 2594.470 1666.580 2594.790 1666.640 ;
        RECT 1416.870 1666.440 2594.790 1666.580 ;
        RECT 1416.870 1666.380 1417.190 1666.440 ;
        RECT 2594.470 1666.380 2594.790 1666.440 ;
      LAYER via ;
        RECT 1416.900 1666.380 1417.160 1666.640 ;
        RECT 2594.500 1666.380 2594.760 1666.640 ;
      LAYER met2 ;
        RECT 1416.800 1700.340 1417.080 1704.000 ;
        RECT 1416.800 1700.000 1417.100 1700.340 ;
        RECT 1416.960 1666.670 1417.100 1700.000 ;
        RECT 1416.900 1666.350 1417.160 1666.670 ;
        RECT 2594.500 1666.350 2594.760 1666.670 ;
        RECT 2594.560 17.410 2594.700 1666.350 ;
        RECT 2594.560 17.270 2595.620 17.410 ;
        RECT 2595.480 2.400 2595.620 17.270 ;
        RECT 2595.270 -4.800 2595.830 2.400 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1418.710 1685.280 1419.030 1685.340 ;
        RECT 1420.090 1685.280 1420.410 1685.340 ;
        RECT 1418.710 1685.140 1420.410 1685.280 ;
        RECT 1418.710 1685.080 1419.030 1685.140 ;
        RECT 1420.090 1685.080 1420.410 1685.140 ;
        RECT 1420.090 1680.520 1420.410 1680.580 ;
        RECT 2608.270 1680.520 2608.590 1680.580 ;
        RECT 1420.090 1680.380 2608.590 1680.520 ;
        RECT 1420.090 1680.320 1420.410 1680.380 ;
        RECT 2608.270 1680.320 2608.590 1680.380 ;
      LAYER via ;
        RECT 1418.740 1685.080 1419.000 1685.340 ;
        RECT 1420.120 1685.080 1420.380 1685.340 ;
        RECT 1420.120 1680.320 1420.380 1680.580 ;
        RECT 2608.300 1680.320 2608.560 1680.580 ;
      LAYER met2 ;
        RECT 1418.640 1700.340 1418.920 1704.000 ;
        RECT 1418.640 1700.000 1418.940 1700.340 ;
        RECT 1418.800 1685.370 1418.940 1700.000 ;
        RECT 1418.740 1685.050 1419.000 1685.370 ;
        RECT 1420.120 1685.050 1420.380 1685.370 ;
        RECT 1420.180 1680.610 1420.320 1685.050 ;
        RECT 1420.120 1680.290 1420.380 1680.610 ;
        RECT 2608.300 1680.290 2608.560 1680.610 ;
        RECT 2608.360 17.410 2608.500 1680.290 ;
        RECT 2608.360 17.270 2613.560 17.410 ;
        RECT 2613.420 2.400 2613.560 17.270 ;
        RECT 2613.210 -4.800 2613.770 2.400 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1455.125 1686.145 1455.295 1689.715 ;
      LAYER mcon ;
        RECT 1455.125 1689.545 1455.295 1689.715 ;
      LAYER met1 ;
        RECT 1455.065 1689.700 1455.355 1689.745 ;
        RECT 1486.790 1689.700 1487.110 1689.760 ;
        RECT 1455.065 1689.560 1487.110 1689.700 ;
        RECT 1455.065 1689.515 1455.355 1689.560 ;
        RECT 1486.790 1689.500 1487.110 1689.560 ;
        RECT 1421.470 1686.300 1421.790 1686.360 ;
        RECT 1455.065 1686.300 1455.355 1686.345 ;
        RECT 1421.470 1686.160 1455.355 1686.300 ;
        RECT 1421.470 1686.100 1421.790 1686.160 ;
        RECT 1455.065 1686.115 1455.355 1686.160 ;
        RECT 1486.790 93.060 1487.110 93.120 ;
        RECT 2628.970 93.060 2629.290 93.120 ;
        RECT 1486.790 92.920 2629.290 93.060 ;
        RECT 1486.790 92.860 1487.110 92.920 ;
        RECT 2628.970 92.860 2629.290 92.920 ;
      LAYER via ;
        RECT 1486.820 1689.500 1487.080 1689.760 ;
        RECT 1421.500 1686.100 1421.760 1686.360 ;
        RECT 1486.820 92.860 1487.080 93.120 ;
        RECT 2629.000 92.860 2629.260 93.120 ;
      LAYER met2 ;
        RECT 1420.480 1700.340 1420.760 1704.000 ;
        RECT 1420.480 1700.000 1420.780 1700.340 ;
        RECT 1420.640 1685.450 1420.780 1700.000 ;
        RECT 1486.820 1689.470 1487.080 1689.790 ;
        RECT 1421.500 1686.070 1421.760 1686.390 ;
        RECT 1421.560 1685.450 1421.700 1686.070 ;
        RECT 1420.640 1685.310 1421.700 1685.450 ;
        RECT 1486.880 93.150 1487.020 1689.470 ;
        RECT 1486.820 92.830 1487.080 93.150 ;
        RECT 2629.000 92.830 2629.260 93.150 ;
        RECT 2629.060 17.410 2629.200 92.830 ;
        RECT 2629.060 17.270 2631.500 17.410 ;
        RECT 2631.360 2.400 2631.500 17.270 ;
        RECT 2631.150 -4.800 2631.710 2.400 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1422.390 1684.940 1422.710 1685.000 ;
        RECT 1427.450 1684.940 1427.770 1685.000 ;
        RECT 1422.390 1684.800 1427.770 1684.940 ;
        RECT 1422.390 1684.740 1422.710 1684.800 ;
        RECT 1427.450 1684.740 1427.770 1684.800 ;
        RECT 1427.450 1673.380 1427.770 1673.440 ;
        RECT 2642.770 1673.380 2643.090 1673.440 ;
        RECT 1427.450 1673.240 2643.090 1673.380 ;
        RECT 1427.450 1673.180 1427.770 1673.240 ;
        RECT 2642.770 1673.180 2643.090 1673.240 ;
        RECT 2642.770 16.900 2643.090 16.960 ;
        RECT 2649.210 16.900 2649.530 16.960 ;
        RECT 2642.770 16.760 2649.530 16.900 ;
        RECT 2642.770 16.700 2643.090 16.760 ;
        RECT 2649.210 16.700 2649.530 16.760 ;
      LAYER via ;
        RECT 1422.420 1684.740 1422.680 1685.000 ;
        RECT 1427.480 1684.740 1427.740 1685.000 ;
        RECT 1427.480 1673.180 1427.740 1673.440 ;
        RECT 2642.800 1673.180 2643.060 1673.440 ;
        RECT 2642.800 16.700 2643.060 16.960 ;
        RECT 2649.240 16.700 2649.500 16.960 ;
      LAYER met2 ;
        RECT 1422.320 1700.340 1422.600 1704.000 ;
        RECT 1422.320 1700.000 1422.620 1700.340 ;
        RECT 1422.480 1685.030 1422.620 1700.000 ;
        RECT 1422.420 1684.710 1422.680 1685.030 ;
        RECT 1427.480 1684.710 1427.740 1685.030 ;
        RECT 1427.540 1673.470 1427.680 1684.710 ;
        RECT 1427.480 1673.150 1427.740 1673.470 ;
        RECT 2642.800 1673.150 2643.060 1673.470 ;
        RECT 2642.860 16.990 2643.000 1673.150 ;
        RECT 2642.800 16.670 2643.060 16.990 ;
        RECT 2649.240 16.670 2649.500 16.990 ;
        RECT 2649.300 2.400 2649.440 16.670 ;
        RECT 2649.090 -4.800 2649.650 2.400 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1424.230 1690.040 1424.550 1690.100 ;
        RECT 1473.450 1690.040 1473.770 1690.100 ;
        RECT 1424.230 1689.900 1473.770 1690.040 ;
        RECT 1424.230 1689.840 1424.550 1689.900 ;
        RECT 1473.450 1689.840 1473.770 1689.900 ;
        RECT 1473.450 99.860 1473.770 99.920 ;
        RECT 2663.470 99.860 2663.790 99.920 ;
        RECT 1473.450 99.720 2663.790 99.860 ;
        RECT 1473.450 99.660 1473.770 99.720 ;
        RECT 2663.470 99.660 2663.790 99.720 ;
      LAYER via ;
        RECT 1424.260 1689.840 1424.520 1690.100 ;
        RECT 1473.480 1689.840 1473.740 1690.100 ;
        RECT 1473.480 99.660 1473.740 99.920 ;
        RECT 2663.500 99.660 2663.760 99.920 ;
      LAYER met2 ;
        RECT 1424.160 1700.340 1424.440 1704.000 ;
        RECT 1424.160 1700.000 1424.460 1700.340 ;
        RECT 1424.320 1690.130 1424.460 1700.000 ;
        RECT 1424.260 1689.810 1424.520 1690.130 ;
        RECT 1473.480 1689.810 1473.740 1690.130 ;
        RECT 1473.540 99.950 1473.680 1689.810 ;
        RECT 1473.480 99.630 1473.740 99.950 ;
        RECT 2663.500 99.630 2663.760 99.950 ;
        RECT 2663.560 17.410 2663.700 99.630 ;
        RECT 2663.560 17.270 2667.380 17.410 ;
        RECT 2667.240 2.400 2667.380 17.270 ;
        RECT 2667.030 -4.800 2667.590 2.400 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1449.145 1658.945 1449.315 1659.795 ;
      LAYER mcon ;
        RECT 1449.145 1659.625 1449.315 1659.795 ;
      LAYER met1 ;
        RECT 1449.085 1659.780 1449.375 1659.825 ;
        RECT 2684.170 1659.780 2684.490 1659.840 ;
        RECT 1449.085 1659.640 2684.490 1659.780 ;
        RECT 1449.085 1659.595 1449.375 1659.640 ;
        RECT 2684.170 1659.580 2684.490 1659.640 ;
        RECT 1426.070 1659.100 1426.390 1659.160 ;
        RECT 1449.085 1659.100 1449.375 1659.145 ;
        RECT 1426.070 1658.960 1449.375 1659.100 ;
        RECT 1426.070 1658.900 1426.390 1658.960 ;
        RECT 1449.085 1658.915 1449.375 1658.960 ;
      LAYER via ;
        RECT 2684.200 1659.580 2684.460 1659.840 ;
        RECT 1426.100 1658.900 1426.360 1659.160 ;
      LAYER met2 ;
        RECT 1426.000 1700.340 1426.280 1704.000 ;
        RECT 1426.000 1700.000 1426.300 1700.340 ;
        RECT 1426.160 1659.190 1426.300 1700.000 ;
        RECT 2684.200 1659.550 2684.460 1659.870 ;
        RECT 1426.100 1658.870 1426.360 1659.190 ;
        RECT 2684.260 17.410 2684.400 1659.550 ;
        RECT 2684.260 17.270 2684.860 17.410 ;
        RECT 2684.720 2.400 2684.860 17.270 ;
        RECT 2684.510 -4.800 2685.070 2.400 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1427.910 1652.980 1428.230 1653.040 ;
        RECT 2697.970 1652.980 2698.290 1653.040 ;
        RECT 1427.910 1652.840 2698.290 1652.980 ;
        RECT 1427.910 1652.780 1428.230 1652.840 ;
        RECT 2697.970 1652.780 2698.290 1652.840 ;
      LAYER via ;
        RECT 1427.940 1652.780 1428.200 1653.040 ;
        RECT 2698.000 1652.780 2698.260 1653.040 ;
      LAYER met2 ;
        RECT 1427.840 1700.340 1428.120 1704.000 ;
        RECT 1427.840 1700.000 1428.140 1700.340 ;
        RECT 1428.000 1653.070 1428.140 1700.000 ;
        RECT 1427.940 1652.750 1428.200 1653.070 ;
        RECT 2698.000 1652.750 2698.260 1653.070 ;
        RECT 2698.060 17.410 2698.200 1652.750 ;
        RECT 2698.060 17.270 2702.800 17.410 ;
        RECT 2702.660 2.400 2702.800 17.270 ;
        RECT 2702.450 -4.800 2703.010 2.400 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1454.665 1688.185 1454.835 1689.715 ;
      LAYER mcon ;
        RECT 1454.665 1689.545 1454.835 1689.715 ;
      LAYER met1 ;
        RECT 1429.750 1689.700 1430.070 1689.760 ;
        RECT 1454.605 1689.700 1454.895 1689.745 ;
        RECT 1429.750 1689.560 1454.895 1689.700 ;
        RECT 1429.750 1689.500 1430.070 1689.560 ;
        RECT 1454.605 1689.515 1454.895 1689.560 ;
        RECT 1454.605 1688.340 1454.895 1688.385 ;
        RECT 1604.090 1688.340 1604.410 1688.400 ;
        RECT 1454.605 1688.200 1604.410 1688.340 ;
        RECT 1454.605 1688.155 1454.895 1688.200 ;
        RECT 1604.090 1688.140 1604.410 1688.200 ;
        RECT 1604.090 107.000 1604.410 107.060 ;
        RECT 2718.670 107.000 2718.990 107.060 ;
        RECT 1604.090 106.860 2718.990 107.000 ;
        RECT 1604.090 106.800 1604.410 106.860 ;
        RECT 2718.670 106.800 2718.990 106.860 ;
      LAYER via ;
        RECT 1429.780 1689.500 1430.040 1689.760 ;
        RECT 1604.120 1688.140 1604.380 1688.400 ;
        RECT 1604.120 106.800 1604.380 107.060 ;
        RECT 2718.700 106.800 2718.960 107.060 ;
      LAYER met2 ;
        RECT 1429.680 1700.340 1429.960 1704.000 ;
        RECT 1429.680 1700.000 1429.980 1700.340 ;
        RECT 1429.840 1689.790 1429.980 1700.000 ;
        RECT 1429.780 1689.470 1430.040 1689.790 ;
        RECT 1604.120 1688.110 1604.380 1688.430 ;
        RECT 1604.180 107.090 1604.320 1688.110 ;
        RECT 1604.120 106.770 1604.380 107.090 ;
        RECT 2718.700 106.770 2718.960 107.090 ;
        RECT 2718.760 17.410 2718.900 106.770 ;
        RECT 2718.760 17.270 2720.740 17.410 ;
        RECT 2720.600 2.400 2720.740 17.270 ;
        RECT 2720.390 -4.800 2720.950 2.400 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1431.590 1688.340 1431.910 1688.400 ;
        RECT 1432.970 1688.340 1433.290 1688.400 ;
        RECT 1431.590 1688.200 1433.290 1688.340 ;
        RECT 1431.590 1688.140 1431.910 1688.200 ;
        RECT 1432.970 1688.140 1433.290 1688.200 ;
        RECT 1432.970 1666.240 1433.290 1666.300 ;
        RECT 2732.470 1666.240 2732.790 1666.300 ;
        RECT 1432.970 1666.100 2732.790 1666.240 ;
        RECT 1432.970 1666.040 1433.290 1666.100 ;
        RECT 2732.470 1666.040 2732.790 1666.100 ;
        RECT 2732.470 18.260 2732.790 18.320 ;
        RECT 2738.450 18.260 2738.770 18.320 ;
        RECT 2732.470 18.120 2738.770 18.260 ;
        RECT 2732.470 18.060 2732.790 18.120 ;
        RECT 2738.450 18.060 2738.770 18.120 ;
      LAYER via ;
        RECT 1431.620 1688.140 1431.880 1688.400 ;
        RECT 1433.000 1688.140 1433.260 1688.400 ;
        RECT 1433.000 1666.040 1433.260 1666.300 ;
        RECT 2732.500 1666.040 2732.760 1666.300 ;
        RECT 2732.500 18.060 2732.760 18.320 ;
        RECT 2738.480 18.060 2738.740 18.320 ;
      LAYER met2 ;
        RECT 1431.520 1700.340 1431.800 1704.000 ;
        RECT 1431.520 1700.000 1431.820 1700.340 ;
        RECT 1431.680 1688.430 1431.820 1700.000 ;
        RECT 1431.620 1688.110 1431.880 1688.430 ;
        RECT 1433.000 1688.110 1433.260 1688.430 ;
        RECT 1433.060 1666.330 1433.200 1688.110 ;
        RECT 1433.000 1666.010 1433.260 1666.330 ;
        RECT 2732.500 1666.010 2732.760 1666.330 ;
        RECT 2732.560 18.350 2732.700 1666.010 ;
        RECT 2732.500 18.030 2732.760 18.350 ;
        RECT 2738.480 18.030 2738.740 18.350 ;
        RECT 2738.540 2.400 2738.680 18.030 ;
        RECT 2738.330 -4.800 2738.890 2.400 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1433.430 1683.920 1433.750 1683.980 ;
        RECT 1434.350 1683.920 1434.670 1683.980 ;
        RECT 1433.430 1683.780 1434.670 1683.920 ;
        RECT 1433.430 1683.720 1433.750 1683.780 ;
        RECT 1434.350 1683.720 1434.670 1683.780 ;
        RECT 1434.350 1645.500 1434.670 1645.560 ;
        RECT 2753.170 1645.500 2753.490 1645.560 ;
        RECT 1434.350 1645.360 2753.490 1645.500 ;
        RECT 1434.350 1645.300 1434.670 1645.360 ;
        RECT 2753.170 1645.300 2753.490 1645.360 ;
      LAYER via ;
        RECT 1433.460 1683.720 1433.720 1683.980 ;
        RECT 1434.380 1683.720 1434.640 1683.980 ;
        RECT 1434.380 1645.300 1434.640 1645.560 ;
        RECT 2753.200 1645.300 2753.460 1645.560 ;
      LAYER met2 ;
        RECT 1433.360 1700.340 1433.640 1704.000 ;
        RECT 1433.360 1700.000 1433.660 1700.340 ;
        RECT 1433.520 1684.010 1433.660 1700.000 ;
        RECT 1433.460 1683.690 1433.720 1684.010 ;
        RECT 1434.380 1683.690 1434.640 1684.010 ;
        RECT 1434.440 1645.590 1434.580 1683.690 ;
        RECT 1434.380 1645.270 1434.640 1645.590 ;
        RECT 2753.200 1645.270 2753.460 1645.590 ;
        RECT 2753.260 17.410 2753.400 1645.270 ;
        RECT 2753.260 17.270 2756.160 17.410 ;
        RECT 2756.020 2.400 2756.160 17.270 ;
        RECT 2755.810 -4.800 2756.370 2.400 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1152.905 1647.385 1153.075 1685.295 ;
        RECT 1160.265 1685.125 1160.435 1686.655 ;
        RECT 1209.025 1686.485 1209.195 1688.695 ;
      LAYER mcon ;
        RECT 1209.025 1688.525 1209.195 1688.695 ;
        RECT 1160.265 1686.485 1160.435 1686.655 ;
        RECT 1152.905 1685.125 1153.075 1685.295 ;
      LAYER met1 ;
        RECT 1208.965 1688.680 1209.255 1688.725 ;
        RECT 1234.710 1688.680 1235.030 1688.740 ;
        RECT 1208.965 1688.540 1235.030 1688.680 ;
        RECT 1208.965 1688.495 1209.255 1688.540 ;
        RECT 1234.710 1688.480 1235.030 1688.540 ;
        RECT 1160.205 1686.640 1160.495 1686.685 ;
        RECT 1208.965 1686.640 1209.255 1686.685 ;
        RECT 1160.205 1686.500 1209.255 1686.640 ;
        RECT 1160.205 1686.455 1160.495 1686.500 ;
        RECT 1208.965 1686.455 1209.255 1686.500 ;
        RECT 1152.845 1685.280 1153.135 1685.325 ;
        RECT 1160.205 1685.280 1160.495 1685.325 ;
        RECT 1152.845 1685.140 1160.495 1685.280 ;
        RECT 1152.845 1685.095 1153.135 1685.140 ;
        RECT 1160.205 1685.095 1160.495 1685.140 ;
        RECT 1134.890 1647.540 1135.210 1647.600 ;
        RECT 1152.845 1647.540 1153.135 1647.585 ;
        RECT 1134.890 1647.400 1153.135 1647.540 ;
        RECT 1134.890 1647.340 1135.210 1647.400 ;
        RECT 1152.845 1647.355 1153.135 1647.400 ;
        RECT 834.510 58.720 834.830 58.780 ;
        RECT 1134.890 58.720 1135.210 58.780 ;
        RECT 834.510 58.580 1135.210 58.720 ;
        RECT 834.510 58.520 834.830 58.580 ;
        RECT 1134.890 58.520 1135.210 58.580 ;
      LAYER via ;
        RECT 1234.740 1688.480 1235.000 1688.740 ;
        RECT 1134.920 1647.340 1135.180 1647.600 ;
        RECT 834.540 58.520 834.800 58.780 ;
        RECT 1134.920 58.520 1135.180 58.780 ;
      LAYER met2 ;
        RECT 1234.640 1700.340 1234.920 1704.000 ;
        RECT 1234.640 1700.000 1234.940 1700.340 ;
        RECT 1234.800 1688.770 1234.940 1700.000 ;
        RECT 1234.740 1688.450 1235.000 1688.770 ;
        RECT 1134.920 1647.310 1135.180 1647.630 ;
        RECT 1134.980 58.810 1135.120 1647.310 ;
        RECT 834.540 58.490 834.800 58.810 ;
        RECT 1134.920 58.490 1135.180 58.810 ;
        RECT 834.600 17.410 834.740 58.490 ;
        RECT 829.540 17.270 834.740 17.410 ;
        RECT 829.540 2.400 829.680 17.270 ;
        RECT 829.330 -4.800 829.890 2.400 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1435.270 1680.180 1435.590 1680.240 ;
        RECT 2773.870 1680.180 2774.190 1680.240 ;
        RECT 1435.270 1680.040 2774.190 1680.180 ;
        RECT 1435.270 1679.980 1435.590 1680.040 ;
        RECT 2773.870 1679.980 2774.190 1680.040 ;
      LAYER via ;
        RECT 1435.300 1679.980 1435.560 1680.240 ;
        RECT 2773.900 1679.980 2774.160 1680.240 ;
      LAYER met2 ;
        RECT 1435.200 1700.340 1435.480 1704.000 ;
        RECT 1435.200 1700.000 1435.500 1700.340 ;
        RECT 1435.360 1680.270 1435.500 1700.000 ;
        RECT 1435.300 1679.950 1435.560 1680.270 ;
        RECT 2773.900 1679.950 2774.160 1680.270 ;
        RECT 2773.960 2.400 2774.100 1679.950 ;
        RECT 2773.750 -4.800 2774.310 2.400 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1437.110 1688.340 1437.430 1688.400 ;
        RECT 1454.130 1688.340 1454.450 1688.400 ;
        RECT 1437.110 1688.200 1454.450 1688.340 ;
        RECT 1437.110 1688.140 1437.430 1688.200 ;
        RECT 1454.130 1688.140 1454.450 1688.200 ;
        RECT 1454.130 1638.700 1454.450 1638.760 ;
        RECT 2787.670 1638.700 2787.990 1638.760 ;
        RECT 1454.130 1638.560 2787.990 1638.700 ;
        RECT 1454.130 1638.500 1454.450 1638.560 ;
        RECT 2787.670 1638.500 2787.990 1638.560 ;
      LAYER via ;
        RECT 1437.140 1688.140 1437.400 1688.400 ;
        RECT 1454.160 1688.140 1454.420 1688.400 ;
        RECT 1454.160 1638.500 1454.420 1638.760 ;
        RECT 2787.700 1638.500 2787.960 1638.760 ;
      LAYER met2 ;
        RECT 1437.040 1700.340 1437.320 1704.000 ;
        RECT 1437.040 1700.000 1437.340 1700.340 ;
        RECT 1437.200 1688.430 1437.340 1700.000 ;
        RECT 1437.140 1688.110 1437.400 1688.430 ;
        RECT 1454.160 1688.110 1454.420 1688.430 ;
        RECT 1454.220 1638.790 1454.360 1688.110 ;
        RECT 1454.160 1638.470 1454.420 1638.790 ;
        RECT 2787.700 1638.470 2787.960 1638.790 ;
        RECT 2787.760 17.410 2787.900 1638.470 ;
        RECT 2787.760 17.270 2792.040 17.410 ;
        RECT 2791.900 2.400 2792.040 17.270 ;
        RECT 2791.690 -4.800 2792.250 2.400 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1438.950 1659.440 1439.270 1659.500 ;
        RECT 2804.690 1659.440 2805.010 1659.500 ;
        RECT 1438.950 1659.300 2805.010 1659.440 ;
        RECT 1438.950 1659.240 1439.270 1659.300 ;
        RECT 2804.690 1659.240 2805.010 1659.300 ;
        RECT 2804.690 16.900 2805.010 16.960 ;
        RECT 2809.750 16.900 2810.070 16.960 ;
        RECT 2804.690 16.760 2810.070 16.900 ;
        RECT 2804.690 16.700 2805.010 16.760 ;
        RECT 2809.750 16.700 2810.070 16.760 ;
      LAYER via ;
        RECT 1438.980 1659.240 1439.240 1659.500 ;
        RECT 2804.720 1659.240 2804.980 1659.500 ;
        RECT 2804.720 16.700 2804.980 16.960 ;
        RECT 2809.780 16.700 2810.040 16.960 ;
      LAYER met2 ;
        RECT 1438.880 1700.340 1439.160 1704.000 ;
        RECT 1438.880 1700.000 1439.180 1700.340 ;
        RECT 1439.040 1659.530 1439.180 1700.000 ;
        RECT 1438.980 1659.210 1439.240 1659.530 ;
        RECT 2804.720 1659.210 2804.980 1659.530 ;
        RECT 2804.780 16.990 2804.920 1659.210 ;
        RECT 2804.720 16.670 2804.980 16.990 ;
        RECT 2809.780 16.670 2810.040 16.990 ;
        RECT 2809.840 2.400 2809.980 16.670 ;
        RECT 2809.630 -4.800 2810.190 2.400 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1437.110 1665.900 1437.430 1665.960 ;
        RECT 1440.790 1665.900 1441.110 1665.960 ;
        RECT 1437.110 1665.760 1441.110 1665.900 ;
        RECT 1437.110 1665.700 1437.430 1665.760 ;
        RECT 1440.790 1665.700 1441.110 1665.760 ;
        RECT 2822.170 1631.900 2822.490 1631.960 ;
        RECT 1446.400 1631.760 2822.490 1631.900 ;
        RECT 1437.110 1631.560 1437.430 1631.620 ;
        RECT 1446.400 1631.560 1446.540 1631.760 ;
        RECT 2822.170 1631.700 2822.490 1631.760 ;
        RECT 1437.110 1631.420 1446.540 1631.560 ;
        RECT 1437.110 1631.360 1437.430 1631.420 ;
      LAYER via ;
        RECT 1437.140 1665.700 1437.400 1665.960 ;
        RECT 1440.820 1665.700 1441.080 1665.960 ;
        RECT 1437.140 1631.360 1437.400 1631.620 ;
        RECT 2822.200 1631.700 2822.460 1631.960 ;
      LAYER met2 ;
        RECT 1440.720 1700.340 1441.000 1704.000 ;
        RECT 1440.720 1700.000 1441.020 1700.340 ;
        RECT 1440.880 1665.990 1441.020 1700.000 ;
        RECT 1437.140 1665.670 1437.400 1665.990 ;
        RECT 1440.820 1665.670 1441.080 1665.990 ;
        RECT 1437.200 1631.650 1437.340 1665.670 ;
        RECT 2822.200 1631.670 2822.460 1631.990 ;
        RECT 1437.140 1631.330 1437.400 1631.650 ;
        RECT 2822.260 16.730 2822.400 1631.670 ;
        RECT 2822.260 16.590 2827.920 16.730 ;
        RECT 2827.780 2.400 2827.920 16.590 ;
        RECT 2827.570 -4.800 2828.130 2.400 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1442.630 1684.940 1442.950 1685.000 ;
        RECT 1453.670 1684.940 1453.990 1685.000 ;
        RECT 1442.630 1684.800 1453.990 1684.940 ;
        RECT 1442.630 1684.740 1442.950 1684.800 ;
        RECT 1453.670 1684.740 1453.990 1684.800 ;
        RECT 1453.670 1624.760 1453.990 1624.820 ;
        RECT 2842.870 1624.760 2843.190 1624.820 ;
        RECT 1453.670 1624.620 2843.190 1624.760 ;
        RECT 1453.670 1624.560 1453.990 1624.620 ;
        RECT 2842.870 1624.560 2843.190 1624.620 ;
      LAYER via ;
        RECT 1442.660 1684.740 1442.920 1685.000 ;
        RECT 1453.700 1684.740 1453.960 1685.000 ;
        RECT 1453.700 1624.560 1453.960 1624.820 ;
        RECT 2842.900 1624.560 2843.160 1624.820 ;
      LAYER met2 ;
        RECT 1442.560 1700.340 1442.840 1704.000 ;
        RECT 1442.560 1700.000 1442.860 1700.340 ;
        RECT 1442.720 1685.030 1442.860 1700.000 ;
        RECT 1442.660 1684.710 1442.920 1685.030 ;
        RECT 1453.700 1684.710 1453.960 1685.030 ;
        RECT 1453.760 1624.850 1453.900 1684.710 ;
        RECT 1453.700 1624.530 1453.960 1624.850 ;
        RECT 2842.900 1624.530 2843.160 1624.850 ;
        RECT 2842.960 16.730 2843.100 1624.530 ;
        RECT 2842.960 16.590 2845.400 16.730 ;
        RECT 2845.260 2.400 2845.400 16.590 ;
        RECT 2845.050 -4.800 2845.610 2.400 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1444.470 1684.260 1444.790 1684.320 ;
        RECT 1453.210 1684.260 1453.530 1684.320 ;
        RECT 1444.470 1684.120 1453.530 1684.260 ;
        RECT 1444.470 1684.060 1444.790 1684.120 ;
        RECT 1453.210 1684.060 1453.530 1684.120 ;
        RECT 1453.210 1617.960 1453.530 1618.020 ;
        RECT 2856.670 1617.960 2856.990 1618.020 ;
        RECT 1453.210 1617.820 2856.990 1617.960 ;
        RECT 1453.210 1617.760 1453.530 1617.820 ;
        RECT 2856.670 1617.760 2856.990 1617.820 ;
        RECT 2856.670 17.920 2856.990 17.980 ;
        RECT 2863.110 17.920 2863.430 17.980 ;
        RECT 2856.670 17.780 2863.430 17.920 ;
        RECT 2856.670 17.720 2856.990 17.780 ;
        RECT 2863.110 17.720 2863.430 17.780 ;
      LAYER via ;
        RECT 1444.500 1684.060 1444.760 1684.320 ;
        RECT 1453.240 1684.060 1453.500 1684.320 ;
        RECT 1453.240 1617.760 1453.500 1618.020 ;
        RECT 2856.700 1617.760 2856.960 1618.020 ;
        RECT 2856.700 17.720 2856.960 17.980 ;
        RECT 2863.140 17.720 2863.400 17.980 ;
      LAYER met2 ;
        RECT 1444.400 1700.340 1444.680 1704.000 ;
        RECT 1444.400 1700.000 1444.700 1700.340 ;
        RECT 1444.560 1684.350 1444.700 1700.000 ;
        RECT 1444.500 1684.030 1444.760 1684.350 ;
        RECT 1453.240 1684.030 1453.500 1684.350 ;
        RECT 1453.300 1618.050 1453.440 1684.030 ;
        RECT 1453.240 1617.730 1453.500 1618.050 ;
        RECT 2856.700 1617.730 2856.960 1618.050 ;
        RECT 2856.760 18.010 2856.900 1617.730 ;
        RECT 2856.700 17.690 2856.960 18.010 ;
        RECT 2863.140 17.690 2863.400 18.010 ;
        RECT 2863.200 2.400 2863.340 17.690 ;
        RECT 2862.990 -4.800 2863.550 2.400 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1446.310 1673.040 1446.630 1673.100 ;
        RECT 2873.690 1673.040 2874.010 1673.100 ;
        RECT 1446.310 1672.900 2874.010 1673.040 ;
        RECT 1446.310 1672.840 1446.630 1672.900 ;
        RECT 2873.690 1672.840 2874.010 1672.900 ;
        RECT 2873.690 15.200 2874.010 15.260 ;
        RECT 2881.050 15.200 2881.370 15.260 ;
        RECT 2873.690 15.060 2881.370 15.200 ;
        RECT 2873.690 15.000 2874.010 15.060 ;
        RECT 2881.050 15.000 2881.370 15.060 ;
      LAYER via ;
        RECT 1446.340 1672.840 1446.600 1673.100 ;
        RECT 2873.720 1672.840 2873.980 1673.100 ;
        RECT 2873.720 15.000 2873.980 15.260 ;
        RECT 2881.080 15.000 2881.340 15.260 ;
      LAYER met2 ;
        RECT 1446.240 1700.340 1446.520 1704.000 ;
        RECT 1446.240 1700.000 1446.540 1700.340 ;
        RECT 1446.400 1673.130 1446.540 1700.000 ;
        RECT 1446.340 1672.810 1446.600 1673.130 ;
        RECT 2873.720 1672.810 2873.980 1673.130 ;
        RECT 2873.780 15.290 2873.920 1672.810 ;
        RECT 2873.720 14.970 2873.980 15.290 ;
        RECT 2881.080 14.970 2881.340 15.290 ;
        RECT 2881.140 2.400 2881.280 14.970 ;
        RECT 2880.930 -4.800 2881.490 2.400 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1448.150 1652.640 1448.470 1652.700 ;
        RECT 2866.790 1652.640 2867.110 1652.700 ;
        RECT 1448.150 1652.500 2867.110 1652.640 ;
        RECT 1448.150 1652.440 1448.470 1652.500 ;
        RECT 2866.790 1652.440 2867.110 1652.500 ;
        RECT 2866.790 18.600 2867.110 18.660 ;
        RECT 2898.990 18.600 2899.310 18.660 ;
        RECT 2866.790 18.460 2899.310 18.600 ;
        RECT 2866.790 18.400 2867.110 18.460 ;
        RECT 2898.990 18.400 2899.310 18.460 ;
      LAYER via ;
        RECT 1448.180 1652.440 1448.440 1652.700 ;
        RECT 2866.820 1652.440 2867.080 1652.700 ;
        RECT 2866.820 18.400 2867.080 18.660 ;
        RECT 2899.020 18.400 2899.280 18.660 ;
      LAYER met2 ;
        RECT 1448.080 1700.340 1448.360 1704.000 ;
        RECT 1448.080 1700.000 1448.380 1700.340 ;
        RECT 1448.240 1652.730 1448.380 1700.000 ;
        RECT 1448.180 1652.410 1448.440 1652.730 ;
        RECT 2866.820 1652.410 2867.080 1652.730 ;
        RECT 2866.880 18.690 2867.020 1652.410 ;
        RECT 2866.820 18.370 2867.080 18.690 ;
        RECT 2899.020 18.370 2899.280 18.690 ;
        RECT 2899.080 2.400 2899.220 18.370 ;
        RECT 2898.870 -4.800 2899.430 2.400 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 848.310 1674.400 848.630 1674.460 ;
        RECT 1236.550 1674.400 1236.870 1674.460 ;
        RECT 848.310 1674.260 1236.870 1674.400 ;
        RECT 848.310 1674.200 848.630 1674.260 ;
        RECT 1236.550 1674.200 1236.870 1674.260 ;
      LAYER via ;
        RECT 848.340 1674.200 848.600 1674.460 ;
        RECT 1236.580 1674.200 1236.840 1674.460 ;
      LAYER met2 ;
        RECT 1236.480 1700.340 1236.760 1704.000 ;
        RECT 1236.480 1700.000 1236.780 1700.340 ;
        RECT 1236.640 1674.490 1236.780 1700.000 ;
        RECT 848.340 1674.170 848.600 1674.490 ;
        RECT 1236.580 1674.170 1236.840 1674.490 ;
        RECT 848.400 17.410 848.540 1674.170 ;
        RECT 847.020 17.270 848.540 17.410 ;
        RECT 847.020 2.400 847.160 17.270 ;
        RECT 846.810 -4.800 847.370 2.400 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 869.010 1667.600 869.330 1667.660 ;
        RECT 1238.850 1667.600 1239.170 1667.660 ;
        RECT 869.010 1667.460 1239.170 1667.600 ;
        RECT 869.010 1667.400 869.330 1667.460 ;
        RECT 1238.850 1667.400 1239.170 1667.460 ;
      LAYER via ;
        RECT 869.040 1667.400 869.300 1667.660 ;
        RECT 1238.880 1667.400 1239.140 1667.660 ;
      LAYER met2 ;
        RECT 1238.320 1700.410 1238.600 1704.000 ;
        RECT 1238.320 1700.270 1239.080 1700.410 ;
        RECT 1238.320 1700.000 1238.600 1700.270 ;
        RECT 1238.940 1667.690 1239.080 1700.270 ;
        RECT 869.040 1667.370 869.300 1667.690 ;
        RECT 1238.880 1667.370 1239.140 1667.690 ;
        RECT 869.100 24.210 869.240 1667.370 ;
        RECT 864.960 24.070 869.240 24.210 ;
        RECT 864.960 2.400 865.100 24.070 ;
        RECT 864.750 -4.800 865.310 2.400 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1055.845 1680.705 1057.395 1680.875 ;
      LAYER mcon ;
        RECT 1057.225 1680.705 1057.395 1680.875 ;
      LAYER met1 ;
        RECT 882.810 1680.860 883.130 1680.920 ;
        RECT 1055.785 1680.860 1056.075 1680.905 ;
        RECT 882.810 1680.720 1056.075 1680.860 ;
        RECT 882.810 1680.660 883.130 1680.720 ;
        RECT 1055.785 1680.675 1056.075 1680.720 ;
        RECT 1057.165 1680.860 1057.455 1680.905 ;
        RECT 1240.230 1680.860 1240.550 1680.920 ;
        RECT 1057.165 1680.720 1240.550 1680.860 ;
        RECT 1057.165 1680.675 1057.455 1680.720 ;
        RECT 1240.230 1680.660 1240.550 1680.720 ;
      LAYER via ;
        RECT 882.840 1680.660 883.100 1680.920 ;
        RECT 1240.260 1680.660 1240.520 1680.920 ;
      LAYER met2 ;
        RECT 1240.160 1700.340 1240.440 1704.000 ;
        RECT 1240.160 1700.000 1240.460 1700.340 ;
        RECT 1240.320 1680.950 1240.460 1700.000 ;
        RECT 882.840 1680.630 883.100 1680.950 ;
        RECT 1240.260 1680.630 1240.520 1680.950 ;
        RECT 882.900 2.400 883.040 1680.630 ;
        RECT 882.690 -4.800 883.250 2.400 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1235.170 1683.920 1235.490 1683.980 ;
        RECT 1242.070 1683.920 1242.390 1683.980 ;
        RECT 1235.170 1683.780 1242.390 1683.920 ;
        RECT 1235.170 1683.720 1235.490 1683.780 ;
        RECT 1242.070 1683.720 1242.390 1683.780 ;
        RECT 903.510 1660.800 903.830 1660.860 ;
        RECT 1235.170 1660.800 1235.490 1660.860 ;
        RECT 903.510 1660.660 1235.490 1660.800 ;
        RECT 903.510 1660.600 903.830 1660.660 ;
        RECT 1235.170 1660.600 1235.490 1660.660 ;
      LAYER via ;
        RECT 1235.200 1683.720 1235.460 1683.980 ;
        RECT 1242.100 1683.720 1242.360 1683.980 ;
        RECT 903.540 1660.600 903.800 1660.860 ;
        RECT 1235.200 1660.600 1235.460 1660.860 ;
      LAYER met2 ;
        RECT 1242.000 1700.340 1242.280 1704.000 ;
        RECT 1242.000 1700.000 1242.300 1700.340 ;
        RECT 1242.160 1684.010 1242.300 1700.000 ;
        RECT 1235.200 1683.690 1235.460 1684.010 ;
        RECT 1242.100 1683.690 1242.360 1684.010 ;
        RECT 1235.260 1660.890 1235.400 1683.690 ;
        RECT 903.540 1660.570 903.800 1660.890 ;
        RECT 1235.200 1660.570 1235.460 1660.890 ;
        RECT 903.600 24.210 903.740 1660.570 ;
        RECT 900.840 24.070 903.740 24.210 ;
        RECT 900.840 2.400 900.980 24.070 ;
        RECT 900.630 -4.800 901.190 2.400 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1242.070 1678.480 1242.390 1678.540 ;
        RECT 1243.910 1678.480 1244.230 1678.540 ;
        RECT 1242.070 1678.340 1244.230 1678.480 ;
        RECT 1242.070 1678.280 1242.390 1678.340 ;
        RECT 1243.910 1678.280 1244.230 1678.340 ;
        RECT 924.210 1667.940 924.530 1668.000 ;
        RECT 1242.070 1667.940 1242.390 1668.000 ;
        RECT 924.210 1667.800 1242.390 1667.940 ;
        RECT 924.210 1667.740 924.530 1667.800 ;
        RECT 1242.070 1667.740 1242.390 1667.800 ;
        RECT 918.690 2.960 919.010 3.020 ;
        RECT 923.750 2.960 924.070 3.020 ;
        RECT 918.690 2.820 924.070 2.960 ;
        RECT 918.690 2.760 919.010 2.820 ;
        RECT 923.750 2.760 924.070 2.820 ;
      LAYER via ;
        RECT 1242.100 1678.280 1242.360 1678.540 ;
        RECT 1243.940 1678.280 1244.200 1678.540 ;
        RECT 924.240 1667.740 924.500 1668.000 ;
        RECT 1242.100 1667.740 1242.360 1668.000 ;
        RECT 918.720 2.760 918.980 3.020 ;
        RECT 923.780 2.760 924.040 3.020 ;
      LAYER met2 ;
        RECT 1243.840 1700.340 1244.120 1704.000 ;
        RECT 1243.840 1700.000 1244.140 1700.340 ;
        RECT 1244.000 1678.570 1244.140 1700.000 ;
        RECT 1242.100 1678.250 1242.360 1678.570 ;
        RECT 1243.940 1678.250 1244.200 1678.570 ;
        RECT 1242.160 1668.030 1242.300 1678.250 ;
        RECT 924.240 1667.710 924.500 1668.030 ;
        RECT 1242.100 1667.710 1242.360 1668.030 ;
        RECT 924.300 33.730 924.440 1667.710 ;
        RECT 923.840 33.590 924.440 33.730 ;
        RECT 923.840 3.050 923.980 33.590 ;
        RECT 918.720 2.730 918.980 3.050 ;
        RECT 923.780 2.730 924.040 3.050 ;
        RECT 918.780 2.400 918.920 2.730 ;
        RECT 918.570 -4.800 919.130 2.400 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1246.210 1678.140 1246.530 1678.200 ;
        RECT 1248.050 1678.140 1248.370 1678.200 ;
        RECT 1246.210 1678.000 1248.370 1678.140 ;
        RECT 1246.210 1677.940 1246.530 1678.000 ;
        RECT 1248.050 1677.940 1248.370 1678.000 ;
        RECT 936.170 26.420 936.490 26.480 ;
        RECT 1248.050 26.420 1248.370 26.480 ;
        RECT 936.170 26.280 1248.370 26.420 ;
        RECT 936.170 26.220 936.490 26.280 ;
        RECT 1248.050 26.220 1248.370 26.280 ;
      LAYER via ;
        RECT 1246.240 1677.940 1246.500 1678.200 ;
        RECT 1248.080 1677.940 1248.340 1678.200 ;
        RECT 936.200 26.220 936.460 26.480 ;
        RECT 1248.080 26.220 1248.340 26.480 ;
      LAYER met2 ;
        RECT 1245.680 1700.410 1245.960 1704.000 ;
        RECT 1245.680 1700.270 1246.440 1700.410 ;
        RECT 1245.680 1700.000 1245.960 1700.270 ;
        RECT 1246.300 1678.230 1246.440 1700.270 ;
        RECT 1246.240 1677.910 1246.500 1678.230 ;
        RECT 1248.080 1677.910 1248.340 1678.230 ;
        RECT 1248.140 26.510 1248.280 1677.910 ;
        RECT 936.200 26.190 936.460 26.510 ;
        RECT 1248.080 26.190 1248.340 26.510 ;
        RECT 936.260 2.400 936.400 26.190 ;
        RECT 936.050 -4.800 936.610 2.400 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1242.530 1679.160 1242.850 1679.220 ;
        RECT 1247.590 1679.160 1247.910 1679.220 ;
        RECT 1242.530 1679.020 1247.910 1679.160 ;
        RECT 1242.530 1678.960 1242.850 1679.020 ;
        RECT 1247.590 1678.960 1247.910 1679.020 ;
        RECT 954.110 26.760 954.430 26.820 ;
        RECT 1242.530 26.760 1242.850 26.820 ;
        RECT 954.110 26.620 1242.850 26.760 ;
        RECT 954.110 26.560 954.430 26.620 ;
        RECT 1242.530 26.560 1242.850 26.620 ;
      LAYER via ;
        RECT 1242.560 1678.960 1242.820 1679.220 ;
        RECT 1247.620 1678.960 1247.880 1679.220 ;
        RECT 954.140 26.560 954.400 26.820 ;
        RECT 1242.560 26.560 1242.820 26.820 ;
      LAYER met2 ;
        RECT 1247.520 1700.340 1247.800 1704.000 ;
        RECT 1247.520 1700.000 1247.820 1700.340 ;
        RECT 1247.680 1679.250 1247.820 1700.000 ;
        RECT 1242.560 1678.930 1242.820 1679.250 ;
        RECT 1247.620 1678.930 1247.880 1679.250 ;
        RECT 1242.620 26.850 1242.760 1678.930 ;
        RECT 954.140 26.530 954.400 26.850 ;
        RECT 1242.560 26.530 1242.820 26.850 ;
        RECT 954.200 2.400 954.340 26.530 ;
        RECT 953.990 -4.800 954.550 2.400 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 972.050 27.100 972.370 27.160 ;
        RECT 1249.890 27.100 1250.210 27.160 ;
        RECT 972.050 26.960 1250.210 27.100 ;
        RECT 972.050 26.900 972.370 26.960 ;
        RECT 1249.890 26.900 1250.210 26.960 ;
      LAYER via ;
        RECT 972.080 26.900 972.340 27.160 ;
        RECT 1249.920 26.900 1250.180 27.160 ;
      LAYER met2 ;
        RECT 1249.360 1700.410 1249.640 1704.000 ;
        RECT 1249.360 1700.270 1250.120 1700.410 ;
        RECT 1249.360 1700.000 1249.640 1700.270 ;
        RECT 1249.980 27.190 1250.120 1700.270 ;
        RECT 972.080 26.870 972.340 27.190 ;
        RECT 1249.920 26.870 1250.180 27.190 ;
        RECT 972.140 2.400 972.280 26.870 ;
        RECT 971.930 -4.800 972.490 2.400 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1216.770 1660.120 1217.090 1660.180 ;
        RECT 1218.150 1660.120 1218.470 1660.180 ;
        RECT 1216.770 1659.980 1218.470 1660.120 ;
        RECT 1216.770 1659.920 1217.090 1659.980 ;
        RECT 1218.150 1659.920 1218.470 1659.980 ;
        RECT 650.970 25.400 651.290 25.460 ;
        RECT 1218.150 25.400 1218.470 25.460 ;
        RECT 650.970 25.260 1218.470 25.400 ;
        RECT 650.970 25.200 651.290 25.260 ;
        RECT 1218.150 25.200 1218.470 25.260 ;
      LAYER via ;
        RECT 1216.800 1659.920 1217.060 1660.180 ;
        RECT 1218.180 1659.920 1218.440 1660.180 ;
        RECT 651.000 25.200 651.260 25.460 ;
        RECT 1218.180 25.200 1218.440 25.460 ;
      LAYER met2 ;
        RECT 1216.700 1700.340 1216.980 1704.000 ;
        RECT 1216.700 1700.000 1217.000 1700.340 ;
        RECT 1216.860 1660.210 1217.000 1700.000 ;
        RECT 1216.800 1659.890 1217.060 1660.210 ;
        RECT 1218.180 1659.890 1218.440 1660.210 ;
        RECT 1218.240 25.490 1218.380 1659.890 ;
        RECT 651.000 25.170 651.260 25.490 ;
        RECT 1218.180 25.170 1218.440 25.490 ;
        RECT 651.060 2.400 651.200 25.170 ;
        RECT 650.850 -4.800 651.410 2.400 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1221.445 25.925 1221.615 27.455 ;
      LAYER mcon ;
        RECT 1221.445 27.285 1221.615 27.455 ;
      LAYER met1 ;
        RECT 1251.730 1678.820 1252.050 1678.880 ;
        RECT 1255.410 1678.820 1255.730 1678.880 ;
        RECT 1251.730 1678.680 1255.730 1678.820 ;
        RECT 1251.730 1678.620 1252.050 1678.680 ;
        RECT 1255.410 1678.620 1255.730 1678.680 ;
        RECT 989.990 27.440 990.310 27.500 ;
        RECT 1221.385 27.440 1221.675 27.485 ;
        RECT 989.990 27.300 1221.675 27.440 ;
        RECT 989.990 27.240 990.310 27.300 ;
        RECT 1221.385 27.255 1221.675 27.300 ;
        RECT 1221.385 26.080 1221.675 26.125 ;
        RECT 1255.410 26.080 1255.730 26.140 ;
        RECT 1221.385 25.940 1255.730 26.080 ;
        RECT 1221.385 25.895 1221.675 25.940 ;
        RECT 1255.410 25.880 1255.730 25.940 ;
      LAYER via ;
        RECT 1251.760 1678.620 1252.020 1678.880 ;
        RECT 1255.440 1678.620 1255.700 1678.880 ;
        RECT 990.020 27.240 990.280 27.500 ;
        RECT 1255.440 25.880 1255.700 26.140 ;
      LAYER met2 ;
        RECT 1251.200 1700.410 1251.480 1704.000 ;
        RECT 1251.200 1700.270 1251.960 1700.410 ;
        RECT 1251.200 1700.000 1251.480 1700.270 ;
        RECT 1251.820 1678.910 1251.960 1700.270 ;
        RECT 1251.760 1678.590 1252.020 1678.910 ;
        RECT 1255.440 1678.590 1255.700 1678.910 ;
        RECT 990.020 27.210 990.280 27.530 ;
        RECT 990.080 2.400 990.220 27.210 ;
        RECT 1255.500 26.170 1255.640 1678.590 ;
        RECT 1255.440 25.850 1255.700 26.170 ;
        RECT 989.870 -4.800 990.430 2.400 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1249.430 1676.440 1249.750 1676.500 ;
        RECT 1253.110 1676.440 1253.430 1676.500 ;
        RECT 1249.430 1676.300 1253.430 1676.440 ;
        RECT 1249.430 1676.240 1249.750 1676.300 ;
        RECT 1253.110 1676.240 1253.430 1676.300 ;
        RECT 1007.470 23.700 1007.790 23.760 ;
        RECT 1249.430 23.700 1249.750 23.760 ;
        RECT 1007.470 23.560 1249.750 23.700 ;
        RECT 1007.470 23.500 1007.790 23.560 ;
        RECT 1249.430 23.500 1249.750 23.560 ;
      LAYER via ;
        RECT 1249.460 1676.240 1249.720 1676.500 ;
        RECT 1253.140 1676.240 1253.400 1676.500 ;
        RECT 1007.500 23.500 1007.760 23.760 ;
        RECT 1249.460 23.500 1249.720 23.760 ;
      LAYER met2 ;
        RECT 1253.040 1700.340 1253.320 1704.000 ;
        RECT 1253.040 1700.000 1253.340 1700.340 ;
        RECT 1253.200 1676.530 1253.340 1700.000 ;
        RECT 1249.460 1676.210 1249.720 1676.530 ;
        RECT 1253.140 1676.210 1253.400 1676.530 ;
        RECT 1249.520 23.790 1249.660 1676.210 ;
        RECT 1007.500 23.470 1007.760 23.790 ;
        RECT 1249.460 23.470 1249.720 23.790 ;
        RECT 1007.560 2.400 1007.700 23.470 ;
        RECT 1007.350 -4.800 1007.910 2.400 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1025.410 23.360 1025.730 23.420 ;
        RECT 1254.950 23.360 1255.270 23.420 ;
        RECT 1025.410 23.220 1255.270 23.360 ;
        RECT 1025.410 23.160 1025.730 23.220 ;
        RECT 1254.950 23.160 1255.270 23.220 ;
      LAYER via ;
        RECT 1025.440 23.160 1025.700 23.420 ;
        RECT 1254.980 23.160 1255.240 23.420 ;
      LAYER met2 ;
        RECT 1254.880 1700.340 1255.160 1704.000 ;
        RECT 1254.880 1700.000 1255.180 1700.340 ;
        RECT 1255.040 23.450 1255.180 1700.000 ;
        RECT 1025.440 23.130 1025.700 23.450 ;
        RECT 1254.980 23.130 1255.240 23.450 ;
        RECT 1025.500 2.400 1025.640 23.130 ;
        RECT 1025.290 -4.800 1025.850 2.400 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1242.530 1684.940 1242.850 1685.000 ;
        RECT 1256.790 1684.940 1257.110 1685.000 ;
        RECT 1242.530 1684.800 1257.110 1684.940 ;
        RECT 1242.530 1684.740 1242.850 1684.800 ;
        RECT 1256.790 1684.740 1257.110 1684.800 ;
        RECT 1048.410 1681.540 1048.730 1681.600 ;
        RECT 1242.530 1681.540 1242.850 1681.600 ;
        RECT 1048.410 1681.400 1242.850 1681.540 ;
        RECT 1048.410 1681.340 1048.730 1681.400 ;
        RECT 1242.530 1681.340 1242.850 1681.400 ;
        RECT 1043.350 2.960 1043.670 3.020 ;
        RECT 1048.410 2.960 1048.730 3.020 ;
        RECT 1043.350 2.820 1048.730 2.960 ;
        RECT 1043.350 2.760 1043.670 2.820 ;
        RECT 1048.410 2.760 1048.730 2.820 ;
      LAYER via ;
        RECT 1242.560 1684.740 1242.820 1685.000 ;
        RECT 1256.820 1684.740 1257.080 1685.000 ;
        RECT 1048.440 1681.340 1048.700 1681.600 ;
        RECT 1242.560 1681.340 1242.820 1681.600 ;
        RECT 1043.380 2.760 1043.640 3.020 ;
        RECT 1048.440 2.760 1048.700 3.020 ;
      LAYER met2 ;
        RECT 1256.720 1700.340 1257.000 1704.000 ;
        RECT 1256.720 1700.000 1257.020 1700.340 ;
        RECT 1256.880 1685.030 1257.020 1700.000 ;
        RECT 1242.560 1684.710 1242.820 1685.030 ;
        RECT 1256.820 1684.710 1257.080 1685.030 ;
        RECT 1242.620 1681.630 1242.760 1684.710 ;
        RECT 1048.440 1681.310 1048.700 1681.630 ;
        RECT 1242.560 1681.310 1242.820 1681.630 ;
        RECT 1048.500 3.050 1048.640 1681.310 ;
        RECT 1043.380 2.730 1043.640 3.050 ;
        RECT 1048.440 2.730 1048.700 3.050 ;
        RECT 1043.440 2.400 1043.580 2.730 ;
        RECT 1043.230 -4.800 1043.790 2.400 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1256.790 1679.500 1257.110 1679.560 ;
        RECT 1258.630 1679.500 1258.950 1679.560 ;
        RECT 1256.790 1679.360 1258.950 1679.500 ;
        RECT 1256.790 1679.300 1257.110 1679.360 ;
        RECT 1258.630 1679.300 1258.950 1679.360 ;
        RECT 1062.210 1674.740 1062.530 1674.800 ;
        RECT 1256.790 1674.740 1257.110 1674.800 ;
        RECT 1062.210 1674.600 1257.110 1674.740 ;
        RECT 1062.210 1674.540 1062.530 1674.600 ;
        RECT 1256.790 1674.540 1257.110 1674.600 ;
      LAYER via ;
        RECT 1256.820 1679.300 1257.080 1679.560 ;
        RECT 1258.660 1679.300 1258.920 1679.560 ;
        RECT 1062.240 1674.540 1062.500 1674.800 ;
        RECT 1256.820 1674.540 1257.080 1674.800 ;
      LAYER met2 ;
        RECT 1258.560 1700.340 1258.840 1704.000 ;
        RECT 1258.560 1700.000 1258.860 1700.340 ;
        RECT 1258.720 1679.590 1258.860 1700.000 ;
        RECT 1256.820 1679.270 1257.080 1679.590 ;
        RECT 1258.660 1679.270 1258.920 1679.590 ;
        RECT 1256.880 1674.830 1257.020 1679.270 ;
        RECT 1062.240 1674.510 1062.500 1674.830 ;
        RECT 1256.820 1674.510 1257.080 1674.830 ;
        RECT 1062.300 18.090 1062.440 1674.510 ;
        RECT 1061.380 17.950 1062.440 18.090 ;
        RECT 1061.380 2.400 1061.520 17.950 ;
        RECT 1061.170 -4.800 1061.730 2.400 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1082.910 1681.880 1083.230 1681.940 ;
        RECT 1260.470 1681.880 1260.790 1681.940 ;
        RECT 1082.910 1681.740 1260.790 1681.880 ;
        RECT 1082.910 1681.680 1083.230 1681.740 ;
        RECT 1260.470 1681.680 1260.790 1681.740 ;
      LAYER via ;
        RECT 1082.940 1681.680 1083.200 1681.940 ;
        RECT 1260.500 1681.680 1260.760 1681.940 ;
      LAYER met2 ;
        RECT 1260.400 1700.340 1260.680 1704.000 ;
        RECT 1260.400 1700.000 1260.700 1700.340 ;
        RECT 1260.560 1681.970 1260.700 1700.000 ;
        RECT 1082.940 1681.650 1083.200 1681.970 ;
        RECT 1260.500 1681.650 1260.760 1681.970 ;
        RECT 1083.000 18.090 1083.140 1681.650 ;
        RECT 1079.320 17.950 1083.140 18.090 ;
        RECT 1079.320 2.400 1079.460 17.950 ;
        RECT 1079.110 -4.800 1079.670 2.400 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1096.710 1668.280 1097.030 1668.340 ;
        RECT 1261.850 1668.280 1262.170 1668.340 ;
        RECT 1096.710 1668.140 1262.170 1668.280 ;
        RECT 1096.710 1668.080 1097.030 1668.140 ;
        RECT 1261.850 1668.080 1262.170 1668.140 ;
      LAYER via ;
        RECT 1096.740 1668.080 1097.000 1668.340 ;
        RECT 1261.880 1668.080 1262.140 1668.340 ;
      LAYER met2 ;
        RECT 1262.240 1700.340 1262.520 1704.000 ;
        RECT 1262.240 1700.000 1262.540 1700.340 ;
        RECT 1262.400 1680.010 1262.540 1700.000 ;
        RECT 1262.400 1679.870 1263.000 1680.010 ;
        RECT 1262.860 1677.290 1263.000 1679.870 ;
        RECT 1261.940 1677.150 1263.000 1677.290 ;
        RECT 1261.940 1668.370 1262.080 1677.150 ;
        RECT 1096.740 1668.050 1097.000 1668.370 ;
        RECT 1261.880 1668.050 1262.140 1668.370 ;
        RECT 1096.800 2.400 1096.940 1668.050 ;
        RECT 1096.590 -4.800 1097.150 2.400 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1248.050 1684.600 1248.370 1684.660 ;
        RECT 1264.150 1684.600 1264.470 1684.660 ;
        RECT 1248.050 1684.460 1264.470 1684.600 ;
        RECT 1248.050 1684.400 1248.370 1684.460 ;
        RECT 1264.150 1684.400 1264.470 1684.460 ;
        RECT 1117.410 1675.420 1117.730 1675.480 ;
        RECT 1247.590 1675.420 1247.910 1675.480 ;
        RECT 1117.410 1675.280 1247.910 1675.420 ;
        RECT 1117.410 1675.220 1117.730 1675.280 ;
        RECT 1247.590 1675.220 1247.910 1675.280 ;
      LAYER via ;
        RECT 1248.080 1684.400 1248.340 1684.660 ;
        RECT 1264.180 1684.400 1264.440 1684.660 ;
        RECT 1117.440 1675.220 1117.700 1675.480 ;
        RECT 1247.620 1675.220 1247.880 1675.480 ;
      LAYER met2 ;
        RECT 1264.080 1700.340 1264.360 1704.000 ;
        RECT 1264.080 1700.000 1264.380 1700.340 ;
        RECT 1264.240 1684.690 1264.380 1700.000 ;
        RECT 1248.080 1684.370 1248.340 1684.690 ;
        RECT 1264.180 1684.370 1264.440 1684.690 ;
        RECT 1248.140 1678.650 1248.280 1684.370 ;
        RECT 1247.680 1678.510 1248.280 1678.650 ;
        RECT 1247.680 1675.510 1247.820 1678.510 ;
        RECT 1117.440 1675.190 1117.700 1675.510 ;
        RECT 1247.620 1675.190 1247.880 1675.510 ;
        RECT 1117.500 16.730 1117.640 1675.190 ;
        RECT 1114.740 16.590 1117.640 16.730 ;
        RECT 1114.740 2.400 1114.880 16.590 ;
        RECT 1114.530 -4.800 1115.090 2.400 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1214.470 1687.320 1214.790 1687.380 ;
        RECT 1266.450 1687.320 1266.770 1687.380 ;
        RECT 1214.470 1687.180 1266.770 1687.320 ;
        RECT 1214.470 1687.120 1214.790 1687.180 ;
        RECT 1266.450 1687.120 1266.770 1687.180 ;
        RECT 1138.110 1682.560 1138.430 1682.620 ;
        RECT 1214.470 1682.560 1214.790 1682.620 ;
        RECT 1138.110 1682.420 1214.790 1682.560 ;
        RECT 1138.110 1682.360 1138.430 1682.420 ;
        RECT 1214.470 1682.360 1214.790 1682.420 ;
      LAYER via ;
        RECT 1214.500 1687.120 1214.760 1687.380 ;
        RECT 1266.480 1687.120 1266.740 1687.380 ;
        RECT 1138.140 1682.360 1138.400 1682.620 ;
        RECT 1214.500 1682.360 1214.760 1682.620 ;
      LAYER met2 ;
        RECT 1265.920 1700.410 1266.200 1704.000 ;
        RECT 1265.920 1700.270 1266.680 1700.410 ;
        RECT 1265.920 1700.000 1266.200 1700.270 ;
        RECT 1266.540 1687.410 1266.680 1700.270 ;
        RECT 1214.500 1687.090 1214.760 1687.410 ;
        RECT 1266.480 1687.090 1266.740 1687.410 ;
        RECT 1214.560 1682.650 1214.700 1687.090 ;
        RECT 1138.140 1682.330 1138.400 1682.650 ;
        RECT 1214.500 1682.330 1214.760 1682.650 ;
        RECT 1138.200 16.730 1138.340 1682.330 ;
        RECT 1132.680 16.590 1138.340 16.730 ;
        RECT 1132.680 2.400 1132.820 16.590 ;
        RECT 1132.470 -4.800 1133.030 2.400 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1258.705 1676.625 1258.875 1684.955 ;
      LAYER mcon ;
        RECT 1258.705 1684.785 1258.875 1684.955 ;
      LAYER met1 ;
        RECT 1258.645 1684.940 1258.935 1684.985 ;
        RECT 1267.830 1684.940 1268.150 1685.000 ;
        RECT 1258.645 1684.800 1268.150 1684.940 ;
        RECT 1258.645 1684.755 1258.935 1684.800 ;
        RECT 1267.830 1684.740 1268.150 1684.800 ;
        RECT 1258.630 1676.780 1258.950 1676.840 ;
        RECT 1258.435 1676.640 1258.950 1676.780 ;
        RECT 1258.630 1676.580 1258.950 1676.640 ;
        RECT 1151.910 1661.480 1152.230 1661.540 ;
        RECT 1258.630 1661.480 1258.950 1661.540 ;
        RECT 1151.910 1661.340 1258.950 1661.480 ;
        RECT 1151.910 1661.280 1152.230 1661.340 ;
        RECT 1258.630 1661.280 1258.950 1661.340 ;
        RECT 1150.530 2.960 1150.850 3.020 ;
        RECT 1151.910 2.960 1152.230 3.020 ;
        RECT 1150.530 2.820 1152.230 2.960 ;
        RECT 1150.530 2.760 1150.850 2.820 ;
        RECT 1151.910 2.760 1152.230 2.820 ;
      LAYER via ;
        RECT 1267.860 1684.740 1268.120 1685.000 ;
        RECT 1258.660 1676.580 1258.920 1676.840 ;
        RECT 1151.940 1661.280 1152.200 1661.540 ;
        RECT 1258.660 1661.280 1258.920 1661.540 ;
        RECT 1150.560 2.760 1150.820 3.020 ;
        RECT 1151.940 2.760 1152.200 3.020 ;
      LAYER met2 ;
        RECT 1267.760 1700.340 1268.040 1704.000 ;
        RECT 1267.760 1700.000 1268.060 1700.340 ;
        RECT 1267.920 1685.030 1268.060 1700.000 ;
        RECT 1267.860 1684.710 1268.120 1685.030 ;
        RECT 1258.660 1676.550 1258.920 1676.870 ;
        RECT 1258.720 1661.570 1258.860 1676.550 ;
        RECT 1151.940 1661.250 1152.200 1661.570 ;
        RECT 1258.660 1661.250 1258.920 1661.570 ;
        RECT 1152.000 3.050 1152.140 1661.250 ;
        RECT 1150.560 2.730 1150.820 3.050 ;
        RECT 1151.940 2.730 1152.200 3.050 ;
        RECT 1150.620 2.400 1150.760 2.730 ;
        RECT 1150.410 -4.800 1150.970 2.400 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 668.910 25.740 669.230 25.800 ;
        RECT 1218.610 25.740 1218.930 25.800 ;
        RECT 668.910 25.600 1218.930 25.740 ;
        RECT 668.910 25.540 669.230 25.600 ;
        RECT 1218.610 25.540 1218.930 25.600 ;
      LAYER via ;
        RECT 668.940 25.540 669.200 25.800 ;
        RECT 1218.640 25.540 1218.900 25.800 ;
      LAYER met2 ;
        RECT 1218.540 1700.340 1218.820 1704.000 ;
        RECT 1218.540 1700.000 1218.840 1700.340 ;
        RECT 1218.700 25.830 1218.840 1700.000 ;
        RECT 668.940 25.510 669.200 25.830 ;
        RECT 1218.640 25.510 1218.900 25.830 ;
        RECT 669.000 2.400 669.140 25.510 ;
        RECT 668.790 -4.800 669.350 2.400 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1270.130 1678.480 1270.450 1678.540 ;
        RECT 1271.970 1678.480 1272.290 1678.540 ;
        RECT 1270.130 1678.340 1272.290 1678.480 ;
        RECT 1270.130 1678.280 1270.450 1678.340 ;
        RECT 1271.970 1678.280 1272.290 1678.340 ;
        RECT 1168.470 24.040 1168.790 24.100 ;
        RECT 1271.970 24.040 1272.290 24.100 ;
        RECT 1168.470 23.900 1272.290 24.040 ;
        RECT 1168.470 23.840 1168.790 23.900 ;
        RECT 1271.970 23.840 1272.290 23.900 ;
      LAYER via ;
        RECT 1270.160 1678.280 1270.420 1678.540 ;
        RECT 1272.000 1678.280 1272.260 1678.540 ;
        RECT 1168.500 23.840 1168.760 24.100 ;
        RECT 1272.000 23.840 1272.260 24.100 ;
      LAYER met2 ;
        RECT 1269.600 1700.410 1269.880 1704.000 ;
        RECT 1269.600 1700.270 1270.360 1700.410 ;
        RECT 1269.600 1700.000 1269.880 1700.270 ;
        RECT 1270.220 1678.570 1270.360 1700.270 ;
        RECT 1270.160 1678.250 1270.420 1678.570 ;
        RECT 1272.000 1678.250 1272.260 1678.570 ;
        RECT 1272.060 24.130 1272.200 1678.250 ;
        RECT 1168.500 23.810 1168.760 24.130 ;
        RECT 1272.000 23.810 1272.260 24.130 ;
        RECT 1168.560 2.400 1168.700 23.810 ;
        RECT 1168.350 -4.800 1168.910 2.400 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1186.410 24.380 1186.730 24.440 ;
        RECT 1271.050 24.380 1271.370 24.440 ;
        RECT 1186.410 24.240 1271.370 24.380 ;
        RECT 1186.410 24.180 1186.730 24.240 ;
        RECT 1271.050 24.180 1271.370 24.240 ;
      LAYER via ;
        RECT 1186.440 24.180 1186.700 24.440 ;
        RECT 1271.080 24.180 1271.340 24.440 ;
      LAYER met2 ;
        RECT 1271.440 1700.340 1271.720 1704.000 ;
        RECT 1271.440 1700.000 1271.740 1700.340 ;
        RECT 1271.600 1678.140 1271.740 1700.000 ;
        RECT 1271.140 1678.000 1271.740 1678.140 ;
        RECT 1271.140 24.470 1271.280 1678.000 ;
        RECT 1186.440 24.150 1186.700 24.470 ;
        RECT 1271.080 24.150 1271.340 24.470 ;
        RECT 1186.500 12.650 1186.640 24.150 ;
        RECT 1186.040 12.510 1186.640 12.650 ;
        RECT 1186.040 2.400 1186.180 12.510 ;
        RECT 1185.830 -4.800 1186.390 2.400 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1271.510 1676.780 1271.830 1676.840 ;
        RECT 1273.350 1676.780 1273.670 1676.840 ;
        RECT 1271.510 1676.640 1273.670 1676.780 ;
        RECT 1271.510 1676.580 1271.830 1676.640 ;
        RECT 1273.350 1676.580 1273.670 1676.640 ;
        RECT 1203.890 24.720 1204.210 24.780 ;
        RECT 1271.510 24.720 1271.830 24.780 ;
        RECT 1203.890 24.580 1271.830 24.720 ;
        RECT 1203.890 24.520 1204.210 24.580 ;
        RECT 1271.510 24.520 1271.830 24.580 ;
      LAYER via ;
        RECT 1271.540 1676.580 1271.800 1676.840 ;
        RECT 1273.380 1676.580 1273.640 1676.840 ;
        RECT 1203.920 24.520 1204.180 24.780 ;
        RECT 1271.540 24.520 1271.800 24.780 ;
      LAYER met2 ;
        RECT 1273.280 1700.340 1273.560 1704.000 ;
        RECT 1273.280 1700.000 1273.580 1700.340 ;
        RECT 1273.440 1676.870 1273.580 1700.000 ;
        RECT 1271.540 1676.550 1271.800 1676.870 ;
        RECT 1273.380 1676.550 1273.640 1676.870 ;
        RECT 1271.600 24.810 1271.740 1676.550 ;
        RECT 1203.920 24.490 1204.180 24.810 ;
        RECT 1271.540 24.490 1271.800 24.810 ;
        RECT 1203.980 2.400 1204.120 24.490 ;
        RECT 1203.770 -4.800 1204.330 2.400 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1238.390 1685.280 1238.710 1685.340 ;
        RECT 1275.190 1685.280 1275.510 1685.340 ;
        RECT 1238.390 1685.140 1275.510 1685.280 ;
        RECT 1238.390 1685.080 1238.710 1685.140 ;
        RECT 1275.190 1685.080 1275.510 1685.140 ;
        RECT 1221.830 27.440 1222.150 27.500 ;
        RECT 1238.390 27.440 1238.710 27.500 ;
        RECT 1221.830 27.300 1238.710 27.440 ;
        RECT 1221.830 27.240 1222.150 27.300 ;
        RECT 1238.390 27.240 1238.710 27.300 ;
      LAYER via ;
        RECT 1238.420 1685.080 1238.680 1685.340 ;
        RECT 1275.220 1685.080 1275.480 1685.340 ;
        RECT 1221.860 27.240 1222.120 27.500 ;
        RECT 1238.420 27.240 1238.680 27.500 ;
      LAYER met2 ;
        RECT 1275.120 1700.340 1275.400 1704.000 ;
        RECT 1275.120 1700.000 1275.420 1700.340 ;
        RECT 1275.280 1685.370 1275.420 1700.000 ;
        RECT 1238.420 1685.050 1238.680 1685.370 ;
        RECT 1275.220 1685.050 1275.480 1685.370 ;
        RECT 1238.480 27.530 1238.620 1685.050 ;
        RECT 1221.860 27.210 1222.120 27.530 ;
        RECT 1238.420 27.210 1238.680 27.530 ;
        RECT 1221.920 2.400 1222.060 27.210 ;
        RECT 1221.710 -4.800 1222.270 2.400 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1273.810 1683.920 1274.130 1683.980 ;
        RECT 1277.030 1683.920 1277.350 1683.980 ;
        RECT 1273.810 1683.780 1277.350 1683.920 ;
        RECT 1273.810 1683.720 1274.130 1683.780 ;
        RECT 1277.030 1683.720 1277.350 1683.780 ;
        RECT 1239.770 18.600 1240.090 18.660 ;
        RECT 1273.350 18.600 1273.670 18.660 ;
        RECT 1239.770 18.460 1273.670 18.600 ;
        RECT 1239.770 18.400 1240.090 18.460 ;
        RECT 1273.350 18.400 1273.670 18.460 ;
      LAYER via ;
        RECT 1273.840 1683.720 1274.100 1683.980 ;
        RECT 1277.060 1683.720 1277.320 1683.980 ;
        RECT 1239.800 18.400 1240.060 18.660 ;
        RECT 1273.380 18.400 1273.640 18.660 ;
      LAYER met2 ;
        RECT 1276.960 1700.340 1277.240 1704.000 ;
        RECT 1276.960 1700.000 1277.260 1700.340 ;
        RECT 1277.120 1684.010 1277.260 1700.000 ;
        RECT 1273.840 1683.690 1274.100 1684.010 ;
        RECT 1277.060 1683.690 1277.320 1684.010 ;
        RECT 1273.900 1675.930 1274.040 1683.690 ;
        RECT 1273.440 1675.790 1274.040 1675.930 ;
        RECT 1273.440 18.690 1273.580 1675.790 ;
        RECT 1239.800 18.370 1240.060 18.690 ;
        RECT 1273.380 18.370 1273.640 18.690 ;
        RECT 1239.860 2.400 1240.000 18.370 ;
        RECT 1239.650 -4.800 1240.210 2.400 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1274.270 1684.260 1274.590 1684.320 ;
        RECT 1278.870 1684.260 1279.190 1684.320 ;
        RECT 1274.270 1684.120 1279.190 1684.260 ;
        RECT 1274.270 1684.060 1274.590 1684.120 ;
        RECT 1278.870 1684.060 1279.190 1684.120 ;
        RECT 1257.250 16.560 1257.570 16.620 ;
        RECT 1273.810 16.560 1274.130 16.620 ;
        RECT 1257.250 16.420 1274.130 16.560 ;
        RECT 1257.250 16.360 1257.570 16.420 ;
        RECT 1273.810 16.360 1274.130 16.420 ;
      LAYER via ;
        RECT 1274.300 1684.060 1274.560 1684.320 ;
        RECT 1278.900 1684.060 1279.160 1684.320 ;
        RECT 1257.280 16.360 1257.540 16.620 ;
        RECT 1273.840 16.360 1274.100 16.620 ;
      LAYER met2 ;
        RECT 1278.800 1700.340 1279.080 1704.000 ;
        RECT 1278.800 1700.000 1279.100 1700.340 ;
        RECT 1278.960 1684.350 1279.100 1700.000 ;
        RECT 1274.300 1684.030 1274.560 1684.350 ;
        RECT 1278.900 1684.030 1279.160 1684.350 ;
        RECT 1274.360 1675.250 1274.500 1684.030 ;
        RECT 1273.900 1675.110 1274.500 1675.250 ;
        RECT 1273.900 16.650 1274.040 1675.110 ;
        RECT 1257.280 16.330 1257.540 16.650 ;
        RECT 1273.840 16.330 1274.100 16.650 ;
        RECT 1257.340 2.400 1257.480 16.330 ;
        RECT 1257.130 -4.800 1257.690 2.400 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1275.190 20.300 1275.510 20.360 ;
        RECT 1279.330 20.300 1279.650 20.360 ;
        RECT 1275.190 20.160 1279.650 20.300 ;
        RECT 1275.190 20.100 1275.510 20.160 ;
        RECT 1279.330 20.100 1279.650 20.160 ;
      LAYER via ;
        RECT 1275.220 20.100 1275.480 20.360 ;
        RECT 1279.360 20.100 1279.620 20.360 ;
      LAYER met2 ;
        RECT 1280.640 1700.340 1280.920 1704.000 ;
        RECT 1280.640 1700.000 1280.940 1700.340 ;
        RECT 1280.800 1677.290 1280.940 1700.000 ;
        RECT 1279.420 1677.150 1280.940 1677.290 ;
        RECT 1279.420 20.390 1279.560 1677.150 ;
        RECT 1275.220 20.070 1275.480 20.390 ;
        RECT 1279.360 20.070 1279.620 20.390 ;
        RECT 1275.280 2.400 1275.420 20.070 ;
        RECT 1275.070 -4.800 1275.630 2.400 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1282.550 1683.920 1282.870 1683.980 ;
        RECT 1286.690 1683.920 1287.010 1683.980 ;
        RECT 1282.550 1683.780 1287.010 1683.920 ;
        RECT 1282.550 1683.720 1282.870 1683.780 ;
        RECT 1286.690 1683.720 1287.010 1683.780 ;
        RECT 1286.690 20.300 1287.010 20.360 ;
        RECT 1293.130 20.300 1293.450 20.360 ;
        RECT 1286.690 20.160 1293.450 20.300 ;
        RECT 1286.690 20.100 1287.010 20.160 ;
        RECT 1293.130 20.100 1293.450 20.160 ;
      LAYER via ;
        RECT 1282.580 1683.720 1282.840 1683.980 ;
        RECT 1286.720 1683.720 1286.980 1683.980 ;
        RECT 1286.720 20.100 1286.980 20.360 ;
        RECT 1293.160 20.100 1293.420 20.360 ;
      LAYER met2 ;
        RECT 1282.480 1700.340 1282.760 1704.000 ;
        RECT 1282.480 1700.000 1282.780 1700.340 ;
        RECT 1282.640 1684.010 1282.780 1700.000 ;
        RECT 1282.580 1683.690 1282.840 1684.010 ;
        RECT 1286.720 1683.690 1286.980 1684.010 ;
        RECT 1286.780 20.390 1286.920 1683.690 ;
        RECT 1286.720 20.070 1286.980 20.390 ;
        RECT 1293.160 20.070 1293.420 20.390 ;
        RECT 1293.220 2.400 1293.360 20.070 ;
        RECT 1293.010 -4.800 1293.570 2.400 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1284.390 1685.280 1284.710 1685.340 ;
        RECT 1290.370 1685.280 1290.690 1685.340 ;
        RECT 1284.390 1685.140 1290.690 1685.280 ;
        RECT 1284.390 1685.080 1284.710 1685.140 ;
        RECT 1290.370 1685.080 1290.690 1685.140 ;
        RECT 1289.910 19.620 1290.230 19.680 ;
        RECT 1311.070 19.620 1311.390 19.680 ;
        RECT 1289.910 19.480 1311.390 19.620 ;
        RECT 1289.910 19.420 1290.230 19.480 ;
        RECT 1311.070 19.420 1311.390 19.480 ;
      LAYER via ;
        RECT 1284.420 1685.080 1284.680 1685.340 ;
        RECT 1290.400 1685.080 1290.660 1685.340 ;
        RECT 1289.940 19.420 1290.200 19.680 ;
        RECT 1311.100 19.420 1311.360 19.680 ;
      LAYER met2 ;
        RECT 1284.320 1700.340 1284.600 1704.000 ;
        RECT 1284.320 1700.000 1284.620 1700.340 ;
        RECT 1284.480 1685.370 1284.620 1700.000 ;
        RECT 1284.420 1685.050 1284.680 1685.370 ;
        RECT 1290.400 1685.050 1290.660 1685.370 ;
        RECT 1290.460 1683.410 1290.600 1685.050 ;
        RECT 1290.000 1683.270 1290.600 1683.410 ;
        RECT 1290.000 19.710 1290.140 1683.270 ;
        RECT 1289.940 19.390 1290.200 19.710 ;
        RECT 1311.100 19.390 1311.360 19.710 ;
        RECT 1311.160 2.400 1311.300 19.390 ;
        RECT 1310.950 -4.800 1311.510 2.400 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1316.205 1684.105 1316.375 1688.355 ;
      LAYER mcon ;
        RECT 1316.205 1688.185 1316.375 1688.355 ;
      LAYER met1 ;
        RECT 1286.230 1688.340 1286.550 1688.400 ;
        RECT 1316.145 1688.340 1316.435 1688.385 ;
        RECT 1286.230 1688.200 1316.435 1688.340 ;
        RECT 1286.230 1688.140 1286.550 1688.200 ;
        RECT 1316.145 1688.155 1316.435 1688.200 ;
        RECT 1324.870 1684.940 1325.190 1685.000 ;
        RECT 1319.440 1684.800 1325.190 1684.940 ;
        RECT 1316.145 1684.260 1316.435 1684.305 ;
        RECT 1319.440 1684.260 1319.580 1684.800 ;
        RECT 1324.870 1684.740 1325.190 1684.800 ;
        RECT 1316.145 1684.120 1319.580 1684.260 ;
        RECT 1316.145 1684.075 1316.435 1684.120 ;
      LAYER via ;
        RECT 1286.260 1688.140 1286.520 1688.400 ;
        RECT 1324.900 1684.740 1325.160 1685.000 ;
      LAYER met2 ;
        RECT 1286.160 1700.340 1286.440 1704.000 ;
        RECT 1286.160 1700.000 1286.460 1700.340 ;
        RECT 1286.320 1688.430 1286.460 1700.000 ;
        RECT 1286.260 1688.110 1286.520 1688.430 ;
        RECT 1324.900 1684.710 1325.160 1685.030 ;
        RECT 1324.960 28.970 1325.100 1684.710 ;
        RECT 1324.960 28.830 1329.240 28.970 ;
        RECT 1329.100 2.400 1329.240 28.830 ;
        RECT 1328.890 -4.800 1329.450 2.400 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 686.390 26.420 686.710 26.480 ;
        RECT 686.390 26.280 719.740 26.420 ;
        RECT 686.390 26.220 686.710 26.280 ;
        RECT 719.600 26.080 719.740 26.280 ;
        RECT 1219.990 26.080 1220.310 26.140 ;
        RECT 719.600 25.940 1220.310 26.080 ;
        RECT 1219.990 25.880 1220.310 25.940 ;
      LAYER via ;
        RECT 686.420 26.220 686.680 26.480 ;
        RECT 1220.020 25.880 1220.280 26.140 ;
      LAYER met2 ;
        RECT 1220.380 1700.410 1220.660 1704.000 ;
        RECT 1220.080 1700.270 1220.660 1700.410 ;
        RECT 686.420 26.190 686.680 26.510 ;
        RECT 686.480 2.400 686.620 26.190 ;
        RECT 1220.080 26.170 1220.220 1700.270 ;
        RECT 1220.380 1700.000 1220.660 1700.270 ;
        RECT 1220.020 25.850 1220.280 26.170 ;
        RECT 686.270 -4.800 686.830 2.400 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1285.310 1684.260 1285.630 1684.320 ;
        RECT 1288.070 1684.260 1288.390 1684.320 ;
        RECT 1285.310 1684.120 1288.390 1684.260 ;
        RECT 1285.310 1684.060 1285.630 1684.120 ;
        RECT 1288.070 1684.060 1288.390 1684.120 ;
        RECT 1285.310 23.700 1285.630 23.760 ;
        RECT 1346.490 23.700 1346.810 23.760 ;
        RECT 1285.310 23.560 1346.810 23.700 ;
        RECT 1285.310 23.500 1285.630 23.560 ;
        RECT 1346.490 23.500 1346.810 23.560 ;
      LAYER via ;
        RECT 1285.340 1684.060 1285.600 1684.320 ;
        RECT 1288.100 1684.060 1288.360 1684.320 ;
        RECT 1285.340 23.500 1285.600 23.760 ;
        RECT 1346.520 23.500 1346.780 23.760 ;
      LAYER met2 ;
        RECT 1288.000 1700.340 1288.280 1704.000 ;
        RECT 1288.000 1700.000 1288.300 1700.340 ;
        RECT 1288.160 1684.350 1288.300 1700.000 ;
        RECT 1285.340 1684.030 1285.600 1684.350 ;
        RECT 1288.100 1684.030 1288.360 1684.350 ;
        RECT 1285.400 23.790 1285.540 1684.030 ;
        RECT 1285.340 23.470 1285.600 23.790 ;
        RECT 1346.520 23.470 1346.780 23.790 ;
        RECT 1346.580 2.400 1346.720 23.470 ;
        RECT 1346.370 -4.800 1346.930 2.400 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1287.610 1683.920 1287.930 1683.980 ;
        RECT 1289.910 1683.920 1290.230 1683.980 ;
        RECT 1287.610 1683.780 1290.230 1683.920 ;
        RECT 1287.610 1683.720 1287.930 1683.780 ;
        RECT 1289.910 1683.720 1290.230 1683.780 ;
        RECT 1287.610 26.760 1287.930 26.820 ;
        RECT 1364.430 26.760 1364.750 26.820 ;
        RECT 1287.610 26.620 1364.750 26.760 ;
        RECT 1287.610 26.560 1287.930 26.620 ;
        RECT 1364.430 26.560 1364.750 26.620 ;
      LAYER via ;
        RECT 1287.640 1683.720 1287.900 1683.980 ;
        RECT 1289.940 1683.720 1290.200 1683.980 ;
        RECT 1287.640 26.560 1287.900 26.820 ;
        RECT 1364.460 26.560 1364.720 26.820 ;
      LAYER met2 ;
        RECT 1289.840 1700.340 1290.120 1704.000 ;
        RECT 1289.840 1700.000 1290.140 1700.340 ;
        RECT 1290.000 1684.010 1290.140 1700.000 ;
        RECT 1287.640 1683.690 1287.900 1684.010 ;
        RECT 1289.940 1683.690 1290.200 1684.010 ;
        RECT 1287.700 26.850 1287.840 1683.690 ;
        RECT 1287.640 26.530 1287.900 26.850 ;
        RECT 1364.460 26.530 1364.720 26.850 ;
        RECT 1364.520 2.400 1364.660 26.530 ;
        RECT 1364.310 -4.800 1364.870 2.400 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1296.885 807.585 1297.055 855.355 ;
        RECT 1296.425 710.685 1296.595 800.275 ;
        RECT 1296.425 372.725 1296.595 420.835 ;
        RECT 1296.425 131.325 1296.595 179.435 ;
      LAYER mcon ;
        RECT 1296.885 855.185 1297.055 855.355 ;
        RECT 1296.425 800.105 1296.595 800.275 ;
        RECT 1296.425 420.665 1296.595 420.835 ;
        RECT 1296.425 179.265 1296.595 179.435 ;
      LAYER met1 ;
        RECT 1291.750 1684.940 1292.070 1685.000 ;
        RECT 1295.890 1684.940 1296.210 1685.000 ;
        RECT 1291.750 1684.800 1296.210 1684.940 ;
        RECT 1291.750 1684.740 1292.070 1684.800 ;
        RECT 1295.890 1684.740 1296.210 1684.800 ;
        RECT 1295.890 1617.280 1296.210 1617.340 ;
        RECT 1296.810 1617.280 1297.130 1617.340 ;
        RECT 1295.890 1617.140 1297.130 1617.280 ;
        RECT 1295.890 1617.080 1296.210 1617.140 ;
        RECT 1296.810 1617.080 1297.130 1617.140 ;
        RECT 1296.810 1221.520 1297.130 1221.580 ;
        RECT 1296.440 1221.380 1297.130 1221.520 ;
        RECT 1296.440 1221.240 1296.580 1221.380 ;
        RECT 1296.810 1221.320 1297.130 1221.380 ;
        RECT 1296.350 1220.980 1296.670 1221.240 ;
        RECT 1295.890 1200.440 1296.210 1200.500 ;
        RECT 1296.350 1200.440 1296.670 1200.500 ;
        RECT 1295.890 1200.300 1296.670 1200.440 ;
        RECT 1295.890 1200.240 1296.210 1200.300 ;
        RECT 1296.350 1200.240 1296.670 1200.300 ;
        RECT 1297.730 1104.220 1298.050 1104.280 ;
        RECT 1298.190 1104.220 1298.510 1104.280 ;
        RECT 1297.730 1104.080 1298.510 1104.220 ;
        RECT 1297.730 1104.020 1298.050 1104.080 ;
        RECT 1298.190 1104.020 1298.510 1104.080 ;
        RECT 1296.810 1062.740 1297.130 1062.800 ;
        RECT 1298.190 1062.740 1298.510 1062.800 ;
        RECT 1296.810 1062.600 1298.510 1062.740 ;
        RECT 1296.810 1062.540 1297.130 1062.600 ;
        RECT 1298.190 1062.540 1298.510 1062.600 ;
        RECT 1296.350 903.960 1296.670 904.020 ;
        RECT 1296.810 903.960 1297.130 904.020 ;
        RECT 1296.350 903.820 1297.130 903.960 ;
        RECT 1296.350 903.760 1296.670 903.820 ;
        RECT 1296.810 903.760 1297.130 903.820 ;
        RECT 1296.810 855.340 1297.130 855.400 ;
        RECT 1296.615 855.200 1297.130 855.340 ;
        RECT 1296.810 855.140 1297.130 855.200 ;
        RECT 1296.810 807.740 1297.130 807.800 ;
        RECT 1296.615 807.600 1297.130 807.740 ;
        RECT 1296.810 807.540 1297.130 807.600 ;
        RECT 1296.365 800.260 1296.655 800.305 ;
        RECT 1296.810 800.260 1297.130 800.320 ;
        RECT 1296.365 800.120 1297.130 800.260 ;
        RECT 1296.365 800.075 1296.655 800.120 ;
        RECT 1296.810 800.060 1297.130 800.120 ;
        RECT 1296.350 710.840 1296.670 710.900 ;
        RECT 1296.155 710.700 1296.670 710.840 ;
        RECT 1296.350 710.640 1296.670 710.700 ;
        RECT 1296.350 613.740 1296.670 614.000 ;
        RECT 1296.440 613.600 1296.580 613.740 ;
        RECT 1296.810 613.600 1297.130 613.660 ;
        RECT 1296.440 613.460 1297.130 613.600 ;
        RECT 1296.810 613.400 1297.130 613.460 ;
        RECT 1296.810 428.980 1297.130 429.040 ;
        RECT 1296.440 428.840 1297.130 428.980 ;
        RECT 1296.440 428.700 1296.580 428.840 ;
        RECT 1296.810 428.780 1297.130 428.840 ;
        RECT 1296.350 428.440 1296.670 428.700 ;
        RECT 1296.350 420.820 1296.670 420.880 ;
        RECT 1296.155 420.680 1296.670 420.820 ;
        RECT 1296.350 420.620 1296.670 420.680 ;
        RECT 1296.365 372.880 1296.655 372.925 ;
        RECT 1296.810 372.880 1297.130 372.940 ;
        RECT 1296.365 372.740 1297.130 372.880 ;
        RECT 1296.365 372.695 1296.655 372.740 ;
        RECT 1296.810 372.680 1297.130 372.740 ;
        RECT 1296.350 331.400 1296.670 331.460 ;
        RECT 1296.810 331.400 1297.130 331.460 ;
        RECT 1296.350 331.260 1297.130 331.400 ;
        RECT 1296.350 331.200 1296.670 331.260 ;
        RECT 1296.810 331.200 1297.130 331.260 ;
        RECT 1296.350 217.500 1296.670 217.560 ;
        RECT 1297.270 217.500 1297.590 217.560 ;
        RECT 1296.350 217.360 1297.590 217.500 ;
        RECT 1296.350 217.300 1296.670 217.360 ;
        RECT 1297.270 217.300 1297.590 217.360 ;
        RECT 1296.365 179.420 1296.655 179.465 ;
        RECT 1297.270 179.420 1297.590 179.480 ;
        RECT 1296.365 179.280 1297.590 179.420 ;
        RECT 1296.365 179.235 1296.655 179.280 ;
        RECT 1297.270 179.220 1297.590 179.280 ;
        RECT 1296.350 131.480 1296.670 131.540 ;
        RECT 1296.155 131.340 1296.670 131.480 ;
        RECT 1296.350 131.280 1296.670 131.340 ;
        RECT 1296.350 26.420 1296.670 26.480 ;
        RECT 1382.370 26.420 1382.690 26.480 ;
        RECT 1296.350 26.280 1382.690 26.420 ;
        RECT 1296.350 26.220 1296.670 26.280 ;
        RECT 1382.370 26.220 1382.690 26.280 ;
      LAYER via ;
        RECT 1291.780 1684.740 1292.040 1685.000 ;
        RECT 1295.920 1684.740 1296.180 1685.000 ;
        RECT 1295.920 1617.080 1296.180 1617.340 ;
        RECT 1296.840 1617.080 1297.100 1617.340 ;
        RECT 1296.840 1221.320 1297.100 1221.580 ;
        RECT 1296.380 1220.980 1296.640 1221.240 ;
        RECT 1295.920 1200.240 1296.180 1200.500 ;
        RECT 1296.380 1200.240 1296.640 1200.500 ;
        RECT 1297.760 1104.020 1298.020 1104.280 ;
        RECT 1298.220 1104.020 1298.480 1104.280 ;
        RECT 1296.840 1062.540 1297.100 1062.800 ;
        RECT 1298.220 1062.540 1298.480 1062.800 ;
        RECT 1296.380 903.760 1296.640 904.020 ;
        RECT 1296.840 903.760 1297.100 904.020 ;
        RECT 1296.840 855.140 1297.100 855.400 ;
        RECT 1296.840 807.540 1297.100 807.800 ;
        RECT 1296.840 800.060 1297.100 800.320 ;
        RECT 1296.380 710.640 1296.640 710.900 ;
        RECT 1296.380 613.740 1296.640 614.000 ;
        RECT 1296.840 613.400 1297.100 613.660 ;
        RECT 1296.840 428.780 1297.100 429.040 ;
        RECT 1296.380 428.440 1296.640 428.700 ;
        RECT 1296.380 420.620 1296.640 420.880 ;
        RECT 1296.840 372.680 1297.100 372.940 ;
        RECT 1296.380 331.200 1296.640 331.460 ;
        RECT 1296.840 331.200 1297.100 331.460 ;
        RECT 1296.380 217.300 1296.640 217.560 ;
        RECT 1297.300 217.300 1297.560 217.560 ;
        RECT 1297.300 179.220 1297.560 179.480 ;
        RECT 1296.380 131.280 1296.640 131.540 ;
        RECT 1296.380 26.220 1296.640 26.480 ;
        RECT 1382.400 26.220 1382.660 26.480 ;
      LAYER met2 ;
        RECT 1291.680 1700.340 1291.960 1704.000 ;
        RECT 1291.680 1700.000 1291.980 1700.340 ;
        RECT 1291.840 1685.030 1291.980 1700.000 ;
        RECT 1291.780 1684.710 1292.040 1685.030 ;
        RECT 1295.920 1684.710 1296.180 1685.030 ;
        RECT 1295.980 1617.370 1296.120 1684.710 ;
        RECT 1295.920 1617.050 1296.180 1617.370 ;
        RECT 1296.840 1617.050 1297.100 1617.370 ;
        RECT 1296.900 1269.970 1297.040 1617.050 ;
        RECT 1296.440 1269.830 1297.040 1269.970 ;
        RECT 1296.440 1269.290 1296.580 1269.830 ;
        RECT 1296.440 1269.150 1297.040 1269.290 ;
        RECT 1296.900 1221.610 1297.040 1269.150 ;
        RECT 1296.840 1221.290 1297.100 1221.610 ;
        RECT 1296.380 1220.950 1296.640 1221.270 ;
        RECT 1296.440 1200.530 1296.580 1220.950 ;
        RECT 1295.920 1200.210 1296.180 1200.530 ;
        RECT 1296.380 1200.210 1296.640 1200.530 ;
        RECT 1295.980 1159.130 1296.120 1200.210 ;
        RECT 1295.980 1158.990 1297.500 1159.130 ;
        RECT 1297.360 1140.770 1297.500 1158.990 ;
        RECT 1297.360 1140.630 1297.960 1140.770 ;
        RECT 1297.820 1104.310 1297.960 1140.630 ;
        RECT 1297.760 1103.990 1298.020 1104.310 ;
        RECT 1298.220 1103.990 1298.480 1104.310 ;
        RECT 1298.280 1062.830 1298.420 1103.990 ;
        RECT 1296.840 1062.510 1297.100 1062.830 ;
        RECT 1298.220 1062.510 1298.480 1062.830 ;
        RECT 1296.900 904.050 1297.040 1062.510 ;
        RECT 1296.380 903.730 1296.640 904.050 ;
        RECT 1296.840 903.730 1297.100 904.050 ;
        RECT 1296.440 855.850 1296.580 903.730 ;
        RECT 1296.440 855.710 1297.040 855.850 ;
        RECT 1296.900 855.430 1297.040 855.710 ;
        RECT 1296.840 855.110 1297.100 855.430 ;
        RECT 1296.840 807.510 1297.100 807.830 ;
        RECT 1296.900 800.350 1297.040 807.510 ;
        RECT 1296.840 800.030 1297.100 800.350 ;
        RECT 1296.380 710.610 1296.640 710.930 ;
        RECT 1296.440 614.030 1296.580 710.610 ;
        RECT 1296.380 613.710 1296.640 614.030 ;
        RECT 1296.840 613.370 1297.100 613.690 ;
        RECT 1296.900 429.070 1297.040 613.370 ;
        RECT 1296.840 428.750 1297.100 429.070 ;
        RECT 1296.380 428.410 1296.640 428.730 ;
        RECT 1296.440 420.910 1296.580 428.410 ;
        RECT 1296.380 420.590 1296.640 420.910 ;
        RECT 1296.840 372.650 1297.100 372.970 ;
        RECT 1296.900 331.490 1297.040 372.650 ;
        RECT 1296.380 331.170 1296.640 331.490 ;
        RECT 1296.840 331.170 1297.100 331.490 ;
        RECT 1296.440 217.590 1296.580 331.170 ;
        RECT 1296.380 217.270 1296.640 217.590 ;
        RECT 1297.300 217.270 1297.560 217.590 ;
        RECT 1297.360 179.510 1297.500 217.270 ;
        RECT 1297.300 179.190 1297.560 179.510 ;
        RECT 1296.380 131.250 1296.640 131.570 ;
        RECT 1296.440 56.170 1296.580 131.250 ;
        RECT 1295.980 56.030 1296.580 56.170 ;
        RECT 1295.980 37.130 1296.120 56.030 ;
        RECT 1295.980 36.990 1296.580 37.130 ;
        RECT 1296.440 26.510 1296.580 36.990 ;
        RECT 1296.380 26.190 1296.640 26.510 ;
        RECT 1382.400 26.190 1382.660 26.510 ;
        RECT 1382.460 2.400 1382.600 26.190 ;
        RECT 1382.250 -4.800 1382.810 2.400 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1292.745 1200.625 1292.915 1222.215 ;
        RECT 1293.205 855.865 1293.375 903.975 ;
        RECT 1293.205 807.245 1293.375 855.355 ;
        RECT 1293.205 710.685 1293.375 758.795 ;
        RECT 1292.745 607.325 1292.915 655.435 ;
        RECT 1293.205 510.765 1293.375 558.875 ;
        RECT 1292.745 421.005 1292.915 486.455 ;
        RECT 1292.745 324.785 1292.915 372.555 ;
        RECT 1293.205 227.885 1293.375 317.475 ;
      LAYER mcon ;
        RECT 1292.745 1222.045 1292.915 1222.215 ;
        RECT 1293.205 903.805 1293.375 903.975 ;
        RECT 1293.205 855.185 1293.375 855.355 ;
        RECT 1293.205 758.625 1293.375 758.795 ;
        RECT 1292.745 655.265 1292.915 655.435 ;
        RECT 1293.205 558.705 1293.375 558.875 ;
        RECT 1292.745 486.285 1292.915 486.455 ;
        RECT 1292.745 372.385 1292.915 372.555 ;
        RECT 1293.205 317.305 1293.375 317.475 ;
      LAYER met1 ;
        RECT 1292.670 1642.100 1292.990 1642.160 ;
        RECT 1293.130 1642.100 1293.450 1642.160 ;
        RECT 1292.670 1641.960 1293.450 1642.100 ;
        RECT 1292.670 1641.900 1292.990 1641.960 ;
        RECT 1293.130 1641.900 1293.450 1641.960 ;
        RECT 1292.685 1222.200 1292.975 1222.245 ;
        RECT 1293.130 1222.200 1293.450 1222.260 ;
        RECT 1292.685 1222.060 1293.450 1222.200 ;
        RECT 1292.685 1222.015 1292.975 1222.060 ;
        RECT 1293.130 1222.000 1293.450 1222.060 ;
        RECT 1292.670 1200.780 1292.990 1200.840 ;
        RECT 1292.475 1200.640 1292.990 1200.780 ;
        RECT 1292.670 1200.580 1292.990 1200.640 ;
        RECT 1292.670 1152.500 1292.990 1152.560 ;
        RECT 1293.130 1152.500 1293.450 1152.560 ;
        RECT 1292.670 1152.360 1293.450 1152.500 ;
        RECT 1292.670 1152.300 1292.990 1152.360 ;
        RECT 1293.130 1152.300 1293.450 1152.360 ;
        RECT 1293.130 1014.460 1293.450 1014.520 ;
        RECT 1293.590 1014.460 1293.910 1014.520 ;
        RECT 1293.130 1014.320 1293.910 1014.460 ;
        RECT 1293.130 1014.260 1293.450 1014.320 ;
        RECT 1293.590 1014.260 1293.910 1014.320 ;
        RECT 1293.130 903.960 1293.450 904.020 ;
        RECT 1292.935 903.820 1293.450 903.960 ;
        RECT 1293.130 903.760 1293.450 903.820 ;
        RECT 1293.130 856.020 1293.450 856.080 ;
        RECT 1292.935 855.880 1293.450 856.020 ;
        RECT 1293.130 855.820 1293.450 855.880 ;
        RECT 1293.130 855.340 1293.450 855.400 ;
        RECT 1292.935 855.200 1293.450 855.340 ;
        RECT 1293.130 855.140 1293.450 855.200 ;
        RECT 1293.130 807.400 1293.450 807.460 ;
        RECT 1292.935 807.260 1293.450 807.400 ;
        RECT 1293.130 807.200 1293.450 807.260 ;
        RECT 1293.130 758.780 1293.450 758.840 ;
        RECT 1292.935 758.640 1293.450 758.780 ;
        RECT 1293.130 758.580 1293.450 758.640 ;
        RECT 1293.130 710.840 1293.450 710.900 ;
        RECT 1292.935 710.700 1293.450 710.840 ;
        RECT 1293.130 710.640 1293.450 710.700 ;
        RECT 1292.670 655.420 1292.990 655.480 ;
        RECT 1292.475 655.280 1292.990 655.420 ;
        RECT 1292.670 655.220 1292.990 655.280 ;
        RECT 1292.685 607.480 1292.975 607.525 ;
        RECT 1293.130 607.480 1293.450 607.540 ;
        RECT 1292.685 607.340 1293.450 607.480 ;
        RECT 1292.685 607.295 1292.975 607.340 ;
        RECT 1293.130 607.280 1293.450 607.340 ;
        RECT 1293.130 558.860 1293.450 558.920 ;
        RECT 1292.935 558.720 1293.450 558.860 ;
        RECT 1293.130 558.660 1293.450 558.720 ;
        RECT 1293.130 510.920 1293.450 510.980 ;
        RECT 1292.935 510.780 1293.450 510.920 ;
        RECT 1293.130 510.720 1293.450 510.780 ;
        RECT 1292.685 486.440 1292.975 486.485 ;
        RECT 1293.130 486.440 1293.450 486.500 ;
        RECT 1292.685 486.300 1293.450 486.440 ;
        RECT 1292.685 486.255 1292.975 486.300 ;
        RECT 1293.130 486.240 1293.450 486.300 ;
        RECT 1292.670 421.160 1292.990 421.220 ;
        RECT 1292.475 421.020 1292.990 421.160 ;
        RECT 1292.670 420.960 1292.990 421.020 ;
        RECT 1292.685 372.540 1292.975 372.585 ;
        RECT 1293.130 372.540 1293.450 372.600 ;
        RECT 1292.685 372.400 1293.450 372.540 ;
        RECT 1292.685 372.355 1292.975 372.400 ;
        RECT 1293.130 372.340 1293.450 372.400 ;
        RECT 1292.670 324.940 1292.990 325.000 ;
        RECT 1292.475 324.800 1292.990 324.940 ;
        RECT 1292.670 324.740 1292.990 324.800 ;
        RECT 1292.670 324.260 1292.990 324.320 ;
        RECT 1293.130 324.260 1293.450 324.320 ;
        RECT 1292.670 324.120 1293.450 324.260 ;
        RECT 1292.670 324.060 1292.990 324.120 ;
        RECT 1293.130 324.060 1293.450 324.120 ;
        RECT 1293.130 317.460 1293.450 317.520 ;
        RECT 1292.935 317.320 1293.450 317.460 ;
        RECT 1293.130 317.260 1293.450 317.320 ;
        RECT 1293.130 228.040 1293.450 228.100 ;
        RECT 1292.935 227.900 1293.450 228.040 ;
        RECT 1293.130 227.840 1293.450 227.900 ;
        RECT 1292.670 90.000 1292.990 90.060 ;
        RECT 1293.130 90.000 1293.450 90.060 ;
        RECT 1292.670 89.860 1293.450 90.000 ;
        RECT 1292.670 89.800 1292.990 89.860 ;
        RECT 1293.130 89.800 1293.450 89.860 ;
        RECT 1292.670 25.740 1292.990 25.800 ;
        RECT 1400.310 25.740 1400.630 25.800 ;
        RECT 1292.670 25.600 1400.630 25.740 ;
        RECT 1292.670 25.540 1292.990 25.600 ;
        RECT 1400.310 25.540 1400.630 25.600 ;
      LAYER via ;
        RECT 1292.700 1641.900 1292.960 1642.160 ;
        RECT 1293.160 1641.900 1293.420 1642.160 ;
        RECT 1293.160 1222.000 1293.420 1222.260 ;
        RECT 1292.700 1200.580 1292.960 1200.840 ;
        RECT 1292.700 1152.300 1292.960 1152.560 ;
        RECT 1293.160 1152.300 1293.420 1152.560 ;
        RECT 1293.160 1014.260 1293.420 1014.520 ;
        RECT 1293.620 1014.260 1293.880 1014.520 ;
        RECT 1293.160 903.760 1293.420 904.020 ;
        RECT 1293.160 855.820 1293.420 856.080 ;
        RECT 1293.160 855.140 1293.420 855.400 ;
        RECT 1293.160 807.200 1293.420 807.460 ;
        RECT 1293.160 758.580 1293.420 758.840 ;
        RECT 1293.160 710.640 1293.420 710.900 ;
        RECT 1292.700 655.220 1292.960 655.480 ;
        RECT 1293.160 607.280 1293.420 607.540 ;
        RECT 1293.160 558.660 1293.420 558.920 ;
        RECT 1293.160 510.720 1293.420 510.980 ;
        RECT 1293.160 486.240 1293.420 486.500 ;
        RECT 1292.700 420.960 1292.960 421.220 ;
        RECT 1293.160 372.340 1293.420 372.600 ;
        RECT 1292.700 324.740 1292.960 325.000 ;
        RECT 1292.700 324.060 1292.960 324.320 ;
        RECT 1293.160 324.060 1293.420 324.320 ;
        RECT 1293.160 317.260 1293.420 317.520 ;
        RECT 1293.160 227.840 1293.420 228.100 ;
        RECT 1292.700 89.800 1292.960 90.060 ;
        RECT 1293.160 89.800 1293.420 90.060 ;
        RECT 1292.700 25.540 1292.960 25.800 ;
        RECT 1400.340 25.540 1400.600 25.800 ;
      LAYER met2 ;
        RECT 1293.520 1700.340 1293.800 1704.000 ;
        RECT 1293.520 1700.000 1293.820 1700.340 ;
        RECT 1293.680 1665.730 1293.820 1700.000 ;
        RECT 1292.760 1665.590 1293.820 1665.730 ;
        RECT 1292.760 1642.190 1292.900 1665.590 ;
        RECT 1292.700 1641.870 1292.960 1642.190 ;
        RECT 1293.160 1641.870 1293.420 1642.190 ;
        RECT 1293.220 1269.970 1293.360 1641.870 ;
        RECT 1292.760 1269.830 1293.360 1269.970 ;
        RECT 1292.760 1269.290 1292.900 1269.830 ;
        RECT 1292.760 1269.150 1293.360 1269.290 ;
        RECT 1293.220 1222.290 1293.360 1269.150 ;
        RECT 1293.160 1221.970 1293.420 1222.290 ;
        RECT 1292.700 1200.550 1292.960 1200.870 ;
        RECT 1292.760 1152.590 1292.900 1200.550 ;
        RECT 1292.700 1152.270 1292.960 1152.590 ;
        RECT 1293.160 1152.270 1293.420 1152.590 ;
        RECT 1293.220 1128.530 1293.360 1152.270 ;
        RECT 1292.760 1128.390 1293.360 1128.530 ;
        RECT 1292.760 1090.450 1292.900 1128.390 ;
        RECT 1292.760 1090.310 1293.820 1090.450 ;
        RECT 1293.680 1014.550 1293.820 1090.310 ;
        RECT 1293.160 1014.230 1293.420 1014.550 ;
        RECT 1293.620 1014.230 1293.880 1014.550 ;
        RECT 1293.220 904.050 1293.360 1014.230 ;
        RECT 1293.160 903.730 1293.420 904.050 ;
        RECT 1293.160 855.790 1293.420 856.110 ;
        RECT 1293.220 855.430 1293.360 855.790 ;
        RECT 1293.160 855.110 1293.420 855.430 ;
        RECT 1293.160 807.170 1293.420 807.490 ;
        RECT 1293.220 758.870 1293.360 807.170 ;
        RECT 1293.160 758.550 1293.420 758.870 ;
        RECT 1293.160 710.610 1293.420 710.930 ;
        RECT 1293.220 662.730 1293.360 710.610 ;
        RECT 1292.760 662.590 1293.360 662.730 ;
        RECT 1292.760 655.510 1292.900 662.590 ;
        RECT 1292.700 655.190 1292.960 655.510 ;
        RECT 1293.160 607.250 1293.420 607.570 ;
        RECT 1293.220 558.950 1293.360 607.250 ;
        RECT 1293.160 558.630 1293.420 558.950 ;
        RECT 1293.160 510.690 1293.420 511.010 ;
        RECT 1293.220 486.530 1293.360 510.690 ;
        RECT 1293.160 486.210 1293.420 486.530 ;
        RECT 1292.700 420.930 1292.960 421.250 ;
        RECT 1292.760 420.765 1292.900 420.930 ;
        RECT 1292.690 420.395 1292.970 420.765 ;
        RECT 1293.610 419.715 1293.890 420.085 ;
        RECT 1293.680 400.250 1293.820 419.715 ;
        RECT 1293.220 400.110 1293.820 400.250 ;
        RECT 1293.220 372.630 1293.360 400.110 ;
        RECT 1293.160 372.310 1293.420 372.630 ;
        RECT 1292.700 324.710 1292.960 325.030 ;
        RECT 1292.760 324.350 1292.900 324.710 ;
        RECT 1292.700 324.030 1292.960 324.350 ;
        RECT 1293.160 324.030 1293.420 324.350 ;
        RECT 1293.220 317.550 1293.360 324.030 ;
        RECT 1293.160 317.230 1293.420 317.550 ;
        RECT 1293.160 227.810 1293.420 228.130 ;
        RECT 1293.220 152.050 1293.360 227.810 ;
        RECT 1292.760 151.910 1293.360 152.050 ;
        RECT 1292.760 90.090 1292.900 151.910 ;
        RECT 1292.700 89.770 1292.960 90.090 ;
        RECT 1293.160 89.770 1293.420 90.090 ;
        RECT 1293.220 48.690 1293.360 89.770 ;
        RECT 1293.220 48.550 1293.820 48.690 ;
        RECT 1293.680 48.010 1293.820 48.550 ;
        RECT 1292.760 47.870 1293.820 48.010 ;
        RECT 1292.760 25.830 1292.900 47.870 ;
        RECT 1292.700 25.510 1292.960 25.830 ;
        RECT 1400.340 25.510 1400.600 25.830 ;
        RECT 1400.400 2.400 1400.540 25.510 ;
        RECT 1400.190 -4.800 1400.750 2.400 ;
      LAYER via2 ;
        RECT 1292.690 420.440 1292.970 420.720 ;
        RECT 1293.610 419.760 1293.890 420.040 ;
      LAYER met3 ;
        RECT 1292.665 420.730 1292.995 420.745 ;
        RECT 1291.990 420.430 1292.995 420.730 ;
        RECT 1291.990 420.050 1292.290 420.430 ;
        RECT 1292.665 420.415 1292.995 420.430 ;
        RECT 1293.585 420.050 1293.915 420.065 ;
        RECT 1291.990 419.750 1293.915 420.050 ;
        RECT 1293.585 419.735 1293.915 419.750 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1291.750 1684.260 1292.070 1684.320 ;
        RECT 1295.430 1684.260 1295.750 1684.320 ;
        RECT 1291.750 1684.120 1295.750 1684.260 ;
        RECT 1291.750 1684.060 1292.070 1684.120 ;
        RECT 1295.430 1684.060 1295.750 1684.120 ;
        RECT 1291.750 25.060 1292.070 25.120 ;
        RECT 1418.250 25.060 1418.570 25.120 ;
        RECT 1291.750 24.920 1418.570 25.060 ;
        RECT 1291.750 24.860 1292.070 24.920 ;
        RECT 1418.250 24.860 1418.570 24.920 ;
      LAYER via ;
        RECT 1291.780 1684.060 1292.040 1684.320 ;
        RECT 1295.460 1684.060 1295.720 1684.320 ;
        RECT 1291.780 24.860 1292.040 25.120 ;
        RECT 1418.280 24.860 1418.540 25.120 ;
      LAYER met2 ;
        RECT 1295.360 1700.340 1295.640 1704.000 ;
        RECT 1295.360 1700.000 1295.660 1700.340 ;
        RECT 1295.520 1684.350 1295.660 1700.000 ;
        RECT 1291.780 1684.030 1292.040 1684.350 ;
        RECT 1295.460 1684.030 1295.720 1684.350 ;
        RECT 1291.840 25.150 1291.980 1684.030 ;
        RECT 1291.780 24.830 1292.040 25.150 ;
        RECT 1418.280 24.830 1418.540 25.150 ;
        RECT 1418.340 2.400 1418.480 24.830 ;
        RECT 1418.130 -4.800 1418.690 2.400 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1301.025 1242.105 1301.195 1290.215 ;
        RECT 1301.485 1152.345 1301.655 1200.455 ;
        RECT 1301.025 959.225 1301.195 1007.335 ;
        RECT 1301.485 893.605 1301.655 917.575 ;
        RECT 1301.485 621.265 1301.655 669.375 ;
        RECT 1301.485 572.645 1301.655 620.755 ;
        RECT 1301.485 379.525 1301.655 432.735 ;
        RECT 1301.485 234.685 1301.655 241.995 ;
        RECT 1301.025 41.565 1301.195 89.335 ;
      LAYER mcon ;
        RECT 1301.025 1290.045 1301.195 1290.215 ;
        RECT 1301.485 1200.285 1301.655 1200.455 ;
        RECT 1301.025 1007.165 1301.195 1007.335 ;
        RECT 1301.485 917.405 1301.655 917.575 ;
        RECT 1301.485 669.205 1301.655 669.375 ;
        RECT 1301.485 620.585 1301.655 620.755 ;
        RECT 1301.485 432.565 1301.655 432.735 ;
        RECT 1301.485 241.825 1301.655 241.995 ;
        RECT 1301.025 89.165 1301.195 89.335 ;
      LAYER met1 ;
        RECT 1297.270 1670.320 1297.590 1670.380 ;
        RECT 1301.870 1670.320 1302.190 1670.380 ;
        RECT 1297.270 1670.180 1302.190 1670.320 ;
        RECT 1297.270 1670.120 1297.590 1670.180 ;
        RECT 1301.870 1670.120 1302.190 1670.180 ;
        RECT 1301.870 1538.740 1302.190 1538.800 ;
        RECT 1302.790 1538.740 1303.110 1538.800 ;
        RECT 1301.870 1538.600 1303.110 1538.740 ;
        RECT 1301.870 1538.540 1302.190 1538.600 ;
        RECT 1302.790 1538.540 1303.110 1538.600 ;
        RECT 1301.410 1401.040 1301.730 1401.100 ;
        RECT 1302.790 1401.040 1303.110 1401.100 ;
        RECT 1301.410 1400.900 1303.110 1401.040 ;
        RECT 1301.410 1400.840 1301.730 1400.900 ;
        RECT 1302.790 1400.840 1303.110 1400.900 ;
        RECT 1301.410 1376.560 1301.730 1376.620 ;
        RECT 1302.790 1376.560 1303.110 1376.620 ;
        RECT 1301.410 1376.420 1303.110 1376.560 ;
        RECT 1301.410 1376.360 1301.730 1376.420 ;
        RECT 1302.790 1376.360 1303.110 1376.420 ;
        RECT 1301.870 1297.340 1302.190 1297.400 ;
        RECT 1302.790 1297.340 1303.110 1297.400 ;
        RECT 1301.870 1297.200 1303.110 1297.340 ;
        RECT 1301.870 1297.140 1302.190 1297.200 ;
        RECT 1302.790 1297.140 1303.110 1297.200 ;
        RECT 1300.965 1290.200 1301.255 1290.245 ;
        RECT 1301.870 1290.200 1302.190 1290.260 ;
        RECT 1300.965 1290.060 1302.190 1290.200 ;
        RECT 1300.965 1290.015 1301.255 1290.060 ;
        RECT 1301.870 1290.000 1302.190 1290.060 ;
        RECT 1300.950 1242.260 1301.270 1242.320 ;
        RECT 1300.755 1242.120 1301.270 1242.260 ;
        RECT 1300.950 1242.060 1301.270 1242.120 ;
        RECT 1300.950 1200.440 1301.270 1200.500 ;
        RECT 1301.425 1200.440 1301.715 1200.485 ;
        RECT 1300.950 1200.300 1301.715 1200.440 ;
        RECT 1300.950 1200.240 1301.270 1200.300 ;
        RECT 1301.425 1200.255 1301.715 1200.300 ;
        RECT 1301.410 1152.500 1301.730 1152.560 ;
        RECT 1301.215 1152.360 1301.730 1152.500 ;
        RECT 1301.410 1152.300 1301.730 1152.360 ;
        RECT 1301.410 1111.500 1301.730 1111.760 ;
        RECT 1301.500 1111.080 1301.640 1111.500 ;
        RECT 1301.410 1110.820 1301.730 1111.080 ;
        RECT 1300.950 1014.460 1301.270 1014.520 ;
        RECT 1301.410 1014.460 1301.730 1014.520 ;
        RECT 1300.950 1014.320 1301.730 1014.460 ;
        RECT 1300.950 1014.260 1301.270 1014.320 ;
        RECT 1301.410 1014.260 1301.730 1014.320 ;
        RECT 1300.965 1007.320 1301.255 1007.365 ;
        RECT 1301.410 1007.320 1301.730 1007.380 ;
        RECT 1300.965 1007.180 1301.730 1007.320 ;
        RECT 1300.965 1007.135 1301.255 1007.180 ;
        RECT 1301.410 1007.120 1301.730 1007.180 ;
        RECT 1300.950 959.380 1301.270 959.440 ;
        RECT 1300.755 959.240 1301.270 959.380 ;
        RECT 1300.950 959.180 1301.270 959.240 ;
        RECT 1301.410 917.560 1301.730 917.620 ;
        RECT 1301.215 917.420 1301.730 917.560 ;
        RECT 1301.410 917.360 1301.730 917.420 ;
        RECT 1301.410 893.760 1301.730 893.820 ;
        RECT 1301.215 893.620 1301.730 893.760 ;
        RECT 1301.410 893.560 1301.730 893.620 ;
        RECT 1301.410 821.000 1301.730 821.060 ;
        RECT 1301.870 821.000 1302.190 821.060 ;
        RECT 1301.410 820.860 1302.190 821.000 ;
        RECT 1301.410 820.800 1301.730 820.860 ;
        RECT 1301.870 820.800 1302.190 820.860 ;
        RECT 1301.870 773.400 1302.190 773.460 ;
        RECT 1301.500 773.260 1302.190 773.400 ;
        RECT 1301.500 772.780 1301.640 773.260 ;
        RECT 1301.870 773.200 1302.190 773.260 ;
        RECT 1301.410 772.520 1301.730 772.780 ;
        RECT 1301.410 724.440 1301.730 724.500 ;
        RECT 1301.870 724.440 1302.190 724.500 ;
        RECT 1301.410 724.300 1302.190 724.440 ;
        RECT 1301.410 724.240 1301.730 724.300 ;
        RECT 1301.870 724.240 1302.190 724.300 ;
        RECT 1300.490 693.500 1300.810 693.560 ;
        RECT 1301.870 693.500 1302.190 693.560 ;
        RECT 1300.490 693.360 1302.190 693.500 ;
        RECT 1300.490 693.300 1300.810 693.360 ;
        RECT 1301.870 693.300 1302.190 693.360 ;
        RECT 1301.410 669.360 1301.730 669.420 ;
        RECT 1301.215 669.220 1301.730 669.360 ;
        RECT 1301.410 669.160 1301.730 669.220 ;
        RECT 1301.410 621.420 1301.730 621.480 ;
        RECT 1301.215 621.280 1301.730 621.420 ;
        RECT 1301.410 621.220 1301.730 621.280 ;
        RECT 1301.410 620.740 1301.730 620.800 ;
        RECT 1301.215 620.600 1301.730 620.740 ;
        RECT 1301.410 620.540 1301.730 620.600 ;
        RECT 1301.425 572.800 1301.715 572.845 ;
        RECT 1301.870 572.800 1302.190 572.860 ;
        RECT 1301.425 572.660 1302.190 572.800 ;
        RECT 1301.425 572.615 1301.715 572.660 ;
        RECT 1301.870 572.600 1302.190 572.660 ;
        RECT 1301.410 496.780 1301.730 497.040 ;
        RECT 1301.500 496.640 1301.640 496.780 ;
        RECT 1301.870 496.640 1302.190 496.700 ;
        RECT 1301.500 496.500 1302.190 496.640 ;
        RECT 1301.870 496.440 1302.190 496.500 ;
        RECT 1301.425 432.720 1301.715 432.765 ;
        RECT 1301.870 432.720 1302.190 432.780 ;
        RECT 1301.425 432.580 1302.190 432.720 ;
        RECT 1301.425 432.535 1301.715 432.580 ;
        RECT 1301.870 432.520 1302.190 432.580 ;
        RECT 1301.425 379.680 1301.715 379.725 ;
        RECT 1301.870 379.680 1302.190 379.740 ;
        RECT 1301.425 379.540 1302.190 379.680 ;
        RECT 1301.425 379.495 1301.715 379.540 ;
        RECT 1301.870 379.480 1302.190 379.540 ;
        RECT 1301.410 289.920 1301.730 289.980 ;
        RECT 1301.870 289.920 1302.190 289.980 ;
        RECT 1301.410 289.780 1302.190 289.920 ;
        RECT 1301.410 289.720 1301.730 289.780 ;
        RECT 1301.870 289.720 1302.190 289.780 ;
        RECT 1301.425 241.980 1301.715 242.025 ;
        RECT 1301.870 241.980 1302.190 242.040 ;
        RECT 1301.425 241.840 1302.190 241.980 ;
        RECT 1301.425 241.795 1301.715 241.840 ;
        RECT 1301.870 241.780 1302.190 241.840 ;
        RECT 1301.410 234.840 1301.730 234.900 ;
        RECT 1301.215 234.700 1301.730 234.840 ;
        RECT 1301.410 234.640 1301.730 234.700 ;
        RECT 1300.490 96.800 1300.810 96.860 ;
        RECT 1301.410 96.800 1301.730 96.860 ;
        RECT 1300.490 96.660 1301.730 96.800 ;
        RECT 1300.490 96.600 1300.810 96.660 ;
        RECT 1301.410 96.600 1301.730 96.660 ;
        RECT 1300.965 89.320 1301.255 89.365 ;
        RECT 1301.870 89.320 1302.190 89.380 ;
        RECT 1300.965 89.180 1302.190 89.320 ;
        RECT 1300.965 89.135 1301.255 89.180 ;
        RECT 1301.870 89.120 1302.190 89.180 ;
        RECT 1300.950 41.720 1301.270 41.780 ;
        RECT 1300.755 41.580 1301.270 41.720 ;
        RECT 1300.950 41.520 1301.270 41.580 ;
        RECT 1300.950 24.380 1301.270 24.440 ;
        RECT 1435.730 24.380 1436.050 24.440 ;
        RECT 1300.950 24.240 1436.050 24.380 ;
        RECT 1300.950 24.180 1301.270 24.240 ;
        RECT 1435.730 24.180 1436.050 24.240 ;
      LAYER via ;
        RECT 1297.300 1670.120 1297.560 1670.380 ;
        RECT 1301.900 1670.120 1302.160 1670.380 ;
        RECT 1301.900 1538.540 1302.160 1538.800 ;
        RECT 1302.820 1538.540 1303.080 1538.800 ;
        RECT 1301.440 1400.840 1301.700 1401.100 ;
        RECT 1302.820 1400.840 1303.080 1401.100 ;
        RECT 1301.440 1376.360 1301.700 1376.620 ;
        RECT 1302.820 1376.360 1303.080 1376.620 ;
        RECT 1301.900 1297.140 1302.160 1297.400 ;
        RECT 1302.820 1297.140 1303.080 1297.400 ;
        RECT 1301.900 1290.000 1302.160 1290.260 ;
        RECT 1300.980 1242.060 1301.240 1242.320 ;
        RECT 1300.980 1200.240 1301.240 1200.500 ;
        RECT 1301.440 1152.300 1301.700 1152.560 ;
        RECT 1301.440 1111.500 1301.700 1111.760 ;
        RECT 1301.440 1110.820 1301.700 1111.080 ;
        RECT 1300.980 1014.260 1301.240 1014.520 ;
        RECT 1301.440 1014.260 1301.700 1014.520 ;
        RECT 1301.440 1007.120 1301.700 1007.380 ;
        RECT 1300.980 959.180 1301.240 959.440 ;
        RECT 1301.440 917.360 1301.700 917.620 ;
        RECT 1301.440 893.560 1301.700 893.820 ;
        RECT 1301.440 820.800 1301.700 821.060 ;
        RECT 1301.900 820.800 1302.160 821.060 ;
        RECT 1301.900 773.200 1302.160 773.460 ;
        RECT 1301.440 772.520 1301.700 772.780 ;
        RECT 1301.440 724.240 1301.700 724.500 ;
        RECT 1301.900 724.240 1302.160 724.500 ;
        RECT 1300.520 693.300 1300.780 693.560 ;
        RECT 1301.900 693.300 1302.160 693.560 ;
        RECT 1301.440 669.160 1301.700 669.420 ;
        RECT 1301.440 621.220 1301.700 621.480 ;
        RECT 1301.440 620.540 1301.700 620.800 ;
        RECT 1301.900 572.600 1302.160 572.860 ;
        RECT 1301.440 496.780 1301.700 497.040 ;
        RECT 1301.900 496.440 1302.160 496.700 ;
        RECT 1301.900 432.520 1302.160 432.780 ;
        RECT 1301.900 379.480 1302.160 379.740 ;
        RECT 1301.440 289.720 1301.700 289.980 ;
        RECT 1301.900 289.720 1302.160 289.980 ;
        RECT 1301.900 241.780 1302.160 242.040 ;
        RECT 1301.440 234.640 1301.700 234.900 ;
        RECT 1300.520 96.600 1300.780 96.860 ;
        RECT 1301.440 96.600 1301.700 96.860 ;
        RECT 1301.900 89.120 1302.160 89.380 ;
        RECT 1300.980 41.520 1301.240 41.780 ;
        RECT 1300.980 24.180 1301.240 24.440 ;
        RECT 1435.760 24.180 1436.020 24.440 ;
      LAYER met2 ;
        RECT 1297.200 1700.340 1297.480 1704.000 ;
        RECT 1297.200 1700.000 1297.500 1700.340 ;
        RECT 1297.360 1670.410 1297.500 1700.000 ;
        RECT 1297.300 1670.090 1297.560 1670.410 ;
        RECT 1301.900 1670.090 1302.160 1670.410 ;
        RECT 1301.960 1538.830 1302.100 1670.090 ;
        RECT 1301.900 1538.510 1302.160 1538.830 ;
        RECT 1302.820 1538.510 1303.080 1538.830 ;
        RECT 1302.880 1401.130 1303.020 1538.510 ;
        RECT 1301.440 1400.810 1301.700 1401.130 ;
        RECT 1302.820 1400.810 1303.080 1401.130 ;
        RECT 1301.500 1376.650 1301.640 1400.810 ;
        RECT 1301.440 1376.330 1301.700 1376.650 ;
        RECT 1302.820 1376.330 1303.080 1376.650 ;
        RECT 1302.880 1297.430 1303.020 1376.330 ;
        RECT 1301.900 1297.110 1302.160 1297.430 ;
        RECT 1302.820 1297.110 1303.080 1297.430 ;
        RECT 1301.960 1290.290 1302.100 1297.110 ;
        RECT 1301.900 1289.970 1302.160 1290.290 ;
        RECT 1300.980 1242.030 1301.240 1242.350 ;
        RECT 1301.040 1200.530 1301.180 1242.030 ;
        RECT 1300.980 1200.210 1301.240 1200.530 ;
        RECT 1301.440 1152.270 1301.700 1152.590 ;
        RECT 1301.500 1111.790 1301.640 1152.270 ;
        RECT 1301.440 1111.470 1301.700 1111.790 ;
        RECT 1301.440 1110.790 1301.700 1111.110 ;
        RECT 1301.500 1104.165 1301.640 1110.790 ;
        RECT 1301.430 1103.795 1301.710 1104.165 ;
        RECT 1302.810 1103.795 1303.090 1104.165 ;
        RECT 1302.880 1055.885 1303.020 1103.795 ;
        RECT 1300.970 1055.515 1301.250 1055.885 ;
        RECT 1302.810 1055.515 1303.090 1055.885 ;
        RECT 1301.040 1014.550 1301.180 1055.515 ;
        RECT 1300.980 1014.230 1301.240 1014.550 ;
        RECT 1301.440 1014.230 1301.700 1014.550 ;
        RECT 1301.500 1007.410 1301.640 1014.230 ;
        RECT 1301.440 1007.090 1301.700 1007.410 ;
        RECT 1300.980 959.150 1301.240 959.470 ;
        RECT 1301.040 942.210 1301.180 959.150 ;
        RECT 1301.040 942.070 1301.640 942.210 ;
        RECT 1301.500 917.650 1301.640 942.070 ;
        RECT 1301.440 917.330 1301.700 917.650 ;
        RECT 1301.440 893.530 1301.700 893.850 ;
        RECT 1301.500 821.090 1301.640 893.530 ;
        RECT 1301.440 820.770 1301.700 821.090 ;
        RECT 1301.900 820.770 1302.160 821.090 ;
        RECT 1301.960 773.490 1302.100 820.770 ;
        RECT 1301.900 773.170 1302.160 773.490 ;
        RECT 1301.440 772.490 1301.700 772.810 ;
        RECT 1301.500 724.530 1301.640 772.490 ;
        RECT 1301.440 724.210 1301.700 724.530 ;
        RECT 1301.900 724.210 1302.160 724.530 ;
        RECT 1301.960 693.590 1302.100 724.210 ;
        RECT 1300.520 693.270 1300.780 693.590 ;
        RECT 1301.900 693.270 1302.160 693.590 ;
        RECT 1300.580 670.325 1300.720 693.270 ;
        RECT 1300.510 669.955 1300.790 670.325 ;
        RECT 1301.430 669.275 1301.710 669.645 ;
        RECT 1301.440 669.130 1301.700 669.275 ;
        RECT 1301.440 621.190 1301.700 621.510 ;
        RECT 1301.500 620.830 1301.640 621.190 ;
        RECT 1301.440 620.510 1301.700 620.830 ;
        RECT 1301.900 572.570 1302.160 572.890 ;
        RECT 1301.960 524.690 1302.100 572.570 ;
        RECT 1301.500 524.550 1302.100 524.690 ;
        RECT 1301.500 497.070 1301.640 524.550 ;
        RECT 1301.440 496.750 1301.700 497.070 ;
        RECT 1301.900 496.410 1302.160 496.730 ;
        RECT 1301.960 432.810 1302.100 496.410 ;
        RECT 1301.900 432.490 1302.160 432.810 ;
        RECT 1301.900 379.450 1302.160 379.770 ;
        RECT 1301.960 362.170 1302.100 379.450 ;
        RECT 1301.040 362.030 1302.100 362.170 ;
        RECT 1301.040 337.690 1301.180 362.030 ;
        RECT 1301.040 337.550 1301.640 337.690 ;
        RECT 1301.500 290.010 1301.640 337.550 ;
        RECT 1301.440 289.690 1301.700 290.010 ;
        RECT 1301.900 289.690 1302.160 290.010 ;
        RECT 1301.960 242.070 1302.100 289.690 ;
        RECT 1301.900 241.750 1302.160 242.070 ;
        RECT 1301.440 234.610 1301.700 234.930 ;
        RECT 1301.500 96.890 1301.640 234.610 ;
        RECT 1300.520 96.570 1300.780 96.890 ;
        RECT 1301.440 96.570 1301.700 96.890 ;
        RECT 1300.580 90.285 1300.720 96.570 ;
        RECT 1300.510 89.915 1300.790 90.285 ;
        RECT 1301.890 89.915 1302.170 90.285 ;
        RECT 1301.960 89.410 1302.100 89.915 ;
        RECT 1301.900 89.090 1302.160 89.410 ;
        RECT 1300.980 41.490 1301.240 41.810 ;
        RECT 1301.040 24.470 1301.180 41.490 ;
        RECT 1300.980 24.150 1301.240 24.470 ;
        RECT 1435.760 24.150 1436.020 24.470 ;
        RECT 1435.820 2.400 1435.960 24.150 ;
        RECT 1435.610 -4.800 1436.170 2.400 ;
      LAYER via2 ;
        RECT 1301.430 1103.840 1301.710 1104.120 ;
        RECT 1302.810 1103.840 1303.090 1104.120 ;
        RECT 1300.970 1055.560 1301.250 1055.840 ;
        RECT 1302.810 1055.560 1303.090 1055.840 ;
        RECT 1300.510 670.000 1300.790 670.280 ;
        RECT 1301.430 669.320 1301.710 669.600 ;
        RECT 1300.510 89.960 1300.790 90.240 ;
        RECT 1301.890 89.960 1302.170 90.240 ;
      LAYER met3 ;
        RECT 1301.405 1104.130 1301.735 1104.145 ;
        RECT 1302.785 1104.130 1303.115 1104.145 ;
        RECT 1301.405 1103.830 1303.115 1104.130 ;
        RECT 1301.405 1103.815 1301.735 1103.830 ;
        RECT 1302.785 1103.815 1303.115 1103.830 ;
        RECT 1300.945 1055.850 1301.275 1055.865 ;
        RECT 1302.785 1055.850 1303.115 1055.865 ;
        RECT 1300.945 1055.550 1303.115 1055.850 ;
        RECT 1300.945 1055.535 1301.275 1055.550 ;
        RECT 1302.785 1055.535 1303.115 1055.550 ;
        RECT 1300.485 670.290 1300.815 670.305 ;
        RECT 1300.485 669.990 1301.490 670.290 ;
        RECT 1300.485 669.975 1300.815 669.990 ;
        RECT 1301.190 669.625 1301.490 669.990 ;
        RECT 1301.190 669.310 1301.735 669.625 ;
        RECT 1301.405 669.295 1301.735 669.310 ;
        RECT 1300.485 90.250 1300.815 90.265 ;
        RECT 1301.865 90.250 1302.195 90.265 ;
        RECT 1300.485 89.950 1302.195 90.250 ;
        RECT 1300.485 89.935 1300.815 89.950 ;
        RECT 1301.865 89.935 1302.195 89.950 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1301.025 1496.765 1301.195 1538.755 ;
        RECT 1299.645 1338.665 1299.815 1393.575 ;
        RECT 1300.565 1248.565 1300.735 1290.215 ;
        RECT 1301.025 766.445 1301.195 814.215 ;
        RECT 1300.565 572.645 1300.735 620.755 ;
        RECT 1300.565 462.485 1300.735 510.595 ;
        RECT 1300.565 234.685 1300.735 241.995 ;
        RECT 1299.645 89.845 1299.815 97.495 ;
      LAYER mcon ;
        RECT 1301.025 1538.585 1301.195 1538.755 ;
        RECT 1299.645 1393.405 1299.815 1393.575 ;
        RECT 1300.565 1290.045 1300.735 1290.215 ;
        RECT 1301.025 814.045 1301.195 814.215 ;
        RECT 1300.565 620.585 1300.735 620.755 ;
        RECT 1300.565 510.425 1300.735 510.595 ;
        RECT 1300.565 241.825 1300.735 241.995 ;
        RECT 1299.645 97.325 1299.815 97.495 ;
      LAYER met1 ;
        RECT 1299.570 1674.060 1299.890 1674.120 ;
        RECT 1300.950 1674.060 1301.270 1674.120 ;
        RECT 1299.570 1673.920 1301.270 1674.060 ;
        RECT 1299.570 1673.860 1299.890 1673.920 ;
        RECT 1300.950 1673.860 1301.270 1673.920 ;
        RECT 1300.950 1538.740 1301.270 1538.800 ;
        RECT 1300.755 1538.600 1301.270 1538.740 ;
        RECT 1300.950 1538.540 1301.270 1538.600 ;
        RECT 1300.965 1496.920 1301.255 1496.965 ;
        RECT 1301.410 1496.920 1301.730 1496.980 ;
        RECT 1300.965 1496.780 1301.730 1496.920 ;
        RECT 1300.965 1496.735 1301.255 1496.780 ;
        RECT 1301.410 1496.720 1301.730 1496.780 ;
        RECT 1300.490 1409.880 1300.810 1409.940 ;
        RECT 1301.410 1409.880 1301.730 1409.940 ;
        RECT 1300.490 1409.740 1301.730 1409.880 ;
        RECT 1300.490 1409.680 1300.810 1409.740 ;
        RECT 1301.410 1409.680 1301.730 1409.740 ;
        RECT 1299.570 1400.700 1299.890 1400.760 ;
        RECT 1300.490 1400.700 1300.810 1400.760 ;
        RECT 1299.570 1400.560 1300.810 1400.700 ;
        RECT 1299.570 1400.500 1299.890 1400.560 ;
        RECT 1300.490 1400.500 1300.810 1400.560 ;
        RECT 1299.570 1393.560 1299.890 1393.620 ;
        RECT 1299.375 1393.420 1299.890 1393.560 ;
        RECT 1299.570 1393.360 1299.890 1393.420 ;
        RECT 1299.585 1338.820 1299.875 1338.865 ;
        RECT 1300.490 1338.820 1300.810 1338.880 ;
        RECT 1299.585 1338.680 1300.810 1338.820 ;
        RECT 1299.585 1338.635 1299.875 1338.680 ;
        RECT 1300.490 1338.620 1300.810 1338.680 ;
        RECT 1300.490 1290.200 1300.810 1290.260 ;
        RECT 1300.295 1290.060 1300.810 1290.200 ;
        RECT 1300.490 1290.000 1300.810 1290.060 ;
        RECT 1300.490 1248.720 1300.810 1248.780 ;
        RECT 1300.295 1248.580 1300.810 1248.720 ;
        RECT 1300.490 1248.520 1300.810 1248.580 ;
        RECT 1299.570 1224.920 1299.890 1224.980 ;
        RECT 1300.490 1224.920 1300.810 1224.980 ;
        RECT 1299.570 1224.780 1300.810 1224.920 ;
        RECT 1299.570 1224.720 1299.890 1224.780 ;
        RECT 1300.490 1224.720 1300.810 1224.780 ;
        RECT 1299.570 1176.640 1299.890 1176.700 ;
        RECT 1300.950 1176.640 1301.270 1176.700 ;
        RECT 1299.570 1176.500 1301.270 1176.640 ;
        RECT 1299.570 1176.440 1299.890 1176.500 ;
        RECT 1300.950 1176.440 1301.270 1176.500 ;
        RECT 1300.490 1111.020 1300.810 1111.080 ;
        RECT 1300.950 1111.020 1301.270 1111.080 ;
        RECT 1300.490 1110.880 1301.270 1111.020 ;
        RECT 1300.490 1110.820 1300.810 1110.880 ;
        RECT 1300.950 1110.820 1301.270 1110.880 ;
        RECT 1299.570 1014.460 1299.890 1014.520 ;
        RECT 1300.490 1014.460 1300.810 1014.520 ;
        RECT 1299.570 1014.320 1300.810 1014.460 ;
        RECT 1299.570 1014.260 1299.890 1014.320 ;
        RECT 1300.490 1014.260 1300.810 1014.320 ;
        RECT 1298.650 1007.320 1298.970 1007.380 ;
        RECT 1300.490 1007.320 1300.810 1007.380 ;
        RECT 1298.650 1007.180 1300.810 1007.320 ;
        RECT 1298.650 1007.120 1298.970 1007.180 ;
        RECT 1300.490 1007.120 1300.810 1007.180 ;
        RECT 1299.570 931.500 1299.890 931.560 ;
        RECT 1300.490 931.500 1300.810 931.560 ;
        RECT 1299.570 931.360 1300.810 931.500 ;
        RECT 1299.570 931.300 1299.890 931.360 ;
        RECT 1300.490 931.300 1300.810 931.360 ;
        RECT 1299.570 893.760 1299.890 893.820 ;
        RECT 1300.490 893.760 1300.810 893.820 ;
        RECT 1299.570 893.620 1300.810 893.760 ;
        RECT 1299.570 893.560 1299.890 893.620 ;
        RECT 1300.490 893.560 1300.810 893.620 ;
        RECT 1300.490 821.000 1300.810 821.060 ;
        RECT 1300.950 821.000 1301.270 821.060 ;
        RECT 1300.490 820.860 1301.270 821.000 ;
        RECT 1300.490 820.800 1300.810 820.860 ;
        RECT 1300.950 820.800 1301.270 820.860 ;
        RECT 1300.950 814.200 1301.270 814.260 ;
        RECT 1300.755 814.060 1301.270 814.200 ;
        RECT 1300.950 814.000 1301.270 814.060 ;
        RECT 1300.950 766.600 1301.270 766.660 ;
        RECT 1300.755 766.460 1301.270 766.600 ;
        RECT 1300.950 766.400 1301.270 766.460 ;
        RECT 1300.490 724.440 1300.810 724.500 ;
        RECT 1300.950 724.440 1301.270 724.500 ;
        RECT 1300.490 724.300 1301.270 724.440 ;
        RECT 1300.490 724.240 1300.810 724.300 ;
        RECT 1300.950 724.240 1301.270 724.300 ;
        RECT 1300.490 628.220 1300.810 628.280 ;
        RECT 1300.950 628.220 1301.270 628.280 ;
        RECT 1300.490 628.080 1301.270 628.220 ;
        RECT 1300.490 628.020 1300.810 628.080 ;
        RECT 1300.950 628.020 1301.270 628.080 ;
        RECT 1300.490 620.740 1300.810 620.800 ;
        RECT 1300.295 620.600 1300.810 620.740 ;
        RECT 1300.490 620.540 1300.810 620.600 ;
        RECT 1300.505 572.800 1300.795 572.845 ;
        RECT 1300.950 572.800 1301.270 572.860 ;
        RECT 1300.505 572.660 1301.270 572.800 ;
        RECT 1300.505 572.615 1300.795 572.660 ;
        RECT 1300.950 572.600 1301.270 572.660 ;
        RECT 1300.490 510.580 1300.810 510.640 ;
        RECT 1300.295 510.440 1300.810 510.580 ;
        RECT 1300.490 510.380 1300.810 510.440 ;
        RECT 1300.505 462.640 1300.795 462.685 ;
        RECT 1300.950 462.640 1301.270 462.700 ;
        RECT 1300.505 462.500 1301.270 462.640 ;
        RECT 1300.505 462.455 1300.795 462.500 ;
        RECT 1300.950 462.440 1301.270 462.500 ;
        RECT 1300.490 337.660 1300.810 337.920 ;
        RECT 1300.580 337.180 1300.720 337.660 ;
        RECT 1300.950 337.180 1301.270 337.240 ;
        RECT 1300.580 337.040 1301.270 337.180 ;
        RECT 1300.950 336.980 1301.270 337.040 ;
        RECT 1300.505 241.980 1300.795 242.025 ;
        RECT 1300.950 241.980 1301.270 242.040 ;
        RECT 1300.505 241.840 1301.270 241.980 ;
        RECT 1300.505 241.795 1300.795 241.840 ;
        RECT 1300.950 241.780 1301.270 241.840 ;
        RECT 1300.490 234.840 1300.810 234.900 ;
        RECT 1300.295 234.700 1300.810 234.840 ;
        RECT 1300.490 234.640 1300.810 234.700 ;
        RECT 1299.585 97.480 1299.875 97.525 ;
        RECT 1300.490 97.480 1300.810 97.540 ;
        RECT 1299.585 97.340 1300.810 97.480 ;
        RECT 1299.585 97.295 1299.875 97.340 ;
        RECT 1300.490 97.280 1300.810 97.340 ;
        RECT 1299.570 90.000 1299.890 90.060 ;
        RECT 1299.375 89.860 1299.890 90.000 ;
        RECT 1299.570 89.800 1299.890 89.860 ;
        RECT 1299.570 89.320 1299.890 89.380 ;
        RECT 1300.490 89.320 1300.810 89.380 ;
        RECT 1299.570 89.180 1300.810 89.320 ;
        RECT 1299.570 89.120 1299.890 89.180 ;
        RECT 1300.490 89.120 1300.810 89.180 ;
        RECT 1300.490 24.040 1300.810 24.100 ;
        RECT 1453.670 24.040 1453.990 24.100 ;
        RECT 1300.490 23.900 1453.990 24.040 ;
        RECT 1300.490 23.840 1300.810 23.900 ;
        RECT 1453.670 23.840 1453.990 23.900 ;
      LAYER via ;
        RECT 1299.600 1673.860 1299.860 1674.120 ;
        RECT 1300.980 1673.860 1301.240 1674.120 ;
        RECT 1300.980 1538.540 1301.240 1538.800 ;
        RECT 1301.440 1496.720 1301.700 1496.980 ;
        RECT 1300.520 1409.680 1300.780 1409.940 ;
        RECT 1301.440 1409.680 1301.700 1409.940 ;
        RECT 1299.600 1400.500 1299.860 1400.760 ;
        RECT 1300.520 1400.500 1300.780 1400.760 ;
        RECT 1299.600 1393.360 1299.860 1393.620 ;
        RECT 1300.520 1338.620 1300.780 1338.880 ;
        RECT 1300.520 1290.000 1300.780 1290.260 ;
        RECT 1300.520 1248.520 1300.780 1248.780 ;
        RECT 1299.600 1224.720 1299.860 1224.980 ;
        RECT 1300.520 1224.720 1300.780 1224.980 ;
        RECT 1299.600 1176.440 1299.860 1176.700 ;
        RECT 1300.980 1176.440 1301.240 1176.700 ;
        RECT 1300.520 1110.820 1300.780 1111.080 ;
        RECT 1300.980 1110.820 1301.240 1111.080 ;
        RECT 1299.600 1014.260 1299.860 1014.520 ;
        RECT 1300.520 1014.260 1300.780 1014.520 ;
        RECT 1298.680 1007.120 1298.940 1007.380 ;
        RECT 1300.520 1007.120 1300.780 1007.380 ;
        RECT 1299.600 931.300 1299.860 931.560 ;
        RECT 1300.520 931.300 1300.780 931.560 ;
        RECT 1299.600 893.560 1299.860 893.820 ;
        RECT 1300.520 893.560 1300.780 893.820 ;
        RECT 1300.520 820.800 1300.780 821.060 ;
        RECT 1300.980 820.800 1301.240 821.060 ;
        RECT 1300.980 814.000 1301.240 814.260 ;
        RECT 1300.980 766.400 1301.240 766.660 ;
        RECT 1300.520 724.240 1300.780 724.500 ;
        RECT 1300.980 724.240 1301.240 724.500 ;
        RECT 1300.520 628.020 1300.780 628.280 ;
        RECT 1300.980 628.020 1301.240 628.280 ;
        RECT 1300.520 620.540 1300.780 620.800 ;
        RECT 1300.980 572.600 1301.240 572.860 ;
        RECT 1300.520 510.380 1300.780 510.640 ;
        RECT 1300.980 462.440 1301.240 462.700 ;
        RECT 1300.520 337.660 1300.780 337.920 ;
        RECT 1300.980 336.980 1301.240 337.240 ;
        RECT 1300.980 241.780 1301.240 242.040 ;
        RECT 1300.520 234.640 1300.780 234.900 ;
        RECT 1300.520 97.280 1300.780 97.540 ;
        RECT 1299.600 89.800 1299.860 90.060 ;
        RECT 1299.600 89.120 1299.860 89.380 ;
        RECT 1300.520 89.120 1300.780 89.380 ;
        RECT 1300.520 23.840 1300.780 24.100 ;
        RECT 1453.700 23.840 1453.960 24.100 ;
      LAYER met2 ;
        RECT 1299.040 1700.410 1299.320 1704.000 ;
        RECT 1299.040 1700.270 1299.800 1700.410 ;
        RECT 1299.040 1700.000 1299.320 1700.270 ;
        RECT 1299.660 1674.150 1299.800 1700.270 ;
        RECT 1299.600 1673.830 1299.860 1674.150 ;
        RECT 1300.980 1673.830 1301.240 1674.150 ;
        RECT 1301.040 1538.830 1301.180 1673.830 ;
        RECT 1300.980 1538.510 1301.240 1538.830 ;
        RECT 1301.440 1496.690 1301.700 1497.010 ;
        RECT 1301.500 1409.970 1301.640 1496.690 ;
        RECT 1300.520 1409.650 1300.780 1409.970 ;
        RECT 1301.440 1409.650 1301.700 1409.970 ;
        RECT 1300.580 1400.790 1300.720 1409.650 ;
        RECT 1299.600 1400.470 1299.860 1400.790 ;
        RECT 1300.520 1400.470 1300.780 1400.790 ;
        RECT 1299.660 1393.650 1299.800 1400.470 ;
        RECT 1299.600 1393.330 1299.860 1393.650 ;
        RECT 1300.520 1338.590 1300.780 1338.910 ;
        RECT 1300.580 1290.290 1300.720 1338.590 ;
        RECT 1300.520 1289.970 1300.780 1290.290 ;
        RECT 1300.520 1248.490 1300.780 1248.810 ;
        RECT 1300.580 1225.010 1300.720 1248.490 ;
        RECT 1299.600 1224.690 1299.860 1225.010 ;
        RECT 1300.520 1224.690 1300.780 1225.010 ;
        RECT 1299.660 1176.730 1299.800 1224.690 ;
        RECT 1299.600 1176.410 1299.860 1176.730 ;
        RECT 1300.980 1176.410 1301.240 1176.730 ;
        RECT 1301.040 1111.110 1301.180 1176.410 ;
        RECT 1300.520 1110.790 1300.780 1111.110 ;
        RECT 1300.980 1110.790 1301.240 1111.110 ;
        RECT 1300.580 1104.165 1300.720 1110.790 ;
        RECT 1298.670 1103.795 1298.950 1104.165 ;
        RECT 1300.510 1103.795 1300.790 1104.165 ;
        RECT 1298.740 1055.885 1298.880 1103.795 ;
        RECT 1298.670 1055.515 1298.950 1055.885 ;
        RECT 1299.590 1055.515 1299.870 1055.885 ;
        RECT 1299.660 1014.550 1299.800 1055.515 ;
        RECT 1299.600 1014.230 1299.860 1014.550 ;
        RECT 1300.520 1014.230 1300.780 1014.550 ;
        RECT 1300.580 1007.410 1300.720 1014.230 ;
        RECT 1298.680 1007.090 1298.940 1007.410 ;
        RECT 1300.520 1007.090 1300.780 1007.410 ;
        RECT 1298.740 959.325 1298.880 1007.090 ;
        RECT 1298.670 958.955 1298.950 959.325 ;
        RECT 1299.590 958.955 1299.870 959.325 ;
        RECT 1299.660 931.590 1299.800 958.955 ;
        RECT 1299.600 931.270 1299.860 931.590 ;
        RECT 1300.520 931.270 1300.780 931.590 ;
        RECT 1300.580 917.845 1300.720 931.270 ;
        RECT 1299.590 917.475 1299.870 917.845 ;
        RECT 1300.510 917.475 1300.790 917.845 ;
        RECT 1299.660 893.850 1299.800 917.475 ;
        RECT 1299.600 893.530 1299.860 893.850 ;
        RECT 1300.520 893.530 1300.780 893.850 ;
        RECT 1300.580 821.090 1300.720 893.530 ;
        RECT 1300.520 820.770 1300.780 821.090 ;
        RECT 1300.980 820.770 1301.240 821.090 ;
        RECT 1301.040 814.290 1301.180 820.770 ;
        RECT 1300.980 813.970 1301.240 814.290 ;
        RECT 1300.980 766.370 1301.240 766.690 ;
        RECT 1301.040 725.405 1301.180 766.370 ;
        RECT 1300.970 725.035 1301.250 725.405 ;
        RECT 1300.510 724.355 1300.790 724.725 ;
        RECT 1300.520 724.210 1300.780 724.355 ;
        RECT 1300.980 724.210 1301.240 724.530 ;
        RECT 1301.040 628.310 1301.180 724.210 ;
        RECT 1300.520 627.990 1300.780 628.310 ;
        RECT 1300.980 627.990 1301.240 628.310 ;
        RECT 1300.580 620.830 1300.720 627.990 ;
        RECT 1300.520 620.510 1300.780 620.830 ;
        RECT 1300.980 572.570 1301.240 572.890 ;
        RECT 1301.040 524.690 1301.180 572.570 ;
        RECT 1300.580 524.550 1301.180 524.690 ;
        RECT 1300.580 510.670 1300.720 524.550 ;
        RECT 1300.520 510.350 1300.780 510.670 ;
        RECT 1300.980 462.410 1301.240 462.730 ;
        RECT 1301.040 362.850 1301.180 462.410 ;
        RECT 1300.580 362.710 1301.180 362.850 ;
        RECT 1300.580 337.950 1300.720 362.710 ;
        RECT 1300.520 337.630 1300.780 337.950 ;
        RECT 1300.980 336.950 1301.240 337.270 ;
        RECT 1301.040 242.070 1301.180 336.950 ;
        RECT 1300.980 241.750 1301.240 242.070 ;
        RECT 1300.520 234.610 1300.780 234.930 ;
        RECT 1300.580 97.570 1300.720 234.610 ;
        RECT 1300.520 97.250 1300.780 97.570 ;
        RECT 1299.600 89.770 1299.860 90.090 ;
        RECT 1299.660 89.410 1299.800 89.770 ;
        RECT 1299.600 89.090 1299.860 89.410 ;
        RECT 1300.520 89.090 1300.780 89.410 ;
        RECT 1300.580 24.130 1300.720 89.090 ;
        RECT 1300.520 23.810 1300.780 24.130 ;
        RECT 1453.700 23.810 1453.960 24.130 ;
        RECT 1453.760 2.400 1453.900 23.810 ;
        RECT 1453.550 -4.800 1454.110 2.400 ;
      LAYER via2 ;
        RECT 1298.670 1103.840 1298.950 1104.120 ;
        RECT 1300.510 1103.840 1300.790 1104.120 ;
        RECT 1298.670 1055.560 1298.950 1055.840 ;
        RECT 1299.590 1055.560 1299.870 1055.840 ;
        RECT 1298.670 959.000 1298.950 959.280 ;
        RECT 1299.590 959.000 1299.870 959.280 ;
        RECT 1299.590 917.520 1299.870 917.800 ;
        RECT 1300.510 917.520 1300.790 917.800 ;
        RECT 1300.970 725.080 1301.250 725.360 ;
        RECT 1300.510 724.400 1300.790 724.680 ;
      LAYER met3 ;
        RECT 1298.645 1104.130 1298.975 1104.145 ;
        RECT 1300.485 1104.130 1300.815 1104.145 ;
        RECT 1298.645 1103.830 1300.815 1104.130 ;
        RECT 1298.645 1103.815 1298.975 1103.830 ;
        RECT 1300.485 1103.815 1300.815 1103.830 ;
        RECT 1298.645 1055.850 1298.975 1055.865 ;
        RECT 1299.565 1055.850 1299.895 1055.865 ;
        RECT 1298.645 1055.550 1299.895 1055.850 ;
        RECT 1298.645 1055.535 1298.975 1055.550 ;
        RECT 1299.565 1055.535 1299.895 1055.550 ;
        RECT 1298.645 959.290 1298.975 959.305 ;
        RECT 1299.565 959.290 1299.895 959.305 ;
        RECT 1298.645 958.990 1299.895 959.290 ;
        RECT 1298.645 958.975 1298.975 958.990 ;
        RECT 1299.565 958.975 1299.895 958.990 ;
        RECT 1299.565 917.810 1299.895 917.825 ;
        RECT 1300.485 917.810 1300.815 917.825 ;
        RECT 1299.565 917.510 1300.815 917.810 ;
        RECT 1299.565 917.495 1299.895 917.510 ;
        RECT 1300.485 917.495 1300.815 917.510 ;
        RECT 1300.945 725.370 1301.275 725.385 ;
        RECT 1300.270 725.070 1301.275 725.370 ;
        RECT 1300.270 724.705 1300.570 725.070 ;
        RECT 1300.945 725.055 1301.275 725.070 ;
        RECT 1300.270 724.390 1300.815 724.705 ;
        RECT 1300.485 724.375 1300.815 724.390 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1388.425 1686.995 1388.595 1687.675 ;
        RECT 1315.745 1684.785 1315.915 1686.995 ;
        RECT 1387.965 1686.825 1388.595 1686.995 ;
      LAYER mcon ;
        RECT 1388.425 1687.505 1388.595 1687.675 ;
        RECT 1315.745 1686.825 1315.915 1686.995 ;
      LAYER met1 ;
        RECT 1388.365 1687.660 1388.655 1687.705 ;
        RECT 1403.530 1687.660 1403.850 1687.720 ;
        RECT 1388.365 1687.520 1403.850 1687.660 ;
        RECT 1388.365 1687.475 1388.655 1687.520 ;
        RECT 1403.530 1687.460 1403.850 1687.520 ;
        RECT 1300.950 1686.980 1301.270 1687.040 ;
        RECT 1315.685 1686.980 1315.975 1687.025 ;
        RECT 1387.905 1686.980 1388.195 1687.025 ;
        RECT 1300.950 1686.840 1315.975 1686.980 ;
        RECT 1300.950 1686.780 1301.270 1686.840 ;
        RECT 1315.685 1686.795 1315.975 1686.840 ;
        RECT 1318.520 1686.840 1388.195 1686.980 ;
        RECT 1315.685 1684.940 1315.975 1684.985 ;
        RECT 1318.520 1684.940 1318.660 1686.840 ;
        RECT 1387.905 1686.795 1388.195 1686.840 ;
        RECT 1315.685 1684.800 1318.660 1684.940 ;
        RECT 1315.685 1684.755 1315.975 1684.800 ;
        RECT 1403.530 1683.240 1403.850 1683.300 ;
        RECT 1469.770 1683.240 1470.090 1683.300 ;
        RECT 1403.530 1683.100 1470.090 1683.240 ;
        RECT 1403.530 1683.040 1403.850 1683.100 ;
        RECT 1469.770 1683.040 1470.090 1683.100 ;
      LAYER via ;
        RECT 1403.560 1687.460 1403.820 1687.720 ;
        RECT 1300.980 1686.780 1301.240 1687.040 ;
        RECT 1403.560 1683.040 1403.820 1683.300 ;
        RECT 1469.800 1683.040 1470.060 1683.300 ;
      LAYER met2 ;
        RECT 1300.880 1700.340 1301.160 1704.000 ;
        RECT 1300.880 1700.000 1301.180 1700.340 ;
        RECT 1301.040 1687.070 1301.180 1700.000 ;
        RECT 1403.560 1687.430 1403.820 1687.750 ;
        RECT 1300.980 1686.750 1301.240 1687.070 ;
        RECT 1403.620 1683.330 1403.760 1687.430 ;
        RECT 1403.560 1683.010 1403.820 1683.330 ;
        RECT 1469.800 1683.010 1470.060 1683.330 ;
        RECT 1469.860 3.130 1470.000 1683.010 ;
        RECT 1469.860 2.990 1471.840 3.130 ;
        RECT 1471.700 2.400 1471.840 2.990 ;
        RECT 1471.490 -4.800 1472.050 2.400 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1318.965 1685.635 1319.135 1688.015 ;
        RECT 1387.045 1687.845 1387.215 1688.695 ;
        RECT 1318.045 1685.465 1319.135 1685.635 ;
      LAYER mcon ;
        RECT 1387.045 1688.525 1387.215 1688.695 ;
        RECT 1318.965 1687.845 1319.135 1688.015 ;
      LAYER met1 ;
        RECT 1386.985 1688.680 1387.275 1688.725 ;
        RECT 1398.010 1688.680 1398.330 1688.740 ;
        RECT 1386.985 1688.540 1398.330 1688.680 ;
        RECT 1386.985 1688.495 1387.275 1688.540 ;
        RECT 1398.010 1688.480 1398.330 1688.540 ;
        RECT 1318.905 1688.000 1319.195 1688.045 ;
        RECT 1386.985 1688.000 1387.275 1688.045 ;
        RECT 1318.905 1687.860 1387.275 1688.000 ;
        RECT 1318.905 1687.815 1319.195 1687.860 ;
        RECT 1386.985 1687.815 1387.275 1687.860 ;
        RECT 1302.790 1686.640 1303.110 1686.700 ;
        RECT 1302.790 1686.500 1311.300 1686.640 ;
        RECT 1302.790 1686.440 1303.110 1686.500 ;
        RECT 1311.160 1685.620 1311.300 1686.500 ;
        RECT 1317.985 1685.620 1318.275 1685.665 ;
        RECT 1311.160 1685.480 1318.275 1685.620 ;
        RECT 1317.985 1685.435 1318.275 1685.480 ;
        RECT 1398.010 1682.900 1398.330 1682.960 ;
        RECT 1483.570 1682.900 1483.890 1682.960 ;
        RECT 1398.010 1682.760 1483.890 1682.900 ;
        RECT 1398.010 1682.700 1398.330 1682.760 ;
        RECT 1483.570 1682.700 1483.890 1682.760 ;
        RECT 1483.570 20.980 1483.890 21.040 ;
        RECT 1489.550 20.980 1489.870 21.040 ;
        RECT 1483.570 20.840 1489.870 20.980 ;
        RECT 1483.570 20.780 1483.890 20.840 ;
        RECT 1489.550 20.780 1489.870 20.840 ;
      LAYER via ;
        RECT 1398.040 1688.480 1398.300 1688.740 ;
        RECT 1302.820 1686.440 1303.080 1686.700 ;
        RECT 1398.040 1682.700 1398.300 1682.960 ;
        RECT 1483.600 1682.700 1483.860 1682.960 ;
        RECT 1483.600 20.780 1483.860 21.040 ;
        RECT 1489.580 20.780 1489.840 21.040 ;
      LAYER met2 ;
        RECT 1302.720 1700.340 1303.000 1704.000 ;
        RECT 1302.720 1700.000 1303.020 1700.340 ;
        RECT 1302.880 1686.730 1303.020 1700.000 ;
        RECT 1398.040 1688.450 1398.300 1688.770 ;
        RECT 1302.820 1686.410 1303.080 1686.730 ;
        RECT 1398.100 1682.990 1398.240 1688.450 ;
        RECT 1398.040 1682.670 1398.300 1682.990 ;
        RECT 1483.600 1682.670 1483.860 1682.990 ;
        RECT 1483.660 21.070 1483.800 1682.670 ;
        RECT 1483.600 20.750 1483.860 21.070 ;
        RECT 1489.580 20.750 1489.840 21.070 ;
        RECT 1489.640 2.400 1489.780 20.750 ;
        RECT 1489.430 -4.800 1489.990 2.400 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1352.545 1683.425 1352.715 1687.675 ;
        RECT 1381.525 1683.765 1381.695 1685.975 ;
        RECT 1412.345 1675.605 1412.515 1685.975 ;
      LAYER mcon ;
        RECT 1352.545 1687.505 1352.715 1687.675 ;
        RECT 1381.525 1685.805 1381.695 1685.975 ;
        RECT 1412.345 1685.805 1412.515 1685.975 ;
      LAYER met1 ;
        RECT 1304.630 1687.660 1304.950 1687.720 ;
        RECT 1352.485 1687.660 1352.775 1687.705 ;
        RECT 1304.630 1687.520 1352.775 1687.660 ;
        RECT 1304.630 1687.460 1304.950 1687.520 ;
        RECT 1352.485 1687.475 1352.775 1687.520 ;
        RECT 1381.465 1685.960 1381.755 1686.005 ;
        RECT 1412.285 1685.960 1412.575 1686.005 ;
        RECT 1381.465 1685.820 1412.575 1685.960 ;
        RECT 1381.465 1685.775 1381.755 1685.820 ;
        RECT 1412.285 1685.775 1412.575 1685.820 ;
        RECT 1381.465 1683.920 1381.755 1683.965 ;
        RECT 1377.400 1683.780 1381.755 1683.920 ;
        RECT 1352.485 1683.580 1352.775 1683.625 ;
        RECT 1377.400 1683.580 1377.540 1683.780 ;
        RECT 1381.465 1683.735 1381.755 1683.780 ;
        RECT 1352.485 1683.440 1377.540 1683.580 ;
        RECT 1352.485 1683.395 1352.775 1683.440 ;
        RECT 1412.285 1675.760 1412.575 1675.805 ;
        RECT 1412.285 1675.620 1413.420 1675.760 ;
        RECT 1412.285 1675.575 1412.575 1675.620 ;
        RECT 1413.280 1675.420 1413.420 1675.620 ;
        RECT 1504.270 1675.420 1504.590 1675.480 ;
        RECT 1413.280 1675.280 1504.590 1675.420 ;
        RECT 1504.270 1675.220 1504.590 1675.280 ;
        RECT 1504.270 2.960 1504.590 3.020 ;
        RECT 1507.030 2.960 1507.350 3.020 ;
        RECT 1504.270 2.820 1507.350 2.960 ;
        RECT 1504.270 2.760 1504.590 2.820 ;
        RECT 1507.030 2.760 1507.350 2.820 ;
      LAYER via ;
        RECT 1304.660 1687.460 1304.920 1687.720 ;
        RECT 1504.300 1675.220 1504.560 1675.480 ;
        RECT 1504.300 2.760 1504.560 3.020 ;
        RECT 1507.060 2.760 1507.320 3.020 ;
      LAYER met2 ;
        RECT 1304.560 1700.340 1304.840 1704.000 ;
        RECT 1304.560 1700.000 1304.860 1700.340 ;
        RECT 1304.720 1687.750 1304.860 1700.000 ;
        RECT 1304.660 1687.430 1304.920 1687.750 ;
        RECT 1504.300 1675.190 1504.560 1675.510 ;
        RECT 1504.360 3.050 1504.500 1675.190 ;
        RECT 1504.300 2.730 1504.560 3.050 ;
        RECT 1507.060 2.730 1507.320 3.050 ;
        RECT 1507.120 2.400 1507.260 2.730 ;
        RECT 1506.910 -4.800 1507.470 2.400 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1222.290 1678.280 1222.610 1678.540 ;
        RECT 1222.380 1677.120 1222.520 1678.280 ;
        RECT 1221.460 1676.980 1222.520 1677.120 ;
        RECT 1221.460 1676.840 1221.600 1676.980 ;
        RECT 1221.370 1676.580 1221.690 1676.840 ;
        RECT 710.310 1660.460 710.630 1660.520 ;
        RECT 1221.370 1660.460 1221.690 1660.520 ;
        RECT 710.310 1660.320 1221.690 1660.460 ;
        RECT 710.310 1660.260 710.630 1660.320 ;
        RECT 1221.370 1660.260 1221.690 1660.320 ;
        RECT 704.330 26.080 704.650 26.140 ;
        RECT 710.310 26.080 710.630 26.140 ;
        RECT 704.330 25.940 710.630 26.080 ;
        RECT 704.330 25.880 704.650 25.940 ;
        RECT 710.310 25.880 710.630 25.940 ;
      LAYER via ;
        RECT 1222.320 1678.280 1222.580 1678.540 ;
        RECT 1221.400 1676.580 1221.660 1676.840 ;
        RECT 710.340 1660.260 710.600 1660.520 ;
        RECT 1221.400 1660.260 1221.660 1660.520 ;
        RECT 704.360 25.880 704.620 26.140 ;
        RECT 710.340 25.880 710.600 26.140 ;
      LAYER met2 ;
        RECT 1222.220 1700.340 1222.500 1704.000 ;
        RECT 1222.220 1700.000 1222.520 1700.340 ;
        RECT 1222.380 1678.570 1222.520 1700.000 ;
        RECT 1222.320 1678.250 1222.580 1678.570 ;
        RECT 1221.400 1676.550 1221.660 1676.870 ;
        RECT 1221.460 1660.550 1221.600 1676.550 ;
        RECT 710.340 1660.230 710.600 1660.550 ;
        RECT 1221.400 1660.230 1221.660 1660.550 ;
        RECT 710.400 26.170 710.540 1660.230 ;
        RECT 704.360 25.850 704.620 26.170 ;
        RECT 710.340 25.850 710.600 26.170 ;
        RECT 704.420 2.400 704.560 25.850 ;
        RECT 704.210 -4.800 704.770 2.400 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1306.470 1685.620 1306.790 1685.680 ;
        RECT 1308.310 1685.620 1308.630 1685.680 ;
        RECT 1306.470 1685.480 1308.630 1685.620 ;
        RECT 1306.470 1685.420 1306.790 1685.480 ;
        RECT 1308.310 1685.420 1308.630 1685.480 ;
        RECT 1308.310 1682.560 1308.630 1682.620 ;
        RECT 1524.970 1682.560 1525.290 1682.620 ;
        RECT 1308.310 1682.420 1525.290 1682.560 ;
        RECT 1308.310 1682.360 1308.630 1682.420 ;
        RECT 1524.970 1682.360 1525.290 1682.420 ;
      LAYER via ;
        RECT 1306.500 1685.420 1306.760 1685.680 ;
        RECT 1308.340 1685.420 1308.600 1685.680 ;
        RECT 1308.340 1682.360 1308.600 1682.620 ;
        RECT 1525.000 1682.360 1525.260 1682.620 ;
      LAYER met2 ;
        RECT 1306.400 1700.340 1306.680 1704.000 ;
        RECT 1306.400 1700.000 1306.700 1700.340 ;
        RECT 1306.560 1685.710 1306.700 1700.000 ;
        RECT 1306.500 1685.390 1306.760 1685.710 ;
        RECT 1308.340 1685.390 1308.600 1685.710 ;
        RECT 1308.400 1682.650 1308.540 1685.390 ;
        RECT 1308.340 1682.330 1308.600 1682.650 ;
        RECT 1525.000 1682.330 1525.260 1682.650 ;
        RECT 1525.060 2.400 1525.200 1682.330 ;
        RECT 1524.850 -4.800 1525.410 2.400 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1307.390 1686.300 1307.710 1686.360 ;
        RECT 1308.310 1686.300 1308.630 1686.360 ;
        RECT 1307.390 1686.160 1308.630 1686.300 ;
        RECT 1307.390 1686.100 1307.710 1686.160 ;
        RECT 1308.310 1686.100 1308.630 1686.160 ;
        RECT 1307.390 1668.280 1307.710 1668.340 ;
        RECT 1538.770 1668.280 1539.090 1668.340 ;
        RECT 1307.390 1668.140 1539.090 1668.280 ;
        RECT 1307.390 1668.080 1307.710 1668.140 ;
        RECT 1538.770 1668.080 1539.090 1668.140 ;
      LAYER via ;
        RECT 1307.420 1686.100 1307.680 1686.360 ;
        RECT 1308.340 1686.100 1308.600 1686.360 ;
        RECT 1307.420 1668.080 1307.680 1668.340 ;
        RECT 1538.800 1668.080 1539.060 1668.340 ;
      LAYER met2 ;
        RECT 1308.240 1700.340 1308.520 1704.000 ;
        RECT 1308.240 1700.000 1308.540 1700.340 ;
        RECT 1308.400 1686.390 1308.540 1700.000 ;
        RECT 1307.420 1686.070 1307.680 1686.390 ;
        RECT 1308.340 1686.070 1308.600 1686.390 ;
        RECT 1307.480 1668.370 1307.620 1686.070 ;
        RECT 1307.420 1668.050 1307.680 1668.370 ;
        RECT 1538.800 1668.050 1539.060 1668.370 ;
        RECT 1538.860 17.410 1539.000 1668.050 ;
        RECT 1538.860 17.270 1543.140 17.410 ;
        RECT 1543.000 2.400 1543.140 17.270 ;
        RECT 1542.790 -4.800 1543.350 2.400 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1310.610 1675.080 1310.930 1675.140 ;
        RECT 1559.470 1675.080 1559.790 1675.140 ;
        RECT 1310.610 1674.940 1559.790 1675.080 ;
        RECT 1310.610 1674.880 1310.930 1674.940 ;
        RECT 1559.470 1674.880 1559.790 1674.940 ;
      LAYER via ;
        RECT 1310.640 1674.880 1310.900 1675.140 ;
        RECT 1559.500 1674.880 1559.760 1675.140 ;
      LAYER met2 ;
        RECT 1310.080 1700.340 1310.360 1704.000 ;
        RECT 1310.080 1700.000 1310.380 1700.340 ;
        RECT 1310.240 1685.450 1310.380 1700.000 ;
        RECT 1310.240 1685.310 1310.840 1685.450 ;
        RECT 1310.700 1675.170 1310.840 1685.310 ;
        RECT 1310.640 1674.850 1310.900 1675.170 ;
        RECT 1559.500 1674.850 1559.760 1675.170 ;
        RECT 1559.560 17.410 1559.700 1674.850 ;
        RECT 1559.560 17.270 1561.080 17.410 ;
        RECT 1560.940 2.400 1561.080 17.270 ;
        RECT 1560.730 -4.800 1561.290 2.400 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1311.990 1689.020 1312.310 1689.080 ;
        RECT 1327.630 1689.020 1327.950 1689.080 ;
        RECT 1311.990 1688.880 1327.950 1689.020 ;
        RECT 1311.990 1688.820 1312.310 1688.880 ;
        RECT 1327.630 1688.820 1327.950 1688.880 ;
        RECT 1327.630 1682.220 1327.950 1682.280 ;
        RECT 1573.270 1682.220 1573.590 1682.280 ;
        RECT 1327.630 1682.080 1573.590 1682.220 ;
        RECT 1327.630 1682.020 1327.950 1682.080 ;
        RECT 1573.270 1682.020 1573.590 1682.080 ;
      LAYER via ;
        RECT 1312.020 1688.820 1312.280 1689.080 ;
        RECT 1327.660 1688.820 1327.920 1689.080 ;
        RECT 1327.660 1682.020 1327.920 1682.280 ;
        RECT 1573.300 1682.020 1573.560 1682.280 ;
      LAYER met2 ;
        RECT 1311.920 1700.340 1312.200 1704.000 ;
        RECT 1311.920 1700.000 1312.220 1700.340 ;
        RECT 1312.080 1689.110 1312.220 1700.000 ;
        RECT 1312.020 1688.790 1312.280 1689.110 ;
        RECT 1327.660 1688.790 1327.920 1689.110 ;
        RECT 1327.720 1682.310 1327.860 1688.790 ;
        RECT 1327.660 1681.990 1327.920 1682.310 ;
        RECT 1573.300 1681.990 1573.560 1682.310 ;
        RECT 1573.360 17.410 1573.500 1681.990 ;
        RECT 1573.360 17.270 1579.020 17.410 ;
        RECT 1578.880 2.400 1579.020 17.270 ;
        RECT 1578.670 -4.800 1579.230 2.400 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1313.830 1685.280 1314.150 1685.340 ;
        RECT 1314.750 1685.280 1315.070 1685.340 ;
        RECT 1313.830 1685.140 1315.070 1685.280 ;
        RECT 1313.830 1685.080 1314.150 1685.140 ;
        RECT 1314.750 1685.080 1315.070 1685.140 ;
        RECT 1314.750 1667.940 1315.070 1668.000 ;
        RECT 1593.970 1667.940 1594.290 1668.000 ;
        RECT 1314.750 1667.800 1594.290 1667.940 ;
        RECT 1314.750 1667.740 1315.070 1667.800 ;
        RECT 1593.970 1667.740 1594.290 1667.800 ;
      LAYER via ;
        RECT 1313.860 1685.080 1314.120 1685.340 ;
        RECT 1314.780 1685.080 1315.040 1685.340 ;
        RECT 1314.780 1667.740 1315.040 1668.000 ;
        RECT 1594.000 1667.740 1594.260 1668.000 ;
      LAYER met2 ;
        RECT 1313.760 1700.340 1314.040 1704.000 ;
        RECT 1313.760 1700.000 1314.060 1700.340 ;
        RECT 1313.920 1685.370 1314.060 1700.000 ;
        RECT 1313.860 1685.050 1314.120 1685.370 ;
        RECT 1314.780 1685.050 1315.040 1685.370 ;
        RECT 1314.840 1668.030 1314.980 1685.050 ;
        RECT 1314.780 1667.710 1315.040 1668.030 ;
        RECT 1594.000 1667.710 1594.260 1668.030 ;
        RECT 1594.060 17.410 1594.200 1667.710 ;
        RECT 1594.060 17.270 1596.500 17.410 ;
        RECT 1596.360 2.400 1596.500 17.270 ;
        RECT 1596.150 -4.800 1596.710 2.400 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1313.370 1684.260 1313.690 1684.320 ;
        RECT 1315.670 1684.260 1315.990 1684.320 ;
        RECT 1313.370 1684.120 1315.990 1684.260 ;
        RECT 1313.370 1684.060 1313.690 1684.120 ;
        RECT 1315.670 1684.060 1315.990 1684.120 ;
        RECT 1313.370 27.780 1313.690 27.840 ;
        RECT 1614.210 27.780 1614.530 27.840 ;
        RECT 1313.370 27.640 1614.530 27.780 ;
        RECT 1313.370 27.580 1313.690 27.640 ;
        RECT 1614.210 27.580 1614.530 27.640 ;
      LAYER via ;
        RECT 1313.400 1684.060 1313.660 1684.320 ;
        RECT 1315.700 1684.060 1315.960 1684.320 ;
        RECT 1313.400 27.580 1313.660 27.840 ;
        RECT 1614.240 27.580 1614.500 27.840 ;
      LAYER met2 ;
        RECT 1315.600 1700.340 1315.880 1704.000 ;
        RECT 1315.600 1700.000 1315.900 1700.340 ;
        RECT 1315.760 1684.350 1315.900 1700.000 ;
        RECT 1313.400 1684.030 1313.660 1684.350 ;
        RECT 1315.700 1684.030 1315.960 1684.350 ;
        RECT 1313.460 27.870 1313.600 1684.030 ;
        RECT 1313.400 27.550 1313.660 27.870 ;
        RECT 1614.240 27.550 1614.500 27.870 ;
        RECT 1614.300 2.400 1614.440 27.550 ;
        RECT 1614.090 -4.800 1614.650 2.400 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1313.830 1684.600 1314.150 1684.660 ;
        RECT 1317.510 1684.600 1317.830 1684.660 ;
        RECT 1313.830 1684.460 1317.830 1684.600 ;
        RECT 1313.830 1684.400 1314.150 1684.460 ;
        RECT 1317.510 1684.400 1317.830 1684.460 ;
        RECT 1313.830 28.120 1314.150 28.180 ;
        RECT 1632.150 28.120 1632.470 28.180 ;
        RECT 1313.830 27.980 1632.470 28.120 ;
        RECT 1313.830 27.920 1314.150 27.980 ;
        RECT 1632.150 27.920 1632.470 27.980 ;
      LAYER via ;
        RECT 1313.860 1684.400 1314.120 1684.660 ;
        RECT 1317.540 1684.400 1317.800 1684.660 ;
        RECT 1313.860 27.920 1314.120 28.180 ;
        RECT 1632.180 27.920 1632.440 28.180 ;
      LAYER met2 ;
        RECT 1317.440 1700.340 1317.720 1704.000 ;
        RECT 1317.440 1700.000 1317.740 1700.340 ;
        RECT 1317.600 1684.690 1317.740 1700.000 ;
        RECT 1313.860 1684.370 1314.120 1684.690 ;
        RECT 1317.540 1684.370 1317.800 1684.690 ;
        RECT 1313.920 28.210 1314.060 1684.370 ;
        RECT 1313.860 27.890 1314.120 28.210 ;
        RECT 1632.180 27.890 1632.440 28.210 ;
        RECT 1632.240 2.400 1632.380 27.890 ;
        RECT 1632.030 -4.800 1632.590 2.400 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1320.270 28.460 1320.590 28.520 ;
        RECT 1650.090 28.460 1650.410 28.520 ;
        RECT 1320.270 28.320 1650.410 28.460 ;
        RECT 1320.270 28.260 1320.590 28.320 ;
        RECT 1650.090 28.260 1650.410 28.320 ;
      LAYER via ;
        RECT 1320.300 28.260 1320.560 28.520 ;
        RECT 1650.120 28.260 1650.380 28.520 ;
      LAYER met2 ;
        RECT 1319.280 1700.340 1319.560 1704.000 ;
        RECT 1319.280 1700.000 1319.580 1700.340 ;
        RECT 1319.440 1684.770 1319.580 1700.000 ;
        RECT 1319.440 1684.630 1320.500 1684.770 ;
        RECT 1320.360 28.550 1320.500 1684.630 ;
        RECT 1320.300 28.230 1320.560 28.550 ;
        RECT 1650.120 28.230 1650.380 28.550 ;
        RECT 1650.180 2.400 1650.320 28.230 ;
        RECT 1649.970 -4.800 1650.530 2.400 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1321.190 28.800 1321.510 28.860 ;
        RECT 1668.030 28.800 1668.350 28.860 ;
        RECT 1321.190 28.660 1668.350 28.800 ;
        RECT 1321.190 28.600 1321.510 28.660 ;
        RECT 1668.030 28.600 1668.350 28.660 ;
      LAYER via ;
        RECT 1321.220 28.600 1321.480 28.860 ;
        RECT 1668.060 28.600 1668.320 28.860 ;
      LAYER met2 ;
        RECT 1321.120 1700.340 1321.400 1704.000 ;
        RECT 1321.120 1700.000 1321.420 1700.340 ;
        RECT 1321.280 28.890 1321.420 1700.000 ;
        RECT 1321.220 28.570 1321.480 28.890 ;
        RECT 1668.060 28.570 1668.320 28.890 ;
        RECT 1668.120 2.400 1668.260 28.570 ;
        RECT 1667.910 -4.800 1668.470 2.400 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1321.650 1683.920 1321.970 1683.980 ;
        RECT 1323.030 1683.920 1323.350 1683.980 ;
        RECT 1321.650 1683.780 1323.350 1683.920 ;
        RECT 1321.650 1683.720 1321.970 1683.780 ;
        RECT 1323.030 1683.720 1323.350 1683.780 ;
        RECT 1321.650 29.140 1321.970 29.200 ;
        RECT 1685.510 29.140 1685.830 29.200 ;
        RECT 1321.650 29.000 1685.830 29.140 ;
        RECT 1321.650 28.940 1321.970 29.000 ;
        RECT 1685.510 28.940 1685.830 29.000 ;
      LAYER via ;
        RECT 1321.680 1683.720 1321.940 1683.980 ;
        RECT 1323.060 1683.720 1323.320 1683.980 ;
        RECT 1321.680 28.940 1321.940 29.200 ;
        RECT 1685.540 28.940 1685.800 29.200 ;
      LAYER met2 ;
        RECT 1322.960 1700.340 1323.240 1704.000 ;
        RECT 1322.960 1700.000 1323.260 1700.340 ;
        RECT 1323.120 1684.010 1323.260 1700.000 ;
        RECT 1321.680 1683.690 1321.940 1684.010 ;
        RECT 1323.060 1683.690 1323.320 1684.010 ;
        RECT 1321.740 29.230 1321.880 1683.690 ;
        RECT 1321.680 28.910 1321.940 29.230 ;
        RECT 1685.540 28.910 1685.800 29.230 ;
        RECT 1685.600 2.400 1685.740 28.910 ;
        RECT 1685.390 -4.800 1685.950 2.400 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1221.370 1679.160 1221.690 1679.220 ;
        RECT 1223.670 1679.160 1223.990 1679.220 ;
        RECT 1221.370 1679.020 1223.990 1679.160 ;
        RECT 1221.370 1678.960 1221.690 1679.020 ;
        RECT 1223.670 1678.960 1223.990 1679.020 ;
        RECT 724.110 1653.660 724.430 1653.720 ;
        RECT 1222.290 1653.660 1222.610 1653.720 ;
        RECT 724.110 1653.520 1222.610 1653.660 ;
        RECT 724.110 1653.460 724.430 1653.520 ;
        RECT 1222.290 1653.460 1222.610 1653.520 ;
      LAYER via ;
        RECT 1221.400 1678.960 1221.660 1679.220 ;
        RECT 1223.700 1678.960 1223.960 1679.220 ;
        RECT 724.140 1653.460 724.400 1653.720 ;
        RECT 1222.320 1653.460 1222.580 1653.720 ;
      LAYER met2 ;
        RECT 1224.060 1700.410 1224.340 1704.000 ;
        RECT 1223.760 1700.270 1224.340 1700.410 ;
        RECT 1223.760 1679.250 1223.900 1700.270 ;
        RECT 1224.060 1700.000 1224.340 1700.270 ;
        RECT 1221.400 1678.930 1221.660 1679.250 ;
        RECT 1223.700 1678.930 1223.960 1679.250 ;
        RECT 1221.460 1677.290 1221.600 1678.930 ;
        RECT 1221.460 1677.150 1222.520 1677.290 ;
        RECT 1222.380 1653.750 1222.520 1677.150 ;
        RECT 724.140 1653.430 724.400 1653.750 ;
        RECT 1222.320 1653.430 1222.580 1653.750 ;
        RECT 724.200 16.730 724.340 1653.430 ;
        RECT 722.360 16.590 724.340 16.730 ;
        RECT 722.360 2.400 722.500 16.590 ;
        RECT 722.150 -4.800 722.710 2.400 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1324.870 1685.620 1325.190 1685.680 ;
        RECT 1329.470 1685.620 1329.790 1685.680 ;
        RECT 1324.870 1685.480 1329.790 1685.620 ;
        RECT 1324.870 1685.420 1325.190 1685.480 ;
        RECT 1329.470 1685.420 1329.790 1685.480 ;
        RECT 1329.930 29.480 1330.250 29.540 ;
        RECT 1703.450 29.480 1703.770 29.540 ;
        RECT 1329.930 29.340 1703.770 29.480 ;
        RECT 1329.930 29.280 1330.250 29.340 ;
        RECT 1703.450 29.280 1703.770 29.340 ;
      LAYER via ;
        RECT 1324.900 1685.420 1325.160 1685.680 ;
        RECT 1329.500 1685.420 1329.760 1685.680 ;
        RECT 1329.960 29.280 1330.220 29.540 ;
        RECT 1703.480 29.280 1703.740 29.540 ;
      LAYER met2 ;
        RECT 1324.800 1700.340 1325.080 1704.000 ;
        RECT 1324.800 1700.000 1325.100 1700.340 ;
        RECT 1324.960 1685.710 1325.100 1700.000 ;
        RECT 1324.900 1685.390 1325.160 1685.710 ;
        RECT 1329.500 1685.390 1329.760 1685.710 ;
        RECT 1329.560 1684.770 1329.700 1685.390 ;
        RECT 1329.560 1684.630 1330.160 1684.770 ;
        RECT 1330.020 29.570 1330.160 1684.630 ;
        RECT 1329.960 29.250 1330.220 29.570 ;
        RECT 1703.480 29.250 1703.740 29.570 ;
        RECT 1703.540 2.400 1703.680 29.250 ;
        RECT 1703.330 -4.800 1703.890 2.400 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1326.710 1681.540 1327.030 1681.600 ;
        RECT 1327.630 1681.540 1327.950 1681.600 ;
        RECT 1326.710 1681.400 1327.950 1681.540 ;
        RECT 1326.710 1681.340 1327.030 1681.400 ;
        RECT 1327.630 1681.340 1327.950 1681.400 ;
        RECT 1326.710 1594.160 1327.030 1594.220 ;
        RECT 1327.630 1594.160 1327.950 1594.220 ;
        RECT 1326.710 1594.020 1327.950 1594.160 ;
        RECT 1326.710 1593.960 1327.030 1594.020 ;
        RECT 1327.630 1593.960 1327.950 1594.020 ;
        RECT 1327.630 29.820 1327.950 29.880 ;
        RECT 1721.390 29.820 1721.710 29.880 ;
        RECT 1327.630 29.680 1721.710 29.820 ;
        RECT 1327.630 29.620 1327.950 29.680 ;
        RECT 1721.390 29.620 1721.710 29.680 ;
      LAYER via ;
        RECT 1326.740 1681.340 1327.000 1681.600 ;
        RECT 1327.660 1681.340 1327.920 1681.600 ;
        RECT 1326.740 1593.960 1327.000 1594.220 ;
        RECT 1327.660 1593.960 1327.920 1594.220 ;
        RECT 1327.660 29.620 1327.920 29.880 ;
        RECT 1721.420 29.620 1721.680 29.880 ;
      LAYER met2 ;
        RECT 1326.640 1700.340 1326.920 1704.000 ;
        RECT 1326.640 1700.000 1326.940 1700.340 ;
        RECT 1326.800 1681.630 1326.940 1700.000 ;
        RECT 1326.740 1681.310 1327.000 1681.630 ;
        RECT 1327.660 1681.310 1327.920 1681.630 ;
        RECT 1327.720 1594.250 1327.860 1681.310 ;
        RECT 1326.740 1593.930 1327.000 1594.250 ;
        RECT 1327.660 1593.930 1327.920 1594.250 ;
        RECT 1326.800 1593.650 1326.940 1593.930 ;
        RECT 1326.800 1593.510 1327.860 1593.650 ;
        RECT 1327.720 29.910 1327.860 1593.510 ;
        RECT 1327.660 29.590 1327.920 29.910 ;
        RECT 1721.420 29.590 1721.680 29.910 ;
        RECT 1721.480 2.400 1721.620 29.590 ;
        RECT 1721.270 -4.800 1721.830 2.400 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1328.550 1683.920 1328.870 1683.980 ;
        RECT 1329.470 1683.920 1329.790 1683.980 ;
        RECT 1328.550 1683.780 1329.790 1683.920 ;
        RECT 1328.550 1683.720 1328.870 1683.780 ;
        RECT 1329.470 1683.720 1329.790 1683.780 ;
        RECT 1329.470 1631.900 1329.790 1631.960 ;
        RECT 1330.390 1631.900 1330.710 1631.960 ;
        RECT 1329.470 1631.760 1330.710 1631.900 ;
        RECT 1329.470 1631.700 1329.790 1631.760 ;
        RECT 1330.390 1631.700 1330.710 1631.760 ;
        RECT 1330.390 30.160 1330.710 30.220 ;
        RECT 1739.330 30.160 1739.650 30.220 ;
        RECT 1330.390 30.020 1739.650 30.160 ;
        RECT 1330.390 29.960 1330.710 30.020 ;
        RECT 1739.330 29.960 1739.650 30.020 ;
      LAYER via ;
        RECT 1328.580 1683.720 1328.840 1683.980 ;
        RECT 1329.500 1683.720 1329.760 1683.980 ;
        RECT 1329.500 1631.700 1329.760 1631.960 ;
        RECT 1330.420 1631.700 1330.680 1631.960 ;
        RECT 1330.420 29.960 1330.680 30.220 ;
        RECT 1739.360 29.960 1739.620 30.220 ;
      LAYER met2 ;
        RECT 1328.480 1700.340 1328.760 1704.000 ;
        RECT 1328.480 1700.000 1328.780 1700.340 ;
        RECT 1328.640 1684.010 1328.780 1700.000 ;
        RECT 1328.580 1683.690 1328.840 1684.010 ;
        RECT 1329.500 1683.690 1329.760 1684.010 ;
        RECT 1329.560 1631.990 1329.700 1683.690 ;
        RECT 1329.500 1631.670 1329.760 1631.990 ;
        RECT 1330.420 1631.670 1330.680 1631.990 ;
        RECT 1330.480 30.250 1330.620 1631.670 ;
        RECT 1330.420 29.930 1330.680 30.250 ;
        RECT 1739.360 29.930 1739.620 30.250 ;
        RECT 1739.420 2.400 1739.560 29.930 ;
        RECT 1739.210 -4.800 1739.770 2.400 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1326.250 1684.940 1326.570 1685.000 ;
        RECT 1330.390 1684.940 1330.710 1685.000 ;
        RECT 1326.250 1684.800 1330.710 1684.940 ;
        RECT 1326.250 1684.740 1326.570 1684.800 ;
        RECT 1330.390 1684.740 1330.710 1684.800 ;
        RECT 1326.710 30.500 1327.030 30.560 ;
        RECT 1756.810 30.500 1757.130 30.560 ;
        RECT 1326.710 30.360 1757.130 30.500 ;
        RECT 1326.710 30.300 1327.030 30.360 ;
        RECT 1756.810 30.300 1757.130 30.360 ;
      LAYER via ;
        RECT 1326.280 1684.740 1326.540 1685.000 ;
        RECT 1330.420 1684.740 1330.680 1685.000 ;
        RECT 1326.740 30.300 1327.000 30.560 ;
        RECT 1756.840 30.300 1757.100 30.560 ;
      LAYER met2 ;
        RECT 1330.320 1700.340 1330.600 1704.000 ;
        RECT 1330.320 1700.000 1330.620 1700.340 ;
        RECT 1330.480 1685.030 1330.620 1700.000 ;
        RECT 1326.280 1684.710 1326.540 1685.030 ;
        RECT 1330.420 1684.710 1330.680 1685.030 ;
        RECT 1326.340 1558.970 1326.480 1684.710 ;
        RECT 1326.340 1558.830 1326.940 1558.970 ;
        RECT 1326.800 30.590 1326.940 1558.830 ;
        RECT 1326.740 30.270 1327.000 30.590 ;
        RECT 1756.840 30.270 1757.100 30.590 ;
        RECT 1756.900 2.400 1757.040 30.270 ;
        RECT 1756.690 -4.800 1757.250 2.400 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1332.230 34.240 1332.550 34.300 ;
        RECT 1774.750 34.240 1775.070 34.300 ;
        RECT 1332.230 34.100 1775.070 34.240 ;
        RECT 1332.230 34.040 1332.550 34.100 ;
        RECT 1774.750 34.040 1775.070 34.100 ;
      LAYER via ;
        RECT 1332.260 34.040 1332.520 34.300 ;
        RECT 1774.780 34.040 1775.040 34.300 ;
      LAYER met2 ;
        RECT 1332.160 1700.340 1332.440 1704.000 ;
        RECT 1332.160 1700.000 1332.460 1700.340 ;
        RECT 1332.320 34.330 1332.460 1700.000 ;
        RECT 1332.260 34.010 1332.520 34.330 ;
        RECT 1774.780 34.010 1775.040 34.330 ;
        RECT 1774.840 2.400 1774.980 34.010 ;
        RECT 1774.630 -4.800 1775.190 2.400 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1334.070 33.900 1334.390 33.960 ;
        RECT 1792.690 33.900 1793.010 33.960 ;
        RECT 1334.070 33.760 1793.010 33.900 ;
        RECT 1334.070 33.700 1334.390 33.760 ;
        RECT 1792.690 33.700 1793.010 33.760 ;
      LAYER via ;
        RECT 1334.100 33.700 1334.360 33.960 ;
        RECT 1792.720 33.700 1792.980 33.960 ;
      LAYER met2 ;
        RECT 1334.000 1700.340 1334.280 1704.000 ;
        RECT 1334.000 1700.000 1334.300 1700.340 ;
        RECT 1334.160 33.990 1334.300 1700.000 ;
        RECT 1334.100 33.670 1334.360 33.990 ;
        RECT 1792.720 33.670 1792.980 33.990 ;
        RECT 1792.780 2.400 1792.920 33.670 ;
        RECT 1792.570 -4.800 1793.130 2.400 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1333.610 1684.600 1333.930 1684.660 ;
        RECT 1335.910 1684.600 1336.230 1684.660 ;
        RECT 1333.610 1684.460 1336.230 1684.600 ;
        RECT 1333.610 1684.400 1333.930 1684.460 ;
        RECT 1335.910 1684.400 1336.230 1684.460 ;
        RECT 1333.610 33.560 1333.930 33.620 ;
        RECT 1810.630 33.560 1810.950 33.620 ;
        RECT 1333.610 33.420 1810.950 33.560 ;
        RECT 1333.610 33.360 1333.930 33.420 ;
        RECT 1810.630 33.360 1810.950 33.420 ;
      LAYER via ;
        RECT 1333.640 1684.400 1333.900 1684.660 ;
        RECT 1335.940 1684.400 1336.200 1684.660 ;
        RECT 1333.640 33.360 1333.900 33.620 ;
        RECT 1810.660 33.360 1810.920 33.620 ;
      LAYER met2 ;
        RECT 1335.840 1700.340 1336.120 1704.000 ;
        RECT 1335.840 1700.000 1336.140 1700.340 ;
        RECT 1336.000 1684.690 1336.140 1700.000 ;
        RECT 1333.640 1684.370 1333.900 1684.690 ;
        RECT 1335.940 1684.370 1336.200 1684.690 ;
        RECT 1333.700 33.650 1333.840 1684.370 ;
        RECT 1333.640 33.330 1333.900 33.650 ;
        RECT 1810.660 33.330 1810.920 33.650 ;
        RECT 1810.720 2.400 1810.860 33.330 ;
        RECT 1810.510 -4.800 1811.070 2.400 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1337.365 1642.285 1337.535 1690.395 ;
      LAYER mcon ;
        RECT 1337.365 1690.225 1337.535 1690.395 ;
      LAYER met1 ;
        RECT 1337.305 1690.380 1337.595 1690.425 ;
        RECT 1337.750 1690.380 1338.070 1690.440 ;
        RECT 1337.305 1690.240 1338.070 1690.380 ;
        RECT 1337.305 1690.195 1337.595 1690.240 ;
        RECT 1337.750 1690.180 1338.070 1690.240 ;
        RECT 1337.290 1642.440 1337.610 1642.500 ;
        RECT 1337.095 1642.300 1337.610 1642.440 ;
        RECT 1337.290 1642.240 1337.610 1642.300 ;
        RECT 1337.290 33.220 1337.610 33.280 ;
        RECT 1829.030 33.220 1829.350 33.280 ;
        RECT 1337.290 33.080 1829.350 33.220 ;
        RECT 1337.290 33.020 1337.610 33.080 ;
        RECT 1829.030 33.020 1829.350 33.080 ;
      LAYER via ;
        RECT 1337.780 1690.180 1338.040 1690.440 ;
        RECT 1337.320 1642.240 1337.580 1642.500 ;
        RECT 1337.320 33.020 1337.580 33.280 ;
        RECT 1829.060 33.020 1829.320 33.280 ;
      LAYER met2 ;
        RECT 1337.680 1700.340 1337.960 1704.000 ;
        RECT 1337.680 1700.000 1337.980 1700.340 ;
        RECT 1337.840 1690.470 1337.980 1700.000 ;
        RECT 1337.780 1690.150 1338.040 1690.470 ;
        RECT 1337.320 1642.210 1337.580 1642.530 ;
        RECT 1337.380 33.310 1337.520 1642.210 ;
        RECT 1337.320 32.990 1337.580 33.310 ;
        RECT 1829.060 32.990 1829.320 33.310 ;
        RECT 1829.120 16.730 1829.260 32.990 ;
        RECT 1828.660 16.590 1829.260 16.730 ;
        RECT 1828.660 2.400 1828.800 16.590 ;
        RECT 1828.450 -4.800 1829.010 2.400 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1339.665 1628.345 1339.835 1689.035 ;
      LAYER mcon ;
        RECT 1339.665 1688.865 1339.835 1689.035 ;
      LAYER met1 ;
        RECT 1339.590 1689.020 1339.910 1689.080 ;
        RECT 1339.395 1688.880 1339.910 1689.020 ;
        RECT 1339.590 1688.820 1339.910 1688.880 ;
        RECT 1339.605 1628.500 1339.895 1628.545 ;
        RECT 1345.110 1628.500 1345.430 1628.560 ;
        RECT 1339.605 1628.360 1345.430 1628.500 ;
        RECT 1339.605 1628.315 1339.895 1628.360 ;
        RECT 1345.110 1628.300 1345.430 1628.360 ;
        RECT 1345.110 1593.480 1345.430 1593.540 ;
        RECT 1346.030 1593.480 1346.350 1593.540 ;
        RECT 1345.110 1593.340 1346.350 1593.480 ;
        RECT 1345.110 1593.280 1345.430 1593.340 ;
        RECT 1346.030 1593.280 1346.350 1593.340 ;
        RECT 1345.110 32.880 1345.430 32.940 ;
        RECT 1846.050 32.880 1846.370 32.940 ;
        RECT 1345.110 32.740 1846.370 32.880 ;
        RECT 1345.110 32.680 1345.430 32.740 ;
        RECT 1846.050 32.680 1846.370 32.740 ;
      LAYER via ;
        RECT 1339.620 1688.820 1339.880 1689.080 ;
        RECT 1345.140 1628.300 1345.400 1628.560 ;
        RECT 1345.140 1593.280 1345.400 1593.540 ;
        RECT 1346.060 1593.280 1346.320 1593.540 ;
        RECT 1345.140 32.680 1345.400 32.940 ;
        RECT 1846.080 32.680 1846.340 32.940 ;
      LAYER met2 ;
        RECT 1339.520 1700.340 1339.800 1704.000 ;
        RECT 1339.520 1700.000 1339.820 1700.340 ;
        RECT 1339.680 1689.110 1339.820 1700.000 ;
        RECT 1339.620 1688.790 1339.880 1689.110 ;
        RECT 1345.140 1628.445 1345.400 1628.590 ;
        RECT 1345.130 1628.075 1345.410 1628.445 ;
        RECT 1346.050 1627.395 1346.330 1627.765 ;
        RECT 1346.120 1593.570 1346.260 1627.395 ;
        RECT 1345.140 1593.250 1345.400 1593.570 ;
        RECT 1346.060 1593.250 1346.320 1593.570 ;
        RECT 1345.200 32.970 1345.340 1593.250 ;
        RECT 1345.140 32.650 1345.400 32.970 ;
        RECT 1846.080 32.650 1846.340 32.970 ;
        RECT 1846.140 2.400 1846.280 32.650 ;
        RECT 1845.930 -4.800 1846.490 2.400 ;
      LAYER via2 ;
        RECT 1345.130 1628.120 1345.410 1628.400 ;
        RECT 1346.050 1627.440 1346.330 1627.720 ;
      LAYER met3 ;
        RECT 1345.105 1628.410 1345.435 1628.425 ;
        RECT 1345.105 1628.095 1345.650 1628.410 ;
        RECT 1345.350 1627.730 1345.650 1628.095 ;
        RECT 1346.025 1627.730 1346.355 1627.745 ;
        RECT 1345.350 1627.430 1346.355 1627.730 ;
        RECT 1346.025 1627.415 1346.355 1627.430 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1341.430 1684.600 1341.750 1684.660 ;
        RECT 1344.190 1684.600 1344.510 1684.660 ;
        RECT 1341.430 1684.460 1344.510 1684.600 ;
        RECT 1341.430 1684.400 1341.750 1684.460 ;
        RECT 1344.190 1684.400 1344.510 1684.460 ;
        RECT 1344.190 32.540 1344.510 32.600 ;
        RECT 1863.990 32.540 1864.310 32.600 ;
        RECT 1344.190 32.400 1864.310 32.540 ;
        RECT 1344.190 32.340 1344.510 32.400 ;
        RECT 1863.990 32.340 1864.310 32.400 ;
      LAYER via ;
        RECT 1341.460 1684.400 1341.720 1684.660 ;
        RECT 1344.220 1684.400 1344.480 1684.660 ;
        RECT 1344.220 32.340 1344.480 32.600 ;
        RECT 1864.020 32.340 1864.280 32.600 ;
      LAYER met2 ;
        RECT 1341.360 1700.340 1341.640 1704.000 ;
        RECT 1341.360 1700.000 1341.660 1700.340 ;
        RECT 1341.520 1684.690 1341.660 1700.000 ;
        RECT 1341.460 1684.370 1341.720 1684.690 ;
        RECT 1344.220 1684.370 1344.480 1684.690 ;
        RECT 1344.280 32.630 1344.420 1684.370 ;
        RECT 1344.220 32.310 1344.480 32.630 ;
        RECT 1864.020 32.310 1864.280 32.630 ;
        RECT 1864.080 2.400 1864.220 32.310 ;
        RECT 1863.870 -4.800 1864.430 2.400 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1180.045 1686.145 1180.215 1689.375 ;
      LAYER mcon ;
        RECT 1180.045 1689.205 1180.215 1689.375 ;
      LAYER met1 ;
        RECT 1179.985 1689.360 1180.275 1689.405 ;
        RECT 1225.510 1689.360 1225.830 1689.420 ;
        RECT 1179.985 1689.220 1225.830 1689.360 ;
        RECT 1179.985 1689.175 1180.275 1689.220 ;
        RECT 1225.510 1689.160 1225.830 1689.220 ;
        RECT 1128.450 1686.300 1128.770 1686.360 ;
        RECT 1179.985 1686.300 1180.275 1686.345 ;
        RECT 1128.450 1686.160 1180.275 1686.300 ;
        RECT 1128.450 1686.100 1128.770 1686.160 ;
        RECT 1179.985 1686.115 1180.275 1686.160 ;
        RECT 744.810 65.520 745.130 65.580 ;
        RECT 1128.450 65.520 1128.770 65.580 ;
        RECT 744.810 65.380 1128.770 65.520 ;
        RECT 744.810 65.320 745.130 65.380 ;
        RECT 1128.450 65.320 1128.770 65.380 ;
      LAYER via ;
        RECT 1225.540 1689.160 1225.800 1689.420 ;
        RECT 1128.480 1686.100 1128.740 1686.360 ;
        RECT 744.840 65.320 745.100 65.580 ;
        RECT 1128.480 65.320 1128.740 65.580 ;
      LAYER met2 ;
        RECT 1225.440 1700.340 1225.720 1704.000 ;
        RECT 1225.440 1700.000 1225.740 1700.340 ;
        RECT 1225.600 1689.450 1225.740 1700.000 ;
        RECT 1225.540 1689.130 1225.800 1689.450 ;
        RECT 1128.480 1686.070 1128.740 1686.390 ;
        RECT 1128.540 65.610 1128.680 1686.070 ;
        RECT 744.840 65.290 745.100 65.610 ;
        RECT 1128.480 65.290 1128.740 65.610 ;
        RECT 744.900 16.730 745.040 65.290 ;
        RECT 740.300 16.590 745.040 16.730 ;
        RECT 740.300 2.400 740.440 16.590 ;
        RECT 740.090 -4.800 740.650 2.400 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1339.590 1684.940 1339.910 1685.000 ;
        RECT 1343.270 1684.940 1343.590 1685.000 ;
        RECT 1339.590 1684.800 1343.590 1684.940 ;
        RECT 1339.590 1684.740 1339.910 1684.800 ;
        RECT 1343.270 1684.740 1343.590 1684.800 ;
        RECT 1339.590 32.200 1339.910 32.260 ;
        RECT 1881.930 32.200 1882.250 32.260 ;
        RECT 1339.590 32.060 1882.250 32.200 ;
        RECT 1339.590 32.000 1339.910 32.060 ;
        RECT 1881.930 32.000 1882.250 32.060 ;
      LAYER via ;
        RECT 1339.620 1684.740 1339.880 1685.000 ;
        RECT 1343.300 1684.740 1343.560 1685.000 ;
        RECT 1339.620 32.000 1339.880 32.260 ;
        RECT 1881.960 32.000 1882.220 32.260 ;
      LAYER met2 ;
        RECT 1343.200 1700.340 1343.480 1704.000 ;
        RECT 1343.200 1700.000 1343.500 1700.340 ;
        RECT 1343.360 1685.030 1343.500 1700.000 ;
        RECT 1339.620 1684.710 1339.880 1685.030 ;
        RECT 1343.300 1684.710 1343.560 1685.030 ;
        RECT 1339.680 32.290 1339.820 1684.710 ;
        RECT 1339.620 31.970 1339.880 32.290 ;
        RECT 1881.960 31.970 1882.220 32.290 ;
        RECT 1882.020 2.400 1882.160 31.970 ;
        RECT 1881.810 -4.800 1882.370 2.400 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1340.050 1645.840 1340.370 1645.900 ;
        RECT 1345.110 1645.840 1345.430 1645.900 ;
        RECT 1340.050 1645.700 1345.430 1645.840 ;
        RECT 1340.050 1645.640 1340.370 1645.700 ;
        RECT 1345.110 1645.640 1345.430 1645.700 ;
        RECT 1340.970 31.860 1341.290 31.920 ;
        RECT 1899.870 31.860 1900.190 31.920 ;
        RECT 1340.970 31.720 1900.190 31.860 ;
        RECT 1340.970 31.660 1341.290 31.720 ;
        RECT 1899.870 31.660 1900.190 31.720 ;
      LAYER via ;
        RECT 1340.080 1645.640 1340.340 1645.900 ;
        RECT 1345.140 1645.640 1345.400 1645.900 ;
        RECT 1341.000 31.660 1341.260 31.920 ;
        RECT 1899.900 31.660 1900.160 31.920 ;
      LAYER met2 ;
        RECT 1345.040 1700.340 1345.320 1704.000 ;
        RECT 1345.040 1700.000 1345.340 1700.340 ;
        RECT 1345.200 1645.930 1345.340 1700.000 ;
        RECT 1340.080 1645.610 1340.340 1645.930 ;
        RECT 1345.140 1645.610 1345.400 1645.930 ;
        RECT 1340.140 1593.650 1340.280 1645.610 ;
        RECT 1340.140 1593.510 1340.740 1593.650 ;
        RECT 1340.600 47.330 1340.740 1593.510 ;
        RECT 1340.600 47.190 1341.200 47.330 ;
        RECT 1341.060 31.950 1341.200 47.190 ;
        RECT 1341.000 31.630 1341.260 31.950 ;
        RECT 1899.900 31.630 1900.160 31.950 ;
        RECT 1899.960 2.400 1900.100 31.630 ;
        RECT 1899.750 -4.800 1900.310 2.400 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1346.950 1677.120 1347.270 1677.180 ;
        RECT 1350.630 1677.120 1350.950 1677.180 ;
        RECT 1346.950 1676.980 1350.950 1677.120 ;
        RECT 1346.950 1676.920 1347.270 1676.980 ;
        RECT 1350.630 1676.920 1350.950 1676.980 ;
        RECT 1350.630 31.520 1350.950 31.580 ;
        RECT 1917.810 31.520 1918.130 31.580 ;
        RECT 1350.630 31.380 1918.130 31.520 ;
        RECT 1350.630 31.320 1350.950 31.380 ;
        RECT 1917.810 31.320 1918.130 31.380 ;
      LAYER via ;
        RECT 1346.980 1676.920 1347.240 1677.180 ;
        RECT 1350.660 1676.920 1350.920 1677.180 ;
        RECT 1350.660 31.320 1350.920 31.580 ;
        RECT 1917.840 31.320 1918.100 31.580 ;
      LAYER met2 ;
        RECT 1346.880 1700.340 1347.160 1704.000 ;
        RECT 1346.880 1700.000 1347.180 1700.340 ;
        RECT 1347.040 1677.210 1347.180 1700.000 ;
        RECT 1346.980 1676.890 1347.240 1677.210 ;
        RECT 1350.660 1676.890 1350.920 1677.210 ;
        RECT 1350.720 31.610 1350.860 1676.890 ;
        RECT 1350.660 31.290 1350.920 31.610 ;
        RECT 1917.840 31.290 1918.100 31.610 ;
        RECT 1917.900 2.400 1918.040 31.290 ;
        RECT 1917.690 -4.800 1918.250 2.400 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1347.410 1683.920 1347.730 1683.980 ;
        RECT 1348.790 1683.920 1349.110 1683.980 ;
        RECT 1347.410 1683.780 1349.110 1683.920 ;
        RECT 1347.410 1683.720 1347.730 1683.780 ;
        RECT 1348.790 1683.720 1349.110 1683.780 ;
        RECT 1347.410 31.180 1347.730 31.240 ;
        RECT 1935.290 31.180 1935.610 31.240 ;
        RECT 1347.410 31.040 1935.610 31.180 ;
        RECT 1347.410 30.980 1347.730 31.040 ;
        RECT 1935.290 30.980 1935.610 31.040 ;
      LAYER via ;
        RECT 1347.440 1683.720 1347.700 1683.980 ;
        RECT 1348.820 1683.720 1349.080 1683.980 ;
        RECT 1347.440 30.980 1347.700 31.240 ;
        RECT 1935.320 30.980 1935.580 31.240 ;
      LAYER met2 ;
        RECT 1348.720 1700.340 1349.000 1704.000 ;
        RECT 1348.720 1700.000 1349.020 1700.340 ;
        RECT 1348.880 1684.010 1349.020 1700.000 ;
        RECT 1347.440 1683.690 1347.700 1684.010 ;
        RECT 1348.820 1683.690 1349.080 1684.010 ;
        RECT 1347.500 31.270 1347.640 1683.690 ;
        RECT 1347.440 30.950 1347.700 31.270 ;
        RECT 1935.320 30.950 1935.580 31.270 ;
        RECT 1935.380 2.400 1935.520 30.950 ;
        RECT 1935.170 -4.800 1935.730 2.400 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1351.090 30.840 1351.410 30.900 ;
        RECT 1953.230 30.840 1953.550 30.900 ;
        RECT 1351.090 30.700 1953.550 30.840 ;
        RECT 1351.090 30.640 1351.410 30.700 ;
        RECT 1953.230 30.640 1953.550 30.700 ;
      LAYER via ;
        RECT 1351.120 30.640 1351.380 30.900 ;
        RECT 1953.260 30.640 1953.520 30.900 ;
      LAYER met2 ;
        RECT 1350.560 1700.340 1350.840 1704.000 ;
        RECT 1350.560 1700.000 1350.860 1700.340 ;
        RECT 1350.720 1677.970 1350.860 1700.000 ;
        RECT 1350.720 1677.830 1351.320 1677.970 ;
        RECT 1351.180 30.930 1351.320 1677.830 ;
        RECT 1351.120 30.610 1351.380 30.930 ;
        RECT 1953.260 30.610 1953.520 30.930 ;
        RECT 1953.320 2.400 1953.460 30.610 ;
        RECT 1953.110 -4.800 1953.670 2.400 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1373.245 1685.465 1373.415 1686.655 ;
        RECT 1388.425 1686.315 1388.595 1686.655 ;
        RECT 1388.425 1686.145 1390.895 1686.315 ;
        RECT 1400.845 1675.945 1401.015 1686.655 ;
      LAYER mcon ;
        RECT 1373.245 1686.485 1373.415 1686.655 ;
        RECT 1388.425 1686.485 1388.595 1686.655 ;
        RECT 1400.845 1686.485 1401.015 1686.655 ;
        RECT 1390.725 1686.145 1390.895 1686.315 ;
      LAYER met1 ;
        RECT 1373.185 1686.640 1373.475 1686.685 ;
        RECT 1388.365 1686.640 1388.655 1686.685 ;
        RECT 1400.785 1686.640 1401.075 1686.685 ;
        RECT 1373.185 1686.500 1388.655 1686.640 ;
        RECT 1373.185 1686.455 1373.475 1686.500 ;
        RECT 1388.365 1686.455 1388.655 1686.500 ;
        RECT 1393.500 1686.500 1401.075 1686.640 ;
        RECT 1390.665 1686.300 1390.955 1686.345 ;
        RECT 1393.500 1686.300 1393.640 1686.500 ;
        RECT 1400.785 1686.455 1401.075 1686.500 ;
        RECT 1390.665 1686.160 1393.640 1686.300 ;
        RECT 1390.665 1686.115 1390.955 1686.160 ;
        RECT 1352.470 1685.620 1352.790 1685.680 ;
        RECT 1373.185 1685.620 1373.475 1685.665 ;
        RECT 1352.470 1685.480 1373.475 1685.620 ;
        RECT 1352.470 1685.420 1352.790 1685.480 ;
        RECT 1373.185 1685.435 1373.475 1685.480 ;
        RECT 1400.770 1676.100 1401.090 1676.160 ;
        RECT 1400.575 1675.960 1401.090 1676.100 ;
        RECT 1400.770 1675.900 1401.090 1675.960 ;
        RECT 1400.770 1646.520 1401.090 1646.580 ;
        RECT 1966.570 1646.520 1966.890 1646.580 ;
        RECT 1400.770 1646.380 1966.890 1646.520 ;
        RECT 1400.770 1646.320 1401.090 1646.380 ;
        RECT 1966.570 1646.320 1966.890 1646.380 ;
      LAYER via ;
        RECT 1352.500 1685.420 1352.760 1685.680 ;
        RECT 1400.800 1675.900 1401.060 1676.160 ;
        RECT 1400.800 1646.320 1401.060 1646.580 ;
        RECT 1966.600 1646.320 1966.860 1646.580 ;
      LAYER met2 ;
        RECT 1352.400 1700.340 1352.680 1704.000 ;
        RECT 1352.400 1700.000 1352.700 1700.340 ;
        RECT 1352.560 1685.710 1352.700 1700.000 ;
        RECT 1352.500 1685.390 1352.760 1685.710 ;
        RECT 1400.800 1675.870 1401.060 1676.190 ;
        RECT 1400.860 1646.610 1401.000 1675.870 ;
        RECT 1400.800 1646.290 1401.060 1646.610 ;
        RECT 1966.600 1646.290 1966.860 1646.610 ;
        RECT 1966.660 17.410 1966.800 1646.290 ;
        RECT 1966.660 17.270 1971.400 17.410 ;
        RECT 1971.260 2.400 1971.400 17.270 ;
        RECT 1971.050 -4.800 1971.610 2.400 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1416.945 1660.305 1417.115 1662.175 ;
      LAYER mcon ;
        RECT 1416.945 1662.005 1417.115 1662.175 ;
      LAYER met1 ;
        RECT 1393.870 1662.160 1394.190 1662.220 ;
        RECT 1416.885 1662.160 1417.175 1662.205 ;
        RECT 1393.870 1662.020 1417.175 1662.160 ;
        RECT 1393.870 1661.960 1394.190 1662.020 ;
        RECT 1416.885 1661.975 1417.175 1662.020 ;
        RECT 1416.885 1660.460 1417.175 1660.505 ;
        RECT 1987.270 1660.460 1987.590 1660.520 ;
        RECT 1416.885 1660.320 1987.590 1660.460 ;
        RECT 1416.885 1660.275 1417.175 1660.320 ;
        RECT 1987.270 1660.260 1987.590 1660.320 ;
      LAYER via ;
        RECT 1393.900 1661.960 1394.160 1662.220 ;
        RECT 1987.300 1660.260 1987.560 1660.520 ;
      LAYER met2 ;
        RECT 1354.240 1700.340 1354.520 1704.000 ;
        RECT 1354.240 1700.000 1354.540 1700.340 ;
        RECT 1354.400 1687.605 1354.540 1700.000 ;
        RECT 1354.330 1687.235 1354.610 1687.605 ;
        RECT 1393.430 1687.235 1393.710 1687.605 ;
        RECT 1393.500 1675.930 1393.640 1687.235 ;
        RECT 1393.500 1675.790 1394.100 1675.930 ;
        RECT 1393.960 1662.250 1394.100 1675.790 ;
        RECT 1393.900 1661.930 1394.160 1662.250 ;
        RECT 1987.300 1660.230 1987.560 1660.550 ;
        RECT 1987.360 17.410 1987.500 1660.230 ;
        RECT 1987.360 17.270 1989.340 17.410 ;
        RECT 1989.200 2.400 1989.340 17.270 ;
        RECT 1988.990 -4.800 1989.550 2.400 ;
      LAYER via2 ;
        RECT 1354.330 1687.280 1354.610 1687.560 ;
        RECT 1393.430 1687.280 1393.710 1687.560 ;
      LAYER met3 ;
        RECT 1354.305 1687.570 1354.635 1687.585 ;
        RECT 1393.405 1687.570 1393.735 1687.585 ;
        RECT 1354.305 1687.270 1393.735 1687.570 ;
        RECT 1354.305 1687.255 1354.635 1687.270 ;
        RECT 1393.405 1687.255 1393.735 1687.270 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1387.505 1684.105 1387.675 1686.315 ;
        RECT 1415.105 1683.425 1415.275 1684.275 ;
      LAYER mcon ;
        RECT 1387.505 1686.145 1387.675 1686.315 ;
        RECT 1415.105 1684.105 1415.275 1684.275 ;
      LAYER met1 ;
        RECT 1356.150 1686.300 1356.470 1686.360 ;
        RECT 1387.445 1686.300 1387.735 1686.345 ;
        RECT 1356.150 1686.160 1387.735 1686.300 ;
        RECT 1356.150 1686.100 1356.470 1686.160 ;
        RECT 1387.445 1686.115 1387.735 1686.160 ;
        RECT 1387.445 1684.260 1387.735 1684.305 ;
        RECT 1415.045 1684.260 1415.335 1684.305 ;
        RECT 1387.445 1684.120 1415.335 1684.260 ;
        RECT 1387.445 1684.075 1387.735 1684.120 ;
        RECT 1415.045 1684.075 1415.335 1684.120 ;
        RECT 1415.045 1683.580 1415.335 1683.625 ;
        RECT 1416.410 1683.580 1416.730 1683.640 ;
        RECT 1415.045 1683.440 1416.730 1683.580 ;
        RECT 1415.045 1683.395 1415.335 1683.440 ;
        RECT 1416.410 1683.380 1416.730 1683.440 ;
        RECT 1416.410 1640.060 1416.730 1640.120 ;
        RECT 2001.530 1640.060 2001.850 1640.120 ;
        RECT 1416.410 1639.920 2001.850 1640.060 ;
        RECT 1416.410 1639.860 1416.730 1639.920 ;
        RECT 2001.530 1639.860 2001.850 1639.920 ;
      LAYER via ;
        RECT 1356.180 1686.100 1356.440 1686.360 ;
        RECT 1416.440 1683.380 1416.700 1683.640 ;
        RECT 1416.440 1639.860 1416.700 1640.120 ;
        RECT 2001.560 1639.860 2001.820 1640.120 ;
      LAYER met2 ;
        RECT 1356.080 1700.340 1356.360 1704.000 ;
        RECT 1356.080 1700.000 1356.380 1700.340 ;
        RECT 1356.240 1686.390 1356.380 1700.000 ;
        RECT 1356.180 1686.070 1356.440 1686.390 ;
        RECT 1416.440 1683.350 1416.700 1683.670 ;
        RECT 1416.500 1640.150 1416.640 1683.350 ;
        RECT 1416.440 1639.830 1416.700 1640.150 ;
        RECT 2001.560 1639.830 2001.820 1640.150 ;
        RECT 2001.620 17.410 2001.760 1639.830 ;
        RECT 2001.620 17.270 2006.820 17.410 ;
        RECT 2006.680 2.400 2006.820 17.270 ;
        RECT 2006.470 -4.800 2007.030 2.400 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1357.990 1667.260 1358.310 1667.320 ;
        RECT 2021.770 1667.260 2022.090 1667.320 ;
        RECT 1357.990 1667.120 2022.090 1667.260 ;
        RECT 1357.990 1667.060 1358.310 1667.120 ;
        RECT 2021.770 1667.060 2022.090 1667.120 ;
      LAYER via ;
        RECT 1358.020 1667.060 1358.280 1667.320 ;
        RECT 2021.800 1667.060 2022.060 1667.320 ;
      LAYER met2 ;
        RECT 1357.920 1700.340 1358.200 1704.000 ;
        RECT 1357.920 1700.000 1358.220 1700.340 ;
        RECT 1358.080 1667.350 1358.220 1700.000 ;
        RECT 1358.020 1667.030 1358.280 1667.350 ;
        RECT 2021.800 1667.030 2022.060 1667.350 ;
        RECT 2021.860 17.410 2022.000 1667.030 ;
        RECT 2021.860 17.270 2024.760 17.410 ;
        RECT 2024.620 2.400 2024.760 17.270 ;
        RECT 2024.410 -4.800 2024.970 2.400 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1402.225 1676.285 1402.395 1689.375 ;
      LAYER mcon ;
        RECT 1402.225 1689.205 1402.395 1689.375 ;
      LAYER met1 ;
        RECT 1359.830 1689.700 1360.150 1689.760 ;
        RECT 1359.830 1689.560 1390.420 1689.700 ;
        RECT 1359.830 1689.500 1360.150 1689.560 ;
        RECT 1390.280 1689.360 1390.420 1689.560 ;
        RECT 1402.165 1689.360 1402.455 1689.405 ;
        RECT 1390.280 1689.220 1402.455 1689.360 ;
        RECT 1402.165 1689.175 1402.455 1689.220 ;
        RECT 1402.150 1676.440 1402.470 1676.500 ;
        RECT 1401.955 1676.300 1402.470 1676.440 ;
        RECT 1402.150 1676.240 1402.470 1676.300 ;
        RECT 1402.150 1632.920 1402.470 1632.980 ;
        RECT 2042.470 1632.920 2042.790 1632.980 ;
        RECT 1402.150 1632.780 2042.790 1632.920 ;
        RECT 1402.150 1632.720 1402.470 1632.780 ;
        RECT 2042.470 1632.720 2042.790 1632.780 ;
      LAYER via ;
        RECT 1359.860 1689.500 1360.120 1689.760 ;
        RECT 1402.180 1676.240 1402.440 1676.500 ;
        RECT 1402.180 1632.720 1402.440 1632.980 ;
        RECT 2042.500 1632.720 2042.760 1632.980 ;
      LAYER met2 ;
        RECT 1359.760 1700.340 1360.040 1704.000 ;
        RECT 1359.760 1700.000 1360.060 1700.340 ;
        RECT 1359.920 1689.790 1360.060 1700.000 ;
        RECT 1359.860 1689.470 1360.120 1689.790 ;
        RECT 1402.180 1676.210 1402.440 1676.530 ;
        RECT 1402.240 1633.010 1402.380 1676.210 ;
        RECT 1402.180 1632.690 1402.440 1633.010 ;
        RECT 2042.500 1632.690 2042.760 1633.010 ;
        RECT 2042.560 2.400 2042.700 1632.690 ;
        RECT 2042.350 -4.800 2042.910 2.400 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1223.670 1659.440 1223.990 1659.500 ;
        RECT 1227.350 1659.440 1227.670 1659.500 ;
        RECT 1223.670 1659.300 1227.670 1659.440 ;
        RECT 1223.670 1659.240 1223.990 1659.300 ;
        RECT 1227.350 1659.240 1227.670 1659.300 ;
        RECT 758.610 1646.180 758.930 1646.240 ;
        RECT 1223.670 1646.180 1223.990 1646.240 ;
        RECT 758.610 1646.040 1223.990 1646.180 ;
        RECT 758.610 1645.980 758.930 1646.040 ;
        RECT 1223.670 1645.980 1223.990 1646.040 ;
      LAYER via ;
        RECT 1223.700 1659.240 1223.960 1659.500 ;
        RECT 1227.380 1659.240 1227.640 1659.500 ;
        RECT 758.640 1645.980 758.900 1646.240 ;
        RECT 1223.700 1645.980 1223.960 1646.240 ;
      LAYER met2 ;
        RECT 1227.280 1700.340 1227.560 1704.000 ;
        RECT 1227.280 1700.000 1227.580 1700.340 ;
        RECT 1227.440 1659.530 1227.580 1700.000 ;
        RECT 1223.700 1659.210 1223.960 1659.530 ;
        RECT 1227.380 1659.210 1227.640 1659.530 ;
        RECT 1223.760 1646.270 1223.900 1659.210 ;
        RECT 758.640 1645.950 758.900 1646.270 ;
        RECT 1223.700 1645.950 1223.960 1646.270 ;
        RECT 758.700 17.410 758.840 1645.950 ;
        RECT 757.780 17.270 758.840 17.410 ;
        RECT 757.780 2.400 757.920 17.270 ;
        RECT 757.570 -4.800 758.130 2.400 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1361.670 1685.280 1361.990 1685.340 ;
        RECT 1365.350 1685.280 1365.670 1685.340 ;
        RECT 1361.670 1685.140 1365.670 1685.280 ;
        RECT 1361.670 1685.080 1361.990 1685.140 ;
        RECT 1365.350 1685.080 1365.670 1685.140 ;
        RECT 1365.350 1653.660 1365.670 1653.720 ;
        RECT 2056.270 1653.660 2056.590 1653.720 ;
        RECT 1365.350 1653.520 2056.590 1653.660 ;
        RECT 1365.350 1653.460 1365.670 1653.520 ;
        RECT 2056.270 1653.460 2056.590 1653.520 ;
      LAYER via ;
        RECT 1361.700 1685.080 1361.960 1685.340 ;
        RECT 1365.380 1685.080 1365.640 1685.340 ;
        RECT 1365.380 1653.460 1365.640 1653.720 ;
        RECT 2056.300 1653.460 2056.560 1653.720 ;
      LAYER met2 ;
        RECT 1361.600 1700.340 1361.880 1704.000 ;
        RECT 1361.600 1700.000 1361.900 1700.340 ;
        RECT 1361.760 1685.370 1361.900 1700.000 ;
        RECT 1361.700 1685.050 1361.960 1685.370 ;
        RECT 1365.380 1685.050 1365.640 1685.370 ;
        RECT 1365.440 1653.750 1365.580 1685.050 ;
        RECT 1365.380 1653.430 1365.640 1653.750 ;
        RECT 2056.300 1653.430 2056.560 1653.750 ;
        RECT 2056.360 17.410 2056.500 1653.430 ;
        RECT 2056.360 17.270 2060.640 17.410 ;
        RECT 2060.500 2.400 2060.640 17.270 ;
        RECT 2060.290 -4.800 2060.850 2.400 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1361.670 1684.600 1361.990 1684.660 ;
        RECT 1363.510 1684.600 1363.830 1684.660 ;
        RECT 1361.670 1684.460 1363.830 1684.600 ;
        RECT 1361.670 1684.400 1361.990 1684.460 ;
        RECT 1363.510 1684.400 1363.830 1684.460 ;
        RECT 1361.670 1646.180 1361.990 1646.240 ;
        RECT 2076.970 1646.180 2077.290 1646.240 ;
        RECT 1361.670 1646.040 2077.290 1646.180 ;
        RECT 1361.670 1645.980 1361.990 1646.040 ;
        RECT 2076.970 1645.980 2077.290 1646.040 ;
      LAYER via ;
        RECT 1361.700 1684.400 1361.960 1684.660 ;
        RECT 1363.540 1684.400 1363.800 1684.660 ;
        RECT 1361.700 1645.980 1361.960 1646.240 ;
        RECT 2077.000 1645.980 2077.260 1646.240 ;
      LAYER met2 ;
        RECT 1363.440 1700.340 1363.720 1704.000 ;
        RECT 1363.440 1700.000 1363.740 1700.340 ;
        RECT 1363.600 1684.690 1363.740 1700.000 ;
        RECT 1361.700 1684.370 1361.960 1684.690 ;
        RECT 1363.540 1684.370 1363.800 1684.690 ;
        RECT 1361.760 1646.270 1361.900 1684.370 ;
        RECT 1361.700 1645.950 1361.960 1646.270 ;
        RECT 2077.000 1645.950 2077.260 1646.270 ;
        RECT 2077.060 17.410 2077.200 1645.950 ;
        RECT 2077.060 17.270 2078.580 17.410 ;
        RECT 2078.440 2.400 2078.580 17.270 ;
        RECT 2078.230 -4.800 2078.790 2.400 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1362.590 1685.960 1362.910 1686.020 ;
        RECT 1365.350 1685.960 1365.670 1686.020 ;
        RECT 1362.590 1685.820 1365.670 1685.960 ;
        RECT 1362.590 1685.760 1362.910 1685.820 ;
        RECT 1365.350 1685.760 1365.670 1685.820 ;
        RECT 1360.750 1677.460 1361.070 1677.520 ;
        RECT 1362.590 1677.460 1362.910 1677.520 ;
        RECT 1360.750 1677.320 1362.910 1677.460 ;
        RECT 1360.750 1677.260 1361.070 1677.320 ;
        RECT 1362.590 1677.260 1362.910 1677.320 ;
        RECT 1360.750 1605.380 1361.070 1605.440 ;
        RECT 2090.770 1605.380 2091.090 1605.440 ;
        RECT 1360.750 1605.240 2091.090 1605.380 ;
        RECT 1360.750 1605.180 1361.070 1605.240 ;
        RECT 2090.770 1605.180 2091.090 1605.240 ;
      LAYER via ;
        RECT 1362.620 1685.760 1362.880 1686.020 ;
        RECT 1365.380 1685.760 1365.640 1686.020 ;
        RECT 1360.780 1677.260 1361.040 1677.520 ;
        RECT 1362.620 1677.260 1362.880 1677.520 ;
        RECT 1360.780 1605.180 1361.040 1605.440 ;
        RECT 2090.800 1605.180 2091.060 1605.440 ;
      LAYER met2 ;
        RECT 1365.280 1700.340 1365.560 1704.000 ;
        RECT 1365.280 1700.000 1365.580 1700.340 ;
        RECT 1365.440 1686.050 1365.580 1700.000 ;
        RECT 1362.620 1685.730 1362.880 1686.050 ;
        RECT 1365.380 1685.730 1365.640 1686.050 ;
        RECT 1362.680 1677.550 1362.820 1685.730 ;
        RECT 1360.780 1677.230 1361.040 1677.550 ;
        RECT 1362.620 1677.230 1362.880 1677.550 ;
        RECT 1360.840 1605.470 1360.980 1677.230 ;
        RECT 1360.780 1605.150 1361.040 1605.470 ;
        RECT 2090.800 1605.150 2091.060 1605.470 ;
        RECT 2090.860 17.410 2091.000 1605.150 ;
        RECT 2090.860 17.270 2096.060 17.410 ;
        RECT 2095.920 2.400 2096.060 17.270 ;
        RECT 2095.710 -4.800 2096.270 2.400 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1367.190 1686.640 1367.510 1686.700 ;
        RECT 1372.710 1686.640 1373.030 1686.700 ;
        RECT 1367.190 1686.500 1373.030 1686.640 ;
        RECT 1367.190 1686.440 1367.510 1686.500 ;
        RECT 1372.710 1686.440 1373.030 1686.500 ;
        RECT 1372.710 1674.060 1373.030 1674.120 ;
        RECT 2111.470 1674.060 2111.790 1674.120 ;
        RECT 1372.710 1673.920 2111.790 1674.060 ;
        RECT 1372.710 1673.860 1373.030 1673.920 ;
        RECT 2111.470 1673.860 2111.790 1673.920 ;
      LAYER via ;
        RECT 1367.220 1686.440 1367.480 1686.700 ;
        RECT 1372.740 1686.440 1373.000 1686.700 ;
        RECT 1372.740 1673.860 1373.000 1674.120 ;
        RECT 2111.500 1673.860 2111.760 1674.120 ;
      LAYER met2 ;
        RECT 1367.120 1700.340 1367.400 1704.000 ;
        RECT 1367.120 1700.000 1367.420 1700.340 ;
        RECT 1367.280 1686.730 1367.420 1700.000 ;
        RECT 1367.220 1686.410 1367.480 1686.730 ;
        RECT 1372.740 1686.410 1373.000 1686.730 ;
        RECT 1372.800 1674.150 1372.940 1686.410 ;
        RECT 1372.740 1673.830 1373.000 1674.150 ;
        RECT 2111.500 1673.830 2111.760 1674.150 ;
        RECT 2111.560 17.410 2111.700 1673.830 ;
        RECT 2111.560 17.270 2114.000 17.410 ;
        RECT 2113.860 2.400 2114.000 17.270 ;
        RECT 2113.650 -4.800 2114.210 2.400 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1366.730 1684.260 1367.050 1684.320 ;
        RECT 1369.030 1684.260 1369.350 1684.320 ;
        RECT 1366.730 1684.120 1369.350 1684.260 ;
        RECT 1366.730 1684.060 1367.050 1684.120 ;
        RECT 1369.030 1684.060 1369.350 1684.120 ;
        RECT 1366.730 1639.720 1367.050 1639.780 ;
        RECT 2125.730 1639.720 2126.050 1639.780 ;
        RECT 1366.730 1639.580 2126.050 1639.720 ;
        RECT 1366.730 1639.520 1367.050 1639.580 ;
        RECT 2125.730 1639.520 2126.050 1639.580 ;
        RECT 2125.730 14.520 2126.050 14.580 ;
        RECT 2131.710 14.520 2132.030 14.580 ;
        RECT 2125.730 14.380 2132.030 14.520 ;
        RECT 2125.730 14.320 2126.050 14.380 ;
        RECT 2131.710 14.320 2132.030 14.380 ;
      LAYER via ;
        RECT 1366.760 1684.060 1367.020 1684.320 ;
        RECT 1369.060 1684.060 1369.320 1684.320 ;
        RECT 1366.760 1639.520 1367.020 1639.780 ;
        RECT 2125.760 1639.520 2126.020 1639.780 ;
        RECT 2125.760 14.320 2126.020 14.580 ;
        RECT 2131.740 14.320 2132.000 14.580 ;
      LAYER met2 ;
        RECT 1368.960 1700.340 1369.240 1704.000 ;
        RECT 1368.960 1700.000 1369.260 1700.340 ;
        RECT 1369.120 1684.350 1369.260 1700.000 ;
        RECT 1366.760 1684.030 1367.020 1684.350 ;
        RECT 1369.060 1684.030 1369.320 1684.350 ;
        RECT 1366.820 1639.810 1366.960 1684.030 ;
        RECT 1366.760 1639.490 1367.020 1639.810 ;
        RECT 2125.760 1639.490 2126.020 1639.810 ;
        RECT 2125.820 14.610 2125.960 1639.490 ;
        RECT 2125.760 14.290 2126.020 14.610 ;
        RECT 2131.740 14.290 2132.000 14.610 ;
        RECT 2131.800 2.400 2131.940 14.290 ;
        RECT 2131.590 -4.800 2132.150 2.400 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1368.110 1683.920 1368.430 1683.980 ;
        RECT 1370.870 1683.920 1371.190 1683.980 ;
        RECT 1368.110 1683.780 1371.190 1683.920 ;
        RECT 1368.110 1683.720 1368.430 1683.780 ;
        RECT 1370.870 1683.720 1371.190 1683.780 ;
        RECT 1368.110 1625.440 1368.430 1625.500 ;
        RECT 2145.970 1625.440 2146.290 1625.500 ;
        RECT 1368.110 1625.300 2146.290 1625.440 ;
        RECT 1368.110 1625.240 1368.430 1625.300 ;
        RECT 2145.970 1625.240 2146.290 1625.300 ;
      LAYER via ;
        RECT 1368.140 1683.720 1368.400 1683.980 ;
        RECT 1370.900 1683.720 1371.160 1683.980 ;
        RECT 1368.140 1625.240 1368.400 1625.500 ;
        RECT 2146.000 1625.240 2146.260 1625.500 ;
      LAYER met2 ;
        RECT 1370.800 1700.340 1371.080 1704.000 ;
        RECT 1370.800 1700.000 1371.100 1700.340 ;
        RECT 1370.960 1684.010 1371.100 1700.000 ;
        RECT 1368.140 1683.690 1368.400 1684.010 ;
        RECT 1370.900 1683.690 1371.160 1684.010 ;
        RECT 1368.200 1625.530 1368.340 1683.690 ;
        RECT 1368.140 1625.210 1368.400 1625.530 ;
        RECT 2146.000 1625.210 2146.260 1625.530 ;
        RECT 2146.060 17.410 2146.200 1625.210 ;
        RECT 2146.060 17.270 2149.880 17.410 ;
        RECT 2149.740 2.400 2149.880 17.270 ;
        RECT 2149.530 -4.800 2150.090 2.400 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1369.490 1689.020 1369.810 1689.080 ;
        RECT 1372.710 1689.020 1373.030 1689.080 ;
        RECT 1369.490 1688.880 1373.030 1689.020 ;
        RECT 1369.490 1688.820 1369.810 1688.880 ;
        RECT 1372.710 1688.820 1373.030 1688.880 ;
        RECT 1369.490 1660.120 1369.810 1660.180 ;
        RECT 2166.670 1660.120 2166.990 1660.180 ;
        RECT 1369.490 1659.980 2166.990 1660.120 ;
        RECT 1369.490 1659.920 1369.810 1659.980 ;
        RECT 2166.670 1659.920 2166.990 1659.980 ;
      LAYER via ;
        RECT 1369.520 1688.820 1369.780 1689.080 ;
        RECT 1372.740 1688.820 1373.000 1689.080 ;
        RECT 1369.520 1659.920 1369.780 1660.180 ;
        RECT 2166.700 1659.920 2166.960 1660.180 ;
      LAYER met2 ;
        RECT 1372.640 1700.340 1372.920 1704.000 ;
        RECT 1372.640 1700.000 1372.940 1700.340 ;
        RECT 1372.800 1689.110 1372.940 1700.000 ;
        RECT 1369.520 1688.790 1369.780 1689.110 ;
        RECT 1372.740 1688.790 1373.000 1689.110 ;
        RECT 1369.580 1660.210 1369.720 1688.790 ;
        RECT 1369.520 1659.890 1369.780 1660.210 ;
        RECT 2166.700 1659.890 2166.960 1660.210 ;
        RECT 2166.760 17.410 2166.900 1659.890 ;
        RECT 2166.760 17.270 2167.820 17.410 ;
        RECT 2167.680 2.400 2167.820 17.270 ;
        RECT 2167.470 -4.800 2168.030 2.400 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1394.865 1675.605 1395.035 1686.315 ;
      LAYER mcon ;
        RECT 1394.865 1686.145 1395.035 1686.315 ;
      LAYER met1 ;
        RECT 1374.550 1690.380 1374.870 1690.440 ;
        RECT 1393.870 1690.380 1394.190 1690.440 ;
        RECT 1374.550 1690.240 1394.190 1690.380 ;
        RECT 1374.550 1690.180 1374.870 1690.240 ;
        RECT 1393.870 1690.180 1394.190 1690.240 ;
        RECT 1393.870 1686.300 1394.190 1686.360 ;
        RECT 1394.805 1686.300 1395.095 1686.345 ;
        RECT 1393.870 1686.160 1395.095 1686.300 ;
        RECT 1393.870 1686.100 1394.190 1686.160 ;
        RECT 1394.805 1686.115 1395.095 1686.160 ;
        RECT 1394.790 1675.760 1395.110 1675.820 ;
        RECT 1394.595 1675.620 1395.110 1675.760 ;
        RECT 1394.790 1675.560 1395.110 1675.620 ;
        RECT 1394.790 1618.640 1395.110 1618.700 ;
        RECT 2180.470 1618.640 2180.790 1618.700 ;
        RECT 1394.790 1618.500 2180.790 1618.640 ;
        RECT 1394.790 1618.440 1395.110 1618.500 ;
        RECT 2180.470 1618.440 2180.790 1618.500 ;
      LAYER via ;
        RECT 1374.580 1690.180 1374.840 1690.440 ;
        RECT 1393.900 1690.180 1394.160 1690.440 ;
        RECT 1393.900 1686.100 1394.160 1686.360 ;
        RECT 1394.820 1675.560 1395.080 1675.820 ;
        RECT 1394.820 1618.440 1395.080 1618.700 ;
        RECT 2180.500 1618.440 2180.760 1618.700 ;
      LAYER met2 ;
        RECT 1374.480 1700.340 1374.760 1704.000 ;
        RECT 1374.480 1700.000 1374.780 1700.340 ;
        RECT 1374.640 1690.470 1374.780 1700.000 ;
        RECT 1374.580 1690.150 1374.840 1690.470 ;
        RECT 1393.900 1690.150 1394.160 1690.470 ;
        RECT 1393.960 1686.390 1394.100 1690.150 ;
        RECT 1393.900 1686.070 1394.160 1686.390 ;
        RECT 1394.820 1675.530 1395.080 1675.850 ;
        RECT 1394.880 1618.730 1395.020 1675.530 ;
        RECT 1394.820 1618.410 1395.080 1618.730 ;
        RECT 2180.500 1618.410 2180.760 1618.730 ;
        RECT 2180.560 17.410 2180.700 1618.410 ;
        RECT 2180.560 17.270 2185.300 17.410 ;
        RECT 2185.160 2.400 2185.300 17.270 ;
        RECT 2184.950 -4.800 2185.510 2.400 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1376.390 1681.200 1376.710 1681.260 ;
        RECT 2201.170 1681.200 2201.490 1681.260 ;
        RECT 1376.390 1681.060 2201.490 1681.200 ;
        RECT 1376.390 1681.000 1376.710 1681.060 ;
        RECT 2201.170 1681.000 2201.490 1681.060 ;
      LAYER via ;
        RECT 1376.420 1681.000 1376.680 1681.260 ;
        RECT 2201.200 1681.000 2201.460 1681.260 ;
      LAYER met2 ;
        RECT 1376.320 1700.340 1376.600 1704.000 ;
        RECT 1376.320 1700.000 1376.620 1700.340 ;
        RECT 1376.480 1681.290 1376.620 1700.000 ;
        RECT 1376.420 1680.970 1376.680 1681.290 ;
        RECT 2201.200 1680.970 2201.460 1681.290 ;
        RECT 2201.260 17.410 2201.400 1680.970 ;
        RECT 2201.260 17.270 2203.240 17.410 ;
        RECT 2203.100 2.400 2203.240 17.270 ;
        RECT 2202.890 -4.800 2203.450 2.400 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1373.630 1685.280 1373.950 1685.340 ;
        RECT 1378.230 1685.280 1378.550 1685.340 ;
        RECT 1373.630 1685.140 1378.550 1685.280 ;
        RECT 1373.630 1685.080 1373.950 1685.140 ;
        RECT 1378.230 1685.080 1378.550 1685.140 ;
        RECT 1373.630 1632.920 1373.950 1632.980 ;
        RECT 1373.630 1632.780 1399.160 1632.920 ;
        RECT 1373.630 1632.720 1373.950 1632.780 ;
        RECT 1399.020 1632.240 1399.160 1632.780 ;
        RECT 2215.430 1632.240 2215.750 1632.300 ;
        RECT 1399.020 1632.100 2215.750 1632.240 ;
        RECT 2215.430 1632.040 2215.750 1632.100 ;
      LAYER via ;
        RECT 1373.660 1685.080 1373.920 1685.340 ;
        RECT 1378.260 1685.080 1378.520 1685.340 ;
        RECT 1373.660 1632.720 1373.920 1632.980 ;
        RECT 2215.460 1632.040 2215.720 1632.300 ;
      LAYER met2 ;
        RECT 1378.160 1700.340 1378.440 1704.000 ;
        RECT 1378.160 1700.000 1378.460 1700.340 ;
        RECT 1378.320 1685.370 1378.460 1700.000 ;
        RECT 1373.660 1685.050 1373.920 1685.370 ;
        RECT 1378.260 1685.050 1378.520 1685.370 ;
        RECT 1373.720 1633.010 1373.860 1685.050 ;
        RECT 1373.660 1632.690 1373.920 1633.010 ;
        RECT 2215.460 1632.010 2215.720 1632.330 ;
        RECT 2215.520 17.410 2215.660 1632.010 ;
        RECT 2215.520 17.270 2221.180 17.410 ;
        RECT 2221.040 2.400 2221.180 17.270 ;
        RECT 2220.830 -4.800 2221.390 2.400 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1226.430 1683.920 1226.750 1683.980 ;
        RECT 1229.190 1683.920 1229.510 1683.980 ;
        RECT 1226.430 1683.780 1229.510 1683.920 ;
        RECT 1226.430 1683.720 1226.750 1683.780 ;
        RECT 1229.190 1683.720 1229.510 1683.780 ;
        RECT 779.310 1667.260 779.630 1667.320 ;
        RECT 1226.430 1667.260 1226.750 1667.320 ;
        RECT 779.310 1667.120 1226.750 1667.260 ;
        RECT 779.310 1667.060 779.630 1667.120 ;
        RECT 1226.430 1667.060 1226.750 1667.120 ;
      LAYER via ;
        RECT 1226.460 1683.720 1226.720 1683.980 ;
        RECT 1229.220 1683.720 1229.480 1683.980 ;
        RECT 779.340 1667.060 779.600 1667.320 ;
        RECT 1226.460 1667.060 1226.720 1667.320 ;
      LAYER met2 ;
        RECT 1229.120 1700.340 1229.400 1704.000 ;
        RECT 1229.120 1700.000 1229.420 1700.340 ;
        RECT 1229.280 1684.010 1229.420 1700.000 ;
        RECT 1226.460 1683.690 1226.720 1684.010 ;
        RECT 1229.220 1683.690 1229.480 1684.010 ;
        RECT 1226.520 1667.350 1226.660 1683.690 ;
        RECT 779.340 1667.030 779.600 1667.350 ;
        RECT 1226.460 1667.030 1226.720 1667.350 ;
        RECT 779.400 18.090 779.540 1667.030 ;
        RECT 775.720 17.950 779.540 18.090 ;
        RECT 775.720 2.400 775.860 17.950 ;
        RECT 775.510 -4.800 776.070 2.400 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1414.185 1685.125 1414.355 1689.035 ;
      LAYER mcon ;
        RECT 1414.185 1688.865 1414.355 1689.035 ;
      LAYER met1 ;
        RECT 1380.070 1689.020 1380.390 1689.080 ;
        RECT 1414.125 1689.020 1414.415 1689.065 ;
        RECT 1380.070 1688.880 1414.415 1689.020 ;
        RECT 1380.070 1688.820 1380.390 1688.880 ;
        RECT 1414.125 1688.835 1414.415 1688.880 ;
        RECT 1414.125 1685.280 1414.415 1685.325 ;
        RECT 1417.330 1685.280 1417.650 1685.340 ;
        RECT 1414.125 1685.140 1417.650 1685.280 ;
        RECT 1414.125 1685.095 1414.415 1685.140 ;
        RECT 1417.330 1685.080 1417.650 1685.140 ;
        RECT 1417.330 1597.900 1417.650 1597.960 ;
        RECT 2235.670 1597.900 2235.990 1597.960 ;
        RECT 1417.330 1597.760 2235.990 1597.900 ;
        RECT 1417.330 1597.700 1417.650 1597.760 ;
        RECT 2235.670 1597.700 2235.990 1597.760 ;
      LAYER via ;
        RECT 1380.100 1688.820 1380.360 1689.080 ;
        RECT 1417.360 1685.080 1417.620 1685.340 ;
        RECT 1417.360 1597.700 1417.620 1597.960 ;
        RECT 2235.700 1597.700 2235.960 1597.960 ;
      LAYER met2 ;
        RECT 1380.000 1700.340 1380.280 1704.000 ;
        RECT 1380.000 1700.000 1380.300 1700.340 ;
        RECT 1380.160 1689.110 1380.300 1700.000 ;
        RECT 1380.100 1688.790 1380.360 1689.110 ;
        RECT 1417.360 1685.050 1417.620 1685.370 ;
        RECT 1417.420 1597.990 1417.560 1685.050 ;
        RECT 1417.360 1597.670 1417.620 1597.990 ;
        RECT 2235.700 1597.670 2235.960 1597.990 ;
        RECT 2235.760 17.410 2235.900 1597.670 ;
        RECT 2235.760 17.270 2239.120 17.410 ;
        RECT 2238.980 2.400 2239.120 17.270 ;
        RECT 2238.770 -4.800 2239.330 2.400 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1381.910 1683.920 1382.230 1683.980 ;
        RECT 1383.290 1683.920 1383.610 1683.980 ;
        RECT 1381.910 1683.780 1383.610 1683.920 ;
        RECT 1381.910 1683.720 1382.230 1683.780 ;
        RECT 1383.290 1683.720 1383.610 1683.780 ;
        RECT 1383.290 1653.320 1383.610 1653.380 ;
        RECT 2256.370 1653.320 2256.690 1653.380 ;
        RECT 1383.290 1653.180 2256.690 1653.320 ;
        RECT 1383.290 1653.120 1383.610 1653.180 ;
        RECT 2256.370 1653.120 2256.690 1653.180 ;
      LAYER via ;
        RECT 1381.940 1683.720 1382.200 1683.980 ;
        RECT 1383.320 1683.720 1383.580 1683.980 ;
        RECT 1383.320 1653.120 1383.580 1653.380 ;
        RECT 2256.400 1653.120 2256.660 1653.380 ;
      LAYER met2 ;
        RECT 1381.840 1700.340 1382.120 1704.000 ;
        RECT 1381.840 1700.000 1382.140 1700.340 ;
        RECT 1382.000 1684.010 1382.140 1700.000 ;
        RECT 1381.940 1683.690 1382.200 1684.010 ;
        RECT 1383.320 1683.690 1383.580 1684.010 ;
        RECT 1383.380 1653.410 1383.520 1683.690 ;
        RECT 1383.320 1653.090 1383.580 1653.410 ;
        RECT 2256.400 1653.090 2256.660 1653.410 ;
        RECT 2256.460 2.400 2256.600 1653.090 ;
        RECT 2256.250 -4.800 2256.810 2.400 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1383.750 1591.100 1384.070 1591.160 ;
        RECT 2270.170 1591.100 2270.490 1591.160 ;
        RECT 1383.750 1590.960 2270.490 1591.100 ;
        RECT 1383.750 1590.900 1384.070 1590.960 ;
        RECT 2270.170 1590.900 2270.490 1590.960 ;
      LAYER via ;
        RECT 1383.780 1590.900 1384.040 1591.160 ;
        RECT 2270.200 1590.900 2270.460 1591.160 ;
      LAYER met2 ;
        RECT 1383.680 1700.340 1383.960 1704.000 ;
        RECT 1383.680 1700.000 1383.980 1700.340 ;
        RECT 1383.840 1591.190 1383.980 1700.000 ;
        RECT 1383.780 1590.870 1384.040 1591.190 ;
        RECT 2270.200 1590.870 2270.460 1591.190 ;
        RECT 2270.260 17.410 2270.400 1590.870 ;
        RECT 2270.260 17.270 2274.540 17.410 ;
        RECT 2274.400 2.400 2274.540 17.270 ;
        RECT 2274.190 -4.800 2274.750 2.400 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1386.510 1611.500 1386.830 1611.560 ;
        RECT 2290.870 1611.500 2291.190 1611.560 ;
        RECT 1386.510 1611.360 2291.190 1611.500 ;
        RECT 1386.510 1611.300 1386.830 1611.360 ;
        RECT 2290.870 1611.300 2291.190 1611.360 ;
      LAYER via ;
        RECT 1386.540 1611.300 1386.800 1611.560 ;
        RECT 2290.900 1611.300 2291.160 1611.560 ;
      LAYER met2 ;
        RECT 1385.520 1700.340 1385.800 1704.000 ;
        RECT 1385.520 1700.000 1385.820 1700.340 ;
        RECT 1385.680 1673.210 1385.820 1700.000 ;
        RECT 1385.680 1673.070 1386.740 1673.210 ;
        RECT 1386.600 1611.590 1386.740 1673.070 ;
        RECT 1386.540 1611.270 1386.800 1611.590 ;
        RECT 2290.900 1611.270 2291.160 1611.590 ;
        RECT 2290.960 17.410 2291.100 1611.270 ;
        RECT 2290.960 17.270 2292.480 17.410 ;
        RECT 2292.340 2.400 2292.480 17.270 ;
        RECT 2292.130 -4.800 2292.690 2.400 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1387.430 1690.040 1387.750 1690.100 ;
        RECT 1392.490 1690.040 1392.810 1690.100 ;
        RECT 1387.430 1689.900 1392.810 1690.040 ;
        RECT 1387.430 1689.840 1387.750 1689.900 ;
        RECT 1392.490 1689.840 1392.810 1689.900 ;
        RECT 1392.490 1683.920 1392.810 1683.980 ;
        RECT 1392.490 1683.780 1397.320 1683.920 ;
        RECT 1392.490 1683.720 1392.810 1683.780 ;
        RECT 1397.180 1683.240 1397.320 1683.780 ;
        RECT 1400.770 1683.240 1401.090 1683.300 ;
        RECT 1397.180 1683.100 1401.090 1683.240 ;
        RECT 1400.770 1683.040 1401.090 1683.100 ;
        RECT 1400.770 1676.780 1401.090 1676.840 ;
        RECT 1402.610 1676.780 1402.930 1676.840 ;
        RECT 1400.770 1676.640 1402.930 1676.780 ;
        RECT 1400.770 1676.580 1401.090 1676.640 ;
        RECT 1402.610 1676.580 1402.930 1676.640 ;
        RECT 1403.070 1583.960 1403.390 1584.020 ;
        RECT 2304.670 1583.960 2304.990 1584.020 ;
        RECT 1403.070 1583.820 2304.990 1583.960 ;
        RECT 1403.070 1583.760 1403.390 1583.820 ;
        RECT 2304.670 1583.760 2304.990 1583.820 ;
      LAYER via ;
        RECT 1387.460 1689.840 1387.720 1690.100 ;
        RECT 1392.520 1689.840 1392.780 1690.100 ;
        RECT 1392.520 1683.720 1392.780 1683.980 ;
        RECT 1400.800 1683.040 1401.060 1683.300 ;
        RECT 1400.800 1676.580 1401.060 1676.840 ;
        RECT 1402.640 1676.580 1402.900 1676.840 ;
        RECT 1403.100 1583.760 1403.360 1584.020 ;
        RECT 2304.700 1583.760 2304.960 1584.020 ;
      LAYER met2 ;
        RECT 1387.360 1700.340 1387.640 1704.000 ;
        RECT 1387.360 1700.000 1387.660 1700.340 ;
        RECT 1387.520 1690.130 1387.660 1700.000 ;
        RECT 1387.460 1689.810 1387.720 1690.130 ;
        RECT 1392.520 1689.810 1392.780 1690.130 ;
        RECT 1392.580 1684.010 1392.720 1689.810 ;
        RECT 1392.520 1683.690 1392.780 1684.010 ;
        RECT 1400.800 1683.010 1401.060 1683.330 ;
        RECT 1400.860 1676.870 1401.000 1683.010 ;
        RECT 1400.800 1676.550 1401.060 1676.870 ;
        RECT 1402.640 1676.550 1402.900 1676.870 ;
        RECT 1402.700 1631.050 1402.840 1676.550 ;
        RECT 1402.700 1630.910 1403.300 1631.050 ;
        RECT 1403.160 1584.050 1403.300 1630.910 ;
        RECT 1403.100 1583.730 1403.360 1584.050 ;
        RECT 2304.700 1583.730 2304.960 1584.050 ;
        RECT 2304.760 17.410 2304.900 1583.730 ;
        RECT 2304.760 17.270 2310.420 17.410 ;
        RECT 2310.280 2.400 2310.420 17.270 ;
        RECT 2310.070 -4.800 2310.630 2.400 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1389.270 1690.720 1389.590 1690.780 ;
        RECT 1390.650 1690.720 1390.970 1690.780 ;
        RECT 1389.270 1690.580 1390.970 1690.720 ;
        RECT 1389.270 1690.520 1389.590 1690.580 ;
        RECT 1390.650 1690.520 1390.970 1690.580 ;
        RECT 1390.650 1685.080 1390.970 1685.340 ;
        RECT 1390.740 1684.940 1390.880 1685.080 ;
        RECT 1392.950 1684.940 1393.270 1685.000 ;
        RECT 1390.740 1684.800 1393.270 1684.940 ;
        RECT 1392.950 1684.740 1393.270 1684.800 ;
        RECT 1392.950 1666.920 1393.270 1666.980 ;
        RECT 2325.370 1666.920 2325.690 1666.980 ;
        RECT 1392.950 1666.780 2325.690 1666.920 ;
        RECT 1392.950 1666.720 1393.270 1666.780 ;
        RECT 2325.370 1666.720 2325.690 1666.780 ;
      LAYER via ;
        RECT 1389.300 1690.520 1389.560 1690.780 ;
        RECT 1390.680 1690.520 1390.940 1690.780 ;
        RECT 1390.680 1685.080 1390.940 1685.340 ;
        RECT 1392.980 1684.740 1393.240 1685.000 ;
        RECT 1392.980 1666.720 1393.240 1666.980 ;
        RECT 2325.400 1666.720 2325.660 1666.980 ;
      LAYER met2 ;
        RECT 1389.200 1700.340 1389.480 1704.000 ;
        RECT 1389.200 1700.000 1389.500 1700.340 ;
        RECT 1389.360 1690.810 1389.500 1700.000 ;
        RECT 1389.300 1690.490 1389.560 1690.810 ;
        RECT 1390.680 1690.490 1390.940 1690.810 ;
        RECT 1390.740 1685.370 1390.880 1690.490 ;
        RECT 1390.680 1685.050 1390.940 1685.370 ;
        RECT 1392.980 1684.710 1393.240 1685.030 ;
        RECT 1393.040 1667.010 1393.180 1684.710 ;
        RECT 1392.980 1666.690 1393.240 1667.010 ;
        RECT 2325.400 1666.690 2325.660 1667.010 ;
        RECT 2325.460 17.410 2325.600 1666.690 ;
        RECT 2325.460 17.270 2328.360 17.410 ;
        RECT 2328.220 2.400 2328.360 17.270 ;
        RECT 2328.010 -4.800 2328.570 2.400 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1391.110 1685.280 1391.430 1685.340 ;
        RECT 1393.870 1685.280 1394.190 1685.340 ;
        RECT 1391.110 1685.140 1394.190 1685.280 ;
        RECT 1391.110 1685.080 1391.430 1685.140 ;
        RECT 1393.870 1685.080 1394.190 1685.140 ;
        RECT 1395.250 1645.840 1395.570 1645.900 ;
        RECT 2339.170 1645.840 2339.490 1645.900 ;
        RECT 1395.250 1645.700 2339.490 1645.840 ;
        RECT 1395.250 1645.640 1395.570 1645.700 ;
        RECT 2339.170 1645.640 2339.490 1645.700 ;
        RECT 2339.170 17.580 2339.490 17.640 ;
        RECT 2345.610 17.580 2345.930 17.640 ;
        RECT 2339.170 17.440 2345.930 17.580 ;
        RECT 2339.170 17.380 2339.490 17.440 ;
        RECT 2345.610 17.380 2345.930 17.440 ;
      LAYER via ;
        RECT 1391.140 1685.080 1391.400 1685.340 ;
        RECT 1393.900 1685.080 1394.160 1685.340 ;
        RECT 1395.280 1645.640 1395.540 1645.900 ;
        RECT 2339.200 1645.640 2339.460 1645.900 ;
        RECT 2339.200 17.380 2339.460 17.640 ;
        RECT 2345.640 17.380 2345.900 17.640 ;
      LAYER met2 ;
        RECT 1391.040 1700.340 1391.320 1704.000 ;
        RECT 1391.040 1700.000 1391.340 1700.340 ;
        RECT 1391.200 1685.370 1391.340 1700.000 ;
        RECT 1391.140 1685.050 1391.400 1685.370 ;
        RECT 1393.900 1685.050 1394.160 1685.370 ;
        RECT 1393.960 1676.610 1394.100 1685.050 ;
        RECT 1393.960 1676.470 1395.480 1676.610 ;
        RECT 1395.340 1645.930 1395.480 1676.470 ;
        RECT 1395.280 1645.610 1395.540 1645.930 ;
        RECT 2339.200 1645.610 2339.460 1645.930 ;
        RECT 2339.260 17.670 2339.400 1645.610 ;
        RECT 2339.200 17.350 2339.460 17.670 ;
        RECT 2345.640 17.350 2345.900 17.670 ;
        RECT 2345.700 2.400 2345.840 17.350 ;
        RECT 2345.490 -4.800 2346.050 2.400 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1389.270 1686.640 1389.590 1686.700 ;
        RECT 1392.950 1686.640 1393.270 1686.700 ;
        RECT 1389.270 1686.500 1393.270 1686.640 ;
        RECT 1389.270 1686.440 1389.590 1686.500 ;
        RECT 1392.950 1686.440 1393.270 1686.500 ;
        RECT 1389.270 1625.100 1389.590 1625.160 ;
        RECT 2359.870 1625.100 2360.190 1625.160 ;
        RECT 1389.270 1624.960 2360.190 1625.100 ;
        RECT 1389.270 1624.900 1389.590 1624.960 ;
        RECT 2359.870 1624.900 2360.190 1624.960 ;
      LAYER via ;
        RECT 1389.300 1686.440 1389.560 1686.700 ;
        RECT 1392.980 1686.440 1393.240 1686.700 ;
        RECT 1389.300 1624.900 1389.560 1625.160 ;
        RECT 2359.900 1624.900 2360.160 1625.160 ;
      LAYER met2 ;
        RECT 1392.880 1700.340 1393.160 1704.000 ;
        RECT 1392.880 1700.000 1393.180 1700.340 ;
        RECT 1393.040 1686.730 1393.180 1700.000 ;
        RECT 1389.300 1686.410 1389.560 1686.730 ;
        RECT 1392.980 1686.410 1393.240 1686.730 ;
        RECT 1389.360 1625.190 1389.500 1686.410 ;
        RECT 1389.300 1624.870 1389.560 1625.190 ;
        RECT 2359.900 1624.870 2360.160 1625.190 ;
        RECT 2359.960 16.730 2360.100 1624.870 ;
        RECT 2359.960 16.590 2363.780 16.730 ;
        RECT 2363.640 2.400 2363.780 16.590 ;
        RECT 2363.430 -4.800 2363.990 2.400 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1396.170 1604.700 1396.490 1604.760 ;
        RECT 2380.570 1604.700 2380.890 1604.760 ;
        RECT 1396.170 1604.560 2380.890 1604.700 ;
        RECT 1396.170 1604.500 1396.490 1604.560 ;
        RECT 2380.570 1604.500 2380.890 1604.560 ;
      LAYER via ;
        RECT 1396.200 1604.500 1396.460 1604.760 ;
        RECT 2380.600 1604.500 2380.860 1604.760 ;
      LAYER met2 ;
        RECT 1394.720 1700.340 1395.000 1704.000 ;
        RECT 1394.720 1700.000 1395.020 1700.340 ;
        RECT 1394.880 1677.970 1395.020 1700.000 ;
        RECT 1394.880 1677.830 1396.400 1677.970 ;
        RECT 1396.260 1604.790 1396.400 1677.830 ;
        RECT 1396.200 1604.470 1396.460 1604.790 ;
        RECT 2380.600 1604.470 2380.860 1604.790 ;
        RECT 2380.660 16.730 2380.800 1604.470 ;
        RECT 2380.660 16.590 2381.720 16.730 ;
        RECT 2381.580 2.400 2381.720 16.590 ;
        RECT 2381.370 -4.800 2381.930 2.400 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1396.630 1684.600 1396.950 1684.660 ;
        RECT 1399.390 1684.600 1399.710 1684.660 ;
        RECT 1396.630 1684.460 1399.710 1684.600 ;
        RECT 1396.630 1684.400 1396.950 1684.460 ;
        RECT 1399.390 1684.400 1399.710 1684.460 ;
        RECT 1398.930 1576.820 1399.250 1576.880 ;
        RECT 2394.370 1576.820 2394.690 1576.880 ;
        RECT 1398.930 1576.680 2394.690 1576.820 ;
        RECT 1398.930 1576.620 1399.250 1576.680 ;
        RECT 2394.370 1576.620 2394.690 1576.680 ;
      LAYER via ;
        RECT 1396.660 1684.400 1396.920 1684.660 ;
        RECT 1399.420 1684.400 1399.680 1684.660 ;
        RECT 1398.960 1576.620 1399.220 1576.880 ;
        RECT 2394.400 1576.620 2394.660 1576.880 ;
      LAYER met2 ;
        RECT 1396.560 1700.340 1396.840 1704.000 ;
        RECT 1396.560 1700.000 1396.860 1700.340 ;
        RECT 1396.720 1684.690 1396.860 1700.000 ;
        RECT 1396.660 1684.370 1396.920 1684.690 ;
        RECT 1399.420 1684.370 1399.680 1684.690 ;
        RECT 1399.480 1650.770 1399.620 1684.370 ;
        RECT 1399.020 1650.630 1399.620 1650.770 ;
        RECT 1399.020 1576.910 1399.160 1650.630 ;
        RECT 1398.960 1576.590 1399.220 1576.910 ;
        RECT 2394.400 1576.590 2394.660 1576.910 ;
        RECT 2394.460 16.730 2394.600 1576.590 ;
        RECT 2394.460 16.590 2399.660 16.730 ;
        RECT 2399.520 2.400 2399.660 16.590 ;
        RECT 2399.310 -4.800 2399.870 2.400 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1231.105 1673.905 1231.275 1679.175 ;
      LAYER mcon ;
        RECT 1231.105 1679.005 1231.275 1679.175 ;
      LAYER met1 ;
        RECT 1231.030 1679.160 1231.350 1679.220 ;
        RECT 1230.835 1679.020 1231.350 1679.160 ;
        RECT 1231.030 1678.960 1231.350 1679.020 ;
        RECT 800.010 1674.060 800.330 1674.120 ;
        RECT 1231.045 1674.060 1231.335 1674.105 ;
        RECT 800.010 1673.920 1231.335 1674.060 ;
        RECT 800.010 1673.860 800.330 1673.920 ;
        RECT 1231.045 1673.875 1231.335 1673.920 ;
        RECT 793.570 20.980 793.890 21.040 ;
        RECT 800.010 20.980 800.330 21.040 ;
        RECT 793.570 20.840 800.330 20.980 ;
        RECT 793.570 20.780 793.890 20.840 ;
        RECT 800.010 20.780 800.330 20.840 ;
      LAYER via ;
        RECT 1231.060 1678.960 1231.320 1679.220 ;
        RECT 800.040 1673.860 800.300 1674.120 ;
        RECT 793.600 20.780 793.860 21.040 ;
        RECT 800.040 20.780 800.300 21.040 ;
      LAYER met2 ;
        RECT 1230.960 1700.340 1231.240 1704.000 ;
        RECT 1230.960 1700.000 1231.260 1700.340 ;
        RECT 1231.120 1679.250 1231.260 1700.000 ;
        RECT 1231.060 1678.930 1231.320 1679.250 ;
        RECT 800.040 1673.830 800.300 1674.150 ;
        RECT 800.100 21.070 800.240 1673.830 ;
        RECT 793.600 20.750 793.860 21.070 ;
        RECT 800.040 20.750 800.300 21.070 ;
        RECT 793.660 2.400 793.800 20.750 ;
        RECT 793.450 -4.800 794.010 2.400 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1215.465 1653.165 1215.635 1690.395 ;
      LAYER mcon ;
        RECT 1215.465 1690.225 1215.635 1690.395 ;
      LAYER met1 ;
        RECT 1215.390 1690.380 1215.710 1690.440 ;
        RECT 1215.195 1690.240 1215.710 1690.380 ;
        RECT 1215.390 1690.180 1215.710 1690.240 ;
        RECT 641.310 1653.320 641.630 1653.380 ;
        RECT 1215.405 1653.320 1215.695 1653.365 ;
        RECT 641.310 1653.180 1215.695 1653.320 ;
        RECT 641.310 1653.120 641.630 1653.180 ;
        RECT 1215.405 1653.135 1215.695 1653.180 ;
      LAYER via ;
        RECT 1215.420 1690.180 1215.680 1690.440 ;
        RECT 641.340 1653.120 641.600 1653.380 ;
      LAYER met2 ;
        RECT 1215.320 1700.340 1215.600 1704.000 ;
        RECT 1215.320 1700.000 1215.620 1700.340 ;
        RECT 1215.480 1690.470 1215.620 1700.000 ;
        RECT 1215.420 1690.150 1215.680 1690.470 ;
        RECT 641.340 1653.090 641.600 1653.410 ;
        RECT 641.400 17.410 641.540 1653.090 ;
        RECT 639.100 17.270 641.540 17.410 ;
        RECT 639.100 2.400 639.240 17.270 ;
        RECT 638.890 -4.800 639.450 2.400 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1397.550 1677.460 1397.870 1677.520 ;
        RECT 1398.930 1677.460 1399.250 1677.520 ;
        RECT 1397.550 1677.320 1399.250 1677.460 ;
        RECT 1397.550 1677.260 1397.870 1677.320 ;
        RECT 1398.930 1677.260 1399.250 1677.320 ;
        RECT 1397.550 1570.020 1397.870 1570.080 ;
        RECT 2421.970 1570.020 2422.290 1570.080 ;
        RECT 1397.550 1569.880 2422.290 1570.020 ;
        RECT 1397.550 1569.820 1397.870 1569.880 ;
        RECT 2421.970 1569.820 2422.290 1569.880 ;
      LAYER via ;
        RECT 1397.580 1677.260 1397.840 1677.520 ;
        RECT 1398.960 1677.260 1399.220 1677.520 ;
        RECT 1397.580 1569.820 1397.840 1570.080 ;
        RECT 2422.000 1569.820 2422.260 1570.080 ;
      LAYER met2 ;
        RECT 1398.860 1700.340 1399.140 1704.000 ;
        RECT 1398.860 1700.000 1399.160 1700.340 ;
        RECT 1399.020 1677.550 1399.160 1700.000 ;
        RECT 1397.580 1677.230 1397.840 1677.550 ;
        RECT 1398.960 1677.230 1399.220 1677.550 ;
        RECT 1397.640 1570.110 1397.780 1677.230 ;
        RECT 1397.580 1569.790 1397.840 1570.110 ;
        RECT 2422.000 1569.790 2422.260 1570.110 ;
        RECT 2422.060 17.410 2422.200 1569.790 ;
        RECT 2422.060 17.270 2423.120 17.410 ;
        RECT 2422.980 2.400 2423.120 17.270 ;
        RECT 2422.770 -4.800 2423.330 2.400 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1400.770 1683.920 1401.090 1683.980 ;
        RECT 1402.150 1683.920 1402.470 1683.980 ;
        RECT 1400.770 1683.780 1402.470 1683.920 ;
        RECT 1400.770 1683.720 1401.090 1683.780 ;
        RECT 1402.150 1683.720 1402.470 1683.780 ;
        RECT 1403.530 1597.560 1403.850 1597.620 ;
        RECT 2435.770 1597.560 2436.090 1597.620 ;
        RECT 1403.530 1597.420 2436.090 1597.560 ;
        RECT 1403.530 1597.360 1403.850 1597.420 ;
        RECT 2435.770 1597.360 2436.090 1597.420 ;
      LAYER via ;
        RECT 1400.800 1683.720 1401.060 1683.980 ;
        RECT 1402.180 1683.720 1402.440 1683.980 ;
        RECT 1403.560 1597.360 1403.820 1597.620 ;
        RECT 2435.800 1597.360 2436.060 1597.620 ;
      LAYER met2 ;
        RECT 1400.700 1700.340 1400.980 1704.000 ;
        RECT 1400.700 1700.000 1401.000 1700.340 ;
        RECT 1400.860 1684.010 1401.000 1700.000 ;
        RECT 1400.800 1683.690 1401.060 1684.010 ;
        RECT 1402.180 1683.690 1402.440 1684.010 ;
        RECT 1402.240 1677.290 1402.380 1683.690 ;
        RECT 1402.240 1677.150 1403.300 1677.290 ;
        RECT 1403.160 1631.730 1403.300 1677.150 ;
        RECT 1403.160 1631.590 1403.760 1631.730 ;
        RECT 1403.620 1597.650 1403.760 1631.590 ;
        RECT 1403.560 1597.330 1403.820 1597.650 ;
        RECT 2435.800 1597.330 2436.060 1597.650 ;
        RECT 2435.860 17.410 2436.000 1597.330 ;
        RECT 2435.860 17.270 2441.060 17.410 ;
        RECT 2440.920 2.400 2441.060 17.270 ;
        RECT 2440.710 -4.800 2441.270 2.400 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1402.610 1683.920 1402.930 1683.980 ;
        RECT 1402.610 1683.780 1403.300 1683.920 ;
        RECT 1402.610 1683.720 1402.930 1683.780 ;
        RECT 1403.160 1683.580 1403.300 1683.780 ;
        RECT 1404.450 1683.580 1404.770 1683.640 ;
        RECT 1403.160 1683.440 1404.770 1683.580 ;
        RECT 1404.450 1683.380 1404.770 1683.440 ;
        RECT 1404.450 1563.220 1404.770 1563.280 ;
        RECT 2456.470 1563.220 2456.790 1563.280 ;
        RECT 1404.450 1563.080 2456.790 1563.220 ;
        RECT 1404.450 1563.020 1404.770 1563.080 ;
        RECT 2456.470 1563.020 2456.790 1563.080 ;
      LAYER via ;
        RECT 1402.640 1683.720 1402.900 1683.980 ;
        RECT 1404.480 1683.380 1404.740 1683.640 ;
        RECT 1404.480 1563.020 1404.740 1563.280 ;
        RECT 2456.500 1563.020 2456.760 1563.280 ;
      LAYER met2 ;
        RECT 1402.540 1700.340 1402.820 1704.000 ;
        RECT 1402.540 1700.000 1402.840 1700.340 ;
        RECT 1402.700 1684.010 1402.840 1700.000 ;
        RECT 1402.640 1683.690 1402.900 1684.010 ;
        RECT 1404.480 1683.350 1404.740 1683.670 ;
        RECT 1404.540 1563.310 1404.680 1683.350 ;
        RECT 1404.480 1562.990 1404.740 1563.310 ;
        RECT 2456.500 1562.990 2456.760 1563.310 ;
        RECT 2456.560 3.130 2456.700 1562.990 ;
        RECT 2456.560 2.990 2459.000 3.130 ;
        RECT 2458.860 2.400 2459.000 2.990 ;
        RECT 2458.650 -4.800 2459.210 2.400 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1401.690 1684.940 1402.010 1685.000 ;
        RECT 1404.450 1684.940 1404.770 1685.000 ;
        RECT 1401.690 1684.800 1404.770 1684.940 ;
        RECT 1401.690 1684.740 1402.010 1684.800 ;
        RECT 1404.450 1684.740 1404.770 1684.800 ;
        RECT 1401.690 1631.900 1402.010 1631.960 ;
        RECT 1404.910 1631.900 1405.230 1631.960 ;
        RECT 1401.690 1631.760 1405.230 1631.900 ;
        RECT 1401.690 1631.700 1402.010 1631.760 ;
        RECT 1404.910 1631.700 1405.230 1631.760 ;
        RECT 1404.910 1549.280 1405.230 1549.340 ;
        RECT 2470.270 1549.280 2470.590 1549.340 ;
        RECT 1404.910 1549.140 2470.590 1549.280 ;
        RECT 1404.910 1549.080 1405.230 1549.140 ;
        RECT 2470.270 1549.080 2470.590 1549.140 ;
        RECT 2470.270 16.900 2470.590 16.960 ;
        RECT 2476.710 16.900 2477.030 16.960 ;
        RECT 2470.270 16.760 2477.030 16.900 ;
        RECT 2470.270 16.700 2470.590 16.760 ;
        RECT 2476.710 16.700 2477.030 16.760 ;
      LAYER via ;
        RECT 1401.720 1684.740 1401.980 1685.000 ;
        RECT 1404.480 1684.740 1404.740 1685.000 ;
        RECT 1401.720 1631.700 1401.980 1631.960 ;
        RECT 1404.940 1631.700 1405.200 1631.960 ;
        RECT 1404.940 1549.080 1405.200 1549.340 ;
        RECT 2470.300 1549.080 2470.560 1549.340 ;
        RECT 2470.300 16.700 2470.560 16.960 ;
        RECT 2476.740 16.700 2477.000 16.960 ;
      LAYER met2 ;
        RECT 1404.380 1700.340 1404.660 1704.000 ;
        RECT 1404.380 1700.000 1404.680 1700.340 ;
        RECT 1404.540 1685.030 1404.680 1700.000 ;
        RECT 1401.720 1684.710 1401.980 1685.030 ;
        RECT 1404.480 1684.710 1404.740 1685.030 ;
        RECT 1401.780 1631.990 1401.920 1684.710 ;
        RECT 1401.720 1631.670 1401.980 1631.990 ;
        RECT 1404.940 1631.670 1405.200 1631.990 ;
        RECT 1405.000 1549.370 1405.140 1631.670 ;
        RECT 1404.940 1549.050 1405.200 1549.370 ;
        RECT 2470.300 1549.050 2470.560 1549.370 ;
        RECT 2470.360 16.990 2470.500 1549.050 ;
        RECT 2470.300 16.670 2470.560 16.990 ;
        RECT 2476.740 16.670 2477.000 16.990 ;
        RECT 2476.800 2.400 2476.940 16.670 ;
        RECT 2476.590 -4.800 2477.150 2.400 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1405.370 1631.900 1405.690 1631.960 ;
        RECT 1406.290 1631.900 1406.610 1631.960 ;
        RECT 1405.370 1631.760 1406.610 1631.900 ;
        RECT 1405.370 1631.700 1405.690 1631.760 ;
        RECT 1406.290 1631.700 1406.610 1631.760 ;
        RECT 1405.370 1542.480 1405.690 1542.540 ;
        RECT 2490.970 1542.480 2491.290 1542.540 ;
        RECT 1405.370 1542.340 2491.290 1542.480 ;
        RECT 1405.370 1542.280 1405.690 1542.340 ;
        RECT 2490.970 1542.280 2491.290 1542.340 ;
        RECT 2490.970 2.960 2491.290 3.020 ;
        RECT 2494.650 2.960 2494.970 3.020 ;
        RECT 2490.970 2.820 2494.970 2.960 ;
        RECT 2490.970 2.760 2491.290 2.820 ;
        RECT 2494.650 2.760 2494.970 2.820 ;
      LAYER via ;
        RECT 1405.400 1631.700 1405.660 1631.960 ;
        RECT 1406.320 1631.700 1406.580 1631.960 ;
        RECT 1405.400 1542.280 1405.660 1542.540 ;
        RECT 2491.000 1542.280 2491.260 1542.540 ;
        RECT 2491.000 2.760 2491.260 3.020 ;
        RECT 2494.680 2.760 2494.940 3.020 ;
      LAYER met2 ;
        RECT 1406.220 1700.340 1406.500 1704.000 ;
        RECT 1406.220 1700.000 1406.520 1700.340 ;
        RECT 1406.380 1631.990 1406.520 1700.000 ;
        RECT 1405.400 1631.670 1405.660 1631.990 ;
        RECT 1406.320 1631.670 1406.580 1631.990 ;
        RECT 1405.460 1542.570 1405.600 1631.670 ;
        RECT 1405.400 1542.250 1405.660 1542.570 ;
        RECT 2491.000 1542.250 2491.260 1542.570 ;
        RECT 2491.060 3.050 2491.200 1542.250 ;
        RECT 2491.000 2.730 2491.260 3.050 ;
        RECT 2494.680 2.730 2494.940 3.050 ;
        RECT 2494.740 2.400 2494.880 2.730 ;
        RECT 2494.530 -4.800 2495.090 2.400 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1408.130 1683.920 1408.450 1683.980 ;
        RECT 1408.130 1683.780 1410.200 1683.920 ;
        RECT 1408.130 1683.720 1408.450 1683.780 ;
        RECT 1410.060 1683.580 1410.200 1683.780 ;
        RECT 1414.110 1683.580 1414.430 1683.640 ;
        RECT 1410.060 1683.440 1414.430 1683.580 ;
        RECT 1414.110 1683.380 1414.430 1683.440 ;
        RECT 1414.110 1639.040 1414.430 1639.100 ;
        RECT 2511.670 1639.040 2511.990 1639.100 ;
        RECT 1414.110 1638.900 2511.990 1639.040 ;
        RECT 1414.110 1638.840 1414.430 1638.900 ;
        RECT 2511.670 1638.840 2511.990 1638.900 ;
      LAYER via ;
        RECT 1408.160 1683.720 1408.420 1683.980 ;
        RECT 1414.140 1683.380 1414.400 1683.640 ;
        RECT 1414.140 1638.840 1414.400 1639.100 ;
        RECT 2511.700 1638.840 2511.960 1639.100 ;
      LAYER met2 ;
        RECT 1408.060 1700.340 1408.340 1704.000 ;
        RECT 1408.060 1700.000 1408.360 1700.340 ;
        RECT 1408.220 1684.010 1408.360 1700.000 ;
        RECT 1408.160 1683.690 1408.420 1684.010 ;
        RECT 1414.140 1683.350 1414.400 1683.670 ;
        RECT 1414.200 1639.130 1414.340 1683.350 ;
        RECT 1414.140 1638.810 1414.400 1639.130 ;
        RECT 2511.700 1638.810 2511.960 1639.130 ;
        RECT 2511.760 17.410 2511.900 1638.810 ;
        RECT 2511.760 17.270 2512.360 17.410 ;
        RECT 2512.220 2.400 2512.360 17.270 ;
        RECT 2512.010 -4.800 2512.570 2.400 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1408.590 1590.760 1408.910 1590.820 ;
        RECT 2525.470 1590.760 2525.790 1590.820 ;
        RECT 1408.590 1590.620 2525.790 1590.760 ;
        RECT 1408.590 1590.560 1408.910 1590.620 ;
        RECT 2525.470 1590.560 2525.790 1590.620 ;
      LAYER via ;
        RECT 1408.620 1590.560 1408.880 1590.820 ;
        RECT 2525.500 1590.560 2525.760 1590.820 ;
      LAYER met2 ;
        RECT 1409.900 1700.340 1410.180 1704.000 ;
        RECT 1409.900 1700.000 1410.200 1700.340 ;
        RECT 1410.060 1677.970 1410.200 1700.000 ;
        RECT 1408.680 1677.830 1410.200 1677.970 ;
        RECT 1408.680 1590.850 1408.820 1677.830 ;
        RECT 1408.620 1590.530 1408.880 1590.850 ;
        RECT 2525.500 1590.530 2525.760 1590.850 ;
        RECT 2525.560 17.410 2525.700 1590.530 ;
        RECT 2525.560 17.270 2530.300 17.410 ;
        RECT 2530.160 2.400 2530.300 17.270 ;
        RECT 2529.950 -4.800 2530.510 2.400 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1409.050 1618.300 1409.370 1618.360 ;
        RECT 2546.170 1618.300 2546.490 1618.360 ;
        RECT 1409.050 1618.160 2546.490 1618.300 ;
        RECT 1409.050 1618.100 1409.370 1618.160 ;
        RECT 2546.170 1618.100 2546.490 1618.160 ;
      LAYER via ;
        RECT 1409.080 1618.100 1409.340 1618.360 ;
        RECT 2546.200 1618.100 2546.460 1618.360 ;
      LAYER met2 ;
        RECT 1411.740 1700.340 1412.020 1704.000 ;
        RECT 1411.740 1700.000 1412.040 1700.340 ;
        RECT 1411.900 1677.290 1412.040 1700.000 ;
        RECT 1409.140 1677.150 1412.040 1677.290 ;
        RECT 1409.140 1618.390 1409.280 1677.150 ;
        RECT 1409.080 1618.070 1409.340 1618.390 ;
        RECT 2546.200 1618.070 2546.460 1618.390 ;
        RECT 2546.260 17.410 2546.400 1618.070 ;
        RECT 2546.260 17.270 2548.240 17.410 ;
        RECT 2548.100 2.400 2548.240 17.270 ;
        RECT 2547.890 -4.800 2548.450 2.400 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1413.650 1535.340 1413.970 1535.400 ;
        RECT 2559.970 1535.340 2560.290 1535.400 ;
        RECT 1413.650 1535.200 2560.290 1535.340 ;
        RECT 1413.650 1535.140 1413.970 1535.200 ;
        RECT 2559.970 1535.140 2560.290 1535.200 ;
        RECT 2559.970 16.900 2560.290 16.960 ;
        RECT 2565.950 16.900 2566.270 16.960 ;
        RECT 2559.970 16.760 2566.270 16.900 ;
        RECT 2559.970 16.700 2560.290 16.760 ;
        RECT 2565.950 16.700 2566.270 16.760 ;
      LAYER via ;
        RECT 1413.680 1535.140 1413.940 1535.400 ;
        RECT 2560.000 1535.140 2560.260 1535.400 ;
        RECT 2560.000 16.700 2560.260 16.960 ;
        RECT 2565.980 16.700 2566.240 16.960 ;
      LAYER met2 ;
        RECT 1413.580 1700.340 1413.860 1704.000 ;
        RECT 1413.580 1700.000 1413.880 1700.340 ;
        RECT 1413.740 1535.430 1413.880 1700.000 ;
        RECT 1413.680 1535.110 1413.940 1535.430 ;
        RECT 2560.000 1535.110 2560.260 1535.430 ;
        RECT 2560.060 16.990 2560.200 1535.110 ;
        RECT 2560.000 16.670 2560.260 16.990 ;
        RECT 2565.980 16.670 2566.240 16.990 ;
        RECT 2566.040 2.400 2566.180 16.670 ;
        RECT 2565.830 -4.800 2566.390 2.400 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1415.950 1655.700 1416.270 1655.760 ;
        RECT 1419.170 1655.700 1419.490 1655.760 ;
        RECT 1415.950 1655.560 1419.490 1655.700 ;
        RECT 1415.950 1655.500 1416.270 1655.560 ;
        RECT 1419.170 1655.500 1419.490 1655.560 ;
        RECT 1419.170 1583.620 1419.490 1583.680 ;
        RECT 2580.670 1583.620 2580.990 1583.680 ;
        RECT 1419.170 1583.480 2580.990 1583.620 ;
        RECT 1419.170 1583.420 1419.490 1583.480 ;
        RECT 2580.670 1583.420 2580.990 1583.480 ;
      LAYER via ;
        RECT 1415.980 1655.500 1416.240 1655.760 ;
        RECT 1419.200 1655.500 1419.460 1655.760 ;
        RECT 1419.200 1583.420 1419.460 1583.680 ;
        RECT 2580.700 1583.420 2580.960 1583.680 ;
      LAYER met2 ;
        RECT 1415.420 1700.340 1415.700 1704.000 ;
        RECT 1415.420 1700.000 1415.720 1700.340 ;
        RECT 1415.580 1666.410 1415.720 1700.000 ;
        RECT 1415.580 1666.270 1416.180 1666.410 ;
        RECT 1416.040 1655.790 1416.180 1666.270 ;
        RECT 1415.980 1655.470 1416.240 1655.790 ;
        RECT 1419.200 1655.470 1419.460 1655.790 ;
        RECT 1419.260 1583.710 1419.400 1655.470 ;
        RECT 1419.200 1583.390 1419.460 1583.710 ;
        RECT 2580.700 1583.390 2580.960 1583.710 ;
        RECT 2580.760 17.410 2580.900 1583.390 ;
        RECT 2580.760 17.270 2584.120 17.410 ;
        RECT 2583.980 2.400 2584.120 17.270 ;
        RECT 2583.770 -4.800 2584.330 2.400 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1141.790 1685.960 1142.110 1686.020 ;
        RECT 1141.790 1685.820 1197.220 1685.960 ;
        RECT 1141.790 1685.760 1142.110 1685.820 ;
        RECT 1197.080 1685.620 1197.220 1685.820 ;
        RECT 1233.790 1685.620 1234.110 1685.680 ;
        RECT 1197.080 1685.480 1234.110 1685.620 ;
        RECT 1233.790 1685.420 1234.110 1685.480 ;
        RECT 820.710 72.320 821.030 72.380 ;
        RECT 1141.790 72.320 1142.110 72.380 ;
        RECT 820.710 72.180 1142.110 72.320 ;
        RECT 820.710 72.120 821.030 72.180 ;
        RECT 1141.790 72.120 1142.110 72.180 ;
      LAYER via ;
        RECT 1141.820 1685.760 1142.080 1686.020 ;
        RECT 1233.820 1685.420 1234.080 1685.680 ;
        RECT 820.740 72.120 821.000 72.380 ;
        RECT 1141.820 72.120 1142.080 72.380 ;
      LAYER met2 ;
        RECT 1233.720 1700.340 1234.000 1704.000 ;
        RECT 1233.720 1700.000 1234.020 1700.340 ;
        RECT 1141.820 1685.730 1142.080 1686.050 ;
        RECT 1141.880 72.410 1142.020 1685.730 ;
        RECT 1233.880 1685.710 1234.020 1700.000 ;
        RECT 1233.820 1685.390 1234.080 1685.710 ;
        RECT 820.740 72.090 821.000 72.410 ;
        RECT 1141.820 72.090 1142.080 72.410 ;
        RECT 820.800 17.410 820.940 72.090 ;
        RECT 817.580 17.270 820.940 17.410 ;
        RECT 817.580 2.400 817.720 17.270 ;
        RECT 817.370 -4.800 817.930 2.400 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1414.570 1685.960 1414.890 1686.020 ;
        RECT 1417.330 1685.960 1417.650 1686.020 ;
        RECT 1414.570 1685.820 1417.650 1685.960 ;
        RECT 1414.570 1685.760 1414.890 1685.820 ;
        RECT 1417.330 1685.760 1417.650 1685.820 ;
        RECT 1414.570 1528.200 1414.890 1528.260 ;
        RECT 2601.370 1528.200 2601.690 1528.260 ;
        RECT 1414.570 1528.060 2601.690 1528.200 ;
        RECT 1414.570 1528.000 1414.890 1528.060 ;
        RECT 2601.370 1528.000 2601.690 1528.060 ;
      LAYER via ;
        RECT 1414.600 1685.760 1414.860 1686.020 ;
        RECT 1417.360 1685.760 1417.620 1686.020 ;
        RECT 1414.600 1528.000 1414.860 1528.260 ;
        RECT 2601.400 1528.000 2601.660 1528.260 ;
      LAYER met2 ;
        RECT 1417.260 1700.340 1417.540 1704.000 ;
        RECT 1417.260 1700.000 1417.560 1700.340 ;
        RECT 1417.420 1686.050 1417.560 1700.000 ;
        RECT 1414.600 1685.730 1414.860 1686.050 ;
        RECT 1417.360 1685.730 1417.620 1686.050 ;
        RECT 1414.660 1528.290 1414.800 1685.730 ;
        RECT 1414.600 1527.970 1414.860 1528.290 ;
        RECT 2601.400 1527.970 2601.660 1528.290 ;
        RECT 2601.460 2.400 2601.600 1527.970 ;
        RECT 2601.250 -4.800 2601.810 2.400 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1419.630 1521.400 1419.950 1521.460 ;
        RECT 2615.170 1521.400 2615.490 1521.460 ;
        RECT 1419.630 1521.260 2615.490 1521.400 ;
        RECT 1419.630 1521.200 1419.950 1521.260 ;
        RECT 2615.170 1521.200 2615.490 1521.260 ;
      LAYER via ;
        RECT 1419.660 1521.200 1419.920 1521.460 ;
        RECT 2615.200 1521.200 2615.460 1521.460 ;
      LAYER met2 ;
        RECT 1419.100 1700.340 1419.380 1704.000 ;
        RECT 1419.100 1700.000 1419.400 1700.340 ;
        RECT 1419.260 1677.970 1419.400 1700.000 ;
        RECT 1419.260 1677.830 1419.860 1677.970 ;
        RECT 1419.720 1521.490 1419.860 1677.830 ;
        RECT 1419.660 1521.170 1419.920 1521.490 ;
        RECT 2615.200 1521.170 2615.460 1521.490 ;
        RECT 2615.260 17.410 2615.400 1521.170 ;
        RECT 2615.260 17.270 2619.540 17.410 ;
        RECT 2619.400 2.400 2619.540 17.270 ;
        RECT 2619.190 -4.800 2619.750 2.400 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1415.105 1514.445 1415.275 1545.215 ;
      LAYER mcon ;
        RECT 1415.105 1545.045 1415.275 1545.215 ;
      LAYER met1 ;
        RECT 1415.030 1686.300 1415.350 1686.360 ;
        RECT 1421.010 1686.300 1421.330 1686.360 ;
        RECT 1415.030 1686.160 1421.330 1686.300 ;
        RECT 1415.030 1686.100 1415.350 1686.160 ;
        RECT 1421.010 1686.100 1421.330 1686.160 ;
        RECT 1415.030 1594.160 1415.350 1594.220 ;
        RECT 1416.870 1594.160 1417.190 1594.220 ;
        RECT 1415.030 1594.020 1417.190 1594.160 ;
        RECT 1415.030 1593.960 1415.350 1594.020 ;
        RECT 1416.870 1593.960 1417.190 1594.020 ;
        RECT 1415.030 1545.200 1415.350 1545.260 ;
        RECT 1414.835 1545.060 1415.350 1545.200 ;
        RECT 1415.030 1545.000 1415.350 1545.060 ;
        RECT 1415.045 1514.600 1415.335 1514.645 ;
        RECT 2635.870 1514.600 2636.190 1514.660 ;
        RECT 1415.045 1514.460 2636.190 1514.600 ;
        RECT 1415.045 1514.415 1415.335 1514.460 ;
        RECT 2635.870 1514.400 2636.190 1514.460 ;
      LAYER via ;
        RECT 1415.060 1686.100 1415.320 1686.360 ;
        RECT 1421.040 1686.100 1421.300 1686.360 ;
        RECT 1415.060 1593.960 1415.320 1594.220 ;
        RECT 1416.900 1593.960 1417.160 1594.220 ;
        RECT 1415.060 1545.000 1415.320 1545.260 ;
        RECT 2635.900 1514.400 2636.160 1514.660 ;
      LAYER met2 ;
        RECT 1420.940 1700.340 1421.220 1704.000 ;
        RECT 1420.940 1700.000 1421.240 1700.340 ;
        RECT 1421.100 1686.390 1421.240 1700.000 ;
        RECT 1415.060 1686.070 1415.320 1686.390 ;
        RECT 1421.040 1686.070 1421.300 1686.390 ;
        RECT 1415.120 1642.725 1415.260 1686.070 ;
        RECT 1415.050 1642.355 1415.330 1642.725 ;
        RECT 1416.890 1641.675 1417.170 1642.045 ;
        RECT 1416.960 1594.250 1417.100 1641.675 ;
        RECT 1415.060 1593.930 1415.320 1594.250 ;
        RECT 1416.900 1593.930 1417.160 1594.250 ;
        RECT 1415.120 1545.290 1415.260 1593.930 ;
        RECT 1415.060 1544.970 1415.320 1545.290 ;
        RECT 2635.900 1514.370 2636.160 1514.690 ;
        RECT 2635.960 17.410 2636.100 1514.370 ;
        RECT 2635.960 17.270 2637.480 17.410 ;
        RECT 2637.340 2.400 2637.480 17.270 ;
        RECT 2637.130 -4.800 2637.690 2.400 ;
      LAYER via2 ;
        RECT 1415.050 1642.400 1415.330 1642.680 ;
        RECT 1416.890 1641.720 1417.170 1642.000 ;
      LAYER met3 ;
        RECT 1415.025 1642.690 1415.355 1642.705 ;
        RECT 1415.025 1642.390 1416.490 1642.690 ;
        RECT 1415.025 1642.375 1415.355 1642.390 ;
        RECT 1416.190 1642.010 1416.490 1642.390 ;
        RECT 1416.865 1642.010 1417.195 1642.025 ;
        RECT 1416.190 1641.710 1417.195 1642.010 ;
        RECT 1416.865 1641.695 1417.195 1641.710 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1421.470 1683.920 1421.790 1683.980 ;
        RECT 1422.850 1683.920 1423.170 1683.980 ;
        RECT 1421.470 1683.780 1423.170 1683.920 ;
        RECT 1421.470 1683.720 1421.790 1683.780 ;
        RECT 1422.850 1683.720 1423.170 1683.780 ;
        RECT 1421.470 1576.480 1421.790 1576.540 ;
        RECT 2649.670 1576.480 2649.990 1576.540 ;
        RECT 1421.470 1576.340 2649.990 1576.480 ;
        RECT 1421.470 1576.280 1421.790 1576.340 ;
        RECT 2649.670 1576.280 2649.990 1576.340 ;
      LAYER via ;
        RECT 1421.500 1683.720 1421.760 1683.980 ;
        RECT 1422.880 1683.720 1423.140 1683.980 ;
        RECT 1421.500 1576.280 1421.760 1576.540 ;
        RECT 2649.700 1576.280 2649.960 1576.540 ;
      LAYER met2 ;
        RECT 1422.780 1700.340 1423.060 1704.000 ;
        RECT 1422.780 1700.000 1423.080 1700.340 ;
        RECT 1422.940 1684.010 1423.080 1700.000 ;
        RECT 1421.500 1683.690 1421.760 1684.010 ;
        RECT 1422.880 1683.690 1423.140 1684.010 ;
        RECT 1421.560 1576.570 1421.700 1683.690 ;
        RECT 1421.500 1576.250 1421.760 1576.570 ;
        RECT 2649.700 1576.250 2649.960 1576.570 ;
        RECT 2649.760 17.410 2649.900 1576.250 ;
        RECT 2649.760 17.270 2655.420 17.410 ;
        RECT 2655.280 2.400 2655.420 17.270 ;
        RECT 2655.070 -4.800 2655.630 2.400 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1422.005 1644.325 1422.175 1678.835 ;
      LAYER mcon ;
        RECT 1422.005 1678.665 1422.175 1678.835 ;
      LAYER met1 ;
        RECT 1421.945 1678.820 1422.235 1678.865 ;
        RECT 1424.690 1678.820 1425.010 1678.880 ;
        RECT 1421.945 1678.680 1425.010 1678.820 ;
        RECT 1421.945 1678.635 1422.235 1678.680 ;
        RECT 1424.690 1678.620 1425.010 1678.680 ;
        RECT 1421.930 1644.480 1422.250 1644.540 ;
        RECT 1421.735 1644.340 1422.250 1644.480 ;
        RECT 1421.930 1644.280 1422.250 1644.340 ;
        RECT 1421.930 1507.460 1422.250 1507.520 ;
        RECT 2670.370 1507.460 2670.690 1507.520 ;
        RECT 1421.930 1507.320 2670.690 1507.460 ;
        RECT 1421.930 1507.260 1422.250 1507.320 ;
        RECT 2670.370 1507.260 2670.690 1507.320 ;
      LAYER via ;
        RECT 1424.720 1678.620 1424.980 1678.880 ;
        RECT 1421.960 1644.280 1422.220 1644.540 ;
        RECT 1421.960 1507.260 1422.220 1507.520 ;
        RECT 2670.400 1507.260 2670.660 1507.520 ;
      LAYER met2 ;
        RECT 1424.620 1700.340 1424.900 1704.000 ;
        RECT 1424.620 1700.000 1424.920 1700.340 ;
        RECT 1424.780 1678.910 1424.920 1700.000 ;
        RECT 1424.720 1678.590 1424.980 1678.910 ;
        RECT 1421.960 1644.250 1422.220 1644.570 ;
        RECT 1422.020 1507.550 1422.160 1644.250 ;
        RECT 1421.960 1507.230 1422.220 1507.550 ;
        RECT 2670.400 1507.230 2670.660 1507.550 ;
        RECT 2670.460 17.410 2670.600 1507.230 ;
        RECT 2670.460 17.270 2672.900 17.410 ;
        RECT 2672.760 2.400 2672.900 17.270 ;
        RECT 2672.550 -4.800 2673.110 2.400 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1426.530 1500.660 1426.850 1500.720 ;
        RECT 2684.630 1500.660 2684.950 1500.720 ;
        RECT 1426.530 1500.520 2684.950 1500.660 ;
        RECT 1426.530 1500.460 1426.850 1500.520 ;
        RECT 2684.630 1500.460 2684.950 1500.520 ;
        RECT 2684.630 18.260 2684.950 18.320 ;
        RECT 2690.610 18.260 2690.930 18.320 ;
        RECT 2684.630 18.120 2690.930 18.260 ;
        RECT 2684.630 18.060 2684.950 18.120 ;
        RECT 2690.610 18.060 2690.930 18.120 ;
      LAYER via ;
        RECT 1426.560 1500.460 1426.820 1500.720 ;
        RECT 2684.660 1500.460 2684.920 1500.720 ;
        RECT 2684.660 18.060 2684.920 18.320 ;
        RECT 2690.640 18.060 2690.900 18.320 ;
      LAYER met2 ;
        RECT 1426.460 1700.340 1426.740 1704.000 ;
        RECT 1426.460 1700.000 1426.760 1700.340 ;
        RECT 1426.620 1500.750 1426.760 1700.000 ;
        RECT 1426.560 1500.430 1426.820 1500.750 ;
        RECT 2684.660 1500.430 2684.920 1500.750 ;
        RECT 2684.720 18.350 2684.860 1500.430 ;
        RECT 2684.660 18.030 2684.920 18.350 ;
        RECT 2690.640 18.030 2690.900 18.350 ;
        RECT 2690.700 2.400 2690.840 18.030 ;
        RECT 2690.490 -4.800 2691.050 2.400 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1428.370 1684.600 1428.690 1684.660 ;
        RECT 1431.590 1684.600 1431.910 1684.660 ;
        RECT 1428.370 1684.460 1431.910 1684.600 ;
        RECT 1428.370 1684.400 1428.690 1684.460 ;
        RECT 1431.590 1684.400 1431.910 1684.460 ;
        RECT 1431.590 1604.360 1431.910 1604.420 ;
        RECT 2704.870 1604.360 2705.190 1604.420 ;
        RECT 1431.590 1604.220 2705.190 1604.360 ;
        RECT 1431.590 1604.160 1431.910 1604.220 ;
        RECT 2704.870 1604.160 2705.190 1604.220 ;
      LAYER via ;
        RECT 1428.400 1684.400 1428.660 1684.660 ;
        RECT 1431.620 1684.400 1431.880 1684.660 ;
        RECT 1431.620 1604.160 1431.880 1604.420 ;
        RECT 2704.900 1604.160 2705.160 1604.420 ;
      LAYER met2 ;
        RECT 1428.300 1700.340 1428.580 1704.000 ;
        RECT 1428.300 1700.000 1428.600 1700.340 ;
        RECT 1428.460 1684.690 1428.600 1700.000 ;
        RECT 1428.400 1684.370 1428.660 1684.690 ;
        RECT 1431.620 1684.370 1431.880 1684.690 ;
        RECT 1431.680 1604.450 1431.820 1684.370 ;
        RECT 1431.620 1604.130 1431.880 1604.450 ;
        RECT 2704.900 1604.130 2705.160 1604.450 ;
        RECT 2704.960 17.410 2705.100 1604.130 ;
        RECT 2704.960 17.270 2708.780 17.410 ;
        RECT 2708.640 2.400 2708.780 17.270 ;
        RECT 2708.430 -4.800 2708.990 2.400 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1430.210 1685.960 1430.530 1686.020 ;
        RECT 1434.810 1685.960 1435.130 1686.020 ;
        RECT 1430.210 1685.820 1435.130 1685.960 ;
        RECT 1430.210 1685.760 1430.530 1685.820 ;
        RECT 1434.810 1685.760 1435.130 1685.820 ;
        RECT 1433.430 1631.900 1433.750 1631.960 ;
        RECT 1434.810 1631.900 1435.130 1631.960 ;
        RECT 1433.430 1631.760 1435.130 1631.900 ;
        RECT 1433.430 1631.700 1433.750 1631.760 ;
        RECT 1434.810 1631.700 1435.130 1631.760 ;
        RECT 1433.430 1569.680 1433.750 1569.740 ;
        RECT 2725.570 1569.680 2725.890 1569.740 ;
        RECT 1433.430 1569.540 2725.890 1569.680 ;
        RECT 1433.430 1569.480 1433.750 1569.540 ;
        RECT 2725.570 1569.480 2725.890 1569.540 ;
      LAYER via ;
        RECT 1430.240 1685.760 1430.500 1686.020 ;
        RECT 1434.840 1685.760 1435.100 1686.020 ;
        RECT 1433.460 1631.700 1433.720 1631.960 ;
        RECT 1434.840 1631.700 1435.100 1631.960 ;
        RECT 1433.460 1569.480 1433.720 1569.740 ;
        RECT 2725.600 1569.480 2725.860 1569.740 ;
      LAYER met2 ;
        RECT 1430.140 1700.340 1430.420 1704.000 ;
        RECT 1430.140 1700.000 1430.440 1700.340 ;
        RECT 1430.300 1686.050 1430.440 1700.000 ;
        RECT 1430.240 1685.730 1430.500 1686.050 ;
        RECT 1434.840 1685.730 1435.100 1686.050 ;
        RECT 1434.900 1631.990 1435.040 1685.730 ;
        RECT 1433.460 1631.670 1433.720 1631.990 ;
        RECT 1434.840 1631.670 1435.100 1631.990 ;
        RECT 1433.520 1569.770 1433.660 1631.670 ;
        RECT 1433.460 1569.450 1433.720 1569.770 ;
        RECT 2725.600 1569.450 2725.860 1569.770 ;
        RECT 2725.660 17.410 2725.800 1569.450 ;
        RECT 2725.660 17.270 2726.720 17.410 ;
        RECT 2726.580 2.400 2726.720 17.270 ;
        RECT 2726.370 -4.800 2726.930 2.400 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1429.750 1684.260 1430.070 1684.320 ;
        RECT 1432.050 1684.260 1432.370 1684.320 ;
        RECT 1429.750 1684.120 1432.370 1684.260 ;
        RECT 1429.750 1684.060 1430.070 1684.120 ;
        RECT 1432.050 1684.060 1432.370 1684.120 ;
        RECT 1429.750 1487.060 1430.070 1487.120 ;
        RECT 2739.370 1487.060 2739.690 1487.120 ;
        RECT 1429.750 1486.920 2739.690 1487.060 ;
        RECT 1429.750 1486.860 1430.070 1486.920 ;
        RECT 2739.370 1486.860 2739.690 1486.920 ;
      LAYER via ;
        RECT 1429.780 1684.060 1430.040 1684.320 ;
        RECT 1432.080 1684.060 1432.340 1684.320 ;
        RECT 1429.780 1486.860 1430.040 1487.120 ;
        RECT 2739.400 1486.860 2739.660 1487.120 ;
      LAYER met2 ;
        RECT 1431.980 1700.340 1432.260 1704.000 ;
        RECT 1431.980 1700.000 1432.280 1700.340 ;
        RECT 1432.140 1684.350 1432.280 1700.000 ;
        RECT 1429.780 1684.030 1430.040 1684.350 ;
        RECT 1432.080 1684.030 1432.340 1684.350 ;
        RECT 1429.840 1487.150 1429.980 1684.030 ;
        RECT 1429.780 1486.830 1430.040 1487.150 ;
        RECT 2739.400 1486.830 2739.660 1487.150 ;
        RECT 2739.460 17.410 2739.600 1486.830 ;
        RECT 2739.460 17.270 2744.660 17.410 ;
        RECT 2744.520 2.400 2744.660 17.270 ;
        RECT 2744.310 -4.800 2744.870 2.400 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1432.970 1562.880 1433.290 1562.940 ;
        RECT 2760.070 1562.880 2760.390 1562.940 ;
        RECT 1432.970 1562.740 2760.390 1562.880 ;
        RECT 1432.970 1562.680 1433.290 1562.740 ;
        RECT 2760.070 1562.680 2760.390 1562.740 ;
      LAYER via ;
        RECT 1433.000 1562.680 1433.260 1562.940 ;
        RECT 2760.100 1562.680 2760.360 1562.940 ;
      LAYER met2 ;
        RECT 1433.820 1700.340 1434.100 1704.000 ;
        RECT 1433.820 1700.000 1434.120 1700.340 ;
        RECT 1433.980 1665.050 1434.120 1700.000 ;
        RECT 1433.060 1664.910 1434.120 1665.050 ;
        RECT 1433.060 1562.970 1433.200 1664.910 ;
        RECT 1433.000 1562.650 1433.260 1562.970 ;
        RECT 2760.100 1562.650 2760.360 1562.970 ;
        RECT 2760.160 17.410 2760.300 1562.650 ;
        RECT 2760.160 17.270 2762.140 17.410 ;
        RECT 2762.000 2.400 2762.140 17.270 ;
        RECT 2761.790 -4.800 2762.350 2.400 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 841.410 1639.720 841.730 1639.780 ;
        RECT 1235.630 1639.720 1235.950 1639.780 ;
        RECT 841.410 1639.580 1235.950 1639.720 ;
        RECT 841.410 1639.520 841.730 1639.580 ;
        RECT 1235.630 1639.520 1235.950 1639.580 ;
        RECT 835.430 20.980 835.750 21.040 ;
        RECT 841.410 20.980 841.730 21.040 ;
        RECT 835.430 20.840 841.730 20.980 ;
        RECT 835.430 20.780 835.750 20.840 ;
        RECT 841.410 20.780 841.730 20.840 ;
      LAYER via ;
        RECT 841.440 1639.520 841.700 1639.780 ;
        RECT 1235.660 1639.520 1235.920 1639.780 ;
        RECT 835.460 20.780 835.720 21.040 ;
        RECT 841.440 20.780 841.700 21.040 ;
      LAYER met2 ;
        RECT 1235.560 1700.340 1235.840 1704.000 ;
        RECT 1235.560 1700.000 1235.860 1700.340 ;
        RECT 1235.720 1639.810 1235.860 1700.000 ;
        RECT 841.440 1639.490 841.700 1639.810 ;
        RECT 1235.660 1639.490 1235.920 1639.810 ;
        RECT 841.500 21.070 841.640 1639.490 ;
        RECT 835.460 20.750 835.720 21.070 ;
        RECT 841.440 20.750 841.700 21.070 ;
        RECT 835.520 2.400 835.660 20.750 ;
        RECT 835.310 -4.800 835.870 2.400 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1435.730 1611.160 1436.050 1611.220 ;
        RECT 2774.330 1611.160 2774.650 1611.220 ;
        RECT 1435.730 1611.020 2774.650 1611.160 ;
        RECT 1435.730 1610.960 1436.050 1611.020 ;
        RECT 2774.330 1610.960 2774.650 1611.020 ;
      LAYER via ;
        RECT 1435.760 1610.960 1436.020 1611.220 ;
        RECT 2774.360 1610.960 2774.620 1611.220 ;
      LAYER met2 ;
        RECT 1435.660 1700.340 1435.940 1704.000 ;
        RECT 1435.660 1700.000 1435.960 1700.340 ;
        RECT 1435.820 1611.250 1435.960 1700.000 ;
        RECT 1435.760 1610.930 1436.020 1611.250 ;
        RECT 2774.360 1610.930 2774.620 1611.250 ;
        RECT 2774.420 17.410 2774.560 1610.930 ;
        RECT 2774.420 17.270 2780.080 17.410 ;
        RECT 2779.940 2.400 2780.080 17.270 ;
        RECT 2779.730 -4.800 2780.290 2.400 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1437.570 1684.260 1437.890 1684.320 ;
        RECT 1440.330 1684.260 1440.650 1684.320 ;
        RECT 1437.570 1684.120 1440.650 1684.260 ;
        RECT 1437.570 1684.060 1437.890 1684.120 ;
        RECT 1440.330 1684.060 1440.650 1684.120 ;
        RECT 1439.870 1597.220 1440.190 1597.280 ;
        RECT 2783.990 1597.220 2784.310 1597.280 ;
        RECT 1439.870 1597.080 2784.310 1597.220 ;
        RECT 1439.870 1597.020 1440.190 1597.080 ;
        RECT 2783.990 1597.020 2784.310 1597.080 ;
        RECT 2783.990 20.640 2784.310 20.700 ;
        RECT 2797.790 20.640 2798.110 20.700 ;
        RECT 2783.990 20.500 2798.110 20.640 ;
        RECT 2783.990 20.440 2784.310 20.500 ;
        RECT 2797.790 20.440 2798.110 20.500 ;
      LAYER via ;
        RECT 1437.600 1684.060 1437.860 1684.320 ;
        RECT 1440.360 1684.060 1440.620 1684.320 ;
        RECT 1439.900 1597.020 1440.160 1597.280 ;
        RECT 2784.020 1597.020 2784.280 1597.280 ;
        RECT 2784.020 20.440 2784.280 20.700 ;
        RECT 2797.820 20.440 2798.080 20.700 ;
      LAYER met2 ;
        RECT 1437.500 1700.340 1437.780 1704.000 ;
        RECT 1437.500 1700.000 1437.800 1700.340 ;
        RECT 1437.660 1684.350 1437.800 1700.000 ;
        RECT 1437.600 1684.030 1437.860 1684.350 ;
        RECT 1440.360 1684.030 1440.620 1684.350 ;
        RECT 1440.420 1677.970 1440.560 1684.030 ;
        RECT 1439.960 1677.830 1440.560 1677.970 ;
        RECT 1439.960 1597.310 1440.100 1677.830 ;
        RECT 1439.900 1596.990 1440.160 1597.310 ;
        RECT 2784.020 1596.990 2784.280 1597.310 ;
        RECT 2784.080 20.730 2784.220 1596.990 ;
        RECT 2784.020 20.410 2784.280 20.730 ;
        RECT 2797.820 20.410 2798.080 20.730 ;
        RECT 2797.880 2.400 2798.020 20.410 ;
        RECT 2797.670 -4.800 2798.230 2.400 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1439.410 1548.940 1439.730 1549.000 ;
        RECT 2815.270 1548.940 2815.590 1549.000 ;
        RECT 1439.410 1548.800 2815.590 1548.940 ;
        RECT 1439.410 1548.740 1439.730 1548.800 ;
        RECT 2815.270 1548.740 2815.590 1548.800 ;
      LAYER via ;
        RECT 1439.440 1548.740 1439.700 1549.000 ;
        RECT 2815.300 1548.740 2815.560 1549.000 ;
      LAYER met2 ;
        RECT 1439.340 1700.340 1439.620 1704.000 ;
        RECT 1439.340 1700.000 1439.640 1700.340 ;
        RECT 1439.500 1549.030 1439.640 1700.000 ;
        RECT 1439.440 1548.710 1439.700 1549.030 ;
        RECT 2815.300 1548.710 2815.560 1549.030 ;
        RECT 2815.360 17.410 2815.500 1548.710 ;
        RECT 2815.360 17.270 2815.960 17.410 ;
        RECT 2815.820 2.400 2815.960 17.270 ;
        RECT 2815.610 -4.800 2816.170 2.400 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1440.330 1479.920 1440.650 1479.980 ;
        RECT 2825.390 1479.920 2825.710 1479.980 ;
        RECT 1440.330 1479.780 2825.710 1479.920 ;
        RECT 1440.330 1479.720 1440.650 1479.780 ;
        RECT 2825.390 1479.720 2825.710 1479.780 ;
        RECT 2825.390 18.260 2825.710 18.320 ;
        RECT 2833.670 18.260 2833.990 18.320 ;
        RECT 2825.390 18.120 2833.990 18.260 ;
        RECT 2825.390 18.060 2825.710 18.120 ;
        RECT 2833.670 18.060 2833.990 18.120 ;
      LAYER via ;
        RECT 1440.360 1479.720 1440.620 1479.980 ;
        RECT 2825.420 1479.720 2825.680 1479.980 ;
        RECT 2825.420 18.060 2825.680 18.320 ;
        RECT 2833.700 18.060 2833.960 18.320 ;
      LAYER met2 ;
        RECT 1441.180 1700.340 1441.460 1704.000 ;
        RECT 1441.180 1700.000 1441.480 1700.340 ;
        RECT 1441.340 1665.050 1441.480 1700.000 ;
        RECT 1440.420 1664.910 1441.480 1665.050 ;
        RECT 1440.420 1480.010 1440.560 1664.910 ;
        RECT 1440.360 1479.690 1440.620 1480.010 ;
        RECT 2825.420 1479.690 2825.680 1480.010 ;
        RECT 2825.480 18.350 2825.620 1479.690 ;
        RECT 2825.420 18.030 2825.680 18.350 ;
        RECT 2833.700 18.030 2833.960 18.350 ;
        RECT 2833.760 2.400 2833.900 18.030 ;
        RECT 2833.550 -4.800 2834.110 2.400 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1443.090 1684.600 1443.410 1684.660 ;
        RECT 1452.750 1684.600 1453.070 1684.660 ;
        RECT 1443.090 1684.460 1453.070 1684.600 ;
        RECT 1443.090 1684.400 1443.410 1684.460 ;
        RECT 1452.750 1684.400 1453.070 1684.460 ;
        RECT 1452.750 1473.120 1453.070 1473.180 ;
        RECT 2849.770 1473.120 2850.090 1473.180 ;
        RECT 1452.750 1472.980 2850.090 1473.120 ;
        RECT 1452.750 1472.920 1453.070 1472.980 ;
        RECT 2849.770 1472.920 2850.090 1472.980 ;
      LAYER via ;
        RECT 1443.120 1684.400 1443.380 1684.660 ;
        RECT 1452.780 1684.400 1453.040 1684.660 ;
        RECT 1452.780 1472.920 1453.040 1473.180 ;
        RECT 2849.800 1472.920 2850.060 1473.180 ;
      LAYER met2 ;
        RECT 1443.020 1700.340 1443.300 1704.000 ;
        RECT 1443.020 1700.000 1443.320 1700.340 ;
        RECT 1443.180 1684.690 1443.320 1700.000 ;
        RECT 1443.120 1684.370 1443.380 1684.690 ;
        RECT 1452.780 1684.370 1453.040 1684.690 ;
        RECT 1452.840 1473.210 1452.980 1684.370 ;
        RECT 1452.780 1472.890 1453.040 1473.210 ;
        RECT 2849.800 1472.890 2850.060 1473.210 ;
        RECT 2849.860 16.730 2850.000 1472.890 ;
        RECT 2849.860 16.590 2851.380 16.730 ;
        RECT 2851.240 2.400 2851.380 16.590 ;
        RECT 2851.030 -4.800 2851.590 2.400 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1446.310 1590.420 1446.630 1590.480 ;
        RECT 2839.190 1590.420 2839.510 1590.480 ;
        RECT 1446.310 1590.280 2839.510 1590.420 ;
        RECT 1446.310 1590.220 1446.630 1590.280 ;
        RECT 2839.190 1590.220 2839.510 1590.280 ;
        RECT 2839.190 18.940 2839.510 19.000 ;
        RECT 2869.090 18.940 2869.410 19.000 ;
        RECT 2839.190 18.800 2869.410 18.940 ;
        RECT 2839.190 18.740 2839.510 18.800 ;
        RECT 2869.090 18.740 2869.410 18.800 ;
      LAYER via ;
        RECT 1446.340 1590.220 1446.600 1590.480 ;
        RECT 2839.220 1590.220 2839.480 1590.480 ;
        RECT 2839.220 18.740 2839.480 19.000 ;
        RECT 2869.120 18.740 2869.380 19.000 ;
      LAYER met2 ;
        RECT 1444.860 1700.340 1445.140 1704.000 ;
        RECT 1444.860 1700.000 1445.160 1700.340 ;
        RECT 1445.020 1660.970 1445.160 1700.000 ;
        RECT 1445.020 1660.830 1446.540 1660.970 ;
        RECT 1446.400 1590.510 1446.540 1660.830 ;
        RECT 1446.340 1590.190 1446.600 1590.510 ;
        RECT 2839.220 1590.190 2839.480 1590.510 ;
        RECT 2839.280 19.030 2839.420 1590.190 ;
        RECT 2839.220 18.710 2839.480 19.030 ;
        RECT 2869.120 18.710 2869.380 19.030 ;
        RECT 2869.180 2.400 2869.320 18.710 ;
        RECT 2868.970 -4.800 2869.530 2.400 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1446.770 1542.140 1447.090 1542.200 ;
        RECT 2874.150 1542.140 2874.470 1542.200 ;
        RECT 1446.770 1542.000 2874.470 1542.140 ;
        RECT 1446.770 1541.940 1447.090 1542.000 ;
        RECT 2874.150 1541.940 2874.470 1542.000 ;
        RECT 2874.150 16.560 2874.470 16.620 ;
        RECT 2887.030 16.560 2887.350 16.620 ;
        RECT 2874.150 16.420 2887.350 16.560 ;
        RECT 2874.150 16.360 2874.470 16.420 ;
        RECT 2887.030 16.360 2887.350 16.420 ;
      LAYER via ;
        RECT 1446.800 1541.940 1447.060 1542.200 ;
        RECT 2874.180 1541.940 2874.440 1542.200 ;
        RECT 2874.180 16.360 2874.440 16.620 ;
        RECT 2887.060 16.360 2887.320 16.620 ;
      LAYER met2 ;
        RECT 1446.700 1700.340 1446.980 1704.000 ;
        RECT 1446.700 1700.000 1447.000 1700.340 ;
        RECT 1446.860 1542.230 1447.000 1700.000 ;
        RECT 1446.800 1541.910 1447.060 1542.230 ;
        RECT 2874.180 1541.910 2874.440 1542.230 ;
        RECT 2874.240 16.650 2874.380 1541.910 ;
        RECT 2874.180 16.330 2874.440 16.650 ;
        RECT 2887.060 16.330 2887.320 16.650 ;
        RECT 2887.120 2.400 2887.260 16.330 ;
        RECT 2886.910 -4.800 2887.470 2.400 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1445.850 1659.780 1446.170 1659.840 ;
        RECT 1448.610 1659.780 1448.930 1659.840 ;
        RECT 1445.850 1659.640 1448.930 1659.780 ;
        RECT 1445.850 1659.580 1446.170 1659.640 ;
        RECT 1448.610 1659.580 1448.930 1659.640 ;
        RECT 1444.470 1631.900 1444.790 1631.960 ;
        RECT 1445.850 1631.900 1446.170 1631.960 ;
        RECT 1444.470 1631.760 1446.170 1631.900 ;
        RECT 1444.470 1631.700 1444.790 1631.760 ;
        RECT 1445.850 1631.700 1446.170 1631.760 ;
        RECT 1445.850 1545.540 1446.170 1545.600 ;
        RECT 1446.310 1545.540 1446.630 1545.600 ;
        RECT 1445.850 1545.400 1446.630 1545.540 ;
        RECT 1445.850 1545.340 1446.170 1545.400 ;
        RECT 1446.310 1545.340 1446.630 1545.400 ;
        RECT 1446.770 1466.320 1447.090 1466.380 ;
        RECT 2867.250 1466.320 2867.570 1466.380 ;
        RECT 1446.770 1466.180 2867.570 1466.320 ;
        RECT 1446.770 1466.120 1447.090 1466.180 ;
        RECT 2867.250 1466.120 2867.570 1466.180 ;
        RECT 2867.250 18.260 2867.570 18.320 ;
        RECT 2904.970 18.260 2905.290 18.320 ;
        RECT 2867.250 18.120 2905.290 18.260 ;
        RECT 2867.250 18.060 2867.570 18.120 ;
        RECT 2904.970 18.060 2905.290 18.120 ;
      LAYER via ;
        RECT 1445.880 1659.580 1446.140 1659.840 ;
        RECT 1448.640 1659.580 1448.900 1659.840 ;
        RECT 1444.500 1631.700 1444.760 1631.960 ;
        RECT 1445.880 1631.700 1446.140 1631.960 ;
        RECT 1445.880 1545.340 1446.140 1545.600 ;
        RECT 1446.340 1545.340 1446.600 1545.600 ;
        RECT 1446.800 1466.120 1447.060 1466.380 ;
        RECT 2867.280 1466.120 2867.540 1466.380 ;
        RECT 2867.280 18.060 2867.540 18.320 ;
        RECT 2905.000 18.060 2905.260 18.320 ;
      LAYER met2 ;
        RECT 1448.540 1700.340 1448.820 1704.000 ;
        RECT 1448.540 1700.000 1448.840 1700.340 ;
        RECT 1448.700 1659.870 1448.840 1700.000 ;
        RECT 1445.880 1659.550 1446.140 1659.870 ;
        RECT 1448.640 1659.550 1448.900 1659.870 ;
        RECT 1445.940 1631.990 1446.080 1659.550 ;
        RECT 1444.500 1631.670 1444.760 1631.990 ;
        RECT 1445.880 1631.670 1446.140 1631.990 ;
        RECT 1444.560 1569.850 1444.700 1631.670 ;
        RECT 1444.560 1569.710 1446.080 1569.850 ;
        RECT 1445.940 1545.630 1446.080 1569.710 ;
        RECT 1445.880 1545.310 1446.140 1545.630 ;
        RECT 1446.340 1545.310 1446.600 1545.630 ;
        RECT 1446.400 1541.290 1446.540 1545.310 ;
        RECT 1446.400 1541.150 1447.000 1541.290 ;
        RECT 1446.860 1466.410 1447.000 1541.150 ;
        RECT 1446.800 1466.090 1447.060 1466.410 ;
        RECT 2867.280 1466.090 2867.540 1466.410 ;
        RECT 2867.340 18.350 2867.480 1466.090 ;
        RECT 2867.280 18.030 2867.540 18.350 ;
        RECT 2905.000 18.030 2905.260 18.350 ;
        RECT 2905.060 2.400 2905.200 18.030 ;
        RECT 2904.850 -4.800 2905.410 2.400 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 855.210 1632.920 855.530 1632.980 ;
        RECT 1237.930 1632.920 1238.250 1632.980 ;
        RECT 855.210 1632.780 1238.250 1632.920 ;
        RECT 855.210 1632.720 855.530 1632.780 ;
        RECT 1237.930 1632.720 1238.250 1632.780 ;
      LAYER via ;
        RECT 855.240 1632.720 855.500 1632.980 ;
        RECT 1237.960 1632.720 1238.220 1632.980 ;
      LAYER met2 ;
        RECT 1237.400 1700.340 1237.680 1704.000 ;
        RECT 1237.400 1700.000 1237.700 1700.340 ;
        RECT 1237.560 1677.290 1237.700 1700.000 ;
        RECT 1237.560 1677.150 1238.160 1677.290 ;
        RECT 1238.020 1633.010 1238.160 1677.150 ;
        RECT 855.240 1632.690 855.500 1633.010 ;
        RECT 1237.960 1632.690 1238.220 1633.010 ;
        RECT 855.300 17.410 855.440 1632.690 ;
        RECT 853.000 17.270 855.440 17.410 ;
        RECT 853.000 2.400 853.140 17.270 ;
        RECT 852.790 -4.800 853.350 2.400 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 870.850 31.860 871.170 31.920 ;
        RECT 1239.310 31.860 1239.630 31.920 ;
        RECT 870.850 31.720 1239.630 31.860 ;
        RECT 870.850 31.660 871.170 31.720 ;
        RECT 1239.310 31.660 1239.630 31.720 ;
      LAYER via ;
        RECT 870.880 31.660 871.140 31.920 ;
        RECT 1239.340 31.660 1239.600 31.920 ;
      LAYER met2 ;
        RECT 1239.240 1700.340 1239.520 1704.000 ;
        RECT 1239.240 1700.000 1239.540 1700.340 ;
        RECT 1239.400 31.950 1239.540 1700.000 ;
        RECT 870.880 31.630 871.140 31.950 ;
        RECT 1239.340 31.630 1239.600 31.950 ;
        RECT 870.940 2.400 871.080 31.630 ;
        RECT 870.730 -4.800 871.290 2.400 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 888.790 32.200 889.110 32.260 ;
        RECT 1240.690 32.200 1241.010 32.260 ;
        RECT 888.790 32.060 1241.010 32.200 ;
        RECT 888.790 32.000 889.110 32.060 ;
        RECT 1240.690 32.000 1241.010 32.060 ;
      LAYER via ;
        RECT 888.820 32.000 889.080 32.260 ;
        RECT 1240.720 32.000 1240.980 32.260 ;
      LAYER met2 ;
        RECT 1241.080 1700.410 1241.360 1704.000 ;
        RECT 1240.780 1700.270 1241.360 1700.410 ;
        RECT 1240.780 32.290 1240.920 1700.270 ;
        RECT 1241.080 1700.000 1241.360 1700.270 ;
        RECT 888.820 31.970 889.080 32.290 ;
        RECT 1240.720 31.970 1240.980 32.290 ;
        RECT 888.880 2.400 889.020 31.970 ;
        RECT 888.670 -4.800 889.230 2.400 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 906.730 32.540 907.050 32.600 ;
        RECT 1242.990 32.540 1243.310 32.600 ;
        RECT 906.730 32.400 1243.310 32.540 ;
        RECT 906.730 32.340 907.050 32.400 ;
        RECT 1242.990 32.340 1243.310 32.400 ;
      LAYER via ;
        RECT 906.760 32.340 907.020 32.600 ;
        RECT 1243.020 32.340 1243.280 32.600 ;
      LAYER met2 ;
        RECT 1242.920 1700.340 1243.200 1704.000 ;
        RECT 1242.920 1700.000 1243.220 1700.340 ;
        RECT 1243.080 32.630 1243.220 1700.000 ;
        RECT 906.760 32.310 907.020 32.630 ;
        RECT 1243.020 32.310 1243.280 32.630 ;
        RECT 906.820 2.400 906.960 32.310 ;
        RECT 906.610 -4.800 907.170 2.400 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 924.210 32.880 924.530 32.940 ;
        RECT 1243.450 32.880 1243.770 32.940 ;
        RECT 924.210 32.740 1243.770 32.880 ;
        RECT 924.210 32.680 924.530 32.740 ;
        RECT 1243.450 32.680 1243.770 32.740 ;
      LAYER via ;
        RECT 924.240 32.680 924.500 32.940 ;
        RECT 1243.480 32.680 1243.740 32.940 ;
      LAYER met2 ;
        RECT 1244.760 1700.410 1245.040 1704.000 ;
        RECT 1244.460 1700.270 1245.040 1700.410 ;
        RECT 1244.460 1677.970 1244.600 1700.270 ;
        RECT 1244.760 1700.000 1245.040 1700.270 ;
        RECT 1243.540 1677.830 1244.600 1677.970 ;
        RECT 1243.540 32.970 1243.680 1677.830 ;
        RECT 924.240 32.650 924.500 32.970 ;
        RECT 1243.480 32.650 1243.740 32.970 ;
        RECT 924.300 2.400 924.440 32.650 ;
        RECT 924.090 -4.800 924.650 2.400 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1244.830 1678.480 1245.150 1678.540 ;
        RECT 1246.670 1678.480 1246.990 1678.540 ;
        RECT 1244.830 1678.340 1246.990 1678.480 ;
        RECT 1244.830 1678.280 1245.150 1678.340 ;
        RECT 1246.670 1678.280 1246.990 1678.340 ;
        RECT 942.150 33.220 942.470 33.280 ;
        RECT 1243.910 33.220 1244.230 33.280 ;
        RECT 942.150 33.080 1244.230 33.220 ;
        RECT 942.150 33.020 942.470 33.080 ;
        RECT 1243.910 33.020 1244.230 33.080 ;
      LAYER via ;
        RECT 1244.860 1678.280 1245.120 1678.540 ;
        RECT 1246.700 1678.280 1246.960 1678.540 ;
        RECT 942.180 33.020 942.440 33.280 ;
        RECT 1243.940 33.020 1244.200 33.280 ;
      LAYER met2 ;
        RECT 1246.600 1700.340 1246.880 1704.000 ;
        RECT 1246.600 1700.000 1246.900 1700.340 ;
        RECT 1246.760 1678.570 1246.900 1700.000 ;
        RECT 1244.860 1678.250 1245.120 1678.570 ;
        RECT 1246.700 1678.250 1246.960 1678.570 ;
        RECT 1244.920 1677.290 1245.060 1678.250 ;
        RECT 1244.000 1677.150 1245.060 1677.290 ;
        RECT 1244.000 33.310 1244.140 1677.150 ;
        RECT 942.180 32.990 942.440 33.310 ;
        RECT 1243.940 32.990 1244.200 33.310 ;
        RECT 942.240 2.400 942.380 32.990 ;
        RECT 942.030 -4.800 942.590 2.400 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1243.985 410.465 1244.155 434.775 ;
      LAYER mcon ;
        RECT 1243.985 434.605 1244.155 434.775 ;
      LAYER met1 ;
        RECT 1244.370 1676.780 1244.690 1676.840 ;
        RECT 1248.510 1676.780 1248.830 1676.840 ;
        RECT 1244.370 1676.640 1248.830 1676.780 ;
        RECT 1244.370 1676.580 1244.690 1676.640 ;
        RECT 1248.510 1676.580 1248.830 1676.640 ;
        RECT 1243.925 434.760 1244.215 434.805 ;
        RECT 1244.370 434.760 1244.690 434.820 ;
        RECT 1243.925 434.620 1244.690 434.760 ;
        RECT 1243.925 434.575 1244.215 434.620 ;
        RECT 1244.370 434.560 1244.690 434.620 ;
        RECT 1243.925 410.620 1244.215 410.665 ;
        RECT 1244.370 410.620 1244.690 410.680 ;
        RECT 1243.925 410.480 1244.690 410.620 ;
        RECT 1243.925 410.435 1244.215 410.480 ;
        RECT 1244.370 410.420 1244.690 410.480 ;
        RECT 960.090 33.560 960.410 33.620 ;
        RECT 1244.370 33.560 1244.690 33.620 ;
        RECT 960.090 33.420 1244.690 33.560 ;
        RECT 960.090 33.360 960.410 33.420 ;
        RECT 1244.370 33.360 1244.690 33.420 ;
      LAYER via ;
        RECT 1244.400 1676.580 1244.660 1676.840 ;
        RECT 1248.540 1676.580 1248.800 1676.840 ;
        RECT 1244.400 434.560 1244.660 434.820 ;
        RECT 1244.400 410.420 1244.660 410.680 ;
        RECT 960.120 33.360 960.380 33.620 ;
        RECT 1244.400 33.360 1244.660 33.620 ;
      LAYER met2 ;
        RECT 1248.440 1700.340 1248.720 1704.000 ;
        RECT 1248.440 1700.000 1248.740 1700.340 ;
        RECT 1248.600 1676.870 1248.740 1700.000 ;
        RECT 1244.400 1676.550 1244.660 1676.870 ;
        RECT 1248.540 1676.550 1248.800 1676.870 ;
        RECT 1244.460 530.925 1244.600 1676.550 ;
        RECT 1244.390 530.555 1244.670 530.925 ;
        RECT 1244.850 529.195 1245.130 529.565 ;
        RECT 1244.920 507.010 1245.060 529.195 ;
        RECT 1244.460 506.870 1245.060 507.010 ;
        RECT 1244.460 434.850 1244.600 506.870 ;
        RECT 1244.400 434.530 1244.660 434.850 ;
        RECT 1244.400 410.390 1244.660 410.710 ;
        RECT 1244.460 33.650 1244.600 410.390 ;
        RECT 960.120 33.330 960.380 33.650 ;
        RECT 1244.400 33.330 1244.660 33.650 ;
        RECT 960.180 2.400 960.320 33.330 ;
        RECT 959.970 -4.800 960.530 2.400 ;
      LAYER via2 ;
        RECT 1244.390 530.600 1244.670 530.880 ;
        RECT 1244.850 529.240 1245.130 529.520 ;
      LAYER met3 ;
        RECT 1244.365 530.890 1244.695 530.905 ;
        RECT 1244.365 530.590 1245.370 530.890 ;
        RECT 1244.365 530.575 1244.695 530.590 ;
        RECT 1245.070 529.545 1245.370 530.590 ;
        RECT 1244.825 529.230 1245.370 529.545 ;
        RECT 1244.825 529.215 1245.155 529.230 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 978.030 33.900 978.350 33.960 ;
        RECT 1251.730 33.900 1252.050 33.960 ;
        RECT 978.030 33.760 1252.050 33.900 ;
        RECT 978.030 33.700 978.350 33.760 ;
        RECT 1251.730 33.700 1252.050 33.760 ;
      LAYER via ;
        RECT 978.060 33.700 978.320 33.960 ;
        RECT 1251.760 33.700 1252.020 33.960 ;
      LAYER met2 ;
        RECT 1250.280 1700.340 1250.560 1704.000 ;
        RECT 1250.280 1700.000 1250.580 1700.340 ;
        RECT 1250.440 1677.970 1250.580 1700.000 ;
        RECT 1250.440 1677.830 1251.960 1677.970 ;
        RECT 1251.820 33.990 1251.960 1677.830 ;
        RECT 978.060 33.670 978.320 33.990 ;
        RECT 1251.760 33.670 1252.020 33.990 ;
        RECT 978.120 2.400 978.260 33.670 ;
        RECT 977.910 -4.800 978.470 2.400 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 656.950 31.180 657.270 31.240 ;
        RECT 1215.850 31.180 1216.170 31.240 ;
        RECT 656.950 31.040 1216.170 31.180 ;
        RECT 656.950 30.980 657.270 31.040 ;
        RECT 1215.850 30.980 1216.170 31.040 ;
      LAYER via ;
        RECT 656.980 30.980 657.240 31.240 ;
        RECT 1215.880 30.980 1216.140 31.240 ;
      LAYER met2 ;
        RECT 1217.160 1700.340 1217.440 1704.000 ;
        RECT 1217.160 1700.000 1217.460 1700.340 ;
        RECT 1217.320 1659.610 1217.460 1700.000 ;
        RECT 1215.940 1659.470 1217.460 1659.610 ;
        RECT 1215.940 31.270 1216.080 1659.470 ;
        RECT 656.980 30.950 657.240 31.270 ;
        RECT 1215.880 30.950 1216.140 31.270 ;
        RECT 657.040 2.400 657.180 30.950 ;
        RECT 656.830 -4.800 657.390 2.400 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1248.970 1676.780 1249.290 1676.840 ;
        RECT 1252.190 1676.780 1252.510 1676.840 ;
        RECT 1248.970 1676.640 1252.510 1676.780 ;
        RECT 1248.970 1676.580 1249.290 1676.640 ;
        RECT 1252.190 1676.580 1252.510 1676.640 ;
        RECT 995.970 34.240 996.290 34.300 ;
        RECT 1248.970 34.240 1249.290 34.300 ;
        RECT 995.970 34.100 1249.290 34.240 ;
        RECT 995.970 34.040 996.290 34.100 ;
        RECT 1248.970 34.040 1249.290 34.100 ;
      LAYER via ;
        RECT 1249.000 1676.580 1249.260 1676.840 ;
        RECT 1252.220 1676.580 1252.480 1676.840 ;
        RECT 996.000 34.040 996.260 34.300 ;
        RECT 1249.000 34.040 1249.260 34.300 ;
      LAYER met2 ;
        RECT 1252.120 1700.340 1252.400 1704.000 ;
        RECT 1252.120 1700.000 1252.420 1700.340 ;
        RECT 1252.280 1676.870 1252.420 1700.000 ;
        RECT 1249.000 1676.550 1249.260 1676.870 ;
        RECT 1252.220 1676.550 1252.480 1676.870 ;
        RECT 1249.060 34.330 1249.200 1676.550 ;
        RECT 996.000 34.010 996.260 34.330 ;
        RECT 1249.000 34.010 1249.260 34.330 ;
        RECT 996.060 2.400 996.200 34.010 ;
        RECT 995.850 -4.800 996.410 2.400 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1013.450 30.500 1013.770 30.560 ;
        RECT 1254.030 30.500 1254.350 30.560 ;
        RECT 1013.450 30.360 1254.350 30.500 ;
        RECT 1013.450 30.300 1013.770 30.360 ;
        RECT 1254.030 30.300 1254.350 30.360 ;
      LAYER via ;
        RECT 1013.480 30.300 1013.740 30.560 ;
        RECT 1254.060 30.300 1254.320 30.560 ;
      LAYER met2 ;
        RECT 1253.960 1700.340 1254.240 1704.000 ;
        RECT 1253.960 1700.000 1254.260 1700.340 ;
        RECT 1254.120 30.590 1254.260 1700.000 ;
        RECT 1013.480 30.270 1013.740 30.590 ;
        RECT 1254.060 30.270 1254.320 30.590 ;
        RECT 1013.540 2.400 1013.680 30.270 ;
        RECT 1013.330 -4.800 1013.890 2.400 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1034.610 1646.860 1034.930 1646.920 ;
        RECT 1255.870 1646.860 1256.190 1646.920 ;
        RECT 1034.610 1646.720 1256.190 1646.860 ;
        RECT 1034.610 1646.660 1034.930 1646.720 ;
        RECT 1255.870 1646.660 1256.190 1646.720 ;
        RECT 1031.390 2.960 1031.710 3.020 ;
        RECT 1034.610 2.960 1034.930 3.020 ;
        RECT 1031.390 2.820 1034.930 2.960 ;
        RECT 1031.390 2.760 1031.710 2.820 ;
        RECT 1034.610 2.760 1034.930 2.820 ;
      LAYER via ;
        RECT 1034.640 1646.660 1034.900 1646.920 ;
        RECT 1255.900 1646.660 1256.160 1646.920 ;
        RECT 1031.420 2.760 1031.680 3.020 ;
        RECT 1034.640 2.760 1034.900 3.020 ;
      LAYER met2 ;
        RECT 1255.800 1700.340 1256.080 1704.000 ;
        RECT 1255.800 1700.000 1256.100 1700.340 ;
        RECT 1255.960 1646.950 1256.100 1700.000 ;
        RECT 1034.640 1646.630 1034.900 1646.950 ;
        RECT 1255.900 1646.630 1256.160 1646.950 ;
        RECT 1034.700 3.050 1034.840 1646.630 ;
        RECT 1031.420 2.730 1031.680 3.050 ;
        RECT 1034.640 2.730 1034.900 3.050 ;
        RECT 1031.480 2.400 1031.620 2.730 ;
        RECT 1031.270 -4.800 1031.830 2.400 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1257.785 1654.185 1257.955 1678.495 ;
      LAYER mcon ;
        RECT 1257.785 1678.325 1257.955 1678.495 ;
      LAYER met1 ;
        RECT 1257.710 1678.480 1258.030 1678.540 ;
        RECT 1257.515 1678.340 1258.030 1678.480 ;
        RECT 1257.710 1678.280 1258.030 1678.340 ;
        RECT 1055.310 1654.340 1055.630 1654.400 ;
        RECT 1257.725 1654.340 1258.015 1654.385 ;
        RECT 1055.310 1654.200 1258.015 1654.340 ;
        RECT 1055.310 1654.140 1055.630 1654.200 ;
        RECT 1257.725 1654.155 1258.015 1654.200 ;
        RECT 1049.330 20.980 1049.650 21.040 ;
        RECT 1055.310 20.980 1055.630 21.040 ;
        RECT 1049.330 20.840 1055.630 20.980 ;
        RECT 1049.330 20.780 1049.650 20.840 ;
        RECT 1055.310 20.780 1055.630 20.840 ;
      LAYER via ;
        RECT 1257.740 1678.280 1258.000 1678.540 ;
        RECT 1055.340 1654.140 1055.600 1654.400 ;
        RECT 1049.360 20.780 1049.620 21.040 ;
        RECT 1055.340 20.780 1055.600 21.040 ;
      LAYER met2 ;
        RECT 1257.640 1700.340 1257.920 1704.000 ;
        RECT 1257.640 1700.000 1257.940 1700.340 ;
        RECT 1257.800 1678.570 1257.940 1700.000 ;
        RECT 1257.740 1678.250 1258.000 1678.570 ;
        RECT 1055.340 1654.110 1055.600 1654.430 ;
        RECT 1055.400 21.070 1055.540 1654.110 ;
        RECT 1049.360 20.750 1049.620 21.070 ;
        RECT 1055.340 20.750 1055.600 21.070 ;
        RECT 1049.420 2.400 1049.560 20.750 ;
        RECT 1049.210 -4.800 1049.770 2.400 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1069.110 1625.780 1069.430 1625.840 ;
        RECT 1257.710 1625.780 1258.030 1625.840 ;
        RECT 1069.110 1625.640 1258.030 1625.780 ;
        RECT 1069.110 1625.580 1069.430 1625.640 ;
        RECT 1257.710 1625.580 1258.030 1625.640 ;
      LAYER via ;
        RECT 1069.140 1625.580 1069.400 1625.840 ;
        RECT 1257.740 1625.580 1258.000 1625.840 ;
      LAYER met2 ;
        RECT 1259.480 1700.410 1259.760 1704.000 ;
        RECT 1259.180 1700.270 1259.760 1700.410 ;
        RECT 1259.180 1677.970 1259.320 1700.270 ;
        RECT 1259.480 1700.000 1259.760 1700.270 ;
        RECT 1257.800 1677.830 1259.320 1677.970 ;
        RECT 1257.800 1625.870 1257.940 1677.830 ;
        RECT 1069.140 1625.550 1069.400 1625.870 ;
        RECT 1257.740 1625.550 1258.000 1625.870 ;
        RECT 1069.200 18.090 1069.340 1625.550 ;
        RECT 1067.360 17.950 1069.340 18.090 ;
        RECT 1067.360 2.400 1067.500 17.950 ;
        RECT 1067.150 -4.800 1067.710 2.400 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1257.250 1678.820 1257.570 1678.880 ;
        RECT 1260.930 1678.820 1261.250 1678.880 ;
        RECT 1257.250 1678.680 1261.250 1678.820 ;
        RECT 1257.250 1678.620 1257.570 1678.680 ;
        RECT 1260.930 1678.620 1261.250 1678.680 ;
        RECT 1089.810 1618.980 1090.130 1619.040 ;
        RECT 1257.250 1618.980 1257.570 1619.040 ;
        RECT 1089.810 1618.840 1257.570 1618.980 ;
        RECT 1089.810 1618.780 1090.130 1618.840 ;
        RECT 1257.250 1618.780 1257.570 1618.840 ;
      LAYER via ;
        RECT 1257.280 1678.620 1257.540 1678.880 ;
        RECT 1260.960 1678.620 1261.220 1678.880 ;
        RECT 1089.840 1618.780 1090.100 1619.040 ;
        RECT 1257.280 1618.780 1257.540 1619.040 ;
      LAYER met2 ;
        RECT 1261.320 1700.410 1261.600 1704.000 ;
        RECT 1261.020 1700.270 1261.600 1700.410 ;
        RECT 1261.020 1678.910 1261.160 1700.270 ;
        RECT 1261.320 1700.000 1261.600 1700.270 ;
        RECT 1257.280 1678.590 1257.540 1678.910 ;
        RECT 1260.960 1678.590 1261.220 1678.910 ;
        RECT 1257.340 1619.070 1257.480 1678.590 ;
        RECT 1089.840 1618.750 1090.100 1619.070 ;
        RECT 1257.280 1618.750 1257.540 1619.070 ;
        RECT 1089.900 18.090 1090.040 1618.750 ;
        RECT 1085.300 17.950 1090.040 18.090 ;
        RECT 1085.300 2.400 1085.440 17.950 ;
        RECT 1085.090 -4.800 1085.650 2.400 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1103.610 1682.220 1103.930 1682.280 ;
        RECT 1263.230 1682.220 1263.550 1682.280 ;
        RECT 1103.610 1682.080 1263.550 1682.220 ;
        RECT 1103.610 1682.020 1103.930 1682.080 ;
        RECT 1263.230 1682.020 1263.550 1682.080 ;
      LAYER via ;
        RECT 1103.640 1682.020 1103.900 1682.280 ;
        RECT 1263.260 1682.020 1263.520 1682.280 ;
      LAYER met2 ;
        RECT 1263.160 1700.340 1263.440 1704.000 ;
        RECT 1263.160 1700.000 1263.460 1700.340 ;
        RECT 1263.320 1682.310 1263.460 1700.000 ;
        RECT 1103.640 1681.990 1103.900 1682.310 ;
        RECT 1263.260 1681.990 1263.520 1682.310 ;
        RECT 1103.700 16.730 1103.840 1681.990 ;
        RECT 1102.780 16.590 1103.840 16.730 ;
        RECT 1102.780 2.400 1102.920 16.590 ;
        RECT 1102.570 -4.800 1103.130 2.400 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1124.310 1661.140 1124.630 1661.200 ;
        RECT 1265.070 1661.140 1265.390 1661.200 ;
        RECT 1124.310 1661.000 1265.390 1661.140 ;
        RECT 1124.310 1660.940 1124.630 1661.000 ;
        RECT 1265.070 1660.940 1265.390 1661.000 ;
      LAYER via ;
        RECT 1124.340 1660.940 1124.600 1661.200 ;
        RECT 1265.100 1660.940 1265.360 1661.200 ;
      LAYER met2 ;
        RECT 1265.000 1700.340 1265.280 1704.000 ;
        RECT 1265.000 1700.000 1265.300 1700.340 ;
        RECT 1265.160 1661.230 1265.300 1700.000 ;
        RECT 1124.340 1660.910 1124.600 1661.230 ;
        RECT 1265.100 1660.910 1265.360 1661.230 ;
        RECT 1124.400 16.730 1124.540 1660.910 ;
        RECT 1120.720 16.590 1124.540 16.730 ;
        RECT 1120.720 2.400 1120.860 16.590 ;
        RECT 1120.510 -4.800 1121.070 2.400 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1145.010 1675.760 1145.330 1675.820 ;
        RECT 1266.910 1675.760 1267.230 1675.820 ;
        RECT 1145.010 1675.620 1267.230 1675.760 ;
        RECT 1145.010 1675.560 1145.330 1675.620 ;
        RECT 1266.910 1675.560 1267.230 1675.620 ;
        RECT 1138.570 20.980 1138.890 21.040 ;
        RECT 1145.010 20.980 1145.330 21.040 ;
        RECT 1138.570 20.840 1145.330 20.980 ;
        RECT 1138.570 20.780 1138.890 20.840 ;
        RECT 1145.010 20.780 1145.330 20.840 ;
      LAYER via ;
        RECT 1145.040 1675.560 1145.300 1675.820 ;
        RECT 1266.940 1675.560 1267.200 1675.820 ;
        RECT 1138.600 20.780 1138.860 21.040 ;
        RECT 1145.040 20.780 1145.300 21.040 ;
      LAYER met2 ;
        RECT 1266.840 1700.340 1267.120 1704.000 ;
        RECT 1266.840 1700.000 1267.140 1700.340 ;
        RECT 1267.000 1675.850 1267.140 1700.000 ;
        RECT 1145.040 1675.530 1145.300 1675.850 ;
        RECT 1266.940 1675.530 1267.200 1675.850 ;
        RECT 1145.100 21.070 1145.240 1675.530 ;
        RECT 1138.600 20.750 1138.860 21.070 ;
        RECT 1145.040 20.750 1145.300 21.070 ;
        RECT 1138.660 2.400 1138.800 20.750 ;
        RECT 1138.450 -4.800 1139.010 2.400 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1261.390 1684.260 1261.710 1684.320 ;
        RECT 1268.750 1684.260 1269.070 1684.320 ;
        RECT 1261.390 1684.120 1269.070 1684.260 ;
        RECT 1261.390 1684.060 1261.710 1684.120 ;
        RECT 1268.750 1684.060 1269.070 1684.120 ;
        RECT 1261.390 1678.280 1261.710 1678.540 ;
        RECT 1259.550 1677.460 1259.870 1677.520 ;
        RECT 1261.480 1677.460 1261.620 1678.280 ;
        RECT 1259.550 1677.320 1261.620 1677.460 ;
        RECT 1259.550 1677.260 1259.870 1677.320 ;
        RECT 1158.810 51.580 1159.130 51.640 ;
        RECT 1259.550 51.580 1259.870 51.640 ;
        RECT 1158.810 51.440 1259.870 51.580 ;
        RECT 1158.810 51.380 1159.130 51.440 ;
        RECT 1259.550 51.380 1259.870 51.440 ;
        RECT 1156.510 17.580 1156.830 17.640 ;
        RECT 1158.810 17.580 1159.130 17.640 ;
        RECT 1156.510 17.440 1159.130 17.580 ;
        RECT 1156.510 17.380 1156.830 17.440 ;
        RECT 1158.810 17.380 1159.130 17.440 ;
      LAYER via ;
        RECT 1261.420 1684.060 1261.680 1684.320 ;
        RECT 1268.780 1684.060 1269.040 1684.320 ;
        RECT 1261.420 1678.280 1261.680 1678.540 ;
        RECT 1259.580 1677.260 1259.840 1677.520 ;
        RECT 1158.840 51.380 1159.100 51.640 ;
        RECT 1259.580 51.380 1259.840 51.640 ;
        RECT 1156.540 17.380 1156.800 17.640 ;
        RECT 1158.840 17.380 1159.100 17.640 ;
      LAYER met2 ;
        RECT 1268.680 1700.340 1268.960 1704.000 ;
        RECT 1268.680 1700.000 1268.980 1700.340 ;
        RECT 1268.840 1684.350 1268.980 1700.000 ;
        RECT 1261.420 1684.030 1261.680 1684.350 ;
        RECT 1268.780 1684.030 1269.040 1684.350 ;
        RECT 1261.480 1678.570 1261.620 1684.030 ;
        RECT 1261.420 1678.250 1261.680 1678.570 ;
        RECT 1259.580 1677.230 1259.840 1677.550 ;
        RECT 1259.640 51.670 1259.780 1677.230 ;
        RECT 1158.840 51.350 1159.100 51.670 ;
        RECT 1259.580 51.350 1259.840 51.670 ;
        RECT 1158.900 17.670 1159.040 51.350 ;
        RECT 1156.540 17.350 1156.800 17.670 ;
        RECT 1158.840 17.350 1159.100 17.670 ;
        RECT 1156.600 2.400 1156.740 17.350 ;
        RECT 1156.390 -4.800 1156.950 2.400 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1216.310 1656.720 1216.630 1656.780 ;
        RECT 1219.070 1656.720 1219.390 1656.780 ;
        RECT 1216.310 1656.580 1219.390 1656.720 ;
        RECT 1216.310 1656.520 1216.630 1656.580 ;
        RECT 1219.070 1656.520 1219.390 1656.580 ;
        RECT 674.430 31.520 674.750 31.580 ;
        RECT 1216.310 31.520 1216.630 31.580 ;
        RECT 674.430 31.380 1216.630 31.520 ;
        RECT 674.430 31.320 674.750 31.380 ;
        RECT 1216.310 31.320 1216.630 31.380 ;
      LAYER via ;
        RECT 1216.340 1656.520 1216.600 1656.780 ;
        RECT 1219.100 1656.520 1219.360 1656.780 ;
        RECT 674.460 31.320 674.720 31.580 ;
        RECT 1216.340 31.320 1216.600 31.580 ;
      LAYER met2 ;
        RECT 1219.000 1700.340 1219.280 1704.000 ;
        RECT 1219.000 1700.000 1219.300 1700.340 ;
        RECT 1219.160 1656.810 1219.300 1700.000 ;
        RECT 1216.340 1656.490 1216.600 1656.810 ;
        RECT 1219.100 1656.490 1219.360 1656.810 ;
        RECT 1216.400 31.610 1216.540 1656.490 ;
        RECT 674.460 31.290 674.720 31.610 ;
        RECT 1216.340 31.290 1216.600 31.610 ;
        RECT 674.520 2.400 674.660 31.290 ;
        RECT 674.310 -4.800 674.870 2.400 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1270.590 1677.600 1270.910 1677.860 ;
        RECT 1270.680 1676.100 1270.820 1677.600 ;
        RECT 1272.430 1676.100 1272.750 1676.160 ;
        RECT 1270.680 1675.960 1272.750 1676.100 ;
        RECT 1272.430 1675.900 1272.750 1675.960 ;
        RECT 1173.990 30.840 1174.310 30.900 ;
        RECT 1272.430 30.840 1272.750 30.900 ;
        RECT 1173.990 30.700 1272.750 30.840 ;
        RECT 1173.990 30.640 1174.310 30.700 ;
        RECT 1272.430 30.640 1272.750 30.700 ;
      LAYER via ;
        RECT 1270.620 1677.600 1270.880 1677.860 ;
        RECT 1272.460 1675.900 1272.720 1676.160 ;
        RECT 1174.020 30.640 1174.280 30.900 ;
        RECT 1272.460 30.640 1272.720 30.900 ;
      LAYER met2 ;
        RECT 1270.520 1700.340 1270.800 1704.000 ;
        RECT 1270.520 1700.000 1270.820 1700.340 ;
        RECT 1270.680 1677.890 1270.820 1700.000 ;
        RECT 1270.620 1677.570 1270.880 1677.890 ;
        RECT 1272.460 1675.870 1272.720 1676.190 ;
        RECT 1272.520 30.930 1272.660 1675.870 ;
        RECT 1174.020 30.610 1174.280 30.930 ;
        RECT 1272.460 30.610 1272.720 30.930 ;
        RECT 1174.080 2.400 1174.220 30.610 ;
        RECT 1173.870 -4.800 1174.430 2.400 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1191.930 30.160 1192.250 30.220 ;
        RECT 1272.890 30.160 1273.210 30.220 ;
        RECT 1191.930 30.020 1273.210 30.160 ;
        RECT 1191.930 29.960 1192.250 30.020 ;
        RECT 1272.890 29.960 1273.210 30.020 ;
      LAYER via ;
        RECT 1191.960 29.960 1192.220 30.220 ;
        RECT 1272.920 29.960 1273.180 30.220 ;
      LAYER met2 ;
        RECT 1272.360 1700.340 1272.640 1704.000 ;
        RECT 1272.360 1700.000 1272.660 1700.340 ;
        RECT 1272.520 1676.610 1272.660 1700.000 ;
        RECT 1272.520 1676.470 1273.120 1676.610 ;
        RECT 1272.980 30.250 1273.120 1676.470 ;
        RECT 1191.960 29.930 1192.220 30.250 ;
        RECT 1272.920 29.930 1273.180 30.250 ;
        RECT 1192.020 2.400 1192.160 29.930 ;
        RECT 1191.810 -4.800 1192.370 2.400 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1258.705 1490.645 1258.875 1538.755 ;
        RECT 1258.245 1435.225 1258.415 1462.595 ;
        RECT 1259.165 1110.865 1259.335 1124.975 ;
        RECT 1258.245 662.405 1258.415 685.695 ;
        RECT 1258.705 503.625 1258.875 552.075 ;
        RECT 1258.705 372.725 1258.875 420.835 ;
      LAYER mcon ;
        RECT 1258.705 1538.585 1258.875 1538.755 ;
        RECT 1258.245 1462.425 1258.415 1462.595 ;
        RECT 1259.165 1124.805 1259.335 1124.975 ;
        RECT 1258.245 685.525 1258.415 685.695 ;
        RECT 1258.705 551.905 1258.875 552.075 ;
        RECT 1258.705 420.665 1258.875 420.835 ;
      LAYER met1 ;
        RECT 1256.330 1685.960 1256.650 1686.020 ;
        RECT 1274.270 1685.960 1274.590 1686.020 ;
        RECT 1256.330 1685.820 1274.590 1685.960 ;
        RECT 1256.330 1685.760 1256.650 1685.820 ;
        RECT 1274.270 1685.760 1274.590 1685.820 ;
        RECT 1256.330 1631.900 1256.650 1631.960 ;
        RECT 1258.630 1631.900 1258.950 1631.960 ;
        RECT 1256.330 1631.760 1258.950 1631.900 ;
        RECT 1256.330 1631.700 1256.650 1631.760 ;
        RECT 1258.630 1631.700 1258.950 1631.760 ;
        RECT 1258.645 1538.740 1258.935 1538.785 ;
        RECT 1259.090 1538.740 1259.410 1538.800 ;
        RECT 1258.645 1538.600 1259.410 1538.740 ;
        RECT 1258.645 1538.555 1258.935 1538.600 ;
        RECT 1259.090 1538.540 1259.410 1538.600 ;
        RECT 1258.630 1490.800 1258.950 1490.860 ;
        RECT 1258.435 1490.660 1258.950 1490.800 ;
        RECT 1258.630 1490.600 1258.950 1490.660 ;
        RECT 1258.185 1462.580 1258.475 1462.625 ;
        RECT 1258.630 1462.580 1258.950 1462.640 ;
        RECT 1258.185 1462.440 1258.950 1462.580 ;
        RECT 1258.185 1462.395 1258.475 1462.440 ;
        RECT 1258.630 1462.380 1258.950 1462.440 ;
        RECT 1258.170 1435.380 1258.490 1435.440 ;
        RECT 1257.975 1435.240 1258.490 1435.380 ;
        RECT 1258.170 1435.180 1258.490 1435.240 ;
        RECT 1256.790 1304.140 1257.110 1304.200 ;
        RECT 1258.170 1304.140 1258.490 1304.200 ;
        RECT 1256.790 1304.000 1258.490 1304.140 ;
        RECT 1256.790 1303.940 1257.110 1304.000 ;
        RECT 1258.170 1303.940 1258.490 1304.000 ;
        RECT 1256.790 1266.060 1257.110 1266.120 ;
        RECT 1257.710 1266.060 1258.030 1266.120 ;
        RECT 1256.790 1265.920 1258.030 1266.060 ;
        RECT 1256.790 1265.860 1257.110 1265.920 ;
        RECT 1257.710 1265.860 1258.030 1265.920 ;
        RECT 1257.710 1224.920 1258.030 1224.980 ;
        RECT 1258.630 1224.920 1258.950 1224.980 ;
        RECT 1257.710 1224.780 1258.950 1224.920 ;
        RECT 1257.710 1224.720 1258.030 1224.780 ;
        RECT 1258.630 1224.720 1258.950 1224.780 ;
        RECT 1259.090 1124.960 1259.410 1125.020 ;
        RECT 1258.895 1124.820 1259.410 1124.960 ;
        RECT 1259.090 1124.760 1259.410 1124.820 ;
        RECT 1259.090 1111.020 1259.410 1111.080 ;
        RECT 1258.895 1110.880 1259.410 1111.020 ;
        RECT 1259.090 1110.820 1259.410 1110.880 ;
        RECT 1257.710 1028.200 1258.030 1028.460 ;
        RECT 1257.800 1027.780 1257.940 1028.200 ;
        RECT 1257.710 1027.520 1258.030 1027.780 ;
        RECT 1258.170 989.640 1258.490 989.700 ;
        RECT 1258.630 989.640 1258.950 989.700 ;
        RECT 1258.170 989.500 1258.950 989.640 ;
        RECT 1258.170 989.440 1258.490 989.500 ;
        RECT 1258.630 989.440 1258.950 989.500 ;
        RECT 1258.170 855.340 1258.490 855.400 ;
        RECT 1259.090 855.340 1259.410 855.400 ;
        RECT 1258.170 855.200 1259.410 855.340 ;
        RECT 1258.170 855.140 1258.490 855.200 ;
        RECT 1259.090 855.140 1259.410 855.200 ;
        RECT 1258.630 759.120 1258.950 759.180 ;
        RECT 1259.090 759.120 1259.410 759.180 ;
        RECT 1258.630 758.980 1259.410 759.120 ;
        RECT 1258.630 758.920 1258.950 758.980 ;
        RECT 1259.090 758.920 1259.410 758.980 ;
        RECT 1258.185 685.680 1258.475 685.725 ;
        RECT 1258.630 685.680 1258.950 685.740 ;
        RECT 1258.185 685.540 1258.950 685.680 ;
        RECT 1258.185 685.495 1258.475 685.540 ;
        RECT 1258.630 685.480 1258.950 685.540 ;
        RECT 1258.170 662.560 1258.490 662.620 ;
        RECT 1257.975 662.420 1258.490 662.560 ;
        RECT 1258.170 662.360 1258.490 662.420 ;
        RECT 1258.170 621.220 1258.490 621.480 ;
        RECT 1258.260 620.400 1258.400 621.220 ;
        RECT 1258.630 620.400 1258.950 620.460 ;
        RECT 1258.260 620.260 1258.950 620.400 ;
        RECT 1258.630 620.200 1258.950 620.260 ;
        RECT 1258.645 552.060 1258.935 552.105 ;
        RECT 1259.090 552.060 1259.410 552.120 ;
        RECT 1258.645 551.920 1259.410 552.060 ;
        RECT 1258.645 551.875 1258.935 551.920 ;
        RECT 1259.090 551.860 1259.410 551.920 ;
        RECT 1258.630 503.780 1258.950 503.840 ;
        RECT 1258.435 503.640 1258.950 503.780 ;
        RECT 1258.630 503.580 1258.950 503.640 ;
        RECT 1258.630 420.820 1258.950 420.880 ;
        RECT 1258.435 420.680 1258.950 420.820 ;
        RECT 1258.630 420.620 1258.950 420.680 ;
        RECT 1258.645 372.880 1258.935 372.925 ;
        RECT 1259.090 372.880 1259.410 372.940 ;
        RECT 1258.645 372.740 1259.410 372.880 ;
        RECT 1258.645 372.695 1258.935 372.740 ;
        RECT 1259.090 372.680 1259.410 372.740 ;
        RECT 1258.170 331.400 1258.490 331.460 ;
        RECT 1259.090 331.400 1259.410 331.460 ;
        RECT 1258.170 331.260 1259.410 331.400 ;
        RECT 1258.170 331.200 1258.490 331.260 ;
        RECT 1259.090 331.200 1259.410 331.260 ;
        RECT 1257.710 241.640 1258.030 241.700 ;
        RECT 1258.170 241.640 1258.490 241.700 ;
        RECT 1257.710 241.500 1258.490 241.640 ;
        RECT 1257.710 241.440 1258.030 241.500 ;
        RECT 1258.170 241.440 1258.490 241.500 ;
        RECT 1257.710 224.980 1258.030 225.040 ;
        RECT 1258.630 224.980 1258.950 225.040 ;
        RECT 1257.710 224.840 1258.950 224.980 ;
        RECT 1257.710 224.780 1258.030 224.840 ;
        RECT 1258.630 224.780 1258.950 224.840 ;
        RECT 1258.170 90.000 1258.490 90.060 ;
        RECT 1258.630 90.000 1258.950 90.060 ;
        RECT 1258.170 89.860 1258.950 90.000 ;
        RECT 1258.170 89.800 1258.490 89.860 ;
        RECT 1258.630 89.800 1258.950 89.860 ;
        RECT 1209.870 44.780 1210.190 44.840 ;
        RECT 1258.170 44.780 1258.490 44.840 ;
        RECT 1209.870 44.640 1258.490 44.780 ;
        RECT 1209.870 44.580 1210.190 44.640 ;
        RECT 1258.170 44.580 1258.490 44.640 ;
      LAYER via ;
        RECT 1256.360 1685.760 1256.620 1686.020 ;
        RECT 1274.300 1685.760 1274.560 1686.020 ;
        RECT 1256.360 1631.700 1256.620 1631.960 ;
        RECT 1258.660 1631.700 1258.920 1631.960 ;
        RECT 1259.120 1538.540 1259.380 1538.800 ;
        RECT 1258.660 1490.600 1258.920 1490.860 ;
        RECT 1258.660 1462.380 1258.920 1462.640 ;
        RECT 1258.200 1435.180 1258.460 1435.440 ;
        RECT 1256.820 1303.940 1257.080 1304.200 ;
        RECT 1258.200 1303.940 1258.460 1304.200 ;
        RECT 1256.820 1265.860 1257.080 1266.120 ;
        RECT 1257.740 1265.860 1258.000 1266.120 ;
        RECT 1257.740 1224.720 1258.000 1224.980 ;
        RECT 1258.660 1224.720 1258.920 1224.980 ;
        RECT 1259.120 1124.760 1259.380 1125.020 ;
        RECT 1259.120 1110.820 1259.380 1111.080 ;
        RECT 1257.740 1028.200 1258.000 1028.460 ;
        RECT 1257.740 1027.520 1258.000 1027.780 ;
        RECT 1258.200 989.440 1258.460 989.700 ;
        RECT 1258.660 989.440 1258.920 989.700 ;
        RECT 1258.200 855.140 1258.460 855.400 ;
        RECT 1259.120 855.140 1259.380 855.400 ;
        RECT 1258.660 758.920 1258.920 759.180 ;
        RECT 1259.120 758.920 1259.380 759.180 ;
        RECT 1258.660 685.480 1258.920 685.740 ;
        RECT 1258.200 662.360 1258.460 662.620 ;
        RECT 1258.200 621.220 1258.460 621.480 ;
        RECT 1258.660 620.200 1258.920 620.460 ;
        RECT 1259.120 551.860 1259.380 552.120 ;
        RECT 1258.660 503.580 1258.920 503.840 ;
        RECT 1258.660 420.620 1258.920 420.880 ;
        RECT 1259.120 372.680 1259.380 372.940 ;
        RECT 1258.200 331.200 1258.460 331.460 ;
        RECT 1259.120 331.200 1259.380 331.460 ;
        RECT 1257.740 241.440 1258.000 241.700 ;
        RECT 1258.200 241.440 1258.460 241.700 ;
        RECT 1257.740 224.780 1258.000 225.040 ;
        RECT 1258.660 224.780 1258.920 225.040 ;
        RECT 1258.200 89.800 1258.460 90.060 ;
        RECT 1258.660 89.800 1258.920 90.060 ;
        RECT 1209.900 44.580 1210.160 44.840 ;
        RECT 1258.200 44.580 1258.460 44.840 ;
      LAYER met2 ;
        RECT 1274.200 1700.340 1274.480 1704.000 ;
        RECT 1274.200 1700.000 1274.500 1700.340 ;
        RECT 1274.360 1686.050 1274.500 1700.000 ;
        RECT 1256.360 1685.730 1256.620 1686.050 ;
        RECT 1274.300 1685.730 1274.560 1686.050 ;
        RECT 1256.420 1631.990 1256.560 1685.730 ;
        RECT 1256.360 1631.670 1256.620 1631.990 ;
        RECT 1258.660 1631.670 1258.920 1631.990 ;
        RECT 1258.720 1569.850 1258.860 1631.670 ;
        RECT 1258.720 1569.710 1259.320 1569.850 ;
        RECT 1259.180 1538.830 1259.320 1569.710 ;
        RECT 1259.120 1538.510 1259.380 1538.830 ;
        RECT 1258.660 1490.570 1258.920 1490.890 ;
        RECT 1258.720 1462.670 1258.860 1490.570 ;
        RECT 1258.660 1462.350 1258.920 1462.670 ;
        RECT 1258.200 1435.150 1258.460 1435.470 ;
        RECT 1258.260 1304.230 1258.400 1435.150 ;
        RECT 1256.820 1303.910 1257.080 1304.230 ;
        RECT 1258.200 1303.910 1258.460 1304.230 ;
        RECT 1256.880 1290.485 1257.020 1303.910 ;
        RECT 1256.810 1290.115 1257.090 1290.485 ;
        RECT 1256.810 1289.435 1257.090 1289.805 ;
        RECT 1256.880 1266.150 1257.020 1289.435 ;
        RECT 1256.820 1265.830 1257.080 1266.150 ;
        RECT 1257.740 1265.830 1258.000 1266.150 ;
        RECT 1257.800 1225.010 1257.940 1265.830 ;
        RECT 1257.740 1224.690 1258.000 1225.010 ;
        RECT 1258.660 1224.690 1258.920 1225.010 ;
        RECT 1258.720 1187.690 1258.860 1224.690 ;
        RECT 1258.720 1187.550 1259.320 1187.690 ;
        RECT 1259.180 1125.050 1259.320 1187.550 ;
        RECT 1259.120 1124.730 1259.380 1125.050 ;
        RECT 1259.120 1110.790 1259.380 1111.110 ;
        RECT 1259.180 1087.050 1259.320 1110.790 ;
        RECT 1257.800 1086.910 1259.320 1087.050 ;
        RECT 1257.800 1028.490 1257.940 1086.910 ;
        RECT 1257.740 1028.170 1258.000 1028.490 ;
        RECT 1257.740 1027.490 1258.000 1027.810 ;
        RECT 1257.800 1014.405 1257.940 1027.490 ;
        RECT 1257.730 1014.035 1258.010 1014.405 ;
        RECT 1258.650 1014.035 1258.930 1014.405 ;
        RECT 1258.720 989.730 1258.860 1014.035 ;
        RECT 1258.200 989.410 1258.460 989.730 ;
        RECT 1258.660 989.410 1258.920 989.730 ;
        RECT 1258.260 855.430 1258.400 989.410 ;
        RECT 1258.200 855.110 1258.460 855.430 ;
        RECT 1259.120 855.110 1259.380 855.430 ;
        RECT 1259.180 759.210 1259.320 855.110 ;
        RECT 1258.660 758.890 1258.920 759.210 ;
        RECT 1259.120 758.890 1259.380 759.210 ;
        RECT 1258.720 685.770 1258.860 758.890 ;
        RECT 1258.660 685.450 1258.920 685.770 ;
        RECT 1258.200 662.330 1258.460 662.650 ;
        RECT 1258.260 621.510 1258.400 662.330 ;
        RECT 1258.200 621.190 1258.460 621.510 ;
        RECT 1258.660 620.170 1258.920 620.490 ;
        RECT 1258.720 552.570 1258.860 620.170 ;
        RECT 1258.720 552.430 1259.320 552.570 ;
        RECT 1259.180 552.150 1259.320 552.430 ;
        RECT 1259.120 551.830 1259.380 552.150 ;
        RECT 1258.720 503.870 1258.860 504.025 ;
        RECT 1258.660 503.610 1258.920 503.870 ;
        RECT 1258.660 503.550 1259.320 503.610 ;
        RECT 1258.720 503.470 1259.320 503.550 ;
        RECT 1259.180 479.810 1259.320 503.470 ;
        RECT 1258.720 479.670 1259.320 479.810 ;
        RECT 1258.720 420.910 1258.860 479.670 ;
        RECT 1258.660 420.590 1258.920 420.910 ;
        RECT 1259.120 372.650 1259.380 372.970 ;
        RECT 1259.180 331.490 1259.320 372.650 ;
        RECT 1258.200 331.170 1258.460 331.490 ;
        RECT 1259.120 331.170 1259.380 331.490 ;
        RECT 1258.260 241.730 1258.400 331.170 ;
        RECT 1257.740 241.410 1258.000 241.730 ;
        RECT 1258.200 241.410 1258.460 241.730 ;
        RECT 1257.800 225.070 1257.940 241.410 ;
        RECT 1257.740 224.750 1258.000 225.070 ;
        RECT 1258.660 224.750 1258.920 225.070 ;
        RECT 1258.720 90.090 1258.860 224.750 ;
        RECT 1258.200 89.770 1258.460 90.090 ;
        RECT 1258.660 89.770 1258.920 90.090 ;
        RECT 1258.260 44.870 1258.400 89.770 ;
        RECT 1209.900 44.550 1210.160 44.870 ;
        RECT 1258.200 44.550 1258.460 44.870 ;
        RECT 1209.960 2.400 1210.100 44.550 ;
        RECT 1209.750 -4.800 1210.310 2.400 ;
      LAYER via2 ;
        RECT 1256.810 1290.160 1257.090 1290.440 ;
        RECT 1256.810 1289.480 1257.090 1289.760 ;
        RECT 1257.730 1014.080 1258.010 1014.360 ;
        RECT 1258.650 1014.080 1258.930 1014.360 ;
      LAYER met3 ;
        RECT 1256.785 1290.450 1257.115 1290.465 ;
        RECT 1256.785 1290.135 1257.330 1290.450 ;
        RECT 1257.030 1289.785 1257.330 1290.135 ;
        RECT 1256.785 1289.470 1257.330 1289.785 ;
        RECT 1256.785 1289.455 1257.115 1289.470 ;
        RECT 1257.705 1014.370 1258.035 1014.385 ;
        RECT 1258.625 1014.370 1258.955 1014.385 ;
        RECT 1257.705 1014.070 1258.955 1014.370 ;
        RECT 1257.705 1014.055 1258.035 1014.070 ;
        RECT 1258.625 1014.055 1258.955 1014.070 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1227.810 18.260 1228.130 18.320 ;
        RECT 1275.650 18.260 1275.970 18.320 ;
        RECT 1227.810 18.120 1275.970 18.260 ;
        RECT 1227.810 18.060 1228.130 18.120 ;
        RECT 1275.650 18.060 1275.970 18.120 ;
      LAYER via ;
        RECT 1227.840 18.060 1228.100 18.320 ;
        RECT 1275.680 18.060 1275.940 18.320 ;
      LAYER met2 ;
        RECT 1276.040 1700.410 1276.320 1704.000 ;
        RECT 1275.740 1700.270 1276.320 1700.410 ;
        RECT 1275.740 18.350 1275.880 1700.270 ;
        RECT 1276.040 1700.000 1276.320 1700.270 ;
        RECT 1227.840 18.030 1228.100 18.350 ;
        RECT 1275.680 18.030 1275.940 18.350 ;
        RECT 1227.900 2.400 1228.040 18.030 ;
        RECT 1227.690 -4.800 1228.250 2.400 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1245.750 16.900 1246.070 16.960 ;
        RECT 1277.950 16.900 1278.270 16.960 ;
        RECT 1245.750 16.760 1278.270 16.900 ;
        RECT 1245.750 16.700 1246.070 16.760 ;
        RECT 1277.950 16.700 1278.270 16.760 ;
      LAYER via ;
        RECT 1245.780 16.700 1246.040 16.960 ;
        RECT 1277.980 16.700 1278.240 16.960 ;
      LAYER met2 ;
        RECT 1277.880 1700.340 1278.160 1704.000 ;
        RECT 1277.880 1700.000 1278.180 1700.340 ;
        RECT 1278.040 16.990 1278.180 1700.000 ;
        RECT 1245.780 16.670 1246.040 16.990 ;
        RECT 1277.980 16.670 1278.240 16.990 ;
        RECT 1245.840 2.400 1245.980 16.670 ;
        RECT 1245.630 -4.800 1246.190 2.400 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1263.230 17.920 1263.550 17.980 ;
        RECT 1278.870 17.920 1279.190 17.980 ;
        RECT 1263.230 17.780 1279.190 17.920 ;
        RECT 1263.230 17.720 1263.550 17.780 ;
        RECT 1278.870 17.720 1279.190 17.780 ;
      LAYER via ;
        RECT 1263.260 17.720 1263.520 17.980 ;
        RECT 1278.900 17.720 1279.160 17.980 ;
      LAYER met2 ;
        RECT 1279.720 1700.410 1280.000 1704.000 ;
        RECT 1279.420 1700.270 1280.000 1700.410 ;
        RECT 1279.420 1678.140 1279.560 1700.270 ;
        RECT 1279.720 1700.000 1280.000 1700.270 ;
        RECT 1278.960 1678.000 1279.560 1678.140 ;
        RECT 1278.960 18.010 1279.100 1678.000 ;
        RECT 1263.260 17.690 1263.520 18.010 ;
        RECT 1278.900 17.690 1279.160 18.010 ;
        RECT 1263.320 2.400 1263.460 17.690 ;
        RECT 1263.110 -4.800 1263.670 2.400 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1277.490 1678.140 1277.810 1678.200 ;
        RECT 1281.170 1678.140 1281.490 1678.200 ;
        RECT 1277.490 1678.000 1281.490 1678.140 ;
        RECT 1277.490 1677.940 1277.810 1678.000 ;
        RECT 1281.170 1677.940 1281.490 1678.000 ;
        RECT 1277.490 20.640 1277.810 20.700 ;
        RECT 1281.170 20.640 1281.490 20.700 ;
        RECT 1277.490 20.500 1281.490 20.640 ;
        RECT 1277.490 20.440 1277.810 20.500 ;
        RECT 1281.170 20.440 1281.490 20.500 ;
      LAYER via ;
        RECT 1277.520 1677.940 1277.780 1678.200 ;
        RECT 1281.200 1677.940 1281.460 1678.200 ;
        RECT 1277.520 20.440 1277.780 20.700 ;
        RECT 1281.200 20.440 1281.460 20.700 ;
      LAYER met2 ;
        RECT 1281.560 1700.410 1281.840 1704.000 ;
        RECT 1281.260 1700.270 1281.840 1700.410 ;
        RECT 1281.260 1678.230 1281.400 1700.270 ;
        RECT 1281.560 1700.000 1281.840 1700.270 ;
        RECT 1277.520 1677.910 1277.780 1678.230 ;
        RECT 1281.200 1677.910 1281.460 1678.230 ;
        RECT 1277.580 20.730 1277.720 1677.910 ;
        RECT 1277.520 20.410 1277.780 20.730 ;
        RECT 1281.200 20.410 1281.460 20.730 ;
        RECT 1281.260 2.400 1281.400 20.410 ;
        RECT 1281.050 -4.800 1281.610 2.400 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1283.470 1685.620 1283.790 1685.680 ;
        RECT 1292.210 1685.620 1292.530 1685.680 ;
        RECT 1283.470 1685.480 1292.530 1685.620 ;
        RECT 1283.470 1685.420 1283.790 1685.480 ;
        RECT 1292.210 1685.420 1292.530 1685.480 ;
        RECT 1292.210 20.640 1292.530 20.700 ;
        RECT 1299.110 20.640 1299.430 20.700 ;
        RECT 1292.210 20.500 1299.430 20.640 ;
        RECT 1292.210 20.440 1292.530 20.500 ;
        RECT 1299.110 20.440 1299.430 20.500 ;
      LAYER via ;
        RECT 1283.500 1685.420 1283.760 1685.680 ;
        RECT 1292.240 1685.420 1292.500 1685.680 ;
        RECT 1292.240 20.440 1292.500 20.700 ;
        RECT 1299.140 20.440 1299.400 20.700 ;
      LAYER met2 ;
        RECT 1283.400 1700.340 1283.680 1704.000 ;
        RECT 1283.400 1700.000 1283.700 1700.340 ;
        RECT 1283.560 1685.710 1283.700 1700.000 ;
        RECT 1283.500 1685.390 1283.760 1685.710 ;
        RECT 1292.240 1685.390 1292.500 1685.710 ;
        RECT 1292.300 20.730 1292.440 1685.390 ;
        RECT 1292.240 20.410 1292.500 20.730 ;
        RECT 1299.140 20.410 1299.400 20.730 ;
        RECT 1299.200 2.400 1299.340 20.410 ;
        RECT 1298.990 -4.800 1299.550 2.400 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1285.310 1684.940 1285.630 1685.000 ;
        RECT 1288.990 1684.940 1289.310 1685.000 ;
        RECT 1285.310 1684.800 1289.310 1684.940 ;
        RECT 1285.310 1684.740 1285.630 1684.800 ;
        RECT 1288.990 1684.740 1289.310 1684.800 ;
        RECT 1289.450 19.280 1289.770 19.340 ;
        RECT 1317.050 19.280 1317.370 19.340 ;
        RECT 1289.450 19.140 1317.370 19.280 ;
        RECT 1289.450 19.080 1289.770 19.140 ;
        RECT 1317.050 19.080 1317.370 19.140 ;
      LAYER via ;
        RECT 1285.340 1684.740 1285.600 1685.000 ;
        RECT 1289.020 1684.740 1289.280 1685.000 ;
        RECT 1289.480 19.080 1289.740 19.340 ;
        RECT 1317.080 19.080 1317.340 19.340 ;
      LAYER met2 ;
        RECT 1285.240 1700.340 1285.520 1704.000 ;
        RECT 1285.240 1700.000 1285.540 1700.340 ;
        RECT 1285.400 1685.030 1285.540 1700.000 ;
        RECT 1285.340 1684.710 1285.600 1685.030 ;
        RECT 1289.020 1684.710 1289.280 1685.030 ;
        RECT 1289.080 1678.140 1289.220 1684.710 ;
        RECT 1289.080 1678.000 1289.680 1678.140 ;
        RECT 1289.540 19.370 1289.680 1678.000 ;
        RECT 1289.480 19.050 1289.740 19.370 ;
        RECT 1317.080 19.050 1317.340 19.370 ;
        RECT 1317.140 2.400 1317.280 19.050 ;
        RECT 1316.930 -4.800 1317.490 2.400 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1306.085 1683.085 1306.255 1686.315 ;
      LAYER mcon ;
        RECT 1306.085 1686.145 1306.255 1686.315 ;
      LAYER met1 ;
        RECT 1287.150 1686.300 1287.470 1686.360 ;
        RECT 1306.025 1686.300 1306.315 1686.345 ;
        RECT 1287.150 1686.160 1306.315 1686.300 ;
        RECT 1287.150 1686.100 1287.470 1686.160 ;
        RECT 1306.025 1686.115 1306.315 1686.160 ;
        RECT 1306.010 1683.240 1306.330 1683.300 ;
        RECT 1305.815 1683.100 1306.330 1683.240 ;
        RECT 1306.010 1683.040 1306.330 1683.100 ;
        RECT 1306.010 1667.600 1306.330 1667.660 ;
        RECT 1307.390 1667.600 1307.710 1667.660 ;
        RECT 1306.010 1667.460 1307.710 1667.600 ;
        RECT 1306.010 1667.400 1306.330 1667.460 ;
        RECT 1307.390 1667.400 1307.710 1667.460 ;
        RECT 1307.390 41.380 1307.710 41.440 ;
        RECT 1334.990 41.380 1335.310 41.440 ;
        RECT 1307.390 41.240 1335.310 41.380 ;
        RECT 1307.390 41.180 1307.710 41.240 ;
        RECT 1334.990 41.180 1335.310 41.240 ;
      LAYER via ;
        RECT 1287.180 1686.100 1287.440 1686.360 ;
        RECT 1306.040 1683.040 1306.300 1683.300 ;
        RECT 1306.040 1667.400 1306.300 1667.660 ;
        RECT 1307.420 1667.400 1307.680 1667.660 ;
        RECT 1307.420 41.180 1307.680 41.440 ;
        RECT 1335.020 41.180 1335.280 41.440 ;
      LAYER met2 ;
        RECT 1287.080 1700.340 1287.360 1704.000 ;
        RECT 1287.080 1700.000 1287.380 1700.340 ;
        RECT 1287.240 1686.390 1287.380 1700.000 ;
        RECT 1287.180 1686.070 1287.440 1686.390 ;
        RECT 1306.040 1683.010 1306.300 1683.330 ;
        RECT 1306.100 1667.690 1306.240 1683.010 ;
        RECT 1306.040 1667.370 1306.300 1667.690 ;
        RECT 1307.420 1667.370 1307.680 1667.690 ;
        RECT 1307.480 41.470 1307.620 1667.370 ;
        RECT 1307.420 41.150 1307.680 41.470 ;
        RECT 1335.020 41.150 1335.280 41.470 ;
        RECT 1335.080 2.400 1335.220 41.150 ;
        RECT 1334.870 -4.800 1335.430 2.400 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 696.510 1660.120 696.830 1660.180 ;
        RECT 696.510 1659.980 1169.620 1660.120 ;
        RECT 696.510 1659.920 696.830 1659.980 ;
        RECT 1169.480 1659.780 1169.620 1659.980 ;
        RECT 1220.910 1659.780 1221.230 1659.840 ;
        RECT 1169.480 1659.640 1221.230 1659.780 ;
        RECT 1220.910 1659.580 1221.230 1659.640 ;
      LAYER via ;
        RECT 696.540 1659.920 696.800 1660.180 ;
        RECT 1220.940 1659.580 1221.200 1659.840 ;
      LAYER met2 ;
        RECT 1220.840 1700.340 1221.120 1704.000 ;
        RECT 1220.840 1700.000 1221.140 1700.340 ;
        RECT 696.540 1659.890 696.800 1660.210 ;
        RECT 696.600 24.210 696.740 1659.890 ;
        RECT 1221.000 1659.870 1221.140 1700.000 ;
        RECT 1220.940 1659.550 1221.200 1659.870 ;
        RECT 692.460 24.070 696.740 24.210 ;
        RECT 692.460 2.400 692.600 24.070 ;
        RECT 692.250 -4.800 692.810 2.400 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1288.530 27.440 1288.850 27.500 ;
        RECT 1352.470 27.440 1352.790 27.500 ;
        RECT 1288.530 27.300 1352.790 27.440 ;
        RECT 1288.530 27.240 1288.850 27.300 ;
        RECT 1352.470 27.240 1352.790 27.300 ;
      LAYER via ;
        RECT 1288.560 27.240 1288.820 27.500 ;
        RECT 1352.500 27.240 1352.760 27.500 ;
      LAYER met2 ;
        RECT 1288.920 1700.410 1289.200 1704.000 ;
        RECT 1288.620 1700.270 1289.200 1700.410 ;
        RECT 1288.620 27.530 1288.760 1700.270 ;
        RECT 1288.920 1700.000 1289.200 1700.270 ;
        RECT 1288.560 27.210 1288.820 27.530 ;
        RECT 1352.500 27.210 1352.760 27.530 ;
        RECT 1352.560 2.400 1352.700 27.210 ;
        RECT 1352.350 -4.800 1352.910 2.400 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1290.830 27.100 1291.150 27.160 ;
        RECT 1370.410 27.100 1370.730 27.160 ;
        RECT 1290.830 26.960 1370.730 27.100 ;
        RECT 1290.830 26.900 1291.150 26.960 ;
        RECT 1370.410 26.900 1370.730 26.960 ;
      LAYER via ;
        RECT 1290.860 26.900 1291.120 27.160 ;
        RECT 1370.440 26.900 1370.700 27.160 ;
      LAYER met2 ;
        RECT 1290.760 1700.340 1291.040 1704.000 ;
        RECT 1290.760 1700.000 1291.060 1700.340 ;
        RECT 1290.920 27.190 1291.060 1700.000 ;
        RECT 1290.860 26.870 1291.120 27.190 ;
        RECT 1370.440 26.870 1370.700 27.190 ;
        RECT 1370.500 2.400 1370.640 26.870 ;
        RECT 1370.290 -4.800 1370.850 2.400 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1292.670 1683.920 1292.990 1683.980 ;
        RECT 1294.510 1683.920 1294.830 1683.980 ;
        RECT 1292.670 1683.780 1294.830 1683.920 ;
        RECT 1292.670 1683.720 1292.990 1683.780 ;
        RECT 1294.510 1683.720 1294.830 1683.780 ;
        RECT 1294.510 26.080 1294.830 26.140 ;
        RECT 1388.350 26.080 1388.670 26.140 ;
        RECT 1294.510 25.940 1388.670 26.080 ;
        RECT 1294.510 25.880 1294.830 25.940 ;
        RECT 1388.350 25.880 1388.670 25.940 ;
      LAYER via ;
        RECT 1292.700 1683.720 1292.960 1683.980 ;
        RECT 1294.540 1683.720 1294.800 1683.980 ;
        RECT 1294.540 25.880 1294.800 26.140 ;
        RECT 1388.380 25.880 1388.640 26.140 ;
      LAYER met2 ;
        RECT 1292.600 1700.340 1292.880 1704.000 ;
        RECT 1292.600 1700.000 1292.900 1700.340 ;
        RECT 1292.760 1684.010 1292.900 1700.000 ;
        RECT 1292.700 1683.690 1292.960 1684.010 ;
        RECT 1294.540 1683.690 1294.800 1684.010 ;
        RECT 1294.600 26.170 1294.740 1683.690 ;
        RECT 1294.540 25.850 1294.800 26.170 ;
        RECT 1388.380 25.850 1388.640 26.170 ;
        RECT 1388.440 2.400 1388.580 25.850 ;
        RECT 1388.230 -4.800 1388.790 2.400 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1294.050 25.400 1294.370 25.460 ;
        RECT 1406.290 25.400 1406.610 25.460 ;
        RECT 1294.050 25.260 1406.610 25.400 ;
        RECT 1294.050 25.200 1294.370 25.260 ;
        RECT 1406.290 25.200 1406.610 25.260 ;
      LAYER via ;
        RECT 1294.080 25.200 1294.340 25.460 ;
        RECT 1406.320 25.200 1406.580 25.460 ;
      LAYER met2 ;
        RECT 1294.440 1700.410 1294.720 1704.000 ;
        RECT 1294.140 1700.270 1294.720 1700.410 ;
        RECT 1294.140 25.490 1294.280 1700.270 ;
        RECT 1294.440 1700.000 1294.720 1700.270 ;
        RECT 1294.080 25.170 1294.340 25.490 ;
        RECT 1406.320 25.170 1406.580 25.490 ;
        RECT 1406.380 2.400 1406.520 25.170 ;
        RECT 1406.170 -4.800 1406.730 2.400 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1291.290 1684.600 1291.610 1684.660 ;
        RECT 1296.350 1684.600 1296.670 1684.660 ;
        RECT 1291.290 1684.460 1296.670 1684.600 ;
        RECT 1291.290 1684.400 1291.610 1684.460 ;
        RECT 1296.350 1684.400 1296.670 1684.460 ;
        RECT 1291.290 24.720 1291.610 24.780 ;
        RECT 1423.770 24.720 1424.090 24.780 ;
        RECT 1291.290 24.580 1424.090 24.720 ;
        RECT 1291.290 24.520 1291.610 24.580 ;
        RECT 1423.770 24.520 1424.090 24.580 ;
      LAYER via ;
        RECT 1291.320 1684.400 1291.580 1684.660 ;
        RECT 1296.380 1684.400 1296.640 1684.660 ;
        RECT 1291.320 24.520 1291.580 24.780 ;
        RECT 1423.800 24.520 1424.060 24.780 ;
      LAYER met2 ;
        RECT 1296.280 1700.340 1296.560 1704.000 ;
        RECT 1296.280 1700.000 1296.580 1700.340 ;
        RECT 1296.440 1684.690 1296.580 1700.000 ;
        RECT 1291.320 1684.370 1291.580 1684.690 ;
        RECT 1296.380 1684.370 1296.640 1684.690 ;
        RECT 1291.380 24.810 1291.520 1684.370 ;
        RECT 1291.320 24.490 1291.580 24.810 ;
        RECT 1423.800 24.490 1424.060 24.810 ;
        RECT 1423.860 2.400 1424.000 24.490 ;
        RECT 1423.650 -4.800 1424.210 2.400 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1304.245 1687.165 1304.415 1689.715 ;
        RECT 1317.585 1688.185 1317.755 1689.715 ;
        RECT 1400.845 1688.525 1401.015 1689.715 ;
      LAYER mcon ;
        RECT 1304.245 1689.545 1304.415 1689.715 ;
        RECT 1317.585 1689.545 1317.755 1689.715 ;
        RECT 1400.845 1689.545 1401.015 1689.715 ;
      LAYER met1 ;
        RECT 1304.185 1689.700 1304.475 1689.745 ;
        RECT 1317.525 1689.700 1317.815 1689.745 ;
        RECT 1304.185 1689.560 1317.815 1689.700 ;
        RECT 1304.185 1689.515 1304.475 1689.560 ;
        RECT 1317.525 1689.515 1317.815 1689.560 ;
        RECT 1396.170 1689.700 1396.490 1689.760 ;
        RECT 1400.785 1689.700 1401.075 1689.745 ;
        RECT 1396.170 1689.560 1401.075 1689.700 ;
        RECT 1396.170 1689.500 1396.490 1689.560 ;
        RECT 1400.785 1689.515 1401.075 1689.560 ;
        RECT 1400.785 1688.680 1401.075 1688.725 ;
        RECT 1400.785 1688.540 1404.680 1688.680 ;
        RECT 1400.785 1688.495 1401.075 1688.540 ;
        RECT 1317.525 1688.340 1317.815 1688.385 ;
        RECT 1375.930 1688.340 1376.250 1688.400 ;
        RECT 1317.525 1688.200 1376.250 1688.340 ;
        RECT 1404.540 1688.340 1404.680 1688.540 ;
        RECT 1417.790 1688.340 1418.110 1688.400 ;
        RECT 1404.540 1688.200 1418.110 1688.340 ;
        RECT 1317.525 1688.155 1317.815 1688.200 ;
        RECT 1375.930 1688.140 1376.250 1688.200 ;
        RECT 1417.790 1688.140 1418.110 1688.200 ;
        RECT 1298.190 1687.320 1298.510 1687.380 ;
        RECT 1304.185 1687.320 1304.475 1687.365 ;
        RECT 1298.190 1687.180 1304.475 1687.320 ;
        RECT 1298.190 1687.120 1298.510 1687.180 ;
        RECT 1304.185 1687.135 1304.475 1687.180 ;
        RECT 1417.790 34.580 1418.110 34.640 ;
        RECT 1441.710 34.580 1442.030 34.640 ;
        RECT 1417.790 34.440 1442.030 34.580 ;
        RECT 1417.790 34.380 1418.110 34.440 ;
        RECT 1441.710 34.380 1442.030 34.440 ;
      LAYER via ;
        RECT 1396.200 1689.500 1396.460 1689.760 ;
        RECT 1375.960 1688.140 1376.220 1688.400 ;
        RECT 1417.820 1688.140 1418.080 1688.400 ;
        RECT 1298.220 1687.120 1298.480 1687.380 ;
        RECT 1417.820 34.380 1418.080 34.640 ;
        RECT 1441.740 34.380 1442.000 34.640 ;
      LAYER met2 ;
        RECT 1298.120 1700.340 1298.400 1704.000 ;
        RECT 1298.120 1700.000 1298.420 1700.340 ;
        RECT 1298.280 1687.410 1298.420 1700.000 ;
        RECT 1396.200 1689.470 1396.460 1689.790 ;
        RECT 1396.260 1688.965 1396.400 1689.470 ;
        RECT 1375.950 1688.595 1376.230 1688.965 ;
        RECT 1396.190 1688.595 1396.470 1688.965 ;
        RECT 1376.020 1688.430 1376.160 1688.595 ;
        RECT 1375.960 1688.110 1376.220 1688.430 ;
        RECT 1417.820 1688.110 1418.080 1688.430 ;
        RECT 1298.220 1687.090 1298.480 1687.410 ;
        RECT 1417.880 34.670 1418.020 1688.110 ;
        RECT 1417.820 34.350 1418.080 34.670 ;
        RECT 1441.740 34.350 1442.000 34.670 ;
        RECT 1441.800 2.400 1441.940 34.350 ;
        RECT 1441.590 -4.800 1442.150 2.400 ;
      LAYER via2 ;
        RECT 1375.950 1688.640 1376.230 1688.920 ;
        RECT 1396.190 1688.640 1396.470 1688.920 ;
      LAYER met3 ;
        RECT 1375.925 1688.930 1376.255 1688.945 ;
        RECT 1396.165 1688.930 1396.495 1688.945 ;
        RECT 1375.925 1688.630 1396.495 1688.930 ;
        RECT 1375.925 1688.615 1376.255 1688.630 ;
        RECT 1396.165 1688.615 1396.495 1688.630 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1300.030 1683.920 1300.350 1683.980 ;
        RECT 1302.330 1683.920 1302.650 1683.980 ;
        RECT 1300.030 1683.780 1302.650 1683.920 ;
        RECT 1300.030 1683.720 1300.350 1683.780 ;
        RECT 1302.330 1683.720 1302.650 1683.780 ;
        RECT 1302.330 46.480 1302.650 46.540 ;
        RECT 1459.650 46.480 1459.970 46.540 ;
        RECT 1302.330 46.340 1459.970 46.480 ;
        RECT 1302.330 46.280 1302.650 46.340 ;
        RECT 1459.650 46.280 1459.970 46.340 ;
      LAYER via ;
        RECT 1300.060 1683.720 1300.320 1683.980 ;
        RECT 1302.360 1683.720 1302.620 1683.980 ;
        RECT 1302.360 46.280 1302.620 46.540 ;
        RECT 1459.680 46.280 1459.940 46.540 ;
      LAYER met2 ;
        RECT 1299.960 1700.340 1300.240 1704.000 ;
        RECT 1299.960 1700.000 1300.260 1700.340 ;
        RECT 1300.120 1684.010 1300.260 1700.000 ;
        RECT 1300.060 1683.690 1300.320 1684.010 ;
        RECT 1302.360 1683.690 1302.620 1684.010 ;
        RECT 1302.420 46.570 1302.560 1683.690 ;
        RECT 1302.360 46.250 1302.620 46.570 ;
        RECT 1459.680 46.250 1459.940 46.570 ;
        RECT 1459.740 2.400 1459.880 46.250 ;
        RECT 1459.530 -4.800 1460.090 2.400 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1300.030 1062.880 1300.350 1063.140 ;
        RECT 1300.120 1062.460 1300.260 1062.880 ;
        RECT 1300.030 1062.200 1300.350 1062.460 ;
        RECT 1300.030 96.940 1300.350 97.200 ;
        RECT 1300.120 96.520 1300.260 96.940 ;
        RECT 1300.030 96.260 1300.350 96.520 ;
        RECT 1300.030 46.140 1300.350 46.200 ;
        RECT 1477.590 46.140 1477.910 46.200 ;
        RECT 1300.030 46.000 1477.910 46.140 ;
        RECT 1300.030 45.940 1300.350 46.000 ;
        RECT 1477.590 45.940 1477.910 46.000 ;
      LAYER via ;
        RECT 1300.060 1062.880 1300.320 1063.140 ;
        RECT 1300.060 1062.200 1300.320 1062.460 ;
        RECT 1300.060 96.940 1300.320 97.200 ;
        RECT 1300.060 96.260 1300.320 96.520 ;
        RECT 1300.060 45.940 1300.320 46.200 ;
        RECT 1477.620 45.940 1477.880 46.200 ;
      LAYER met2 ;
        RECT 1301.340 1700.340 1301.620 1704.000 ;
        RECT 1301.340 1700.000 1301.640 1700.340 ;
        RECT 1301.500 1678.650 1301.640 1700.000 ;
        RECT 1300.120 1678.510 1301.640 1678.650 ;
        RECT 1300.120 1063.170 1300.260 1678.510 ;
        RECT 1300.060 1062.850 1300.320 1063.170 ;
        RECT 1300.060 1062.170 1300.320 1062.490 ;
        RECT 1300.120 97.230 1300.260 1062.170 ;
        RECT 1300.060 96.910 1300.320 97.230 ;
        RECT 1300.060 96.230 1300.320 96.550 ;
        RECT 1300.120 46.230 1300.260 96.230 ;
        RECT 1300.060 45.910 1300.320 46.230 ;
        RECT 1477.620 45.910 1477.880 46.230 ;
        RECT 1477.680 2.400 1477.820 45.910 ;
        RECT 1477.470 -4.800 1478.030 2.400 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1299.110 1684.600 1299.430 1684.660 ;
        RECT 1303.250 1684.600 1303.570 1684.660 ;
        RECT 1299.110 1684.460 1303.570 1684.600 ;
        RECT 1299.110 1684.400 1299.430 1684.460 ;
        RECT 1303.250 1684.400 1303.570 1684.460 ;
        RECT 1299.110 45.800 1299.430 45.860 ;
        RECT 1495.530 45.800 1495.850 45.860 ;
        RECT 1299.110 45.660 1495.850 45.800 ;
        RECT 1299.110 45.600 1299.430 45.660 ;
        RECT 1495.530 45.600 1495.850 45.660 ;
      LAYER via ;
        RECT 1299.140 1684.400 1299.400 1684.660 ;
        RECT 1303.280 1684.400 1303.540 1684.660 ;
        RECT 1299.140 45.600 1299.400 45.860 ;
        RECT 1495.560 45.600 1495.820 45.860 ;
      LAYER met2 ;
        RECT 1303.180 1700.340 1303.460 1704.000 ;
        RECT 1303.180 1700.000 1303.480 1700.340 ;
        RECT 1303.340 1684.690 1303.480 1700.000 ;
        RECT 1299.140 1684.370 1299.400 1684.690 ;
        RECT 1303.280 1684.370 1303.540 1684.690 ;
        RECT 1299.200 45.890 1299.340 1684.370 ;
        RECT 1299.140 45.570 1299.400 45.890 ;
        RECT 1495.560 45.570 1495.820 45.890 ;
        RECT 1495.620 2.400 1495.760 45.570 ;
        RECT 1495.410 -4.800 1495.970 2.400 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1306.010 44.780 1306.330 44.840 ;
        RECT 1513.010 44.780 1513.330 44.840 ;
        RECT 1306.010 44.640 1513.330 44.780 ;
        RECT 1306.010 44.580 1306.330 44.640 ;
        RECT 1513.010 44.580 1513.330 44.640 ;
      LAYER via ;
        RECT 1306.040 44.580 1306.300 44.840 ;
        RECT 1513.040 44.580 1513.300 44.840 ;
      LAYER met2 ;
        RECT 1305.020 1700.410 1305.300 1704.000 ;
        RECT 1305.020 1700.270 1305.780 1700.410 ;
        RECT 1305.020 1700.000 1305.300 1700.270 ;
        RECT 1305.640 1667.090 1305.780 1700.270 ;
        RECT 1305.640 1666.950 1306.240 1667.090 ;
        RECT 1306.100 44.870 1306.240 1666.950 ;
        RECT 1306.040 44.550 1306.300 44.870 ;
        RECT 1513.040 44.550 1513.300 44.870 ;
        RECT 1513.100 2.400 1513.240 44.550 ;
        RECT 1512.890 -4.800 1513.450 2.400 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 709.850 1625.440 710.170 1625.500 ;
        RECT 1224.130 1625.440 1224.450 1625.500 ;
        RECT 709.850 1625.300 1224.450 1625.440 ;
        RECT 709.850 1625.240 710.170 1625.300 ;
        RECT 1224.130 1625.240 1224.450 1625.300 ;
      LAYER via ;
        RECT 709.880 1625.240 710.140 1625.500 ;
        RECT 1224.160 1625.240 1224.420 1625.500 ;
      LAYER met2 ;
        RECT 1222.680 1700.340 1222.960 1704.000 ;
        RECT 1222.680 1700.000 1222.980 1700.340 ;
        RECT 1222.840 1678.650 1222.980 1700.000 ;
        RECT 1222.840 1678.510 1224.360 1678.650 ;
        RECT 1224.220 1625.530 1224.360 1678.510 ;
        RECT 709.880 1625.210 710.140 1625.530 ;
        RECT 1224.160 1625.210 1224.420 1625.530 ;
        RECT 709.940 24.210 710.080 1625.210 ;
        RECT 709.940 24.070 710.540 24.210 ;
        RECT 710.400 2.400 710.540 24.070 ;
        RECT 710.190 -4.800 710.750 2.400 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1306.930 45.460 1307.250 45.520 ;
        RECT 1530.950 45.460 1531.270 45.520 ;
        RECT 1306.930 45.320 1531.270 45.460 ;
        RECT 1306.930 45.260 1307.250 45.320 ;
        RECT 1530.950 45.260 1531.270 45.320 ;
      LAYER via ;
        RECT 1306.960 45.260 1307.220 45.520 ;
        RECT 1530.980 45.260 1531.240 45.520 ;
      LAYER met2 ;
        RECT 1306.860 1700.340 1307.140 1704.000 ;
        RECT 1306.860 1700.000 1307.160 1700.340 ;
        RECT 1307.020 45.550 1307.160 1700.000 ;
        RECT 1306.960 45.230 1307.220 45.550 ;
        RECT 1530.980 45.230 1531.240 45.550 ;
        RECT 1531.040 2.400 1531.180 45.230 ;
        RECT 1530.830 -4.800 1531.390 2.400 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1306.470 1683.920 1306.790 1683.980 ;
        RECT 1308.770 1683.920 1309.090 1683.980 ;
        RECT 1306.470 1683.780 1309.090 1683.920 ;
        RECT 1306.470 1683.720 1306.790 1683.780 ;
        RECT 1308.770 1683.720 1309.090 1683.780 ;
        RECT 1306.470 45.120 1306.790 45.180 ;
        RECT 1548.890 45.120 1549.210 45.180 ;
        RECT 1306.470 44.980 1549.210 45.120 ;
        RECT 1306.470 44.920 1306.790 44.980 ;
        RECT 1548.890 44.920 1549.210 44.980 ;
      LAYER via ;
        RECT 1306.500 1683.720 1306.760 1683.980 ;
        RECT 1308.800 1683.720 1309.060 1683.980 ;
        RECT 1306.500 44.920 1306.760 45.180 ;
        RECT 1548.920 44.920 1549.180 45.180 ;
      LAYER met2 ;
        RECT 1308.700 1700.340 1308.980 1704.000 ;
        RECT 1308.700 1700.000 1309.000 1700.340 ;
        RECT 1308.860 1684.010 1309.000 1700.000 ;
        RECT 1306.500 1683.690 1306.760 1684.010 ;
        RECT 1308.800 1683.690 1309.060 1684.010 ;
        RECT 1306.560 45.210 1306.700 1683.690 ;
        RECT 1306.500 44.890 1306.760 45.210 ;
        RECT 1548.920 44.890 1549.180 45.210 ;
        RECT 1548.980 2.400 1549.120 44.890 ;
        RECT 1548.770 -4.800 1549.330 2.400 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1310.610 1685.760 1310.930 1686.020 ;
        RECT 1309.690 1684.260 1310.010 1684.320 ;
        RECT 1310.700 1684.260 1310.840 1685.760 ;
        RECT 1309.690 1684.120 1310.840 1684.260 ;
        RECT 1309.690 1684.060 1310.010 1684.120 ;
        RECT 1309.690 1661.480 1310.010 1661.540 ;
        RECT 1566.370 1661.480 1566.690 1661.540 ;
        RECT 1309.690 1661.340 1566.690 1661.480 ;
        RECT 1309.690 1661.280 1310.010 1661.340 ;
        RECT 1566.370 1661.280 1566.690 1661.340 ;
      LAYER via ;
        RECT 1310.640 1685.760 1310.900 1686.020 ;
        RECT 1309.720 1684.060 1309.980 1684.320 ;
        RECT 1309.720 1661.280 1309.980 1661.540 ;
        RECT 1566.400 1661.280 1566.660 1661.540 ;
      LAYER met2 ;
        RECT 1310.540 1700.340 1310.820 1704.000 ;
        RECT 1310.540 1700.000 1310.840 1700.340 ;
        RECT 1310.700 1686.050 1310.840 1700.000 ;
        RECT 1310.640 1685.730 1310.900 1686.050 ;
        RECT 1309.720 1684.030 1309.980 1684.350 ;
        RECT 1309.780 1661.570 1309.920 1684.030 ;
        RECT 1309.720 1661.250 1309.980 1661.570 ;
        RECT 1566.400 1661.250 1566.660 1661.570 ;
        RECT 1566.460 17.410 1566.600 1661.250 ;
        RECT 1566.460 17.270 1567.060 17.410 ;
        RECT 1566.920 2.400 1567.060 17.270 ;
        RECT 1566.710 -4.800 1567.270 2.400 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1311.530 1674.740 1311.850 1674.800 ;
        RECT 1580.170 1674.740 1580.490 1674.800 ;
        RECT 1311.530 1674.600 1580.490 1674.740 ;
        RECT 1311.530 1674.540 1311.850 1674.600 ;
        RECT 1580.170 1674.540 1580.490 1674.600 ;
      LAYER via ;
        RECT 1311.560 1674.540 1311.820 1674.800 ;
        RECT 1580.200 1674.540 1580.460 1674.800 ;
      LAYER met2 ;
        RECT 1312.380 1700.340 1312.660 1704.000 ;
        RECT 1312.380 1700.000 1312.680 1700.340 ;
        RECT 1312.540 1686.300 1312.680 1700.000 ;
        RECT 1311.620 1686.160 1312.680 1686.300 ;
        RECT 1311.620 1674.830 1311.760 1686.160 ;
        RECT 1311.560 1674.510 1311.820 1674.830 ;
        RECT 1580.200 1674.510 1580.460 1674.830 ;
        RECT 1580.260 18.090 1580.400 1674.510 ;
        RECT 1580.260 17.950 1585.000 18.090 ;
        RECT 1584.860 2.400 1585.000 17.950 ;
        RECT 1584.650 -4.800 1585.210 2.400 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1312.450 1683.920 1312.770 1683.980 ;
        RECT 1314.290 1683.920 1314.610 1683.980 ;
        RECT 1312.450 1683.780 1314.610 1683.920 ;
        RECT 1312.450 1683.720 1312.770 1683.780 ;
        RECT 1314.290 1683.720 1314.610 1683.780 ;
        RECT 1312.450 1654.680 1312.770 1654.740 ;
        RECT 1600.870 1654.680 1601.190 1654.740 ;
        RECT 1312.450 1654.540 1601.190 1654.680 ;
        RECT 1312.450 1654.480 1312.770 1654.540 ;
        RECT 1600.870 1654.480 1601.190 1654.540 ;
      LAYER via ;
        RECT 1312.480 1683.720 1312.740 1683.980 ;
        RECT 1314.320 1683.720 1314.580 1683.980 ;
        RECT 1312.480 1654.480 1312.740 1654.740 ;
        RECT 1600.900 1654.480 1601.160 1654.740 ;
      LAYER met2 ;
        RECT 1314.220 1700.340 1314.500 1704.000 ;
        RECT 1314.220 1700.000 1314.520 1700.340 ;
        RECT 1314.380 1684.010 1314.520 1700.000 ;
        RECT 1312.480 1683.690 1312.740 1684.010 ;
        RECT 1314.320 1683.690 1314.580 1684.010 ;
        RECT 1312.540 1654.770 1312.680 1683.690 ;
        RECT 1312.480 1654.450 1312.740 1654.770 ;
        RECT 1600.900 1654.450 1601.160 1654.770 ;
        RECT 1600.960 17.410 1601.100 1654.450 ;
        RECT 1600.960 17.270 1602.480 17.410 ;
        RECT 1602.340 2.400 1602.480 17.270 ;
        RECT 1602.130 -4.800 1602.690 2.400 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1316.130 1633.600 1316.450 1633.660 ;
        RECT 1614.670 1633.600 1614.990 1633.660 ;
        RECT 1316.130 1633.460 1614.990 1633.600 ;
        RECT 1316.130 1633.400 1316.450 1633.460 ;
        RECT 1614.670 1633.400 1614.990 1633.460 ;
      LAYER via ;
        RECT 1316.160 1633.400 1316.420 1633.660 ;
        RECT 1614.700 1633.400 1614.960 1633.660 ;
      LAYER met2 ;
        RECT 1316.060 1700.340 1316.340 1704.000 ;
        RECT 1316.060 1700.000 1316.360 1700.340 ;
        RECT 1316.220 1633.690 1316.360 1700.000 ;
        RECT 1316.160 1633.370 1316.420 1633.690 ;
        RECT 1614.700 1633.370 1614.960 1633.690 ;
        RECT 1614.760 17.410 1614.900 1633.370 ;
        RECT 1614.760 17.270 1620.420 17.410 ;
        RECT 1620.280 2.400 1620.420 17.270 ;
        RECT 1620.070 -4.800 1620.630 2.400 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1317.970 1689.700 1318.290 1689.760 ;
        RECT 1338.670 1689.700 1338.990 1689.760 ;
        RECT 1317.970 1689.560 1338.990 1689.700 ;
        RECT 1317.970 1689.500 1318.290 1689.560 ;
        RECT 1338.670 1689.500 1338.990 1689.560 ;
        RECT 1338.670 1681.880 1338.990 1681.940 ;
        RECT 1635.370 1681.880 1635.690 1681.940 ;
        RECT 1338.670 1681.740 1635.690 1681.880 ;
        RECT 1338.670 1681.680 1338.990 1681.740 ;
        RECT 1635.370 1681.680 1635.690 1681.740 ;
      LAYER via ;
        RECT 1318.000 1689.500 1318.260 1689.760 ;
        RECT 1338.700 1689.500 1338.960 1689.760 ;
        RECT 1338.700 1681.680 1338.960 1681.940 ;
        RECT 1635.400 1681.680 1635.660 1681.940 ;
      LAYER met2 ;
        RECT 1317.900 1700.340 1318.180 1704.000 ;
        RECT 1317.900 1700.000 1318.200 1700.340 ;
        RECT 1318.060 1689.790 1318.200 1700.000 ;
        RECT 1318.000 1689.470 1318.260 1689.790 ;
        RECT 1338.700 1689.470 1338.960 1689.790 ;
        RECT 1338.760 1681.970 1338.900 1689.470 ;
        RECT 1338.700 1681.650 1338.960 1681.970 ;
        RECT 1635.400 1681.650 1635.660 1681.970 ;
        RECT 1635.460 17.410 1635.600 1681.650 ;
        RECT 1635.460 17.270 1638.360 17.410 ;
        RECT 1638.220 2.400 1638.360 17.270 ;
        RECT 1638.010 -4.800 1638.570 2.400 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1319.810 1686.640 1320.130 1686.700 ;
        RECT 1356.610 1686.640 1356.930 1686.700 ;
        RECT 1319.810 1686.500 1356.930 1686.640 ;
        RECT 1319.810 1686.440 1320.130 1686.500 ;
        RECT 1356.610 1686.440 1356.930 1686.500 ;
        RECT 1356.610 1661.140 1356.930 1661.200 ;
        RECT 1656.070 1661.140 1656.390 1661.200 ;
        RECT 1356.610 1661.000 1656.390 1661.140 ;
        RECT 1356.610 1660.940 1356.930 1661.000 ;
        RECT 1656.070 1660.940 1656.390 1661.000 ;
      LAYER via ;
        RECT 1319.840 1686.440 1320.100 1686.700 ;
        RECT 1356.640 1686.440 1356.900 1686.700 ;
        RECT 1356.640 1660.940 1356.900 1661.200 ;
        RECT 1656.100 1660.940 1656.360 1661.200 ;
      LAYER met2 ;
        RECT 1319.740 1700.340 1320.020 1704.000 ;
        RECT 1319.740 1700.000 1320.040 1700.340 ;
        RECT 1319.900 1686.730 1320.040 1700.000 ;
        RECT 1319.840 1686.410 1320.100 1686.730 ;
        RECT 1356.640 1686.410 1356.900 1686.730 ;
        RECT 1356.700 1661.230 1356.840 1686.410 ;
        RECT 1356.640 1660.910 1356.900 1661.230 ;
        RECT 1656.100 1660.910 1656.360 1661.230 ;
        RECT 1656.160 2.400 1656.300 1660.910 ;
        RECT 1655.950 -4.800 1656.510 2.400 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1322.110 1674.400 1322.430 1674.460 ;
        RECT 1669.870 1674.400 1670.190 1674.460 ;
        RECT 1322.110 1674.260 1670.190 1674.400 ;
        RECT 1322.110 1674.200 1322.430 1674.260 ;
        RECT 1669.870 1674.200 1670.190 1674.260 ;
      LAYER via ;
        RECT 1322.140 1674.200 1322.400 1674.460 ;
        RECT 1669.900 1674.200 1670.160 1674.460 ;
      LAYER met2 ;
        RECT 1321.580 1700.410 1321.860 1704.000 ;
        RECT 1321.580 1700.270 1322.340 1700.410 ;
        RECT 1321.580 1700.000 1321.860 1700.270 ;
        RECT 1322.200 1674.490 1322.340 1700.270 ;
        RECT 1322.140 1674.170 1322.400 1674.490 ;
        RECT 1669.900 1674.170 1670.160 1674.490 ;
        RECT 1669.960 17.410 1670.100 1674.170 ;
        RECT 1669.960 17.270 1673.780 17.410 ;
        RECT 1673.640 2.400 1673.780 17.270 ;
        RECT 1673.430 -4.800 1673.990 2.400 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1324.410 1647.200 1324.730 1647.260 ;
        RECT 1690.570 1647.200 1690.890 1647.260 ;
        RECT 1324.410 1647.060 1690.890 1647.200 ;
        RECT 1324.410 1647.000 1324.730 1647.060 ;
        RECT 1690.570 1647.000 1690.890 1647.060 ;
      LAYER via ;
        RECT 1324.440 1647.000 1324.700 1647.260 ;
        RECT 1690.600 1647.000 1690.860 1647.260 ;
      LAYER met2 ;
        RECT 1323.420 1700.410 1323.700 1704.000 ;
        RECT 1323.420 1700.270 1324.180 1700.410 ;
        RECT 1323.420 1700.000 1323.700 1700.270 ;
        RECT 1324.040 1677.970 1324.180 1700.270 ;
        RECT 1324.040 1677.830 1324.640 1677.970 ;
        RECT 1324.500 1647.290 1324.640 1677.830 ;
        RECT 1324.440 1646.970 1324.700 1647.290 ;
        RECT 1690.600 1646.970 1690.860 1647.290 ;
        RECT 1690.660 17.410 1690.800 1646.970 ;
        RECT 1690.660 17.270 1691.720 17.410 ;
        RECT 1691.580 2.400 1691.720 17.270 ;
        RECT 1691.370 -4.800 1691.930 2.400 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1223.210 1678.140 1223.530 1678.200 ;
        RECT 1224.590 1678.140 1224.910 1678.200 ;
        RECT 1223.210 1678.000 1224.910 1678.140 ;
        RECT 1223.210 1677.940 1223.530 1678.000 ;
        RECT 1224.590 1677.940 1224.910 1678.000 ;
        RECT 731.010 1611.840 731.330 1611.900 ;
        RECT 1223.210 1611.840 1223.530 1611.900 ;
        RECT 731.010 1611.700 1223.530 1611.840 ;
        RECT 731.010 1611.640 731.330 1611.700 ;
        RECT 1223.210 1611.640 1223.530 1611.700 ;
      LAYER via ;
        RECT 1223.240 1677.940 1223.500 1678.200 ;
        RECT 1224.620 1677.940 1224.880 1678.200 ;
        RECT 731.040 1611.640 731.300 1611.900 ;
        RECT 1223.240 1611.640 1223.500 1611.900 ;
      LAYER met2 ;
        RECT 1224.520 1700.340 1224.800 1704.000 ;
        RECT 1224.520 1700.000 1224.820 1700.340 ;
        RECT 1224.680 1678.230 1224.820 1700.000 ;
        RECT 1223.240 1677.910 1223.500 1678.230 ;
        RECT 1224.620 1677.910 1224.880 1678.230 ;
        RECT 1223.300 1611.930 1223.440 1677.910 ;
        RECT 731.040 1611.610 731.300 1611.930 ;
        RECT 1223.240 1611.610 1223.500 1611.930 ;
        RECT 731.100 16.730 731.240 1611.610 ;
        RECT 728.340 16.590 731.240 16.730 ;
        RECT 728.340 2.400 728.480 16.590 ;
        RECT 728.130 -4.800 728.690 2.400 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1325.330 50.220 1325.650 50.280 ;
        RECT 1704.370 50.220 1704.690 50.280 ;
        RECT 1325.330 50.080 1704.690 50.220 ;
        RECT 1325.330 50.020 1325.650 50.080 ;
        RECT 1704.370 50.020 1704.690 50.080 ;
      LAYER via ;
        RECT 1325.360 50.020 1325.620 50.280 ;
        RECT 1704.400 50.020 1704.660 50.280 ;
      LAYER met2 ;
        RECT 1325.260 1700.340 1325.540 1704.000 ;
        RECT 1325.260 1700.000 1325.560 1700.340 ;
        RECT 1325.420 50.310 1325.560 1700.000 ;
        RECT 1325.360 49.990 1325.620 50.310 ;
        RECT 1704.400 49.990 1704.660 50.310 ;
        RECT 1704.460 17.410 1704.600 49.990 ;
        RECT 1704.460 17.270 1709.660 17.410 ;
        RECT 1709.520 2.400 1709.660 17.270 ;
        RECT 1709.310 -4.800 1709.870 2.400 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1327.170 1684.600 1327.490 1684.660 ;
        RECT 1331.310 1684.600 1331.630 1684.660 ;
        RECT 1327.170 1684.460 1331.630 1684.600 ;
        RECT 1327.170 1684.400 1327.490 1684.460 ;
        RECT 1331.310 1684.400 1331.630 1684.460 ;
        RECT 1329.470 1631.220 1329.790 1631.280 ;
        RECT 1331.310 1631.220 1331.630 1631.280 ;
        RECT 1329.470 1631.080 1331.630 1631.220 ;
        RECT 1329.470 1631.020 1329.790 1631.080 ;
        RECT 1331.310 1631.020 1331.630 1631.080 ;
        RECT 1329.470 50.560 1329.790 50.620 ;
        RECT 1725.070 50.560 1725.390 50.620 ;
        RECT 1329.470 50.420 1725.390 50.560 ;
        RECT 1329.470 50.360 1329.790 50.420 ;
        RECT 1725.070 50.360 1725.390 50.420 ;
      LAYER via ;
        RECT 1327.200 1684.400 1327.460 1684.660 ;
        RECT 1331.340 1684.400 1331.600 1684.660 ;
        RECT 1329.500 1631.020 1329.760 1631.280 ;
        RECT 1331.340 1631.020 1331.600 1631.280 ;
        RECT 1329.500 50.360 1329.760 50.620 ;
        RECT 1725.100 50.360 1725.360 50.620 ;
      LAYER met2 ;
        RECT 1327.100 1700.340 1327.380 1704.000 ;
        RECT 1327.100 1700.000 1327.400 1700.340 ;
        RECT 1327.260 1684.690 1327.400 1700.000 ;
        RECT 1327.200 1684.370 1327.460 1684.690 ;
        RECT 1331.340 1684.370 1331.600 1684.690 ;
        RECT 1331.400 1631.310 1331.540 1684.370 ;
        RECT 1329.500 1630.990 1329.760 1631.310 ;
        RECT 1331.340 1630.990 1331.600 1631.310 ;
        RECT 1329.560 50.650 1329.700 1630.990 ;
        RECT 1329.500 50.330 1329.760 50.650 ;
        RECT 1725.100 50.330 1725.360 50.650 ;
        RECT 1725.160 17.410 1725.300 50.330 ;
        RECT 1725.160 17.270 1727.600 17.410 ;
        RECT 1727.460 2.400 1727.600 17.270 ;
        RECT 1727.250 -4.800 1727.810 2.400 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1328.550 50.900 1328.870 50.960 ;
        RECT 1738.870 50.900 1739.190 50.960 ;
        RECT 1328.550 50.760 1739.190 50.900 ;
        RECT 1328.550 50.700 1328.870 50.760 ;
        RECT 1738.870 50.700 1739.190 50.760 ;
        RECT 1738.870 20.980 1739.190 21.040 ;
        RECT 1745.310 20.980 1745.630 21.040 ;
        RECT 1738.870 20.840 1745.630 20.980 ;
        RECT 1738.870 20.780 1739.190 20.840 ;
        RECT 1745.310 20.780 1745.630 20.840 ;
      LAYER via ;
        RECT 1328.580 50.700 1328.840 50.960 ;
        RECT 1738.900 50.700 1739.160 50.960 ;
        RECT 1738.900 20.780 1739.160 21.040 ;
        RECT 1745.340 20.780 1745.600 21.040 ;
      LAYER met2 ;
        RECT 1328.940 1700.340 1329.220 1704.000 ;
        RECT 1328.940 1700.000 1329.240 1700.340 ;
        RECT 1329.100 1666.410 1329.240 1700.000 ;
        RECT 1328.640 1666.270 1329.240 1666.410 ;
        RECT 1328.640 50.990 1328.780 1666.270 ;
        RECT 1328.580 50.670 1328.840 50.990 ;
        RECT 1738.900 50.670 1739.160 50.990 ;
        RECT 1738.960 21.070 1739.100 50.670 ;
        RECT 1738.900 20.750 1739.160 21.070 ;
        RECT 1745.340 20.750 1745.600 21.070 ;
        RECT 1745.400 2.400 1745.540 20.750 ;
        RECT 1745.190 -4.800 1745.750 2.400 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1328.090 1684.260 1328.410 1684.320 ;
        RECT 1330.850 1684.260 1331.170 1684.320 ;
        RECT 1328.090 1684.120 1331.170 1684.260 ;
        RECT 1328.090 1684.060 1328.410 1684.120 ;
        RECT 1330.850 1684.060 1331.170 1684.120 ;
        RECT 1328.090 51.240 1328.410 51.300 ;
        RECT 1759.570 51.240 1759.890 51.300 ;
        RECT 1328.090 51.100 1759.890 51.240 ;
        RECT 1328.090 51.040 1328.410 51.100 ;
        RECT 1759.570 51.040 1759.890 51.100 ;
      LAYER via ;
        RECT 1328.120 1684.060 1328.380 1684.320 ;
        RECT 1330.880 1684.060 1331.140 1684.320 ;
        RECT 1328.120 51.040 1328.380 51.300 ;
        RECT 1759.600 51.040 1759.860 51.300 ;
      LAYER met2 ;
        RECT 1330.780 1700.340 1331.060 1704.000 ;
        RECT 1330.780 1700.000 1331.080 1700.340 ;
        RECT 1330.940 1684.350 1331.080 1700.000 ;
        RECT 1328.120 1684.030 1328.380 1684.350 ;
        RECT 1330.880 1684.030 1331.140 1684.350 ;
        RECT 1328.180 51.330 1328.320 1684.030 ;
        RECT 1328.120 51.010 1328.380 51.330 ;
        RECT 1759.600 51.010 1759.860 51.330 ;
        RECT 1759.660 17.410 1759.800 51.010 ;
        RECT 1759.660 17.270 1763.020 17.410 ;
        RECT 1762.880 2.400 1763.020 17.270 ;
        RECT 1762.670 -4.800 1763.230 2.400 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1332.690 54.980 1333.010 55.040 ;
        RECT 1780.730 54.980 1781.050 55.040 ;
        RECT 1332.690 54.840 1781.050 54.980 ;
        RECT 1332.690 54.780 1333.010 54.840 ;
        RECT 1780.730 54.780 1781.050 54.840 ;
      LAYER via ;
        RECT 1332.720 54.780 1332.980 55.040 ;
        RECT 1780.760 54.780 1781.020 55.040 ;
      LAYER met2 ;
        RECT 1332.620 1700.340 1332.900 1704.000 ;
        RECT 1332.620 1700.000 1332.920 1700.340 ;
        RECT 1332.780 55.070 1332.920 1700.000 ;
        RECT 1332.720 54.750 1332.980 55.070 ;
        RECT 1780.760 54.750 1781.020 55.070 ;
        RECT 1780.820 2.400 1780.960 54.750 ;
        RECT 1780.610 -4.800 1781.170 2.400 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1334.530 1684.260 1334.850 1684.320 ;
        RECT 1336.830 1684.260 1337.150 1684.320 ;
        RECT 1334.530 1684.120 1337.150 1684.260 ;
        RECT 1334.530 1684.060 1334.850 1684.120 ;
        RECT 1336.830 1684.060 1337.150 1684.120 ;
        RECT 1336.830 54.640 1337.150 54.700 ;
        RECT 1794.070 54.640 1794.390 54.700 ;
        RECT 1336.830 54.500 1794.390 54.640 ;
        RECT 1336.830 54.440 1337.150 54.500 ;
        RECT 1794.070 54.440 1794.390 54.500 ;
      LAYER via ;
        RECT 1334.560 1684.060 1334.820 1684.320 ;
        RECT 1336.860 1684.060 1337.120 1684.320 ;
        RECT 1336.860 54.440 1337.120 54.700 ;
        RECT 1794.100 54.440 1794.360 54.700 ;
      LAYER met2 ;
        RECT 1334.460 1700.340 1334.740 1704.000 ;
        RECT 1334.460 1700.000 1334.760 1700.340 ;
        RECT 1334.620 1684.350 1334.760 1700.000 ;
        RECT 1334.560 1684.030 1334.820 1684.350 ;
        RECT 1336.860 1684.030 1337.120 1684.350 ;
        RECT 1336.920 54.730 1337.060 1684.030 ;
        RECT 1336.860 54.410 1337.120 54.730 ;
        RECT 1794.100 54.410 1794.360 54.730 ;
        RECT 1794.160 17.410 1794.300 54.410 ;
        RECT 1794.160 17.270 1798.900 17.410 ;
        RECT 1798.760 2.400 1798.900 17.270 ;
        RECT 1798.550 -4.800 1799.110 2.400 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1336.370 54.300 1336.690 54.360 ;
        RECT 1814.770 54.300 1815.090 54.360 ;
        RECT 1336.370 54.160 1815.090 54.300 ;
        RECT 1336.370 54.100 1336.690 54.160 ;
        RECT 1814.770 54.100 1815.090 54.160 ;
      LAYER via ;
        RECT 1336.400 54.100 1336.660 54.360 ;
        RECT 1814.800 54.100 1815.060 54.360 ;
      LAYER met2 ;
        RECT 1336.300 1700.340 1336.580 1704.000 ;
        RECT 1336.300 1700.000 1336.600 1700.340 ;
        RECT 1336.460 54.390 1336.600 1700.000 ;
        RECT 1336.400 54.070 1336.660 54.390 ;
        RECT 1814.800 54.070 1815.060 54.390 ;
        RECT 1814.860 17.410 1815.000 54.070 ;
        RECT 1814.860 17.270 1816.840 17.410 ;
        RECT 1816.700 2.400 1816.840 17.270 ;
        RECT 1816.490 -4.800 1817.050 2.400 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1331.770 1684.940 1332.090 1685.000 ;
        RECT 1338.210 1684.940 1338.530 1685.000 ;
        RECT 1331.770 1684.800 1338.530 1684.940 ;
        RECT 1331.770 1684.740 1332.090 1684.800 ;
        RECT 1338.210 1684.740 1338.530 1684.800 ;
        RECT 1331.770 53.960 1332.090 54.020 ;
        RECT 1828.570 53.960 1828.890 54.020 ;
        RECT 1331.770 53.820 1828.890 53.960 ;
        RECT 1331.770 53.760 1332.090 53.820 ;
        RECT 1828.570 53.760 1828.890 53.820 ;
        RECT 1828.570 20.980 1828.890 21.040 ;
        RECT 1834.550 20.980 1834.870 21.040 ;
        RECT 1828.570 20.840 1834.870 20.980 ;
        RECT 1828.570 20.780 1828.890 20.840 ;
        RECT 1834.550 20.780 1834.870 20.840 ;
      LAYER via ;
        RECT 1331.800 1684.740 1332.060 1685.000 ;
        RECT 1338.240 1684.740 1338.500 1685.000 ;
        RECT 1331.800 53.760 1332.060 54.020 ;
        RECT 1828.600 53.760 1828.860 54.020 ;
        RECT 1828.600 20.780 1828.860 21.040 ;
        RECT 1834.580 20.780 1834.840 21.040 ;
      LAYER met2 ;
        RECT 1338.140 1700.340 1338.420 1704.000 ;
        RECT 1338.140 1700.000 1338.440 1700.340 ;
        RECT 1338.300 1685.030 1338.440 1700.000 ;
        RECT 1331.800 1684.710 1332.060 1685.030 ;
        RECT 1338.240 1684.710 1338.500 1685.030 ;
        RECT 1331.860 54.050 1332.000 1684.710 ;
        RECT 1331.800 53.730 1332.060 54.050 ;
        RECT 1828.600 53.730 1828.860 54.050 ;
        RECT 1828.660 21.070 1828.800 53.730 ;
        RECT 1828.600 20.750 1828.860 21.070 ;
        RECT 1834.580 20.750 1834.840 21.070 ;
        RECT 1834.640 2.400 1834.780 20.750 ;
        RECT 1834.430 -4.800 1834.990 2.400 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1340.050 1656.180 1340.370 1656.440 ;
        RECT 1340.140 1656.040 1340.280 1656.180 ;
        RECT 1342.350 1656.040 1342.670 1656.100 ;
        RECT 1340.140 1655.900 1342.670 1656.040 ;
        RECT 1342.350 1655.840 1342.670 1655.900 ;
        RECT 1342.350 53.620 1342.670 53.680 ;
        RECT 1849.270 53.620 1849.590 53.680 ;
        RECT 1342.350 53.480 1849.590 53.620 ;
        RECT 1342.350 53.420 1342.670 53.480 ;
        RECT 1849.270 53.420 1849.590 53.480 ;
      LAYER via ;
        RECT 1340.080 1656.180 1340.340 1656.440 ;
        RECT 1342.380 1655.840 1342.640 1656.100 ;
        RECT 1342.380 53.420 1342.640 53.680 ;
        RECT 1849.300 53.420 1849.560 53.680 ;
      LAYER met2 ;
        RECT 1339.980 1700.340 1340.260 1704.000 ;
        RECT 1339.980 1700.000 1340.280 1700.340 ;
        RECT 1340.140 1656.470 1340.280 1700.000 ;
        RECT 1340.080 1656.150 1340.340 1656.470 ;
        RECT 1342.380 1655.810 1342.640 1656.130 ;
        RECT 1342.440 53.710 1342.580 1655.810 ;
        RECT 1342.380 53.390 1342.640 53.710 ;
        RECT 1849.300 53.390 1849.560 53.710 ;
        RECT 1849.360 17.410 1849.500 53.390 ;
        RECT 1849.360 17.270 1852.260 17.410 ;
        RECT 1852.120 2.400 1852.260 17.270 ;
        RECT 1851.910 -4.800 1852.470 2.400 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1342.810 53.280 1343.130 53.340 ;
        RECT 1870.430 53.280 1870.750 53.340 ;
        RECT 1342.810 53.140 1870.750 53.280 ;
        RECT 1342.810 53.080 1343.130 53.140 ;
        RECT 1870.430 53.080 1870.750 53.140 ;
      LAYER via ;
        RECT 1342.840 53.080 1343.100 53.340 ;
        RECT 1870.460 53.080 1870.720 53.340 ;
      LAYER met2 ;
        RECT 1341.820 1700.410 1342.100 1704.000 ;
        RECT 1341.820 1700.270 1342.580 1700.410 ;
        RECT 1341.820 1700.000 1342.100 1700.270 ;
        RECT 1342.440 1677.970 1342.580 1700.270 ;
        RECT 1342.440 1677.830 1343.040 1677.970 ;
        RECT 1342.900 53.370 1343.040 1677.830 ;
        RECT 1342.840 53.050 1343.100 53.370 ;
        RECT 1870.460 53.050 1870.720 53.370 ;
        RECT 1870.520 7.210 1870.660 53.050 ;
        RECT 1870.060 7.070 1870.660 7.210 ;
        RECT 1870.060 2.400 1870.200 7.070 ;
        RECT 1869.850 -4.800 1870.410 2.400 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1221.830 1676.780 1222.150 1676.840 ;
        RECT 1225.970 1676.780 1226.290 1676.840 ;
        RECT 1221.830 1676.640 1226.290 1676.780 ;
        RECT 1221.830 1676.580 1222.150 1676.640 ;
        RECT 1225.970 1676.580 1226.290 1676.640 ;
        RECT 751.710 1639.380 752.030 1639.440 ;
        RECT 1221.830 1639.380 1222.150 1639.440 ;
        RECT 751.710 1639.240 1222.150 1639.380 ;
        RECT 751.710 1639.180 752.030 1639.240 ;
        RECT 1221.830 1639.180 1222.150 1639.240 ;
      LAYER via ;
        RECT 1221.860 1676.580 1222.120 1676.840 ;
        RECT 1226.000 1676.580 1226.260 1676.840 ;
        RECT 751.740 1639.180 752.000 1639.440 ;
        RECT 1221.860 1639.180 1222.120 1639.440 ;
      LAYER met2 ;
        RECT 1226.360 1700.410 1226.640 1704.000 ;
        RECT 1226.060 1700.270 1226.640 1700.410 ;
        RECT 1226.060 1676.870 1226.200 1700.270 ;
        RECT 1226.360 1700.000 1226.640 1700.270 ;
        RECT 1221.860 1676.550 1222.120 1676.870 ;
        RECT 1226.000 1676.550 1226.260 1676.870 ;
        RECT 1221.920 1639.470 1222.060 1676.550 ;
        RECT 751.740 1639.150 752.000 1639.470 ;
        RECT 1221.860 1639.150 1222.120 1639.470 ;
        RECT 751.800 16.730 751.940 1639.150 ;
        RECT 746.280 16.590 751.940 16.730 ;
        RECT 746.280 2.400 746.420 16.590 ;
        RECT 746.070 -4.800 746.630 2.400 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1343.730 52.940 1344.050 53.000 ;
        RECT 1883.770 52.940 1884.090 53.000 ;
        RECT 1343.730 52.800 1884.090 52.940 ;
        RECT 1343.730 52.740 1344.050 52.800 ;
        RECT 1883.770 52.740 1884.090 52.800 ;
      LAYER via ;
        RECT 1343.760 52.740 1344.020 53.000 ;
        RECT 1883.800 52.740 1884.060 53.000 ;
      LAYER met2 ;
        RECT 1343.660 1700.340 1343.940 1704.000 ;
        RECT 1343.660 1700.000 1343.960 1700.340 ;
        RECT 1343.820 53.030 1343.960 1700.000 ;
        RECT 1343.760 52.710 1344.020 53.030 ;
        RECT 1883.800 52.710 1884.060 53.030 ;
        RECT 1883.860 17.410 1884.000 52.710 ;
        RECT 1883.860 17.270 1888.140 17.410 ;
        RECT 1888.000 2.400 1888.140 17.270 ;
        RECT 1887.790 -4.800 1888.350 2.400 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1345.570 1628.500 1345.890 1628.560 ;
        RECT 1346.030 1628.500 1346.350 1628.560 ;
        RECT 1345.570 1628.360 1346.350 1628.500 ;
        RECT 1345.570 1628.300 1345.890 1628.360 ;
        RECT 1346.030 1628.300 1346.350 1628.360 ;
        RECT 1345.570 52.600 1345.890 52.660 ;
        RECT 1904.470 52.600 1904.790 52.660 ;
        RECT 1345.570 52.460 1904.790 52.600 ;
        RECT 1345.570 52.400 1345.890 52.460 ;
        RECT 1904.470 52.400 1904.790 52.460 ;
      LAYER via ;
        RECT 1345.600 1628.300 1345.860 1628.560 ;
        RECT 1346.060 1628.300 1346.320 1628.560 ;
        RECT 1345.600 52.400 1345.860 52.660 ;
        RECT 1904.500 52.400 1904.760 52.660 ;
      LAYER met2 ;
        RECT 1345.500 1700.340 1345.780 1704.000 ;
        RECT 1345.500 1700.000 1345.800 1700.340 ;
        RECT 1345.660 1629.690 1345.800 1700.000 ;
        RECT 1345.660 1629.550 1346.260 1629.690 ;
        RECT 1346.120 1628.590 1346.260 1629.550 ;
        RECT 1345.600 1628.270 1345.860 1628.590 ;
        RECT 1346.060 1628.270 1346.320 1628.590 ;
        RECT 1345.660 52.690 1345.800 1628.270 ;
        RECT 1345.600 52.370 1345.860 52.690 ;
        RECT 1904.500 52.370 1904.760 52.690 ;
        RECT 1904.560 17.410 1904.700 52.370 ;
        RECT 1904.560 17.270 1906.080 17.410 ;
        RECT 1905.940 2.400 1906.080 17.270 ;
        RECT 1905.730 -4.800 1906.290 2.400 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1347.870 1677.460 1348.190 1677.520 ;
        RECT 1349.710 1677.460 1350.030 1677.520 ;
        RECT 1347.870 1677.320 1350.030 1677.460 ;
        RECT 1347.870 1677.260 1348.190 1677.320 ;
        RECT 1349.710 1677.260 1350.030 1677.320 ;
        RECT 1349.710 52.260 1350.030 52.320 ;
        RECT 1918.270 52.260 1918.590 52.320 ;
        RECT 1349.710 52.120 1918.590 52.260 ;
        RECT 1349.710 52.060 1350.030 52.120 ;
        RECT 1918.270 52.060 1918.590 52.120 ;
      LAYER via ;
        RECT 1347.900 1677.260 1348.160 1677.520 ;
        RECT 1349.740 1677.260 1350.000 1677.520 ;
        RECT 1349.740 52.060 1350.000 52.320 ;
        RECT 1918.300 52.060 1918.560 52.320 ;
      LAYER met2 ;
        RECT 1347.340 1700.410 1347.620 1704.000 ;
        RECT 1347.340 1700.270 1348.100 1700.410 ;
        RECT 1347.340 1700.000 1347.620 1700.270 ;
        RECT 1347.960 1677.550 1348.100 1700.270 ;
        RECT 1347.900 1677.230 1348.160 1677.550 ;
        RECT 1349.740 1677.230 1350.000 1677.550 ;
        RECT 1349.800 52.350 1349.940 1677.230 ;
        RECT 1349.740 52.030 1350.000 52.350 ;
        RECT 1918.300 52.030 1918.560 52.350 ;
        RECT 1918.360 17.410 1918.500 52.030 ;
        RECT 1918.360 17.270 1923.560 17.410 ;
        RECT 1923.420 2.400 1923.560 17.270 ;
        RECT 1923.210 -4.800 1923.770 2.400 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1346.490 1678.480 1346.810 1678.540 ;
        RECT 1349.250 1678.480 1349.570 1678.540 ;
        RECT 1346.490 1678.340 1349.570 1678.480 ;
        RECT 1346.490 1678.280 1346.810 1678.340 ;
        RECT 1349.250 1678.280 1349.570 1678.340 ;
        RECT 1346.490 51.920 1346.810 51.980 ;
        RECT 1938.970 51.920 1939.290 51.980 ;
        RECT 1346.490 51.780 1939.290 51.920 ;
        RECT 1346.490 51.720 1346.810 51.780 ;
        RECT 1938.970 51.720 1939.290 51.780 ;
      LAYER via ;
        RECT 1346.520 1678.280 1346.780 1678.540 ;
        RECT 1349.280 1678.280 1349.540 1678.540 ;
        RECT 1346.520 51.720 1346.780 51.980 ;
        RECT 1939.000 51.720 1939.260 51.980 ;
      LAYER met2 ;
        RECT 1349.180 1700.340 1349.460 1704.000 ;
        RECT 1349.180 1700.000 1349.480 1700.340 ;
        RECT 1349.340 1678.570 1349.480 1700.000 ;
        RECT 1346.520 1678.250 1346.780 1678.570 ;
        RECT 1349.280 1678.250 1349.540 1678.570 ;
        RECT 1346.580 52.010 1346.720 1678.250 ;
        RECT 1346.520 51.690 1346.780 52.010 ;
        RECT 1939.000 51.690 1939.260 52.010 ;
        RECT 1939.060 17.410 1939.200 51.690 ;
        RECT 1939.060 17.270 1941.500 17.410 ;
        RECT 1941.360 2.400 1941.500 17.270 ;
        RECT 1941.150 -4.800 1941.710 2.400 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1350.170 1683.920 1350.490 1683.980 ;
        RECT 1351.090 1683.920 1351.410 1683.980 ;
        RECT 1350.170 1683.780 1351.410 1683.920 ;
        RECT 1350.170 1683.720 1350.490 1683.780 ;
        RECT 1351.090 1683.720 1351.410 1683.780 ;
        RECT 1350.170 51.580 1350.490 51.640 ;
        RECT 1952.770 51.580 1953.090 51.640 ;
        RECT 1350.170 51.440 1953.090 51.580 ;
        RECT 1350.170 51.380 1350.490 51.440 ;
        RECT 1952.770 51.380 1953.090 51.440 ;
        RECT 1952.770 14.180 1953.090 14.240 ;
        RECT 1959.210 14.180 1959.530 14.240 ;
        RECT 1952.770 14.040 1959.530 14.180 ;
        RECT 1952.770 13.980 1953.090 14.040 ;
        RECT 1959.210 13.980 1959.530 14.040 ;
      LAYER via ;
        RECT 1350.200 1683.720 1350.460 1683.980 ;
        RECT 1351.120 1683.720 1351.380 1683.980 ;
        RECT 1350.200 51.380 1350.460 51.640 ;
        RECT 1952.800 51.380 1953.060 51.640 ;
        RECT 1952.800 13.980 1953.060 14.240 ;
        RECT 1959.240 13.980 1959.500 14.240 ;
      LAYER met2 ;
        RECT 1351.020 1700.340 1351.300 1704.000 ;
        RECT 1351.020 1700.000 1351.320 1700.340 ;
        RECT 1351.180 1684.010 1351.320 1700.000 ;
        RECT 1350.200 1683.690 1350.460 1684.010 ;
        RECT 1351.120 1683.690 1351.380 1684.010 ;
        RECT 1350.260 51.670 1350.400 1683.690 ;
        RECT 1350.200 51.350 1350.460 51.670 ;
        RECT 1952.800 51.350 1953.060 51.670 ;
        RECT 1952.860 14.270 1953.000 51.350 ;
        RECT 1952.800 13.950 1953.060 14.270 ;
        RECT 1959.240 13.950 1959.500 14.270 ;
        RECT 1959.300 2.400 1959.440 13.950 ;
        RECT 1959.090 -4.800 1959.650 2.400 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1352.930 1684.600 1353.250 1684.660 ;
        RECT 1356.150 1684.600 1356.470 1684.660 ;
        RECT 1352.930 1684.460 1356.470 1684.600 ;
        RECT 1352.930 1684.400 1353.250 1684.460 ;
        RECT 1356.150 1684.400 1356.470 1684.460 ;
        RECT 1356.150 1625.780 1356.470 1625.840 ;
        RECT 1973.470 1625.780 1973.790 1625.840 ;
        RECT 1356.150 1625.640 1973.790 1625.780 ;
        RECT 1356.150 1625.580 1356.470 1625.640 ;
        RECT 1973.470 1625.580 1973.790 1625.640 ;
      LAYER via ;
        RECT 1352.960 1684.400 1353.220 1684.660 ;
        RECT 1356.180 1684.400 1356.440 1684.660 ;
        RECT 1356.180 1625.580 1356.440 1625.840 ;
        RECT 1973.500 1625.580 1973.760 1625.840 ;
      LAYER met2 ;
        RECT 1352.860 1700.340 1353.140 1704.000 ;
        RECT 1352.860 1700.000 1353.160 1700.340 ;
        RECT 1353.020 1684.690 1353.160 1700.000 ;
        RECT 1352.960 1684.370 1353.220 1684.690 ;
        RECT 1356.180 1684.370 1356.440 1684.690 ;
        RECT 1356.240 1625.870 1356.380 1684.370 ;
        RECT 1356.180 1625.550 1356.440 1625.870 ;
        RECT 1973.500 1625.550 1973.760 1625.870 ;
        RECT 1973.560 17.410 1973.700 1625.550 ;
        RECT 1973.560 17.270 1977.380 17.410 ;
        RECT 1977.240 2.400 1977.380 17.270 ;
        RECT 1977.030 -4.800 1977.590 2.400 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1354.770 1618.980 1355.090 1619.040 ;
        RECT 1994.170 1618.980 1994.490 1619.040 ;
        RECT 1354.770 1618.840 1994.490 1618.980 ;
        RECT 1354.770 1618.780 1355.090 1618.840 ;
        RECT 1994.170 1618.780 1994.490 1618.840 ;
      LAYER via ;
        RECT 1354.800 1618.780 1355.060 1619.040 ;
        RECT 1994.200 1618.780 1994.460 1619.040 ;
      LAYER met2 ;
        RECT 1354.700 1700.340 1354.980 1704.000 ;
        RECT 1354.700 1700.000 1355.000 1700.340 ;
        RECT 1354.860 1619.070 1355.000 1700.000 ;
        RECT 1354.800 1618.750 1355.060 1619.070 ;
        RECT 1994.200 1618.750 1994.460 1619.070 ;
        RECT 1994.260 17.410 1994.400 1618.750 ;
        RECT 1994.260 17.270 1995.320 17.410 ;
        RECT 1995.180 2.400 1995.320 17.270 ;
        RECT 1994.970 -4.800 1995.530 2.400 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1357.070 1556.080 1357.390 1556.140 ;
        RECT 2007.970 1556.080 2008.290 1556.140 ;
        RECT 1357.070 1555.940 2008.290 1556.080 ;
        RECT 1357.070 1555.880 1357.390 1555.940 ;
        RECT 2007.970 1555.880 2008.290 1555.940 ;
      LAYER via ;
        RECT 1357.100 1555.880 1357.360 1556.140 ;
        RECT 2008.000 1555.880 2008.260 1556.140 ;
      LAYER met2 ;
        RECT 1356.540 1700.410 1356.820 1704.000 ;
        RECT 1356.540 1700.270 1357.300 1700.410 ;
        RECT 1356.540 1700.000 1356.820 1700.270 ;
        RECT 1357.160 1556.170 1357.300 1700.270 ;
        RECT 1357.100 1555.850 1357.360 1556.170 ;
        RECT 2008.000 1555.850 2008.260 1556.170 ;
        RECT 2008.060 17.410 2008.200 1555.850 ;
        RECT 2008.060 17.270 2012.800 17.410 ;
        RECT 2012.660 2.400 2012.800 17.270 ;
        RECT 2012.450 -4.800 2013.010 2.400 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1358.450 1584.300 1358.770 1584.360 ;
        RECT 2028.670 1584.300 2028.990 1584.360 ;
        RECT 1358.450 1584.160 2028.990 1584.300 ;
        RECT 1358.450 1584.100 1358.770 1584.160 ;
        RECT 2028.670 1584.100 2028.990 1584.160 ;
      LAYER via ;
        RECT 1358.480 1584.100 1358.740 1584.360 ;
        RECT 2028.700 1584.100 2028.960 1584.360 ;
      LAYER met2 ;
        RECT 1358.380 1700.340 1358.660 1704.000 ;
        RECT 1358.380 1700.000 1358.680 1700.340 ;
        RECT 1358.540 1584.390 1358.680 1700.000 ;
        RECT 1358.480 1584.070 1358.740 1584.390 ;
        RECT 2028.700 1584.070 2028.960 1584.390 ;
        RECT 2028.760 17.410 2028.900 1584.070 ;
        RECT 2028.760 17.270 2030.740 17.410 ;
        RECT 2030.600 2.400 2030.740 17.270 ;
        RECT 2030.390 -4.800 2030.950 2.400 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1360.290 1577.160 1360.610 1577.220 ;
        RECT 2042.930 1577.160 2043.250 1577.220 ;
        RECT 1360.290 1577.020 2043.250 1577.160 ;
        RECT 1360.290 1576.960 1360.610 1577.020 ;
        RECT 2042.930 1576.960 2043.250 1577.020 ;
      LAYER via ;
        RECT 1360.320 1576.960 1360.580 1577.220 ;
        RECT 2042.960 1576.960 2043.220 1577.220 ;
      LAYER met2 ;
        RECT 1360.220 1700.340 1360.500 1704.000 ;
        RECT 1360.220 1700.000 1360.520 1700.340 ;
        RECT 1360.380 1577.250 1360.520 1700.000 ;
        RECT 1360.320 1576.930 1360.580 1577.250 ;
        RECT 2042.960 1576.930 2043.220 1577.250 ;
        RECT 2043.020 17.410 2043.160 1576.930 ;
        RECT 2043.020 17.270 2048.680 17.410 ;
        RECT 2048.540 2.400 2048.680 17.270 ;
        RECT 2048.330 -4.800 2048.890 2.400 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 765.510 1646.520 765.830 1646.580 ;
        RECT 1230.110 1646.520 1230.430 1646.580 ;
        RECT 765.510 1646.380 1230.430 1646.520 ;
        RECT 765.510 1646.320 765.830 1646.380 ;
        RECT 1230.110 1646.320 1230.430 1646.380 ;
      LAYER via ;
        RECT 765.540 1646.320 765.800 1646.580 ;
        RECT 1230.140 1646.320 1230.400 1646.580 ;
      LAYER met2 ;
        RECT 1228.200 1700.340 1228.480 1704.000 ;
        RECT 1228.200 1700.000 1228.500 1700.340 ;
        RECT 1228.360 1677.970 1228.500 1700.000 ;
        RECT 1228.360 1677.830 1230.340 1677.970 ;
        RECT 1230.200 1646.610 1230.340 1677.830 ;
        RECT 765.540 1646.290 765.800 1646.610 ;
        RECT 1230.140 1646.290 1230.400 1646.610 ;
        RECT 765.600 18.090 765.740 1646.290 ;
        RECT 763.760 17.950 765.740 18.090 ;
        RECT 763.760 2.400 763.900 17.950 ;
        RECT 763.550 -4.800 764.110 2.400 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1362.130 1683.920 1362.450 1683.980 ;
        RECT 1363.510 1683.920 1363.830 1683.980 ;
        RECT 1362.130 1683.780 1363.830 1683.920 ;
        RECT 1362.130 1683.720 1362.450 1683.780 ;
        RECT 1363.510 1683.720 1363.830 1683.780 ;
        RECT 1363.510 1536.020 1363.830 1536.080 ;
        RECT 2063.170 1536.020 2063.490 1536.080 ;
        RECT 1363.510 1535.880 2063.490 1536.020 ;
        RECT 1363.510 1535.820 1363.830 1535.880 ;
        RECT 2063.170 1535.820 2063.490 1535.880 ;
      LAYER via ;
        RECT 1362.160 1683.720 1362.420 1683.980 ;
        RECT 1363.540 1683.720 1363.800 1683.980 ;
        RECT 1363.540 1535.820 1363.800 1536.080 ;
        RECT 2063.200 1535.820 2063.460 1536.080 ;
      LAYER met2 ;
        RECT 1362.060 1700.340 1362.340 1704.000 ;
        RECT 1362.060 1700.000 1362.360 1700.340 ;
        RECT 1362.220 1684.010 1362.360 1700.000 ;
        RECT 1362.160 1683.690 1362.420 1684.010 ;
        RECT 1363.540 1683.690 1363.800 1684.010 ;
        RECT 1363.600 1536.110 1363.740 1683.690 ;
        RECT 1363.540 1535.790 1363.800 1536.110 ;
        RECT 2063.200 1535.790 2063.460 1536.110 ;
        RECT 2063.260 17.410 2063.400 1535.790 ;
        RECT 2063.260 17.270 2066.620 17.410 ;
        RECT 2066.480 2.400 2066.620 17.270 ;
        RECT 2066.270 -4.800 2066.830 2.400 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1363.970 1528.540 1364.290 1528.600 ;
        RECT 2084.330 1528.540 2084.650 1528.600 ;
        RECT 1363.970 1528.400 2084.650 1528.540 ;
        RECT 1363.970 1528.340 1364.290 1528.400 ;
        RECT 2084.330 1528.340 2084.650 1528.400 ;
      LAYER via ;
        RECT 1364.000 1528.340 1364.260 1528.600 ;
        RECT 2084.360 1528.340 2084.620 1528.600 ;
      LAYER met2 ;
        RECT 1363.900 1700.340 1364.180 1704.000 ;
        RECT 1363.900 1700.000 1364.200 1700.340 ;
        RECT 1364.060 1528.630 1364.200 1700.000 ;
        RECT 1364.000 1528.310 1364.260 1528.630 ;
        RECT 2084.360 1528.310 2084.620 1528.630 ;
        RECT 2084.420 2.400 2084.560 1528.310 ;
        RECT 2084.210 -4.800 2084.770 2.400 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1364.430 1683.920 1364.750 1683.980 ;
        RECT 1365.810 1683.920 1366.130 1683.980 ;
        RECT 1364.430 1683.780 1366.130 1683.920 ;
        RECT 1364.430 1683.720 1364.750 1683.780 ;
        RECT 1365.810 1683.720 1366.130 1683.780 ;
        RECT 1364.430 1459.520 1364.750 1459.580 ;
        RECT 2097.670 1459.520 2097.990 1459.580 ;
        RECT 1364.430 1459.380 2097.990 1459.520 ;
        RECT 1364.430 1459.320 1364.750 1459.380 ;
        RECT 2097.670 1459.320 2097.990 1459.380 ;
      LAYER via ;
        RECT 1364.460 1683.720 1364.720 1683.980 ;
        RECT 1365.840 1683.720 1366.100 1683.980 ;
        RECT 1364.460 1459.320 1364.720 1459.580 ;
        RECT 2097.700 1459.320 2097.960 1459.580 ;
      LAYER met2 ;
        RECT 1365.740 1700.340 1366.020 1704.000 ;
        RECT 1365.740 1700.000 1366.040 1700.340 ;
        RECT 1365.900 1684.010 1366.040 1700.000 ;
        RECT 1364.460 1683.690 1364.720 1684.010 ;
        RECT 1365.840 1683.690 1366.100 1684.010 ;
        RECT 1364.520 1459.610 1364.660 1683.690 ;
        RECT 1364.460 1459.290 1364.720 1459.610 ;
        RECT 2097.700 1459.290 2097.960 1459.610 ;
        RECT 2097.760 17.410 2097.900 1459.290 ;
        RECT 2097.760 17.270 2102.040 17.410 ;
        RECT 2101.900 2.400 2102.040 17.270 ;
        RECT 2101.690 -4.800 2102.250 2.400 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1367.650 1570.360 1367.970 1570.420 ;
        RECT 2118.370 1570.360 2118.690 1570.420 ;
        RECT 1367.650 1570.220 2118.690 1570.360 ;
        RECT 1367.650 1570.160 1367.970 1570.220 ;
        RECT 2118.370 1570.160 2118.690 1570.220 ;
      LAYER via ;
        RECT 1367.680 1570.160 1367.940 1570.420 ;
        RECT 2118.400 1570.160 2118.660 1570.420 ;
      LAYER met2 ;
        RECT 1367.580 1700.340 1367.860 1704.000 ;
        RECT 1367.580 1700.000 1367.880 1700.340 ;
        RECT 1367.740 1570.450 1367.880 1700.000 ;
        RECT 1367.680 1570.130 1367.940 1570.450 ;
        RECT 2118.400 1570.130 2118.660 1570.450 ;
        RECT 2118.460 17.410 2118.600 1570.130 ;
        RECT 2118.460 17.270 2119.980 17.410 ;
        RECT 2119.840 2.400 2119.980 17.270 ;
        RECT 2119.630 -4.800 2120.190 2.400 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1370.410 1521.740 1370.730 1521.800 ;
        RECT 2132.170 1521.740 2132.490 1521.800 ;
        RECT 1370.410 1521.600 2132.490 1521.740 ;
        RECT 1370.410 1521.540 1370.730 1521.600 ;
        RECT 2132.170 1521.540 2132.490 1521.600 ;
      LAYER via ;
        RECT 1370.440 1521.540 1370.700 1521.800 ;
        RECT 2132.200 1521.540 2132.460 1521.800 ;
      LAYER met2 ;
        RECT 1369.420 1700.410 1369.700 1704.000 ;
        RECT 1369.420 1700.270 1370.180 1700.410 ;
        RECT 1369.420 1700.000 1369.700 1700.270 ;
        RECT 1370.040 1618.130 1370.180 1700.270 ;
        RECT 1370.040 1617.990 1370.640 1618.130 ;
        RECT 1370.500 1521.830 1370.640 1617.990 ;
        RECT 1370.440 1521.510 1370.700 1521.830 ;
        RECT 2132.200 1521.510 2132.460 1521.830 ;
        RECT 2132.260 17.410 2132.400 1521.510 ;
        RECT 2132.260 17.270 2137.920 17.410 ;
        RECT 2137.780 2.400 2137.920 17.270 ;
        RECT 2137.570 -4.800 2138.130 2.400 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1370.870 1452.720 1371.190 1452.780 ;
        RECT 2152.870 1452.720 2153.190 1452.780 ;
        RECT 1370.870 1452.580 2153.190 1452.720 ;
        RECT 1370.870 1452.520 1371.190 1452.580 ;
        RECT 2152.870 1452.520 2153.190 1452.580 ;
      LAYER via ;
        RECT 1370.900 1452.520 1371.160 1452.780 ;
        RECT 2152.900 1452.520 2153.160 1452.780 ;
      LAYER met2 ;
        RECT 1371.260 1700.340 1371.540 1704.000 ;
        RECT 1371.260 1700.000 1371.560 1700.340 ;
        RECT 1371.420 1666.410 1371.560 1700.000 ;
        RECT 1370.960 1666.270 1371.560 1666.410 ;
        RECT 1370.960 1452.810 1371.100 1666.270 ;
        RECT 1370.900 1452.490 1371.160 1452.810 ;
        RECT 2152.900 1452.490 2153.160 1452.810 ;
        RECT 2152.960 17.410 2153.100 1452.490 ;
        RECT 2152.960 17.270 2155.860 17.410 ;
        RECT 2155.720 2.400 2155.860 17.270 ;
        RECT 2155.510 -4.800 2156.070 2.400 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1399.465 1632.425 1399.635 1633.955 ;
      LAYER mcon ;
        RECT 1399.465 1633.785 1399.635 1633.955 ;
      LAYER met1 ;
        RECT 1373.170 1633.940 1373.490 1634.000 ;
        RECT 1399.405 1633.940 1399.695 1633.985 ;
        RECT 1373.170 1633.800 1399.695 1633.940 ;
        RECT 1373.170 1633.740 1373.490 1633.800 ;
        RECT 1399.405 1633.755 1399.695 1633.800 ;
        RECT 1399.405 1632.580 1399.695 1632.625 ;
        RECT 2167.130 1632.580 2167.450 1632.640 ;
        RECT 1399.405 1632.440 2167.450 1632.580 ;
        RECT 1399.405 1632.395 1399.695 1632.440 ;
        RECT 2167.130 1632.380 2167.450 1632.440 ;
        RECT 2167.130 19.280 2167.450 19.340 ;
        RECT 2173.110 19.280 2173.430 19.340 ;
        RECT 2167.130 19.140 2173.430 19.280 ;
        RECT 2167.130 19.080 2167.450 19.140 ;
        RECT 2173.110 19.080 2173.430 19.140 ;
      LAYER via ;
        RECT 1373.200 1633.740 1373.460 1634.000 ;
        RECT 2167.160 1632.380 2167.420 1632.640 ;
        RECT 2167.160 19.080 2167.420 19.340 ;
        RECT 2173.140 19.080 2173.400 19.340 ;
      LAYER met2 ;
        RECT 1373.100 1700.340 1373.380 1704.000 ;
        RECT 1373.100 1700.000 1373.400 1700.340 ;
        RECT 1373.260 1634.030 1373.400 1700.000 ;
        RECT 1373.200 1633.710 1373.460 1634.030 ;
        RECT 2167.160 1632.350 2167.420 1632.670 ;
        RECT 2167.220 19.370 2167.360 1632.350 ;
        RECT 2167.160 19.050 2167.420 19.370 ;
        RECT 2173.140 19.050 2173.400 19.370 ;
        RECT 2173.200 2.400 2173.340 19.050 ;
        RECT 2172.990 -4.800 2173.550 2.400 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1375.010 1683.920 1375.330 1683.980 ;
        RECT 1376.850 1683.920 1377.170 1683.980 ;
        RECT 1375.010 1683.780 1377.170 1683.920 ;
        RECT 1375.010 1683.720 1375.330 1683.780 ;
        RECT 1376.850 1683.720 1377.170 1683.780 ;
        RECT 1376.850 1563.560 1377.170 1563.620 ;
        RECT 2187.370 1563.560 2187.690 1563.620 ;
        RECT 1376.850 1563.420 2187.690 1563.560 ;
        RECT 1376.850 1563.360 1377.170 1563.420 ;
        RECT 2187.370 1563.360 2187.690 1563.420 ;
      LAYER via ;
        RECT 1375.040 1683.720 1375.300 1683.980 ;
        RECT 1376.880 1683.720 1377.140 1683.980 ;
        RECT 1376.880 1563.360 1377.140 1563.620 ;
        RECT 2187.400 1563.360 2187.660 1563.620 ;
      LAYER met2 ;
        RECT 1374.940 1700.340 1375.220 1704.000 ;
        RECT 1374.940 1700.000 1375.240 1700.340 ;
        RECT 1375.100 1684.010 1375.240 1700.000 ;
        RECT 1375.040 1683.690 1375.300 1684.010 ;
        RECT 1376.880 1683.690 1377.140 1684.010 ;
        RECT 1376.940 1563.650 1377.080 1683.690 ;
        RECT 1376.880 1563.330 1377.140 1563.650 ;
        RECT 2187.400 1563.330 2187.660 1563.650 ;
        RECT 2187.460 17.410 2187.600 1563.330 ;
        RECT 2187.460 17.270 2191.280 17.410 ;
        RECT 2191.140 2.400 2191.280 17.270 ;
        RECT 2190.930 -4.800 2191.490 2.400 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1374.090 1684.600 1374.410 1684.660 ;
        RECT 1376.850 1684.600 1377.170 1684.660 ;
        RECT 1374.090 1684.460 1377.170 1684.600 ;
        RECT 1374.090 1684.400 1374.410 1684.460 ;
        RECT 1376.850 1684.400 1377.170 1684.460 ;
        RECT 1374.550 1555.740 1374.870 1555.800 ;
        RECT 2208.070 1555.740 2208.390 1555.800 ;
        RECT 1374.550 1555.600 2208.390 1555.740 ;
        RECT 1374.550 1555.540 1374.870 1555.600 ;
        RECT 2208.070 1555.540 2208.390 1555.600 ;
      LAYER via ;
        RECT 1374.120 1684.400 1374.380 1684.660 ;
        RECT 1376.880 1684.400 1377.140 1684.660 ;
        RECT 1374.580 1555.540 1374.840 1555.800 ;
        RECT 2208.100 1555.540 2208.360 1555.800 ;
      LAYER met2 ;
        RECT 1376.780 1700.340 1377.060 1704.000 ;
        RECT 1376.780 1700.000 1377.080 1700.340 ;
        RECT 1376.940 1684.690 1377.080 1700.000 ;
        RECT 1374.120 1684.370 1374.380 1684.690 ;
        RECT 1376.880 1684.370 1377.140 1684.690 ;
        RECT 1374.180 1666.410 1374.320 1684.370 ;
        RECT 1374.180 1666.270 1374.780 1666.410 ;
        RECT 1374.640 1555.830 1374.780 1666.270 ;
        RECT 1374.580 1555.510 1374.840 1555.830 ;
        RECT 2208.100 1555.510 2208.360 1555.830 ;
        RECT 2208.160 17.410 2208.300 1555.510 ;
        RECT 2208.160 17.270 2209.220 17.410 ;
        RECT 2209.080 2.400 2209.220 17.270 ;
        RECT 2208.870 -4.800 2209.430 2.400 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1377.770 1514.940 1378.090 1515.000 ;
        RECT 2221.870 1514.940 2222.190 1515.000 ;
        RECT 1377.770 1514.800 2222.190 1514.940 ;
        RECT 1377.770 1514.740 1378.090 1514.800 ;
        RECT 2221.870 1514.740 2222.190 1514.800 ;
      LAYER via ;
        RECT 1377.800 1514.740 1378.060 1515.000 ;
        RECT 2221.900 1514.740 2222.160 1515.000 ;
      LAYER met2 ;
        RECT 1378.620 1700.340 1378.900 1704.000 ;
        RECT 1378.620 1700.000 1378.920 1700.340 ;
        RECT 1378.780 1674.570 1378.920 1700.000 ;
        RECT 1377.860 1674.430 1378.920 1674.570 ;
        RECT 1377.860 1515.030 1378.000 1674.430 ;
        RECT 1377.800 1514.710 1378.060 1515.030 ;
        RECT 2221.900 1514.710 2222.160 1515.030 ;
        RECT 2221.960 17.410 2222.100 1514.710 ;
        RECT 2221.960 17.270 2227.160 17.410 ;
        RECT 2227.020 2.400 2227.160 17.270 ;
        RECT 2226.810 -4.800 2227.370 2.400 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1230.110 1678.480 1230.430 1678.540 ;
        RECT 1233.330 1678.480 1233.650 1678.540 ;
        RECT 1230.110 1678.340 1233.650 1678.480 ;
        RECT 1230.110 1678.280 1230.430 1678.340 ;
        RECT 1233.330 1678.280 1233.650 1678.340 ;
        RECT 786.210 1632.580 786.530 1632.640 ;
        RECT 1233.330 1632.580 1233.650 1632.640 ;
        RECT 786.210 1632.440 1233.650 1632.580 ;
        RECT 786.210 1632.380 786.530 1632.440 ;
        RECT 1233.330 1632.380 1233.650 1632.440 ;
      LAYER via ;
        RECT 1230.140 1678.280 1230.400 1678.540 ;
        RECT 1233.360 1678.280 1233.620 1678.540 ;
        RECT 786.240 1632.380 786.500 1632.640 ;
        RECT 1233.360 1632.380 1233.620 1632.640 ;
      LAYER met2 ;
        RECT 1230.040 1700.340 1230.320 1704.000 ;
        RECT 1230.040 1700.000 1230.340 1700.340 ;
        RECT 1230.200 1678.570 1230.340 1700.000 ;
        RECT 1230.140 1678.250 1230.400 1678.570 ;
        RECT 1233.360 1678.250 1233.620 1678.570 ;
        RECT 1233.420 1632.670 1233.560 1678.250 ;
        RECT 786.240 1632.350 786.500 1632.670 ;
        RECT 1233.360 1632.350 1233.620 1632.670 ;
        RECT 786.300 18.090 786.440 1632.350 ;
        RECT 781.700 17.950 786.440 18.090 ;
        RECT 781.700 2.400 781.840 17.950 ;
        RECT 781.490 -4.800 782.050 2.400 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1380.530 1684.940 1380.850 1685.000 ;
        RECT 1385.130 1684.940 1385.450 1685.000 ;
        RECT 1380.530 1684.800 1385.450 1684.940 ;
        RECT 1380.530 1684.740 1380.850 1684.800 ;
        RECT 1385.130 1684.740 1385.450 1684.800 ;
        RECT 1385.130 1507.800 1385.450 1507.860 ;
        RECT 2242.570 1507.800 2242.890 1507.860 ;
        RECT 1385.130 1507.660 2242.890 1507.800 ;
        RECT 1385.130 1507.600 1385.450 1507.660 ;
        RECT 2242.570 1507.600 2242.890 1507.660 ;
      LAYER via ;
        RECT 1380.560 1684.740 1380.820 1685.000 ;
        RECT 1385.160 1684.740 1385.420 1685.000 ;
        RECT 1385.160 1507.600 1385.420 1507.860 ;
        RECT 2242.600 1507.600 2242.860 1507.860 ;
      LAYER met2 ;
        RECT 1380.460 1700.340 1380.740 1704.000 ;
        RECT 1380.460 1700.000 1380.760 1700.340 ;
        RECT 1380.620 1685.030 1380.760 1700.000 ;
        RECT 1380.560 1684.710 1380.820 1685.030 ;
        RECT 1385.160 1684.710 1385.420 1685.030 ;
        RECT 1385.220 1507.890 1385.360 1684.710 ;
        RECT 1385.160 1507.570 1385.420 1507.890 ;
        RECT 2242.600 1507.570 2242.860 1507.890 ;
        RECT 2242.660 17.410 2242.800 1507.570 ;
        RECT 2242.660 17.270 2245.100 17.410 ;
        RECT 2244.960 2.400 2245.100 17.270 ;
        RECT 2244.750 -4.800 2245.310 2.400 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1380.070 1684.260 1380.390 1684.320 ;
        RECT 1382.370 1684.260 1382.690 1684.320 ;
        RECT 1380.070 1684.120 1382.690 1684.260 ;
        RECT 1380.070 1684.060 1380.390 1684.120 ;
        RECT 1382.370 1684.060 1382.690 1684.120 ;
        RECT 1380.070 1445.920 1380.390 1445.980 ;
        RECT 2256.830 1445.920 2257.150 1445.980 ;
        RECT 1380.070 1445.780 2257.150 1445.920 ;
        RECT 1380.070 1445.720 1380.390 1445.780 ;
        RECT 2256.830 1445.720 2257.150 1445.780 ;
      LAYER via ;
        RECT 1380.100 1684.060 1380.360 1684.320 ;
        RECT 1382.400 1684.060 1382.660 1684.320 ;
        RECT 1380.100 1445.720 1380.360 1445.980 ;
        RECT 2256.860 1445.720 2257.120 1445.980 ;
      LAYER met2 ;
        RECT 1382.300 1700.340 1382.580 1704.000 ;
        RECT 1382.300 1700.000 1382.600 1700.340 ;
        RECT 1382.460 1684.350 1382.600 1700.000 ;
        RECT 1380.100 1684.030 1380.360 1684.350 ;
        RECT 1382.400 1684.030 1382.660 1684.350 ;
        RECT 1380.160 1446.010 1380.300 1684.030 ;
        RECT 1380.100 1445.690 1380.360 1446.010 ;
        RECT 2256.860 1445.690 2257.120 1446.010 ;
        RECT 2256.920 17.410 2257.060 1445.690 ;
        RECT 2256.920 17.270 2262.580 17.410 ;
        RECT 2262.440 2.400 2262.580 17.270 ;
        RECT 2262.230 -4.800 2262.790 2.400 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1384.210 1501.000 1384.530 1501.060 ;
        RECT 2277.070 1501.000 2277.390 1501.060 ;
        RECT 1384.210 1500.860 2277.390 1501.000 ;
        RECT 1384.210 1500.800 1384.530 1500.860 ;
        RECT 2277.070 1500.800 2277.390 1500.860 ;
      LAYER via ;
        RECT 1384.240 1500.800 1384.500 1501.060 ;
        RECT 2277.100 1500.800 2277.360 1501.060 ;
      LAYER met2 ;
        RECT 1384.140 1700.340 1384.420 1704.000 ;
        RECT 1384.140 1700.000 1384.440 1700.340 ;
        RECT 1384.300 1501.090 1384.440 1700.000 ;
        RECT 1384.240 1500.770 1384.500 1501.090 ;
        RECT 2277.100 1500.770 2277.360 1501.090 ;
        RECT 2277.160 17.410 2277.300 1500.770 ;
        RECT 2277.160 17.270 2280.520 17.410 ;
        RECT 2280.380 2.400 2280.520 17.270 ;
        RECT 2280.170 -4.800 2280.730 2.400 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1384.670 1683.920 1384.990 1683.980 ;
        RECT 1386.050 1683.920 1386.370 1683.980 ;
        RECT 1384.670 1683.780 1386.370 1683.920 ;
        RECT 1384.670 1683.720 1384.990 1683.780 ;
        RECT 1386.050 1683.720 1386.370 1683.780 ;
        RECT 1381.450 1631.900 1381.770 1631.960 ;
        RECT 1384.670 1631.900 1384.990 1631.960 ;
        RECT 1381.450 1631.760 1384.990 1631.900 ;
        RECT 1381.450 1631.700 1381.770 1631.760 ;
        RECT 1384.670 1631.700 1384.990 1631.760 ;
        RECT 1381.450 1438.780 1381.770 1438.840 ;
        RECT 2298.230 1438.780 2298.550 1438.840 ;
        RECT 1381.450 1438.640 2298.550 1438.780 ;
        RECT 1381.450 1438.580 1381.770 1438.640 ;
        RECT 2298.230 1438.580 2298.550 1438.640 ;
      LAYER via ;
        RECT 1384.700 1683.720 1384.960 1683.980 ;
        RECT 1386.080 1683.720 1386.340 1683.980 ;
        RECT 1381.480 1631.700 1381.740 1631.960 ;
        RECT 1384.700 1631.700 1384.960 1631.960 ;
        RECT 1381.480 1438.580 1381.740 1438.840 ;
        RECT 2298.260 1438.580 2298.520 1438.840 ;
      LAYER met2 ;
        RECT 1385.980 1700.340 1386.260 1704.000 ;
        RECT 1385.980 1700.000 1386.280 1700.340 ;
        RECT 1386.140 1684.010 1386.280 1700.000 ;
        RECT 1384.700 1683.690 1384.960 1684.010 ;
        RECT 1386.080 1683.690 1386.340 1684.010 ;
        RECT 1384.760 1631.990 1384.900 1683.690 ;
        RECT 1381.480 1631.670 1381.740 1631.990 ;
        RECT 1384.700 1631.670 1384.960 1631.990 ;
        RECT 1381.540 1438.870 1381.680 1631.670 ;
        RECT 1381.480 1438.550 1381.740 1438.870 ;
        RECT 2298.260 1438.550 2298.520 1438.870 ;
        RECT 2298.320 2.400 2298.460 1438.550 ;
        RECT 2298.110 -4.800 2298.670 2.400 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1386.970 1639.380 1387.290 1639.440 ;
        RECT 2311.570 1639.380 2311.890 1639.440 ;
        RECT 1386.970 1639.240 2311.890 1639.380 ;
        RECT 1386.970 1639.180 1387.290 1639.240 ;
        RECT 2311.570 1639.180 2311.890 1639.240 ;
      LAYER via ;
        RECT 1387.000 1639.180 1387.260 1639.440 ;
        RECT 2311.600 1639.180 2311.860 1639.440 ;
      LAYER met2 ;
        RECT 1387.820 1700.340 1388.100 1704.000 ;
        RECT 1387.820 1700.000 1388.120 1700.340 ;
        RECT 1387.980 1688.850 1388.120 1700.000 ;
        RECT 1387.060 1688.710 1388.120 1688.850 ;
        RECT 1387.060 1639.470 1387.200 1688.710 ;
        RECT 1387.000 1639.150 1387.260 1639.470 ;
        RECT 2311.600 1639.150 2311.860 1639.470 ;
        RECT 2311.660 17.410 2311.800 1639.150 ;
        RECT 2311.660 17.270 2316.400 17.410 ;
        RECT 2316.260 2.400 2316.400 17.270 ;
        RECT 2316.050 -4.800 2316.610 2.400 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1389.730 1683.920 1390.050 1683.980 ;
        RECT 1391.110 1683.920 1391.430 1683.980 ;
        RECT 1389.730 1683.780 1391.430 1683.920 ;
        RECT 1389.730 1683.720 1390.050 1683.780 ;
        RECT 1391.110 1683.720 1391.430 1683.780 ;
        RECT 1391.110 1605.040 1391.430 1605.100 ;
        RECT 2332.270 1605.040 2332.590 1605.100 ;
        RECT 1391.110 1604.900 2332.590 1605.040 ;
        RECT 1391.110 1604.840 1391.430 1604.900 ;
        RECT 2332.270 1604.840 2332.590 1604.900 ;
      LAYER via ;
        RECT 1389.760 1683.720 1390.020 1683.980 ;
        RECT 1391.140 1683.720 1391.400 1683.980 ;
        RECT 1391.140 1604.840 1391.400 1605.100 ;
        RECT 2332.300 1604.840 2332.560 1605.100 ;
      LAYER met2 ;
        RECT 1389.660 1700.340 1389.940 1704.000 ;
        RECT 1389.660 1700.000 1389.960 1700.340 ;
        RECT 1389.820 1684.010 1389.960 1700.000 ;
        RECT 1389.760 1683.690 1390.020 1684.010 ;
        RECT 1391.140 1683.690 1391.400 1684.010 ;
        RECT 1391.200 1605.130 1391.340 1683.690 ;
        RECT 1391.140 1604.810 1391.400 1605.130 ;
        RECT 2332.300 1604.810 2332.560 1605.130 ;
        RECT 2332.360 17.410 2332.500 1604.810 ;
        RECT 2332.360 17.270 2334.340 17.410 ;
        RECT 2334.200 2.400 2334.340 17.270 ;
        RECT 2333.990 -4.800 2334.550 2.400 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1388.810 1686.980 1389.130 1687.040 ;
        RECT 1391.570 1686.980 1391.890 1687.040 ;
        RECT 1388.810 1686.840 1391.890 1686.980 ;
        RECT 1388.810 1686.780 1389.130 1686.840 ;
        RECT 1391.570 1686.780 1391.890 1686.840 ;
        RECT 1387.890 1683.920 1388.210 1683.980 ;
        RECT 1388.810 1683.920 1389.130 1683.980 ;
        RECT 1387.890 1683.780 1389.130 1683.920 ;
        RECT 1387.890 1683.720 1388.210 1683.780 ;
        RECT 1388.810 1683.720 1389.130 1683.780 ;
        RECT 1387.890 1493.860 1388.210 1493.920 ;
        RECT 2346.070 1493.860 2346.390 1493.920 ;
        RECT 1387.890 1493.720 2346.390 1493.860 ;
        RECT 1387.890 1493.660 1388.210 1493.720 ;
        RECT 2346.070 1493.660 2346.390 1493.720 ;
      LAYER via ;
        RECT 1388.840 1686.780 1389.100 1687.040 ;
        RECT 1391.600 1686.780 1391.860 1687.040 ;
        RECT 1387.920 1683.720 1388.180 1683.980 ;
        RECT 1388.840 1683.720 1389.100 1683.980 ;
        RECT 1387.920 1493.660 1388.180 1493.920 ;
        RECT 2346.100 1493.660 2346.360 1493.920 ;
      LAYER met2 ;
        RECT 1391.500 1700.340 1391.780 1704.000 ;
        RECT 1391.500 1700.000 1391.800 1700.340 ;
        RECT 1391.660 1687.070 1391.800 1700.000 ;
        RECT 1388.840 1686.750 1389.100 1687.070 ;
        RECT 1391.600 1686.750 1391.860 1687.070 ;
        RECT 1388.900 1684.010 1389.040 1686.750 ;
        RECT 1387.920 1683.690 1388.180 1684.010 ;
        RECT 1388.840 1683.690 1389.100 1684.010 ;
        RECT 1387.980 1493.950 1388.120 1683.690 ;
        RECT 1387.920 1493.630 1388.180 1493.950 ;
        RECT 2346.100 1493.630 2346.360 1493.950 ;
        RECT 2346.160 17.410 2346.300 1493.630 ;
        RECT 2346.160 17.270 2351.820 17.410 ;
        RECT 2351.680 2.400 2351.820 17.270 ;
        RECT 2351.470 -4.800 2352.030 2.400 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1387.430 1688.000 1387.750 1688.060 ;
        RECT 1393.410 1688.000 1393.730 1688.060 ;
        RECT 1387.430 1687.860 1393.730 1688.000 ;
        RECT 1387.430 1687.800 1387.750 1687.860 ;
        RECT 1393.410 1687.800 1393.730 1687.860 ;
        RECT 1387.430 1535.680 1387.750 1535.740 ;
        RECT 2366.770 1535.680 2367.090 1535.740 ;
        RECT 1387.430 1535.540 2367.090 1535.680 ;
        RECT 1387.430 1535.480 1387.750 1535.540 ;
        RECT 2366.770 1535.480 2367.090 1535.540 ;
      LAYER via ;
        RECT 1387.460 1687.800 1387.720 1688.060 ;
        RECT 1393.440 1687.800 1393.700 1688.060 ;
        RECT 1387.460 1535.480 1387.720 1535.740 ;
        RECT 2366.800 1535.480 2367.060 1535.740 ;
      LAYER met2 ;
        RECT 1393.340 1700.340 1393.620 1704.000 ;
        RECT 1393.340 1700.000 1393.640 1700.340 ;
        RECT 1393.500 1688.090 1393.640 1700.000 ;
        RECT 1387.460 1687.770 1387.720 1688.090 ;
        RECT 1393.440 1687.770 1393.700 1688.090 ;
        RECT 1387.520 1535.770 1387.660 1687.770 ;
        RECT 1387.460 1535.450 1387.720 1535.770 ;
        RECT 2366.800 1535.450 2367.060 1535.770 ;
        RECT 2366.860 16.730 2367.000 1535.450 ;
        RECT 2366.860 16.590 2369.760 16.730 ;
        RECT 2369.620 2.400 2369.760 16.590 ;
        RECT 2369.410 -4.800 2369.970 2.400 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1395.250 1684.940 1395.570 1685.000 ;
        RECT 1398.470 1684.940 1398.790 1685.000 ;
        RECT 1395.250 1684.800 1398.790 1684.940 ;
        RECT 1395.250 1684.740 1395.570 1684.800 ;
        RECT 1398.470 1684.740 1398.790 1684.800 ;
        RECT 1398.010 1431.640 1398.330 1431.700 ;
        RECT 2387.470 1431.640 2387.790 1431.700 ;
        RECT 1398.010 1431.500 2387.790 1431.640 ;
        RECT 1398.010 1431.440 1398.330 1431.500 ;
        RECT 2387.470 1431.440 2387.790 1431.500 ;
      LAYER via ;
        RECT 1395.280 1684.740 1395.540 1685.000 ;
        RECT 1398.500 1684.740 1398.760 1685.000 ;
        RECT 1398.040 1431.440 1398.300 1431.700 ;
        RECT 2387.500 1431.440 2387.760 1431.700 ;
      LAYER met2 ;
        RECT 1395.180 1700.340 1395.460 1704.000 ;
        RECT 1395.180 1700.000 1395.480 1700.340 ;
        RECT 1395.340 1685.030 1395.480 1700.000 ;
        RECT 1395.280 1684.710 1395.540 1685.030 ;
        RECT 1398.500 1684.710 1398.760 1685.030 ;
        RECT 1398.560 1631.730 1398.700 1684.710 ;
        RECT 1398.100 1631.590 1398.700 1631.730 ;
        RECT 1398.100 1431.730 1398.240 1631.590 ;
        RECT 1398.040 1431.410 1398.300 1431.730 ;
        RECT 2387.500 1431.410 2387.760 1431.730 ;
        RECT 2387.560 2.400 2387.700 1431.410 ;
        RECT 2387.350 -4.800 2387.910 2.400 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1398.010 1632.240 1398.330 1632.300 ;
        RECT 1398.010 1632.100 1398.700 1632.240 ;
        RECT 1398.010 1632.040 1398.330 1632.100 ;
        RECT 1398.560 1631.280 1398.700 1632.100 ;
        RECT 1398.470 1631.020 1398.790 1631.280 ;
        RECT 1398.470 1424.840 1398.790 1424.900 ;
        RECT 2401.270 1424.840 2401.590 1424.900 ;
        RECT 1398.470 1424.700 2401.590 1424.840 ;
        RECT 1398.470 1424.640 1398.790 1424.700 ;
        RECT 2401.270 1424.640 2401.590 1424.700 ;
      LAYER via ;
        RECT 1398.040 1632.040 1398.300 1632.300 ;
        RECT 1398.500 1631.020 1398.760 1631.280 ;
        RECT 1398.500 1424.640 1398.760 1424.900 ;
        RECT 2401.300 1424.640 2401.560 1424.900 ;
      LAYER met2 ;
        RECT 1397.020 1700.340 1397.300 1704.000 ;
        RECT 1397.020 1700.000 1397.320 1700.340 ;
        RECT 1397.180 1677.970 1397.320 1700.000 ;
        RECT 1397.180 1677.830 1398.240 1677.970 ;
        RECT 1398.100 1632.330 1398.240 1677.830 ;
        RECT 1398.040 1632.010 1398.300 1632.330 ;
        RECT 1398.500 1630.990 1398.760 1631.310 ;
        RECT 1398.560 1424.930 1398.700 1630.990 ;
        RECT 1398.500 1424.610 1398.760 1424.930 ;
        RECT 2401.300 1424.610 2401.560 1424.930 ;
        RECT 2401.360 17.410 2401.500 1424.610 ;
        RECT 2401.360 17.270 2405.640 17.410 ;
        RECT 2405.500 2.400 2405.640 17.270 ;
        RECT 2405.290 -4.800 2405.850 2.400 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1229.650 1677.460 1229.970 1677.520 ;
        RECT 1231.030 1677.460 1231.350 1677.520 ;
        RECT 1229.650 1677.320 1231.350 1677.460 ;
        RECT 1229.650 1677.260 1229.970 1677.320 ;
        RECT 1231.030 1677.260 1231.350 1677.320 ;
        RECT 799.550 1618.640 799.870 1618.700 ;
        RECT 1229.650 1618.640 1229.970 1618.700 ;
        RECT 799.550 1618.500 1229.970 1618.640 ;
        RECT 799.550 1618.440 799.870 1618.500 ;
        RECT 1229.650 1618.440 1229.970 1618.500 ;
      LAYER via ;
        RECT 1229.680 1677.260 1229.940 1677.520 ;
        RECT 1231.060 1677.260 1231.320 1677.520 ;
        RECT 799.580 1618.440 799.840 1618.700 ;
        RECT 1229.680 1618.440 1229.940 1618.700 ;
      LAYER met2 ;
        RECT 1231.880 1700.410 1232.160 1704.000 ;
        RECT 1231.580 1700.270 1232.160 1700.410 ;
        RECT 1231.580 1678.650 1231.720 1700.270 ;
        RECT 1231.880 1700.000 1232.160 1700.270 ;
        RECT 1231.120 1678.510 1231.720 1678.650 ;
        RECT 1231.120 1677.550 1231.260 1678.510 ;
        RECT 1229.680 1677.230 1229.940 1677.550 ;
        RECT 1231.060 1677.230 1231.320 1677.550 ;
        RECT 1229.740 1618.730 1229.880 1677.230 ;
        RECT 799.580 1618.410 799.840 1618.730 ;
        RECT 1229.680 1618.410 1229.940 1618.730 ;
        RECT 799.640 2.400 799.780 1618.410 ;
        RECT 799.430 -4.800 799.990 2.400 ;
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 648.210 1666.920 648.530 1666.980 ;
        RECT 1215.850 1666.920 1216.170 1666.980 ;
        RECT 648.210 1666.780 1216.170 1666.920 ;
        RECT 648.210 1666.720 648.530 1666.780 ;
        RECT 1215.850 1666.720 1216.170 1666.780 ;
      LAYER via ;
        RECT 648.240 1666.720 648.500 1666.980 ;
        RECT 1215.880 1666.720 1216.140 1666.980 ;
      LAYER met2 ;
        RECT 1215.780 1700.340 1216.060 1704.000 ;
        RECT 1215.780 1700.000 1216.080 1700.340 ;
        RECT 1215.940 1667.010 1216.080 1700.000 ;
        RECT 648.240 1666.690 648.500 1667.010 ;
        RECT 1215.880 1666.690 1216.140 1667.010 ;
        RECT 648.300 17.410 648.440 1666.690 ;
        RECT 645.080 17.270 648.440 17.410 ;
        RECT 645.080 2.400 645.220 17.270 ;
        RECT 644.870 -4.800 645.430 2.400 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1396.170 1685.620 1396.490 1685.680 ;
        RECT 1399.390 1685.620 1399.710 1685.680 ;
        RECT 1396.170 1685.480 1399.710 1685.620 ;
        RECT 1396.170 1685.420 1396.490 1685.480 ;
        RECT 1399.390 1685.420 1399.710 1685.480 ;
        RECT 1394.330 1676.100 1394.650 1676.160 ;
        RECT 1396.630 1676.100 1396.950 1676.160 ;
        RECT 1394.330 1675.960 1396.950 1676.100 ;
        RECT 1394.330 1675.900 1394.650 1675.960 ;
        RECT 1396.630 1675.900 1396.950 1675.960 ;
        RECT 1394.330 1418.040 1394.650 1418.100 ;
        RECT 2428.870 1418.040 2429.190 1418.100 ;
        RECT 1394.330 1417.900 2429.190 1418.040 ;
        RECT 1394.330 1417.840 1394.650 1417.900 ;
        RECT 2428.870 1417.840 2429.190 1417.900 ;
      LAYER via ;
        RECT 1396.200 1685.420 1396.460 1685.680 ;
        RECT 1399.420 1685.420 1399.680 1685.680 ;
        RECT 1394.360 1675.900 1394.620 1676.160 ;
        RECT 1396.660 1675.900 1396.920 1676.160 ;
        RECT 1394.360 1417.840 1394.620 1418.100 ;
        RECT 2428.900 1417.840 2429.160 1418.100 ;
      LAYER met2 ;
        RECT 1399.320 1700.340 1399.600 1704.000 ;
        RECT 1399.320 1700.000 1399.620 1700.340 ;
        RECT 1399.480 1685.710 1399.620 1700.000 ;
        RECT 1396.200 1685.390 1396.460 1685.710 ;
        RECT 1399.420 1685.390 1399.680 1685.710 ;
        RECT 1396.260 1678.650 1396.400 1685.390 ;
        RECT 1396.260 1678.510 1396.860 1678.650 ;
        RECT 1396.720 1676.190 1396.860 1678.510 ;
        RECT 1394.360 1675.870 1394.620 1676.190 ;
        RECT 1396.660 1675.870 1396.920 1676.190 ;
        RECT 1394.420 1418.130 1394.560 1675.870 ;
        RECT 1394.360 1417.810 1394.620 1418.130 ;
        RECT 2428.900 1417.810 2429.160 1418.130 ;
        RECT 2428.960 2.400 2429.100 1417.810 ;
        RECT 2428.750 -4.800 2429.310 2.400 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1401.230 1410.900 1401.550 1410.960 ;
        RECT 2442.670 1410.900 2442.990 1410.960 ;
        RECT 1401.230 1410.760 2442.990 1410.900 ;
        RECT 1401.230 1410.700 1401.550 1410.760 ;
        RECT 2442.670 1410.700 2442.990 1410.760 ;
      LAYER via ;
        RECT 1401.260 1410.700 1401.520 1410.960 ;
        RECT 2442.700 1410.700 2442.960 1410.960 ;
      LAYER met2 ;
        RECT 1401.160 1700.340 1401.440 1704.000 ;
        RECT 1401.160 1700.000 1401.460 1700.340 ;
        RECT 1401.320 1410.990 1401.460 1700.000 ;
        RECT 1401.260 1410.670 1401.520 1410.990 ;
        RECT 2442.700 1410.670 2442.960 1410.990 ;
        RECT 2442.760 18.090 2442.900 1410.670 ;
        RECT 2442.760 17.950 2447.040 18.090 ;
        RECT 2446.900 2.400 2447.040 17.950 ;
        RECT 2446.690 -4.800 2447.250 2.400 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1403.070 1684.600 1403.390 1684.660 ;
        RECT 1405.830 1684.600 1406.150 1684.660 ;
        RECT 1403.070 1684.460 1406.150 1684.600 ;
        RECT 1403.070 1684.400 1403.390 1684.460 ;
        RECT 1405.830 1684.400 1406.150 1684.460 ;
        RECT 1406.290 1404.100 1406.610 1404.160 ;
        RECT 2463.370 1404.100 2463.690 1404.160 ;
        RECT 1406.290 1403.960 2463.690 1404.100 ;
        RECT 1406.290 1403.900 1406.610 1403.960 ;
        RECT 2463.370 1403.900 2463.690 1403.960 ;
        RECT 2463.370 2.960 2463.690 3.020 ;
        RECT 2464.750 2.960 2465.070 3.020 ;
        RECT 2463.370 2.820 2465.070 2.960 ;
        RECT 2463.370 2.760 2463.690 2.820 ;
        RECT 2464.750 2.760 2465.070 2.820 ;
      LAYER via ;
        RECT 1403.100 1684.400 1403.360 1684.660 ;
        RECT 1405.860 1684.400 1406.120 1684.660 ;
        RECT 1406.320 1403.900 1406.580 1404.160 ;
        RECT 2463.400 1403.900 2463.660 1404.160 ;
        RECT 2463.400 2.760 2463.660 3.020 ;
        RECT 2464.780 2.760 2465.040 3.020 ;
      LAYER met2 ;
        RECT 1403.000 1700.340 1403.280 1704.000 ;
        RECT 1403.000 1700.000 1403.300 1700.340 ;
        RECT 1403.160 1684.690 1403.300 1700.000 ;
        RECT 1403.100 1684.370 1403.360 1684.690 ;
        RECT 1405.860 1684.370 1406.120 1684.690 ;
        RECT 1405.920 1631.050 1406.060 1684.370 ;
        RECT 1405.920 1630.910 1406.520 1631.050 ;
        RECT 1406.380 1404.190 1406.520 1630.910 ;
        RECT 1406.320 1403.870 1406.580 1404.190 ;
        RECT 2463.400 1403.870 2463.660 1404.190 ;
        RECT 2463.460 3.050 2463.600 1403.870 ;
        RECT 2463.400 2.730 2463.660 3.050 ;
        RECT 2464.780 2.730 2465.040 3.050 ;
        RECT 2464.840 2.400 2464.980 2.730 ;
        RECT 2464.630 -4.800 2465.190 2.400 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1404.910 1683.920 1405.230 1683.980 ;
        RECT 1407.210 1683.920 1407.530 1683.980 ;
        RECT 1404.910 1683.780 1407.530 1683.920 ;
        RECT 1404.910 1683.720 1405.230 1683.780 ;
        RECT 1407.210 1683.720 1407.530 1683.780 ;
        RECT 1407.210 672.760 1407.530 672.820 ;
        RECT 2477.170 672.760 2477.490 672.820 ;
        RECT 1407.210 672.620 2477.490 672.760 ;
        RECT 1407.210 672.560 1407.530 672.620 ;
        RECT 2477.170 672.560 2477.490 672.620 ;
        RECT 2477.170 2.960 2477.490 3.020 ;
        RECT 2482.690 2.960 2483.010 3.020 ;
        RECT 2477.170 2.820 2483.010 2.960 ;
        RECT 2477.170 2.760 2477.490 2.820 ;
        RECT 2482.690 2.760 2483.010 2.820 ;
      LAYER via ;
        RECT 1404.940 1683.720 1405.200 1683.980 ;
        RECT 1407.240 1683.720 1407.500 1683.980 ;
        RECT 1407.240 672.560 1407.500 672.820 ;
        RECT 2477.200 672.560 2477.460 672.820 ;
        RECT 2477.200 2.760 2477.460 3.020 ;
        RECT 2482.720 2.760 2482.980 3.020 ;
      LAYER met2 ;
        RECT 1404.840 1700.340 1405.120 1704.000 ;
        RECT 1404.840 1700.000 1405.140 1700.340 ;
        RECT 1405.000 1684.010 1405.140 1700.000 ;
        RECT 1404.940 1683.690 1405.200 1684.010 ;
        RECT 1407.240 1683.690 1407.500 1684.010 ;
        RECT 1407.300 672.850 1407.440 1683.690 ;
        RECT 1407.240 672.530 1407.500 672.850 ;
        RECT 2477.200 672.530 2477.460 672.850 ;
        RECT 2477.260 3.050 2477.400 672.530 ;
        RECT 2477.200 2.730 2477.460 3.050 ;
        RECT 2482.720 2.730 2482.980 3.050 ;
        RECT 2482.780 2.400 2482.920 2.730 ;
        RECT 2482.570 -4.800 2483.130 2.400 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1406.750 1397.300 1407.070 1397.360 ;
        RECT 2497.870 1397.300 2498.190 1397.360 ;
        RECT 1406.750 1397.160 2498.190 1397.300 ;
        RECT 1406.750 1397.100 1407.070 1397.160 ;
        RECT 2497.870 1397.100 2498.190 1397.160 ;
      LAYER via ;
        RECT 1406.780 1397.100 1407.040 1397.360 ;
        RECT 2497.900 1397.100 2498.160 1397.360 ;
      LAYER met2 ;
        RECT 1406.680 1700.340 1406.960 1704.000 ;
        RECT 1406.680 1700.000 1406.980 1700.340 ;
        RECT 1406.840 1397.390 1406.980 1700.000 ;
        RECT 1406.780 1397.070 1407.040 1397.390 ;
        RECT 2497.900 1397.070 2498.160 1397.390 ;
        RECT 2497.960 17.410 2498.100 1397.070 ;
        RECT 2497.960 17.270 2500.860 17.410 ;
        RECT 2500.720 2.400 2500.860 17.270 ;
        RECT 2500.510 -4.800 2501.070 2.400 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1408.130 1675.420 1408.450 1675.480 ;
        RECT 1412.730 1675.420 1413.050 1675.480 ;
        RECT 1408.130 1675.280 1413.050 1675.420 ;
        RECT 1408.130 1675.220 1408.450 1675.280 ;
        RECT 1412.730 1675.220 1413.050 1675.280 ;
        RECT 1412.730 1487.400 1413.050 1487.460 ;
        RECT 2512.130 1487.400 2512.450 1487.460 ;
        RECT 1412.730 1487.260 2512.450 1487.400 ;
        RECT 1412.730 1487.200 1413.050 1487.260 ;
        RECT 2512.130 1487.200 2512.450 1487.260 ;
        RECT 2512.130 18.260 2512.450 18.320 ;
        RECT 2518.110 18.260 2518.430 18.320 ;
        RECT 2512.130 18.120 2518.430 18.260 ;
        RECT 2512.130 18.060 2512.450 18.120 ;
        RECT 2518.110 18.060 2518.430 18.120 ;
      LAYER via ;
        RECT 1408.160 1675.220 1408.420 1675.480 ;
        RECT 1412.760 1675.220 1413.020 1675.480 ;
        RECT 1412.760 1487.200 1413.020 1487.460 ;
        RECT 2512.160 1487.200 2512.420 1487.460 ;
        RECT 2512.160 18.060 2512.420 18.320 ;
        RECT 2518.140 18.060 2518.400 18.320 ;
      LAYER met2 ;
        RECT 1408.520 1700.340 1408.800 1704.000 ;
        RECT 1408.520 1700.000 1408.820 1700.340 ;
        RECT 1408.680 1678.650 1408.820 1700.000 ;
        RECT 1408.220 1678.510 1408.820 1678.650 ;
        RECT 1408.220 1675.510 1408.360 1678.510 ;
        RECT 1408.160 1675.190 1408.420 1675.510 ;
        RECT 1412.760 1675.190 1413.020 1675.510 ;
        RECT 1412.820 1487.490 1412.960 1675.190 ;
        RECT 1412.760 1487.170 1413.020 1487.490 ;
        RECT 2512.160 1487.170 2512.420 1487.490 ;
        RECT 2512.220 18.350 2512.360 1487.170 ;
        RECT 2512.160 18.030 2512.420 18.350 ;
        RECT 2518.140 18.030 2518.400 18.350 ;
        RECT 2518.200 2.400 2518.340 18.030 ;
        RECT 2517.990 -4.800 2518.550 2.400 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1410.430 1683.920 1410.750 1683.980 ;
        RECT 1413.190 1683.920 1413.510 1683.980 ;
        RECT 1410.430 1683.780 1413.510 1683.920 ;
        RECT 1410.430 1683.720 1410.750 1683.780 ;
        RECT 1413.190 1683.720 1413.510 1683.780 ;
        RECT 1413.190 1459.180 1413.510 1459.240 ;
        RECT 2532.370 1459.180 2532.690 1459.240 ;
        RECT 1413.190 1459.040 2532.690 1459.180 ;
        RECT 1413.190 1458.980 1413.510 1459.040 ;
        RECT 2532.370 1458.980 2532.690 1459.040 ;
      LAYER via ;
        RECT 1410.460 1683.720 1410.720 1683.980 ;
        RECT 1413.220 1683.720 1413.480 1683.980 ;
        RECT 1413.220 1458.980 1413.480 1459.240 ;
        RECT 2532.400 1458.980 2532.660 1459.240 ;
      LAYER met2 ;
        RECT 1410.360 1700.340 1410.640 1704.000 ;
        RECT 1410.360 1700.000 1410.660 1700.340 ;
        RECT 1410.520 1684.010 1410.660 1700.000 ;
        RECT 1410.460 1683.690 1410.720 1684.010 ;
        RECT 1413.220 1683.690 1413.480 1684.010 ;
        RECT 1413.280 1459.270 1413.420 1683.690 ;
        RECT 1413.220 1458.950 1413.480 1459.270 ;
        RECT 2532.400 1458.950 2532.660 1459.270 ;
        RECT 2532.460 17.410 2532.600 1458.950 ;
        RECT 2532.460 17.270 2536.280 17.410 ;
        RECT 2536.140 2.400 2536.280 17.270 ;
        RECT 2535.930 -4.800 2536.490 2.400 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1409.510 1390.160 1409.830 1390.220 ;
        RECT 2553.070 1390.160 2553.390 1390.220 ;
        RECT 1409.510 1390.020 2553.390 1390.160 ;
        RECT 1409.510 1389.960 1409.830 1390.020 ;
        RECT 2553.070 1389.960 2553.390 1390.020 ;
      LAYER via ;
        RECT 1409.540 1389.960 1409.800 1390.220 ;
        RECT 2553.100 1389.960 2553.360 1390.220 ;
      LAYER met2 ;
        RECT 1412.200 1700.340 1412.480 1704.000 ;
        RECT 1412.200 1700.000 1412.500 1700.340 ;
        RECT 1412.360 1676.610 1412.500 1700.000 ;
        RECT 1409.600 1676.470 1412.500 1676.610 ;
        RECT 1409.600 1390.250 1409.740 1676.470 ;
        RECT 1409.540 1389.930 1409.800 1390.250 ;
        RECT 2553.100 1389.930 2553.360 1390.250 ;
        RECT 2553.160 17.410 2553.300 1389.930 ;
        RECT 2553.160 17.270 2554.220 17.410 ;
        RECT 2554.080 2.400 2554.220 17.270 ;
        RECT 2553.870 -4.800 2554.430 2.400 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1412.730 1685.960 1413.050 1686.020 ;
        RECT 1414.110 1685.960 1414.430 1686.020 ;
        RECT 1412.730 1685.820 1414.430 1685.960 ;
        RECT 1412.730 1685.760 1413.050 1685.820 ;
        RECT 1414.110 1685.760 1414.430 1685.820 ;
        RECT 1410.430 1383.360 1410.750 1383.420 ;
        RECT 2566.870 1383.360 2567.190 1383.420 ;
        RECT 1410.430 1383.220 2567.190 1383.360 ;
        RECT 1410.430 1383.160 1410.750 1383.220 ;
        RECT 2566.870 1383.160 2567.190 1383.220 ;
      LAYER via ;
        RECT 1412.760 1685.760 1413.020 1686.020 ;
        RECT 1414.140 1685.760 1414.400 1686.020 ;
        RECT 1410.460 1383.160 1410.720 1383.420 ;
        RECT 2566.900 1383.160 2567.160 1383.420 ;
      LAYER met2 ;
        RECT 1414.040 1700.340 1414.320 1704.000 ;
        RECT 1414.040 1700.000 1414.340 1700.340 ;
        RECT 1414.200 1686.050 1414.340 1700.000 ;
        RECT 1412.760 1685.730 1413.020 1686.050 ;
        RECT 1414.140 1685.730 1414.400 1686.050 ;
        RECT 1412.820 1675.930 1412.960 1685.730 ;
        RECT 1410.520 1675.790 1412.960 1675.930 ;
        RECT 1410.520 1383.450 1410.660 1675.790 ;
        RECT 1410.460 1383.130 1410.720 1383.450 ;
        RECT 2566.900 1383.130 2567.160 1383.450 ;
        RECT 2566.960 17.410 2567.100 1383.130 ;
        RECT 2566.960 17.270 2572.160 17.410 ;
        RECT 2572.020 2.400 2572.160 17.270 ;
        RECT 2571.810 -4.800 2572.370 2.400 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1415.950 1684.940 1416.270 1685.000 ;
        RECT 1420.550 1684.940 1420.870 1685.000 ;
        RECT 1415.950 1684.800 1420.870 1684.940 ;
        RECT 1415.950 1684.740 1416.270 1684.800 ;
        RECT 1420.550 1684.740 1420.870 1684.800 ;
        RECT 1420.550 1369.760 1420.870 1369.820 ;
        RECT 2587.570 1369.760 2587.890 1369.820 ;
        RECT 1420.550 1369.620 2587.890 1369.760 ;
        RECT 1420.550 1369.560 1420.870 1369.620 ;
        RECT 2587.570 1369.560 2587.890 1369.620 ;
      LAYER via ;
        RECT 1415.980 1684.740 1416.240 1685.000 ;
        RECT 1420.580 1684.740 1420.840 1685.000 ;
        RECT 1420.580 1369.560 1420.840 1369.820 ;
        RECT 2587.600 1369.560 2587.860 1369.820 ;
      LAYER met2 ;
        RECT 1415.880 1700.340 1416.160 1704.000 ;
        RECT 1415.880 1700.000 1416.180 1700.340 ;
        RECT 1416.040 1685.030 1416.180 1700.000 ;
        RECT 1415.980 1684.710 1416.240 1685.030 ;
        RECT 1420.580 1684.710 1420.840 1685.030 ;
        RECT 1420.640 1369.850 1420.780 1684.710 ;
        RECT 1420.580 1369.530 1420.840 1369.850 ;
        RECT 2587.600 1369.530 2587.860 1369.850 ;
        RECT 2587.660 17.410 2587.800 1369.530 ;
        RECT 2587.660 17.270 2589.640 17.410 ;
        RECT 2589.500 2.400 2589.640 17.270 ;
        RECT 2589.290 -4.800 2589.850 2.400 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 827.610 1654.000 827.930 1654.060 ;
        RECT 1234.250 1654.000 1234.570 1654.060 ;
        RECT 827.610 1653.860 1234.570 1654.000 ;
        RECT 827.610 1653.800 827.930 1653.860 ;
        RECT 1234.250 1653.800 1234.570 1653.860 ;
      LAYER via ;
        RECT 827.640 1653.800 827.900 1654.060 ;
        RECT 1234.280 1653.800 1234.540 1654.060 ;
      LAYER met2 ;
        RECT 1234.180 1700.340 1234.460 1704.000 ;
        RECT 1234.180 1700.000 1234.480 1700.340 ;
        RECT 1234.340 1654.090 1234.480 1700.000 ;
        RECT 827.640 1653.770 827.900 1654.090 ;
        RECT 1234.280 1653.770 1234.540 1654.090 ;
        RECT 827.700 17.410 827.840 1653.770 ;
        RECT 823.560 17.270 827.840 17.410 ;
        RECT 823.560 2.400 823.700 17.270 ;
        RECT 823.350 -4.800 823.910 2.400 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1418.325 1642.625 1418.495 1689.715 ;
        RECT 1418.785 1497.785 1418.955 1587.035 ;
        RECT 1418.785 1442.025 1418.955 1490.475 ;
      LAYER mcon ;
        RECT 1418.325 1689.545 1418.495 1689.715 ;
        RECT 1418.785 1586.865 1418.955 1587.035 ;
        RECT 1418.785 1490.305 1418.955 1490.475 ;
      LAYER met1 ;
        RECT 1417.790 1689.700 1418.110 1689.760 ;
        RECT 1418.265 1689.700 1418.555 1689.745 ;
        RECT 1417.790 1689.560 1418.555 1689.700 ;
        RECT 1417.790 1689.500 1418.110 1689.560 ;
        RECT 1418.265 1689.515 1418.555 1689.560 ;
        RECT 1418.250 1642.780 1418.570 1642.840 ;
        RECT 1418.055 1642.640 1418.570 1642.780 ;
        RECT 1418.250 1642.580 1418.570 1642.640 ;
        RECT 1418.710 1587.020 1419.030 1587.080 ;
        RECT 1418.515 1586.880 1419.030 1587.020 ;
        RECT 1418.710 1586.820 1419.030 1586.880 ;
        RECT 1418.710 1497.940 1419.030 1498.000 ;
        RECT 1418.515 1497.800 1419.030 1497.940 ;
        RECT 1418.710 1497.740 1419.030 1497.800 ;
        RECT 1418.710 1490.460 1419.030 1490.520 ;
        RECT 1418.515 1490.320 1419.030 1490.460 ;
        RECT 1418.710 1490.260 1419.030 1490.320 ;
        RECT 1418.725 1442.180 1419.015 1442.225 ;
        RECT 1419.170 1442.180 1419.490 1442.240 ;
        RECT 1418.725 1442.040 1419.490 1442.180 ;
        RECT 1418.725 1441.995 1419.015 1442.040 ;
        RECT 1419.170 1441.980 1419.490 1442.040 ;
        RECT 1418.710 1362.620 1419.030 1362.680 ;
        RECT 2601.830 1362.620 2602.150 1362.680 ;
        RECT 1418.710 1362.480 2602.150 1362.620 ;
        RECT 1418.710 1362.420 1419.030 1362.480 ;
        RECT 2601.830 1362.420 2602.150 1362.480 ;
      LAYER via ;
        RECT 1417.820 1689.500 1418.080 1689.760 ;
        RECT 1418.280 1642.580 1418.540 1642.840 ;
        RECT 1418.740 1586.820 1419.000 1587.080 ;
        RECT 1418.740 1497.740 1419.000 1498.000 ;
        RECT 1418.740 1490.260 1419.000 1490.520 ;
        RECT 1419.200 1441.980 1419.460 1442.240 ;
        RECT 1418.740 1362.420 1419.000 1362.680 ;
        RECT 2601.860 1362.420 2602.120 1362.680 ;
      LAYER met2 ;
        RECT 1417.720 1700.340 1418.000 1704.000 ;
        RECT 1417.720 1700.000 1418.020 1700.340 ;
        RECT 1417.880 1689.790 1418.020 1700.000 ;
        RECT 1417.820 1689.470 1418.080 1689.790 ;
        RECT 1418.280 1642.550 1418.540 1642.870 ;
        RECT 1418.340 1618.130 1418.480 1642.550 ;
        RECT 1418.340 1617.990 1418.940 1618.130 ;
        RECT 1418.800 1587.110 1418.940 1617.990 ;
        RECT 1418.740 1586.790 1419.000 1587.110 ;
        RECT 1418.740 1497.710 1419.000 1498.030 ;
        RECT 1418.800 1490.550 1418.940 1497.710 ;
        RECT 1418.740 1490.230 1419.000 1490.550 ;
        RECT 1419.200 1441.950 1419.460 1442.270 ;
        RECT 1419.260 1400.530 1419.400 1441.950 ;
        RECT 1418.800 1400.390 1419.400 1400.530 ;
        RECT 1418.800 1362.710 1418.940 1400.390 ;
        RECT 1418.740 1362.390 1419.000 1362.710 ;
        RECT 2601.860 1362.390 2602.120 1362.710 ;
        RECT 2601.920 17.410 2602.060 1362.390 ;
        RECT 2601.920 17.270 2607.580 17.410 ;
        RECT 2607.440 2.400 2607.580 17.270 ;
        RECT 2607.230 -4.800 2607.790 2.400 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1420.090 1666.240 1420.410 1666.300 ;
        RECT 1424.690 1666.240 1425.010 1666.300 ;
        RECT 1420.090 1666.100 1425.010 1666.240 ;
        RECT 1420.090 1666.040 1420.410 1666.100 ;
        RECT 1424.690 1666.040 1425.010 1666.100 ;
        RECT 1424.690 1452.380 1425.010 1452.440 ;
        RECT 2622.070 1452.380 2622.390 1452.440 ;
        RECT 1424.690 1452.240 2622.390 1452.380 ;
        RECT 1424.690 1452.180 1425.010 1452.240 ;
        RECT 2622.070 1452.180 2622.390 1452.240 ;
      LAYER via ;
        RECT 1420.120 1666.040 1420.380 1666.300 ;
        RECT 1424.720 1666.040 1424.980 1666.300 ;
        RECT 1424.720 1452.180 1424.980 1452.440 ;
        RECT 2622.100 1452.180 2622.360 1452.440 ;
      LAYER met2 ;
        RECT 1419.560 1700.340 1419.840 1704.000 ;
        RECT 1419.560 1700.000 1419.860 1700.340 ;
        RECT 1419.720 1678.650 1419.860 1700.000 ;
        RECT 1419.720 1678.510 1420.320 1678.650 ;
        RECT 1420.180 1666.330 1420.320 1678.510 ;
        RECT 1420.120 1666.010 1420.380 1666.330 ;
        RECT 1424.720 1666.010 1424.980 1666.330 ;
        RECT 1424.780 1452.470 1424.920 1666.010 ;
        RECT 1424.720 1452.150 1424.980 1452.470 ;
        RECT 2622.100 1452.150 2622.360 1452.470 ;
        RECT 2622.160 17.410 2622.300 1452.150 ;
        RECT 2622.160 17.270 2625.520 17.410 ;
        RECT 2625.380 2.400 2625.520 17.270 ;
        RECT 2625.170 -4.800 2625.730 2.400 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1422.390 1355.820 1422.710 1355.880 ;
        RECT 2643.230 1355.820 2643.550 1355.880 ;
        RECT 1422.390 1355.680 2643.550 1355.820 ;
        RECT 1422.390 1355.620 1422.710 1355.680 ;
        RECT 2643.230 1355.620 2643.550 1355.680 ;
      LAYER via ;
        RECT 1422.420 1355.620 1422.680 1355.880 ;
        RECT 2643.260 1355.620 2643.520 1355.880 ;
      LAYER met2 ;
        RECT 1421.400 1700.410 1421.680 1704.000 ;
        RECT 1421.400 1700.270 1422.160 1700.410 ;
        RECT 1421.400 1700.000 1421.680 1700.270 ;
        RECT 1422.020 1666.410 1422.160 1700.270 ;
        RECT 1422.020 1666.270 1422.620 1666.410 ;
        RECT 1422.480 1355.910 1422.620 1666.270 ;
        RECT 1422.420 1355.590 1422.680 1355.910 ;
        RECT 2643.260 1355.590 2643.520 1355.910 ;
        RECT 2643.320 2.400 2643.460 1355.590 ;
        RECT 2643.110 -4.800 2643.670 2.400 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1422.925 1594.005 1423.095 1642.115 ;
        RECT 1423.385 1510.705 1423.555 1545.555 ;
      LAYER mcon ;
        RECT 1422.925 1641.945 1423.095 1642.115 ;
        RECT 1423.385 1545.385 1423.555 1545.555 ;
      LAYER met1 ;
        RECT 1422.850 1642.100 1423.170 1642.160 ;
        RECT 1422.655 1641.960 1423.170 1642.100 ;
        RECT 1422.850 1641.900 1423.170 1641.960 ;
        RECT 1422.850 1594.160 1423.170 1594.220 ;
        RECT 1422.655 1594.020 1423.170 1594.160 ;
        RECT 1422.850 1593.960 1423.170 1594.020 ;
        RECT 1423.310 1545.540 1423.630 1545.600 ;
        RECT 1423.115 1545.400 1423.630 1545.540 ;
        RECT 1423.310 1545.340 1423.630 1545.400 ;
        RECT 1423.310 1510.860 1423.630 1510.920 ;
        RECT 1423.115 1510.720 1423.630 1510.860 ;
        RECT 1423.310 1510.660 1423.630 1510.720 ;
        RECT 1421.930 1448.980 1422.250 1449.040 ;
        RECT 1423.310 1448.980 1423.630 1449.040 ;
        RECT 1421.930 1448.840 1423.630 1448.980 ;
        RECT 1421.930 1448.780 1422.250 1448.840 ;
        RECT 1423.310 1448.780 1423.630 1448.840 ;
        RECT 1421.930 1395.940 1422.250 1396.000 ;
        RECT 1424.690 1395.940 1425.010 1396.000 ;
        RECT 1421.930 1395.800 1425.010 1395.940 ;
        RECT 1421.930 1395.740 1422.250 1395.800 ;
        RECT 1424.690 1395.740 1425.010 1395.800 ;
        RECT 1424.690 1349.020 1425.010 1349.080 ;
        RECT 2656.570 1349.020 2656.890 1349.080 ;
        RECT 1424.690 1348.880 2656.890 1349.020 ;
        RECT 1424.690 1348.820 1425.010 1348.880 ;
        RECT 2656.570 1348.820 2656.890 1348.880 ;
      LAYER via ;
        RECT 1422.880 1641.900 1423.140 1642.160 ;
        RECT 1422.880 1593.960 1423.140 1594.220 ;
        RECT 1423.340 1545.340 1423.600 1545.600 ;
        RECT 1423.340 1510.660 1423.600 1510.920 ;
        RECT 1421.960 1448.780 1422.220 1449.040 ;
        RECT 1423.340 1448.780 1423.600 1449.040 ;
        RECT 1421.960 1395.740 1422.220 1396.000 ;
        RECT 1424.720 1395.740 1424.980 1396.000 ;
        RECT 1424.720 1348.820 1424.980 1349.080 ;
        RECT 2656.600 1348.820 2656.860 1349.080 ;
      LAYER met2 ;
        RECT 1423.240 1700.340 1423.520 1704.000 ;
        RECT 1423.240 1700.000 1423.540 1700.340 ;
        RECT 1423.400 1666.410 1423.540 1700.000 ;
        RECT 1422.940 1666.270 1423.540 1666.410 ;
        RECT 1422.940 1642.190 1423.080 1666.270 ;
        RECT 1422.880 1641.870 1423.140 1642.190 ;
        RECT 1422.880 1593.930 1423.140 1594.250 ;
        RECT 1422.940 1569.850 1423.080 1593.930 ;
        RECT 1422.940 1569.710 1423.540 1569.850 ;
        RECT 1423.400 1545.630 1423.540 1569.710 ;
        RECT 1423.340 1545.310 1423.600 1545.630 ;
        RECT 1423.340 1510.630 1423.600 1510.950 ;
        RECT 1423.400 1449.070 1423.540 1510.630 ;
        RECT 1421.960 1448.750 1422.220 1449.070 ;
        RECT 1423.340 1448.750 1423.600 1449.070 ;
        RECT 1422.020 1396.030 1422.160 1448.750 ;
        RECT 1421.960 1395.710 1422.220 1396.030 ;
        RECT 1424.720 1395.710 1424.980 1396.030 ;
        RECT 1424.780 1349.110 1424.920 1395.710 ;
        RECT 1424.720 1348.790 1424.980 1349.110 ;
        RECT 2656.600 1348.790 2656.860 1349.110 ;
        RECT 2656.660 17.410 2656.800 1348.790 ;
        RECT 2656.660 17.270 2661.400 17.410 ;
        RECT 2661.260 2.400 2661.400 17.270 ;
        RECT 2661.050 -4.800 2661.610 2.400 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1423.770 1341.880 1424.090 1341.940 ;
        RECT 2677.270 1341.880 2677.590 1341.940 ;
        RECT 1423.770 1341.740 2677.590 1341.880 ;
        RECT 1423.770 1341.680 1424.090 1341.740 ;
        RECT 2677.270 1341.680 2677.590 1341.740 ;
      LAYER via ;
        RECT 1423.800 1341.680 1424.060 1341.940 ;
        RECT 2677.300 1341.680 2677.560 1341.940 ;
      LAYER met2 ;
        RECT 1425.080 1700.340 1425.360 1704.000 ;
        RECT 1425.080 1700.000 1425.380 1700.340 ;
        RECT 1425.240 1677.970 1425.380 1700.000 ;
        RECT 1423.860 1677.830 1425.380 1677.970 ;
        RECT 1423.860 1341.970 1424.000 1677.830 ;
        RECT 1423.800 1341.650 1424.060 1341.970 ;
        RECT 2677.300 1341.650 2677.560 1341.970 ;
        RECT 2677.360 17.410 2677.500 1341.650 ;
        RECT 2677.360 17.270 2678.880 17.410 ;
        RECT 2678.740 2.400 2678.880 17.270 ;
        RECT 2678.530 -4.800 2679.090 2.400 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1424.230 1621.360 1424.550 1621.420 ;
        RECT 1426.990 1621.360 1427.310 1621.420 ;
        RECT 1424.230 1621.220 1427.310 1621.360 ;
        RECT 1424.230 1621.160 1424.550 1621.220 ;
        RECT 1426.990 1621.160 1427.310 1621.220 ;
        RECT 1424.230 1335.080 1424.550 1335.140 ;
        RECT 2691.070 1335.080 2691.390 1335.140 ;
        RECT 1424.230 1334.940 2691.390 1335.080 ;
        RECT 1424.230 1334.880 1424.550 1334.940 ;
        RECT 2691.070 1334.880 2691.390 1334.940 ;
      LAYER via ;
        RECT 1424.260 1621.160 1424.520 1621.420 ;
        RECT 1427.020 1621.160 1427.280 1621.420 ;
        RECT 1424.260 1334.880 1424.520 1335.140 ;
        RECT 2691.100 1334.880 2691.360 1335.140 ;
      LAYER met2 ;
        RECT 1426.920 1700.340 1427.200 1704.000 ;
        RECT 1426.920 1700.000 1427.220 1700.340 ;
        RECT 1427.080 1621.450 1427.220 1700.000 ;
        RECT 1424.260 1621.130 1424.520 1621.450 ;
        RECT 1427.020 1621.130 1427.280 1621.450 ;
        RECT 1424.320 1335.170 1424.460 1621.130 ;
        RECT 1424.260 1334.850 1424.520 1335.170 ;
        RECT 2691.100 1334.850 2691.360 1335.170 ;
        RECT 2691.160 17.410 2691.300 1334.850 ;
        RECT 2691.160 17.270 2696.820 17.410 ;
        RECT 2696.680 2.400 2696.820 17.270 ;
        RECT 2696.470 -4.800 2697.030 2.400 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1429.290 1664.540 1429.610 1664.600 ;
        RECT 1433.890 1664.540 1434.210 1664.600 ;
        RECT 1429.290 1664.400 1434.210 1664.540 ;
        RECT 1429.290 1664.340 1429.610 1664.400 ;
        RECT 1433.890 1664.340 1434.210 1664.400 ;
        RECT 1433.890 1328.280 1434.210 1328.340 ;
        RECT 2711.770 1328.280 2712.090 1328.340 ;
        RECT 1433.890 1328.140 2712.090 1328.280 ;
        RECT 1433.890 1328.080 1434.210 1328.140 ;
        RECT 2711.770 1328.080 2712.090 1328.140 ;
      LAYER via ;
        RECT 1429.320 1664.340 1429.580 1664.600 ;
        RECT 1433.920 1664.340 1434.180 1664.600 ;
        RECT 1433.920 1328.080 1434.180 1328.340 ;
        RECT 2711.800 1328.080 2712.060 1328.340 ;
      LAYER met2 ;
        RECT 1428.760 1700.410 1429.040 1704.000 ;
        RECT 1428.760 1700.270 1429.520 1700.410 ;
        RECT 1428.760 1700.000 1429.040 1700.270 ;
        RECT 1429.380 1664.630 1429.520 1700.270 ;
        RECT 1429.320 1664.310 1429.580 1664.630 ;
        RECT 1433.920 1664.310 1434.180 1664.630 ;
        RECT 1433.980 1328.370 1434.120 1664.310 ;
        RECT 1433.920 1328.050 1434.180 1328.370 ;
        RECT 2711.800 1328.050 2712.060 1328.370 ;
        RECT 2711.860 17.410 2712.000 1328.050 ;
        RECT 2711.860 17.270 2714.760 17.410 ;
        RECT 2714.620 2.400 2714.760 17.270 ;
        RECT 2714.410 -4.800 2714.970 2.400 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1430.670 1314.340 1430.990 1314.400 ;
        RECT 2732.930 1314.340 2733.250 1314.400 ;
        RECT 1430.670 1314.200 2733.250 1314.340 ;
        RECT 1430.670 1314.140 1430.990 1314.200 ;
        RECT 2732.930 1314.140 2733.250 1314.200 ;
      LAYER via ;
        RECT 1430.700 1314.140 1430.960 1314.400 ;
        RECT 2732.960 1314.140 2733.220 1314.400 ;
      LAYER met2 ;
        RECT 1430.600 1700.340 1430.880 1704.000 ;
        RECT 1430.600 1700.000 1430.900 1700.340 ;
        RECT 1430.760 1314.430 1430.900 1700.000 ;
        RECT 1430.700 1314.110 1430.960 1314.430 ;
        RECT 2732.960 1314.110 2733.220 1314.430 ;
        RECT 2733.020 17.410 2733.160 1314.110 ;
        RECT 2732.560 17.270 2733.160 17.410 ;
        RECT 2732.560 2.400 2732.700 17.270 ;
        RECT 2732.350 -4.800 2732.910 2.400 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1430.210 1683.920 1430.530 1683.980 ;
        RECT 1432.510 1683.920 1432.830 1683.980 ;
        RECT 1430.210 1683.780 1432.830 1683.920 ;
        RECT 1430.210 1683.720 1430.530 1683.780 ;
        RECT 1432.510 1683.720 1432.830 1683.780 ;
        RECT 1430.210 1445.580 1430.530 1445.640 ;
        RECT 2746.270 1445.580 2746.590 1445.640 ;
        RECT 1430.210 1445.440 2746.590 1445.580 ;
        RECT 1430.210 1445.380 1430.530 1445.440 ;
        RECT 2746.270 1445.380 2746.590 1445.440 ;
      LAYER via ;
        RECT 1430.240 1683.720 1430.500 1683.980 ;
        RECT 1432.540 1683.720 1432.800 1683.980 ;
        RECT 1430.240 1445.380 1430.500 1445.640 ;
        RECT 2746.300 1445.380 2746.560 1445.640 ;
      LAYER met2 ;
        RECT 1432.440 1700.340 1432.720 1704.000 ;
        RECT 1432.440 1700.000 1432.740 1700.340 ;
        RECT 1432.600 1684.010 1432.740 1700.000 ;
        RECT 1430.240 1683.690 1430.500 1684.010 ;
        RECT 1432.540 1683.690 1432.800 1684.010 ;
        RECT 1430.300 1445.670 1430.440 1683.690 ;
        RECT 1430.240 1445.350 1430.500 1445.670 ;
        RECT 2746.300 1445.350 2746.560 1445.670 ;
        RECT 2746.360 17.410 2746.500 1445.350 ;
        RECT 2746.360 17.270 2750.640 17.410 ;
        RECT 2750.500 2.400 2750.640 17.270 ;
        RECT 2750.290 -4.800 2750.850 2.400 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1431.130 1684.940 1431.450 1685.000 ;
        RECT 1434.350 1684.940 1434.670 1685.000 ;
        RECT 1431.130 1684.800 1434.670 1684.940 ;
        RECT 1431.130 1684.740 1431.450 1684.800 ;
        RECT 1434.350 1684.740 1434.670 1684.800 ;
        RECT 1431.130 1307.540 1431.450 1307.600 ;
        RECT 2766.970 1307.540 2767.290 1307.600 ;
        RECT 1431.130 1307.400 2767.290 1307.540 ;
        RECT 1431.130 1307.340 1431.450 1307.400 ;
        RECT 2766.970 1307.340 2767.290 1307.400 ;
      LAYER via ;
        RECT 1431.160 1684.740 1431.420 1685.000 ;
        RECT 1434.380 1684.740 1434.640 1685.000 ;
        RECT 1431.160 1307.340 1431.420 1307.600 ;
        RECT 2767.000 1307.340 2767.260 1307.600 ;
      LAYER met2 ;
        RECT 1434.280 1700.340 1434.560 1704.000 ;
        RECT 1434.280 1700.000 1434.580 1700.340 ;
        RECT 1434.440 1685.030 1434.580 1700.000 ;
        RECT 1431.160 1684.710 1431.420 1685.030 ;
        RECT 1434.380 1684.710 1434.640 1685.030 ;
        RECT 1431.220 1307.630 1431.360 1684.710 ;
        RECT 1431.160 1307.310 1431.420 1307.630 ;
        RECT 2767.000 1307.310 2767.260 1307.630 ;
        RECT 2767.060 17.410 2767.200 1307.310 ;
        RECT 2767.060 17.270 2768.120 17.410 ;
        RECT 2767.980 2.400 2768.120 17.270 ;
        RECT 2767.770 -4.800 2768.330 2.400 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 840.950 38.320 841.270 38.380 ;
        RECT 1236.550 38.320 1236.870 38.380 ;
        RECT 840.950 38.180 1236.870 38.320 ;
        RECT 840.950 38.120 841.270 38.180 ;
        RECT 1236.550 38.120 1236.870 38.180 ;
      LAYER via ;
        RECT 840.980 38.120 841.240 38.380 ;
        RECT 1236.580 38.120 1236.840 38.380 ;
      LAYER met2 ;
        RECT 1236.020 1700.340 1236.300 1704.000 ;
        RECT 1236.020 1700.000 1236.320 1700.340 ;
        RECT 1236.180 1673.890 1236.320 1700.000 ;
        RECT 1236.180 1673.750 1236.780 1673.890 ;
        RECT 1236.640 38.410 1236.780 1673.750 ;
        RECT 840.980 38.090 841.240 38.410 ;
        RECT 1236.580 38.090 1236.840 38.410 ;
        RECT 841.040 2.400 841.180 38.090 ;
        RECT 840.830 -4.800 841.390 2.400 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1436.190 1300.740 1436.510 1300.800 ;
        RECT 2780.770 1300.740 2781.090 1300.800 ;
        RECT 1436.190 1300.600 2781.090 1300.740 ;
        RECT 1436.190 1300.540 1436.510 1300.600 ;
        RECT 2780.770 1300.540 2781.090 1300.600 ;
      LAYER via ;
        RECT 1436.220 1300.540 1436.480 1300.800 ;
        RECT 2780.800 1300.540 2781.060 1300.800 ;
      LAYER met2 ;
        RECT 1436.120 1700.340 1436.400 1704.000 ;
        RECT 1436.120 1700.000 1436.420 1700.340 ;
        RECT 1436.280 1300.830 1436.420 1700.000 ;
        RECT 1436.220 1300.510 1436.480 1300.830 ;
        RECT 2780.800 1300.510 2781.060 1300.830 ;
        RECT 2780.860 18.090 2781.000 1300.510 ;
        RECT 2780.860 17.950 2786.060 18.090 ;
        RECT 2785.920 2.400 2786.060 17.950 ;
        RECT 2785.710 -4.800 2786.270 2.400 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1438.105 1635.485 1438.275 1678.495 ;
        RECT 1440.865 1538.925 1441.035 1587.035 ;
        RECT 1440.865 1442.025 1441.035 1490.475 ;
      LAYER mcon ;
        RECT 1438.105 1678.325 1438.275 1678.495 ;
        RECT 1440.865 1586.865 1441.035 1587.035 ;
        RECT 1440.865 1490.305 1441.035 1490.475 ;
      LAYER met1 ;
        RECT 1438.030 1678.480 1438.350 1678.540 ;
        RECT 1437.835 1678.340 1438.350 1678.480 ;
        RECT 1438.030 1678.280 1438.350 1678.340 ;
        RECT 1438.045 1635.640 1438.335 1635.685 ;
        RECT 1440.790 1635.640 1441.110 1635.700 ;
        RECT 1438.045 1635.500 1441.110 1635.640 ;
        RECT 1438.045 1635.455 1438.335 1635.500 ;
        RECT 1440.790 1635.440 1441.110 1635.500 ;
        RECT 1440.790 1587.020 1441.110 1587.080 ;
        RECT 1440.595 1586.880 1441.110 1587.020 ;
        RECT 1440.790 1586.820 1441.110 1586.880 ;
        RECT 1440.790 1539.080 1441.110 1539.140 ;
        RECT 1440.595 1538.940 1441.110 1539.080 ;
        RECT 1440.790 1538.880 1441.110 1538.940 ;
        RECT 1440.790 1490.460 1441.110 1490.520 ;
        RECT 1440.595 1490.320 1441.110 1490.460 ;
        RECT 1440.790 1490.260 1441.110 1490.320 ;
        RECT 1440.790 1442.180 1441.110 1442.240 ;
        RECT 1440.595 1442.040 1441.110 1442.180 ;
        RECT 1440.790 1441.980 1441.110 1442.040 ;
        RECT 1440.330 1345.620 1440.650 1345.680 ;
        RECT 1440.790 1345.620 1441.110 1345.680 ;
        RECT 1440.330 1345.480 1441.110 1345.620 ;
        RECT 1440.330 1345.420 1440.650 1345.480 ;
        RECT 1440.790 1345.420 1441.110 1345.480 ;
        RECT 1440.790 1293.600 1441.110 1293.660 ;
        RECT 2801.470 1293.600 2801.790 1293.660 ;
        RECT 1440.790 1293.460 2801.790 1293.600 ;
        RECT 1440.790 1293.400 1441.110 1293.460 ;
        RECT 2801.470 1293.400 2801.790 1293.460 ;
      LAYER via ;
        RECT 1438.060 1678.280 1438.320 1678.540 ;
        RECT 1440.820 1635.440 1441.080 1635.700 ;
        RECT 1440.820 1586.820 1441.080 1587.080 ;
        RECT 1440.820 1538.880 1441.080 1539.140 ;
        RECT 1440.820 1490.260 1441.080 1490.520 ;
        RECT 1440.820 1441.980 1441.080 1442.240 ;
        RECT 1440.360 1345.420 1440.620 1345.680 ;
        RECT 1440.820 1345.420 1441.080 1345.680 ;
        RECT 1440.820 1293.400 1441.080 1293.660 ;
        RECT 2801.500 1293.400 2801.760 1293.660 ;
      LAYER met2 ;
        RECT 1437.960 1700.340 1438.240 1704.000 ;
        RECT 1437.960 1700.000 1438.260 1700.340 ;
        RECT 1438.120 1678.570 1438.260 1700.000 ;
        RECT 1438.060 1678.250 1438.320 1678.570 ;
        RECT 1440.820 1635.410 1441.080 1635.730 ;
        RECT 1440.880 1587.110 1441.020 1635.410 ;
        RECT 1440.820 1586.790 1441.080 1587.110 ;
        RECT 1440.820 1538.850 1441.080 1539.170 ;
        RECT 1440.880 1490.550 1441.020 1538.850 ;
        RECT 1440.820 1490.230 1441.080 1490.550 ;
        RECT 1440.820 1441.950 1441.080 1442.270 ;
        RECT 1440.880 1424.840 1441.020 1441.950 ;
        RECT 1440.880 1424.700 1441.480 1424.840 ;
        RECT 1441.340 1393.845 1441.480 1424.700 ;
        RECT 1440.350 1393.475 1440.630 1393.845 ;
        RECT 1441.270 1393.475 1441.550 1393.845 ;
        RECT 1440.420 1345.710 1440.560 1393.475 ;
        RECT 1440.360 1345.390 1440.620 1345.710 ;
        RECT 1440.820 1345.390 1441.080 1345.710 ;
        RECT 1440.880 1293.690 1441.020 1345.390 ;
        RECT 1440.820 1293.370 1441.080 1293.690 ;
        RECT 2801.500 1293.370 2801.760 1293.690 ;
        RECT 2801.560 17.410 2801.700 1293.370 ;
        RECT 2801.560 17.270 2804.000 17.410 ;
        RECT 2803.860 2.400 2804.000 17.270 ;
        RECT 2803.650 -4.800 2804.210 2.400 ;
      LAYER via2 ;
        RECT 1440.350 1393.520 1440.630 1393.800 ;
        RECT 1441.270 1393.520 1441.550 1393.800 ;
      LAYER met3 ;
        RECT 1440.325 1393.810 1440.655 1393.825 ;
        RECT 1441.245 1393.810 1441.575 1393.825 ;
        RECT 1440.325 1393.510 1441.575 1393.810 ;
        RECT 1440.325 1393.495 1440.655 1393.510 ;
        RECT 1441.245 1393.495 1441.575 1393.510 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1438.490 1683.920 1438.810 1683.980 ;
        RECT 1439.870 1683.920 1440.190 1683.980 ;
        RECT 1438.490 1683.780 1440.190 1683.920 ;
        RECT 1438.490 1683.720 1438.810 1683.780 ;
        RECT 1439.870 1683.720 1440.190 1683.780 ;
        RECT 1437.570 1608.100 1437.890 1608.160 ;
        RECT 1438.490 1608.100 1438.810 1608.160 ;
        RECT 1437.570 1607.960 1438.810 1608.100 ;
        RECT 1437.570 1607.900 1437.890 1607.960 ;
        RECT 1438.490 1607.900 1438.810 1607.960 ;
        RECT 1437.570 1286.800 1437.890 1286.860 ;
        RECT 2815.730 1286.800 2816.050 1286.860 ;
        RECT 1437.570 1286.660 2816.050 1286.800 ;
        RECT 1437.570 1286.600 1437.890 1286.660 ;
        RECT 2815.730 1286.600 2816.050 1286.660 ;
        RECT 2815.730 18.260 2816.050 18.320 ;
        RECT 2821.710 18.260 2822.030 18.320 ;
        RECT 2815.730 18.120 2822.030 18.260 ;
        RECT 2815.730 18.060 2816.050 18.120 ;
        RECT 2821.710 18.060 2822.030 18.120 ;
      LAYER via ;
        RECT 1438.520 1683.720 1438.780 1683.980 ;
        RECT 1439.900 1683.720 1440.160 1683.980 ;
        RECT 1437.600 1607.900 1437.860 1608.160 ;
        RECT 1438.520 1607.900 1438.780 1608.160 ;
        RECT 1437.600 1286.600 1437.860 1286.860 ;
        RECT 2815.760 1286.600 2816.020 1286.860 ;
        RECT 2815.760 18.060 2816.020 18.320 ;
        RECT 2821.740 18.060 2822.000 18.320 ;
      LAYER met2 ;
        RECT 1439.800 1700.340 1440.080 1704.000 ;
        RECT 1439.800 1700.000 1440.100 1700.340 ;
        RECT 1439.960 1684.010 1440.100 1700.000 ;
        RECT 1438.520 1683.690 1438.780 1684.010 ;
        RECT 1439.900 1683.690 1440.160 1684.010 ;
        RECT 1438.580 1608.190 1438.720 1683.690 ;
        RECT 1437.600 1607.870 1437.860 1608.190 ;
        RECT 1438.520 1607.870 1438.780 1608.190 ;
        RECT 1437.660 1286.890 1437.800 1607.870 ;
        RECT 1437.600 1286.570 1437.860 1286.890 ;
        RECT 2815.760 1286.570 2816.020 1286.890 ;
        RECT 2815.820 18.350 2815.960 1286.570 ;
        RECT 2815.760 18.030 2816.020 18.350 ;
        RECT 2821.740 18.030 2822.000 18.350 ;
        RECT 2821.800 2.400 2821.940 18.030 ;
        RECT 2821.590 -4.800 2822.150 2.400 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1437.110 1685.960 1437.430 1686.020 ;
        RECT 1441.710 1685.960 1442.030 1686.020 ;
        RECT 1437.110 1685.820 1442.030 1685.960 ;
        RECT 1437.110 1685.760 1437.430 1685.820 ;
        RECT 1441.710 1685.760 1442.030 1685.820 ;
        RECT 1438.030 113.800 1438.350 113.860 ;
        RECT 2835.970 113.800 2836.290 113.860 ;
        RECT 1438.030 113.660 2836.290 113.800 ;
        RECT 1438.030 113.600 1438.350 113.660 ;
        RECT 2835.970 113.600 2836.290 113.660 ;
      LAYER via ;
        RECT 1437.140 1685.760 1437.400 1686.020 ;
        RECT 1441.740 1685.760 1442.000 1686.020 ;
        RECT 1438.060 113.600 1438.320 113.860 ;
        RECT 2836.000 113.600 2836.260 113.860 ;
      LAYER met2 ;
        RECT 1441.640 1700.340 1441.920 1704.000 ;
        RECT 1441.640 1700.000 1441.940 1700.340 ;
        RECT 1441.800 1686.050 1441.940 1700.000 ;
        RECT 1437.140 1685.730 1437.400 1686.050 ;
        RECT 1441.740 1685.730 1442.000 1686.050 ;
        RECT 1437.200 1677.970 1437.340 1685.730 ;
        RECT 1437.200 1677.830 1438.260 1677.970 ;
        RECT 1438.120 113.890 1438.260 1677.830 ;
        RECT 1438.060 113.570 1438.320 113.890 ;
        RECT 2836.000 113.570 2836.260 113.890 ;
        RECT 2836.060 16.730 2836.200 113.570 ;
        RECT 2836.060 16.590 2839.420 16.730 ;
        RECT 2839.280 2.400 2839.420 16.590 ;
        RECT 2839.070 -4.800 2839.630 2.400 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1444.930 1559.140 1445.250 1559.200 ;
        RECT 1446.310 1559.140 1446.630 1559.200 ;
        RECT 1444.930 1559.000 1446.630 1559.140 ;
        RECT 1444.930 1558.940 1445.250 1559.000 ;
        RECT 1446.310 1558.940 1446.630 1559.000 ;
        RECT 1446.770 1438.440 1447.090 1438.500 ;
        RECT 2857.130 1438.440 2857.450 1438.500 ;
        RECT 1446.770 1438.300 2857.450 1438.440 ;
        RECT 1446.770 1438.240 1447.090 1438.300 ;
        RECT 2857.130 1438.240 2857.450 1438.300 ;
      LAYER via ;
        RECT 1444.960 1558.940 1445.220 1559.200 ;
        RECT 1446.340 1558.940 1446.600 1559.200 ;
        RECT 1446.800 1438.240 1447.060 1438.500 ;
        RECT 2857.160 1438.240 2857.420 1438.500 ;
      LAYER met2 ;
        RECT 1443.480 1700.410 1443.760 1704.000 ;
        RECT 1443.480 1700.270 1444.240 1700.410 ;
        RECT 1443.480 1700.000 1443.760 1700.270 ;
        RECT 1444.100 1660.290 1444.240 1700.270 ;
        RECT 1444.100 1660.150 1445.160 1660.290 ;
        RECT 1445.020 1631.050 1445.160 1660.150 ;
        RECT 1445.020 1630.910 1446.080 1631.050 ;
        RECT 1445.940 1583.450 1446.080 1630.910 ;
        RECT 1445.940 1583.310 1446.540 1583.450 ;
        RECT 1446.400 1559.230 1446.540 1583.310 ;
        RECT 1444.960 1558.910 1445.220 1559.230 ;
        RECT 1446.340 1558.910 1446.600 1559.230 ;
        RECT 1445.020 1465.810 1445.160 1558.910 ;
        RECT 1445.020 1465.670 1447.000 1465.810 ;
        RECT 1446.860 1438.530 1447.000 1465.670 ;
        RECT 1446.800 1438.210 1447.060 1438.530 ;
        RECT 2857.160 1438.210 2857.420 1438.530 ;
        RECT 2857.220 2.400 2857.360 1438.210 ;
        RECT 2857.010 -4.800 2857.570 2.400 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2855.365 16.065 2855.535 17.935 ;
      LAYER mcon ;
        RECT 2855.365 17.765 2855.535 17.935 ;
      LAYER met1 ;
        RECT 1445.390 1683.920 1445.710 1683.980 ;
        RECT 1447.230 1683.920 1447.550 1683.980 ;
        RECT 1445.390 1683.780 1447.550 1683.920 ;
        RECT 1445.390 1683.720 1445.710 1683.780 ;
        RECT 1447.230 1683.720 1447.550 1683.780 ;
        RECT 1447.230 1480.260 1447.550 1480.320 ;
        RECT 2411.390 1480.260 2411.710 1480.320 ;
        RECT 1447.230 1480.120 2411.710 1480.260 ;
        RECT 1447.230 1480.060 1447.550 1480.120 ;
        RECT 2411.390 1480.060 2411.710 1480.120 ;
        RECT 2411.390 17.920 2411.710 17.980 ;
        RECT 2855.305 17.920 2855.595 17.965 ;
        RECT 2411.390 17.780 2855.595 17.920 ;
        RECT 2411.390 17.720 2411.710 17.780 ;
        RECT 2855.305 17.735 2855.595 17.780 ;
        RECT 2855.305 16.220 2855.595 16.265 ;
        RECT 2875.070 16.220 2875.390 16.280 ;
        RECT 2855.305 16.080 2875.390 16.220 ;
        RECT 2855.305 16.035 2855.595 16.080 ;
        RECT 2875.070 16.020 2875.390 16.080 ;
      LAYER via ;
        RECT 1445.420 1683.720 1445.680 1683.980 ;
        RECT 1447.260 1683.720 1447.520 1683.980 ;
        RECT 1447.260 1480.060 1447.520 1480.320 ;
        RECT 2411.420 1480.060 2411.680 1480.320 ;
        RECT 2411.420 17.720 2411.680 17.980 ;
        RECT 2875.100 16.020 2875.360 16.280 ;
      LAYER met2 ;
        RECT 1445.320 1700.340 1445.600 1704.000 ;
        RECT 1445.320 1700.000 1445.620 1700.340 ;
        RECT 1445.480 1684.010 1445.620 1700.000 ;
        RECT 1445.420 1683.690 1445.680 1684.010 ;
        RECT 1447.260 1683.690 1447.520 1684.010 ;
        RECT 1447.320 1480.350 1447.460 1683.690 ;
        RECT 1447.260 1480.030 1447.520 1480.350 ;
        RECT 2411.420 1480.030 2411.680 1480.350 ;
        RECT 2411.480 18.010 2411.620 1480.030 ;
        RECT 2411.420 17.690 2411.680 18.010 ;
        RECT 2875.100 15.990 2875.360 16.310 ;
        RECT 2875.160 2.400 2875.300 15.990 ;
        RECT 2874.950 -4.800 2875.510 2.400 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2859.965 16.745 2860.135 17.595 ;
      LAYER mcon ;
        RECT 2859.965 17.425 2860.135 17.595 ;
      LAYER met1 ;
        RECT 1447.690 1473.460 1448.010 1473.520 ;
        RECT 2376.890 1473.460 2377.210 1473.520 ;
        RECT 1447.690 1473.320 2377.210 1473.460 ;
        RECT 1447.690 1473.260 1448.010 1473.320 ;
        RECT 2376.890 1473.260 2377.210 1473.320 ;
        RECT 2376.890 17.580 2377.210 17.640 ;
        RECT 2859.905 17.580 2860.195 17.625 ;
        RECT 2376.890 17.440 2860.195 17.580 ;
        RECT 2376.890 17.380 2377.210 17.440 ;
        RECT 2859.905 17.395 2860.195 17.440 ;
        RECT 2859.905 16.900 2860.195 16.945 ;
        RECT 2893.010 16.900 2893.330 16.960 ;
        RECT 2859.905 16.760 2893.330 16.900 ;
        RECT 2859.905 16.715 2860.195 16.760 ;
        RECT 2893.010 16.700 2893.330 16.760 ;
      LAYER via ;
        RECT 1447.720 1473.260 1447.980 1473.520 ;
        RECT 2376.920 1473.260 2377.180 1473.520 ;
        RECT 2376.920 17.380 2377.180 17.640 ;
        RECT 2893.040 16.700 2893.300 16.960 ;
      LAYER met2 ;
        RECT 1447.160 1700.410 1447.440 1704.000 ;
        RECT 1447.160 1700.270 1447.920 1700.410 ;
        RECT 1447.160 1700.000 1447.440 1700.270 ;
        RECT 1447.780 1473.550 1447.920 1700.270 ;
        RECT 1447.720 1473.230 1447.980 1473.550 ;
        RECT 2376.920 1473.230 2377.180 1473.550 ;
        RECT 2376.980 17.670 2377.120 1473.230 ;
        RECT 2376.920 17.350 2377.180 17.670 ;
        RECT 2893.040 16.670 2893.300 16.990 ;
        RECT 2893.100 2.400 2893.240 16.670 ;
        RECT 2892.890 -4.800 2893.450 2.400 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1449.070 1683.920 1449.390 1683.980 ;
        RECT 1455.510 1683.920 1455.830 1683.980 ;
        RECT 1449.070 1683.780 1455.830 1683.920 ;
        RECT 1449.070 1683.720 1449.390 1683.780 ;
        RECT 1455.510 1683.720 1455.830 1683.780 ;
        RECT 1455.510 1280.000 1455.830 1280.060 ;
        RECT 2356.190 1280.000 2356.510 1280.060 ;
        RECT 1455.510 1279.860 2356.510 1280.000 ;
        RECT 1455.510 1279.800 1455.830 1279.860 ;
        RECT 2356.190 1279.800 2356.510 1279.860 ;
        RECT 2356.190 17.240 2356.510 17.300 ;
        RECT 2910.950 17.240 2911.270 17.300 ;
        RECT 2356.190 17.100 2911.270 17.240 ;
        RECT 2356.190 17.040 2356.510 17.100 ;
        RECT 2910.950 17.040 2911.270 17.100 ;
      LAYER via ;
        RECT 1449.100 1683.720 1449.360 1683.980 ;
        RECT 1455.540 1683.720 1455.800 1683.980 ;
        RECT 1455.540 1279.800 1455.800 1280.060 ;
        RECT 2356.220 1279.800 2356.480 1280.060 ;
        RECT 2356.220 17.040 2356.480 17.300 ;
        RECT 2910.980 17.040 2911.240 17.300 ;
      LAYER met2 ;
        RECT 1449.000 1700.340 1449.280 1704.000 ;
        RECT 1449.000 1700.000 1449.300 1700.340 ;
        RECT 1449.160 1684.010 1449.300 1700.000 ;
        RECT 1449.100 1683.690 1449.360 1684.010 ;
        RECT 1455.540 1683.690 1455.800 1684.010 ;
        RECT 1455.600 1280.090 1455.740 1683.690 ;
        RECT 1455.540 1279.770 1455.800 1280.090 ;
        RECT 2356.220 1279.770 2356.480 1280.090 ;
        RECT 2356.280 17.330 2356.420 1279.770 ;
        RECT 2356.220 17.010 2356.480 17.330 ;
        RECT 2910.980 17.010 2911.240 17.330 ;
        RECT 2911.040 2.400 2911.180 17.010 ;
        RECT 2910.830 -4.800 2911.390 2.400 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1237.010 1678.140 1237.330 1678.200 ;
        RECT 1237.930 1678.140 1238.250 1678.200 ;
        RECT 1237.010 1678.000 1238.250 1678.140 ;
        RECT 1237.010 1677.940 1237.330 1678.000 ;
        RECT 1237.930 1677.940 1238.250 1678.000 ;
        RECT 858.890 38.660 859.210 38.720 ;
        RECT 1237.010 38.660 1237.330 38.720 ;
        RECT 858.890 38.520 1237.330 38.660 ;
        RECT 858.890 38.460 859.210 38.520 ;
        RECT 1237.010 38.460 1237.330 38.520 ;
      LAYER via ;
        RECT 1237.040 1677.940 1237.300 1678.200 ;
        RECT 1237.960 1677.940 1238.220 1678.200 ;
        RECT 858.920 38.460 859.180 38.720 ;
        RECT 1237.040 38.460 1237.300 38.720 ;
      LAYER met2 ;
        RECT 1237.860 1700.340 1238.140 1704.000 ;
        RECT 1237.860 1700.000 1238.160 1700.340 ;
        RECT 1238.020 1678.230 1238.160 1700.000 ;
        RECT 1237.040 1677.910 1237.300 1678.230 ;
        RECT 1237.960 1677.910 1238.220 1678.230 ;
        RECT 1237.100 38.750 1237.240 1677.910 ;
        RECT 858.920 38.430 859.180 38.750 ;
        RECT 1237.040 38.430 1237.300 38.750 ;
        RECT 858.980 2.400 859.120 38.430 ;
        RECT 858.770 -4.800 859.330 2.400 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 876.830 39.000 877.150 39.060 ;
        RECT 1239.770 39.000 1240.090 39.060 ;
        RECT 876.830 38.860 1240.090 39.000 ;
        RECT 876.830 38.800 877.150 38.860 ;
        RECT 1239.770 38.800 1240.090 38.860 ;
      LAYER via ;
        RECT 876.860 38.800 877.120 39.060 ;
        RECT 1239.800 38.800 1240.060 39.060 ;
      LAYER met2 ;
        RECT 1239.700 1700.340 1239.980 1704.000 ;
        RECT 1239.700 1700.000 1240.000 1700.340 ;
        RECT 1239.860 39.090 1240.000 1700.000 ;
        RECT 876.860 38.770 877.120 39.090 ;
        RECT 1239.800 38.770 1240.060 39.090 ;
        RECT 876.920 2.400 877.060 38.770 ;
        RECT 876.710 -4.800 877.270 2.400 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 894.770 39.340 895.090 39.400 ;
        RECT 1241.610 39.340 1241.930 39.400 ;
        RECT 894.770 39.200 1241.930 39.340 ;
        RECT 894.770 39.140 895.090 39.200 ;
        RECT 1241.610 39.140 1241.930 39.200 ;
      LAYER via ;
        RECT 894.800 39.140 895.060 39.400 ;
        RECT 1241.640 39.140 1241.900 39.400 ;
      LAYER met2 ;
        RECT 1241.540 1700.340 1241.820 1704.000 ;
        RECT 1241.540 1700.000 1241.840 1700.340 ;
        RECT 1241.700 39.430 1241.840 1700.000 ;
        RECT 894.800 39.110 895.060 39.430 ;
        RECT 1241.640 39.110 1241.900 39.430 ;
        RECT 894.860 2.400 895.000 39.110 ;
        RECT 894.650 -4.800 895.210 2.400 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1243.525 1642.285 1243.695 1680.535 ;
        RECT 1245.825 1545.725 1245.995 1593.835 ;
        RECT 1245.825 386.325 1245.995 434.775 ;
      LAYER mcon ;
        RECT 1243.525 1680.365 1243.695 1680.535 ;
        RECT 1245.825 1593.665 1245.995 1593.835 ;
        RECT 1245.825 434.605 1245.995 434.775 ;
      LAYER met1 ;
        RECT 1243.450 1680.520 1243.770 1680.580 ;
        RECT 1243.255 1680.380 1243.770 1680.520 ;
        RECT 1243.450 1680.320 1243.770 1680.380 ;
        RECT 1243.465 1642.440 1243.755 1642.485 ;
        RECT 1245.750 1642.440 1246.070 1642.500 ;
        RECT 1243.465 1642.300 1246.070 1642.440 ;
        RECT 1243.465 1642.255 1243.755 1642.300 ;
        RECT 1245.750 1642.240 1246.070 1642.300 ;
        RECT 1245.750 1593.820 1246.070 1593.880 ;
        RECT 1245.555 1593.680 1246.070 1593.820 ;
        RECT 1245.750 1593.620 1246.070 1593.680 ;
        RECT 1245.750 1545.880 1246.070 1545.940 ;
        RECT 1245.555 1545.740 1246.070 1545.880 ;
        RECT 1245.750 1545.680 1246.070 1545.740 ;
        RECT 1245.750 530.780 1246.070 531.040 ;
        RECT 1245.840 530.360 1245.980 530.780 ;
        RECT 1245.750 530.100 1246.070 530.360 ;
        RECT 1245.750 434.760 1246.070 434.820 ;
        RECT 1245.555 434.620 1246.070 434.760 ;
        RECT 1245.750 434.560 1246.070 434.620 ;
        RECT 1245.750 386.480 1246.070 386.540 ;
        RECT 1245.555 386.340 1246.070 386.480 ;
        RECT 1245.750 386.280 1246.070 386.340 ;
        RECT 1245.750 193.360 1246.070 193.420 ;
        RECT 1246.210 193.360 1246.530 193.420 ;
        RECT 1245.750 193.220 1246.530 193.360 ;
        RECT 1245.750 193.160 1246.070 193.220 ;
        RECT 1246.210 193.160 1246.530 193.220 ;
        RECT 912.710 39.680 913.030 39.740 ;
        RECT 1245.750 39.680 1246.070 39.740 ;
        RECT 912.710 39.540 1246.070 39.680 ;
        RECT 912.710 39.480 913.030 39.540 ;
        RECT 1245.750 39.480 1246.070 39.540 ;
      LAYER via ;
        RECT 1243.480 1680.320 1243.740 1680.580 ;
        RECT 1245.780 1642.240 1246.040 1642.500 ;
        RECT 1245.780 1593.620 1246.040 1593.880 ;
        RECT 1245.780 1545.680 1246.040 1545.940 ;
        RECT 1245.780 530.780 1246.040 531.040 ;
        RECT 1245.780 530.100 1246.040 530.360 ;
        RECT 1245.780 434.560 1246.040 434.820 ;
        RECT 1245.780 386.280 1246.040 386.540 ;
        RECT 1245.780 193.160 1246.040 193.420 ;
        RECT 1246.240 193.160 1246.500 193.420 ;
        RECT 912.740 39.480 913.000 39.740 ;
        RECT 1245.780 39.480 1246.040 39.740 ;
      LAYER met2 ;
        RECT 1243.380 1700.340 1243.660 1704.000 ;
        RECT 1243.380 1700.000 1243.680 1700.340 ;
        RECT 1243.540 1680.610 1243.680 1700.000 ;
        RECT 1243.480 1680.290 1243.740 1680.610 ;
        RECT 1245.780 1642.210 1246.040 1642.530 ;
        RECT 1245.840 1593.910 1245.980 1642.210 ;
        RECT 1245.780 1593.590 1246.040 1593.910 ;
        RECT 1245.780 1545.650 1246.040 1545.970 ;
        RECT 1245.840 531.070 1245.980 1545.650 ;
        RECT 1245.780 530.750 1246.040 531.070 ;
        RECT 1245.780 530.070 1246.040 530.390 ;
        RECT 1245.840 434.850 1245.980 530.070 ;
        RECT 1245.780 434.530 1246.040 434.850 ;
        RECT 1245.780 386.250 1246.040 386.570 ;
        RECT 1245.840 241.130 1245.980 386.250 ;
        RECT 1245.840 240.990 1246.440 241.130 ;
        RECT 1246.300 193.450 1246.440 240.990 ;
        RECT 1245.780 193.130 1246.040 193.450 ;
        RECT 1246.240 193.130 1246.500 193.450 ;
        RECT 1245.840 39.770 1245.980 193.130 ;
        RECT 912.740 39.450 913.000 39.770 ;
        RECT 1245.780 39.450 1246.040 39.770 ;
        RECT 912.800 2.400 912.940 39.450 ;
        RECT 912.590 -4.800 913.150 2.400 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1244.905 489.005 1245.075 530.995 ;
        RECT 1244.905 392.105 1245.075 434.435 ;
      LAYER mcon ;
        RECT 1244.905 530.825 1245.075 530.995 ;
        RECT 1244.905 434.265 1245.075 434.435 ;
      LAYER met1 ;
        RECT 1244.830 530.980 1245.150 531.040 ;
        RECT 1244.635 530.840 1245.150 530.980 ;
        RECT 1244.830 530.780 1245.150 530.840 ;
        RECT 1244.830 489.160 1245.150 489.220 ;
        RECT 1244.635 489.020 1245.150 489.160 ;
        RECT 1244.830 488.960 1245.150 489.020 ;
        RECT 1244.830 434.420 1245.150 434.480 ;
        RECT 1244.635 434.280 1245.150 434.420 ;
        RECT 1244.830 434.220 1245.150 434.280 ;
        RECT 1244.830 392.260 1245.150 392.320 ;
        RECT 1244.635 392.120 1245.150 392.260 ;
        RECT 1244.830 392.060 1245.150 392.120 ;
        RECT 930.190 40.020 930.510 40.080 ;
        RECT 1244.830 40.020 1245.150 40.080 ;
        RECT 930.190 39.880 1245.150 40.020 ;
        RECT 930.190 39.820 930.510 39.880 ;
        RECT 1244.830 39.820 1245.150 39.880 ;
      LAYER via ;
        RECT 1244.860 530.780 1245.120 531.040 ;
        RECT 1244.860 488.960 1245.120 489.220 ;
        RECT 1244.860 434.220 1245.120 434.480 ;
        RECT 1244.860 392.060 1245.120 392.320 ;
        RECT 930.220 39.820 930.480 40.080 ;
        RECT 1244.860 39.820 1245.120 40.080 ;
      LAYER met2 ;
        RECT 1245.220 1700.340 1245.500 1704.000 ;
        RECT 1245.220 1700.000 1245.520 1700.340 ;
        RECT 1245.380 1668.450 1245.520 1700.000 ;
        RECT 1244.920 1668.310 1245.520 1668.450 ;
        RECT 1244.920 531.070 1245.060 1668.310 ;
        RECT 1244.860 530.750 1245.120 531.070 ;
        RECT 1244.860 488.930 1245.120 489.250 ;
        RECT 1244.920 434.510 1245.060 488.930 ;
        RECT 1244.860 434.190 1245.120 434.510 ;
        RECT 1244.860 392.030 1245.120 392.350 ;
        RECT 1244.920 40.110 1245.060 392.030 ;
        RECT 930.220 39.790 930.480 40.110 ;
        RECT 1244.860 39.790 1245.120 40.110 ;
        RECT 930.280 2.400 930.420 39.790 ;
        RECT 930.070 -4.800 930.630 2.400 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1245.290 1645.160 1245.610 1645.220 ;
        RECT 1247.130 1645.160 1247.450 1645.220 ;
        RECT 1245.290 1645.020 1247.450 1645.160 ;
        RECT 1245.290 1644.960 1245.610 1645.020 ;
        RECT 1247.130 1644.960 1247.450 1645.020 ;
        RECT 1245.290 531.120 1245.610 531.380 ;
        RECT 1245.380 530.700 1245.520 531.120 ;
        RECT 1245.290 530.440 1245.610 530.700 ;
        RECT 1245.290 434.220 1245.610 434.480 ;
        RECT 1245.380 433.800 1245.520 434.220 ;
        RECT 1245.290 433.540 1245.610 433.800 ;
        RECT 948.130 40.360 948.450 40.420 ;
        RECT 1245.290 40.360 1245.610 40.420 ;
        RECT 948.130 40.220 1245.610 40.360 ;
        RECT 948.130 40.160 948.450 40.220 ;
        RECT 1245.290 40.160 1245.610 40.220 ;
      LAYER via ;
        RECT 1245.320 1644.960 1245.580 1645.220 ;
        RECT 1247.160 1644.960 1247.420 1645.220 ;
        RECT 1245.320 531.120 1245.580 531.380 ;
        RECT 1245.320 530.440 1245.580 530.700 ;
        RECT 1245.320 434.220 1245.580 434.480 ;
        RECT 1245.320 433.540 1245.580 433.800 ;
        RECT 948.160 40.160 948.420 40.420 ;
        RECT 1245.320 40.160 1245.580 40.420 ;
      LAYER met2 ;
        RECT 1247.060 1700.340 1247.340 1704.000 ;
        RECT 1247.060 1700.000 1247.360 1700.340 ;
        RECT 1247.220 1645.250 1247.360 1700.000 ;
        RECT 1245.320 1644.930 1245.580 1645.250 ;
        RECT 1247.160 1644.930 1247.420 1645.250 ;
        RECT 1245.380 531.410 1245.520 1644.930 ;
        RECT 1245.320 531.090 1245.580 531.410 ;
        RECT 1245.320 530.410 1245.580 530.730 ;
        RECT 1245.380 434.510 1245.520 530.410 ;
        RECT 1245.320 434.190 1245.580 434.510 ;
        RECT 1245.320 433.510 1245.580 433.830 ;
        RECT 1245.380 40.450 1245.520 433.510 ;
        RECT 948.160 40.130 948.420 40.450 ;
        RECT 1245.320 40.130 1245.580 40.450 ;
        RECT 948.220 2.400 948.360 40.130 ;
        RECT 948.010 -4.800 948.570 2.400 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1248.970 1677.460 1249.290 1677.520 ;
        RECT 1250.350 1677.460 1250.670 1677.520 ;
        RECT 1248.970 1677.320 1250.670 1677.460 ;
        RECT 1248.970 1677.260 1249.290 1677.320 ;
        RECT 1250.350 1677.260 1250.670 1677.320 ;
        RECT 966.070 40.700 966.390 40.760 ;
        RECT 1250.350 40.700 1250.670 40.760 ;
        RECT 966.070 40.560 1250.670 40.700 ;
        RECT 966.070 40.500 966.390 40.560 ;
        RECT 1250.350 40.500 1250.670 40.560 ;
      LAYER via ;
        RECT 1249.000 1677.260 1249.260 1677.520 ;
        RECT 1250.380 1677.260 1250.640 1677.520 ;
        RECT 966.100 40.500 966.360 40.760 ;
        RECT 1250.380 40.500 1250.640 40.760 ;
      LAYER met2 ;
        RECT 1248.900 1700.340 1249.180 1704.000 ;
        RECT 1248.900 1700.000 1249.200 1700.340 ;
        RECT 1249.060 1677.550 1249.200 1700.000 ;
        RECT 1249.000 1677.230 1249.260 1677.550 ;
        RECT 1250.380 1677.230 1250.640 1677.550 ;
        RECT 1250.440 40.790 1250.580 1677.230 ;
        RECT 966.100 40.470 966.360 40.790 ;
        RECT 1250.380 40.470 1250.640 40.790 ;
        RECT 966.160 2.400 966.300 40.470 ;
        RECT 965.950 -4.800 966.510 2.400 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1250.810 1678.480 1251.130 1678.540 ;
        RECT 1253.570 1678.480 1253.890 1678.540 ;
        RECT 1250.810 1678.340 1253.890 1678.480 ;
        RECT 1250.810 1678.280 1251.130 1678.340 ;
        RECT 1253.570 1678.280 1253.890 1678.340 ;
        RECT 984.010 41.040 984.330 41.100 ;
        RECT 1253.570 41.040 1253.890 41.100 ;
        RECT 984.010 40.900 1253.890 41.040 ;
        RECT 984.010 40.840 984.330 40.900 ;
        RECT 1253.570 40.840 1253.890 40.900 ;
      LAYER via ;
        RECT 1250.840 1678.280 1251.100 1678.540 ;
        RECT 1253.600 1678.280 1253.860 1678.540 ;
        RECT 984.040 40.840 984.300 41.100 ;
        RECT 1253.600 40.840 1253.860 41.100 ;
      LAYER met2 ;
        RECT 1250.740 1700.340 1251.020 1704.000 ;
        RECT 1250.740 1700.000 1251.040 1700.340 ;
        RECT 1250.900 1678.570 1251.040 1700.000 ;
        RECT 1250.840 1678.250 1251.100 1678.570 ;
        RECT 1253.600 1678.250 1253.860 1678.570 ;
        RECT 1253.660 41.130 1253.800 1678.250 ;
        RECT 984.040 40.810 984.300 41.130 ;
        RECT 1253.600 40.810 1253.860 41.130 ;
        RECT 984.100 2.400 984.240 40.810 ;
        RECT 983.890 -4.800 984.450 2.400 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1217.305 1400.885 1217.475 1448.995 ;
        RECT 1217.305 1283.585 1217.475 1393.575 ;
        RECT 1217.305 1200.965 1217.475 1276.275 ;
        RECT 1217.305 1097.265 1217.475 1186.855 ;
        RECT 1217.305 1014.305 1217.475 1096.755 ;
        RECT 1216.845 931.345 1217.015 959.055 ;
        RECT 1217.305 871.845 1217.475 910.435 ;
        RECT 1217.305 766.445 1217.475 787.015 ;
        RECT 1217.305 620.925 1217.475 710.515 ;
        RECT 1217.765 544.765 1217.935 594.575 ;
        RECT 1217.765 386.325 1217.935 434.775 ;
        RECT 1217.305 138.125 1217.475 241.315 ;
        RECT 1217.305 110.245 1217.475 137.615 ;
      LAYER mcon ;
        RECT 1217.305 1448.825 1217.475 1448.995 ;
        RECT 1217.305 1393.405 1217.475 1393.575 ;
        RECT 1217.305 1276.105 1217.475 1276.275 ;
        RECT 1217.305 1186.685 1217.475 1186.855 ;
        RECT 1217.305 1096.585 1217.475 1096.755 ;
        RECT 1216.845 958.885 1217.015 959.055 ;
        RECT 1217.305 910.265 1217.475 910.435 ;
        RECT 1217.305 786.845 1217.475 787.015 ;
        RECT 1217.305 710.345 1217.475 710.515 ;
        RECT 1217.765 594.405 1217.935 594.575 ;
        RECT 1217.765 434.605 1217.935 434.775 ;
        RECT 1217.305 241.145 1217.475 241.315 ;
        RECT 1217.305 137.445 1217.475 137.615 ;
      LAYER met1 ;
        RECT 1216.770 1594.160 1217.090 1594.220 ;
        RECT 1217.690 1594.160 1218.010 1594.220 ;
        RECT 1216.770 1594.020 1218.010 1594.160 ;
        RECT 1216.770 1593.960 1217.090 1594.020 ;
        RECT 1217.690 1593.960 1218.010 1594.020 ;
        RECT 1216.770 1545.880 1217.090 1545.940 ;
        RECT 1217.690 1545.880 1218.010 1545.940 ;
        RECT 1216.770 1545.740 1218.010 1545.880 ;
        RECT 1216.770 1545.680 1217.090 1545.740 ;
        RECT 1217.690 1545.680 1218.010 1545.740 ;
        RECT 1217.230 1448.980 1217.550 1449.040 ;
        RECT 1217.035 1448.840 1217.550 1448.980 ;
        RECT 1217.230 1448.780 1217.550 1448.840 ;
        RECT 1217.245 1401.040 1217.535 1401.085 ;
        RECT 1217.690 1401.040 1218.010 1401.100 ;
        RECT 1217.245 1400.900 1218.010 1401.040 ;
        RECT 1217.245 1400.855 1217.535 1400.900 ;
        RECT 1217.690 1400.840 1218.010 1400.900 ;
        RECT 1217.245 1393.560 1217.535 1393.605 ;
        RECT 1217.690 1393.560 1218.010 1393.620 ;
        RECT 1217.245 1393.420 1218.010 1393.560 ;
        RECT 1217.245 1393.375 1217.535 1393.420 ;
        RECT 1217.690 1393.360 1218.010 1393.420 ;
        RECT 1217.245 1283.740 1217.535 1283.785 ;
        RECT 1217.690 1283.740 1218.010 1283.800 ;
        RECT 1217.245 1283.600 1218.010 1283.740 ;
        RECT 1217.245 1283.555 1217.535 1283.600 ;
        RECT 1217.690 1283.540 1218.010 1283.600 ;
        RECT 1217.245 1276.260 1217.535 1276.305 ;
        RECT 1217.690 1276.260 1218.010 1276.320 ;
        RECT 1217.245 1276.120 1218.010 1276.260 ;
        RECT 1217.245 1276.075 1217.535 1276.120 ;
        RECT 1217.690 1276.060 1218.010 1276.120 ;
        RECT 1217.245 1201.120 1217.535 1201.165 ;
        RECT 1217.690 1201.120 1218.010 1201.180 ;
        RECT 1217.245 1200.980 1218.010 1201.120 ;
        RECT 1217.245 1200.935 1217.535 1200.980 ;
        RECT 1217.690 1200.920 1218.010 1200.980 ;
        RECT 1217.245 1186.840 1217.535 1186.885 ;
        RECT 1217.690 1186.840 1218.010 1186.900 ;
        RECT 1217.245 1186.700 1218.010 1186.840 ;
        RECT 1217.245 1186.655 1217.535 1186.700 ;
        RECT 1217.690 1186.640 1218.010 1186.700 ;
        RECT 1217.230 1097.420 1217.550 1097.480 ;
        RECT 1217.035 1097.280 1217.550 1097.420 ;
        RECT 1217.230 1097.220 1217.550 1097.280 ;
        RECT 1217.230 1096.740 1217.550 1096.800 ;
        RECT 1217.035 1096.600 1217.550 1096.740 ;
        RECT 1217.230 1096.540 1217.550 1096.600 ;
        RECT 1217.245 1014.460 1217.535 1014.505 ;
        RECT 1217.690 1014.460 1218.010 1014.520 ;
        RECT 1217.245 1014.320 1218.010 1014.460 ;
        RECT 1217.245 1014.275 1217.535 1014.320 ;
        RECT 1217.690 1014.260 1218.010 1014.320 ;
        RECT 1216.770 959.040 1217.090 959.100 ;
        RECT 1216.575 958.900 1217.090 959.040 ;
        RECT 1216.770 958.840 1217.090 958.900 ;
        RECT 1216.785 931.500 1217.075 931.545 ;
        RECT 1217.230 931.500 1217.550 931.560 ;
        RECT 1216.785 931.360 1217.550 931.500 ;
        RECT 1216.785 931.315 1217.075 931.360 ;
        RECT 1217.230 931.300 1217.550 931.360 ;
        RECT 1217.245 910.420 1217.535 910.465 ;
        RECT 1217.690 910.420 1218.010 910.480 ;
        RECT 1217.245 910.280 1218.010 910.420 ;
        RECT 1217.245 910.235 1217.535 910.280 ;
        RECT 1217.690 910.220 1218.010 910.280 ;
        RECT 1217.230 872.000 1217.550 872.060 ;
        RECT 1217.035 871.860 1217.550 872.000 ;
        RECT 1217.230 871.800 1217.550 871.860 ;
        RECT 1217.230 835.080 1217.550 835.340 ;
        RECT 1217.320 834.600 1217.460 835.080 ;
        RECT 1217.690 834.600 1218.010 834.660 ;
        RECT 1217.320 834.460 1218.010 834.600 ;
        RECT 1217.690 834.400 1218.010 834.460 ;
        RECT 1217.245 787.000 1217.535 787.045 ;
        RECT 1217.690 787.000 1218.010 787.060 ;
        RECT 1217.245 786.860 1218.010 787.000 ;
        RECT 1217.245 786.815 1217.535 786.860 ;
        RECT 1217.690 786.800 1218.010 786.860 ;
        RECT 1217.230 766.600 1217.550 766.660 ;
        RECT 1217.035 766.460 1217.550 766.600 ;
        RECT 1217.230 766.400 1217.550 766.460 ;
        RECT 1217.230 738.520 1217.550 738.780 ;
        RECT 1217.320 738.100 1217.460 738.520 ;
        RECT 1217.230 737.840 1217.550 738.100 ;
        RECT 1217.245 710.500 1217.535 710.545 ;
        RECT 1217.690 710.500 1218.010 710.560 ;
        RECT 1217.245 710.360 1218.010 710.500 ;
        RECT 1217.245 710.315 1217.535 710.360 ;
        RECT 1217.690 710.300 1218.010 710.360 ;
        RECT 1217.230 621.080 1217.550 621.140 ;
        RECT 1217.035 620.940 1217.550 621.080 ;
        RECT 1217.230 620.880 1217.550 620.940 ;
        RECT 1217.230 594.560 1217.550 594.620 ;
        RECT 1217.705 594.560 1217.995 594.605 ;
        RECT 1217.230 594.420 1217.995 594.560 ;
        RECT 1217.230 594.360 1217.550 594.420 ;
        RECT 1217.705 594.375 1217.995 594.420 ;
        RECT 1217.690 544.920 1218.010 544.980 ;
        RECT 1217.495 544.780 1218.010 544.920 ;
        RECT 1217.690 544.720 1218.010 544.780 ;
        RECT 1217.690 506.980 1218.010 507.240 ;
        RECT 1217.780 506.560 1217.920 506.980 ;
        RECT 1217.690 506.300 1218.010 506.560 ;
        RECT 1217.690 434.760 1218.010 434.820 ;
        RECT 1217.495 434.620 1218.010 434.760 ;
        RECT 1217.690 434.560 1218.010 434.620 ;
        RECT 1217.690 386.480 1218.010 386.540 ;
        RECT 1217.495 386.340 1218.010 386.480 ;
        RECT 1217.690 386.280 1218.010 386.340 ;
        RECT 1217.230 255.720 1217.550 255.980 ;
        RECT 1217.320 255.300 1217.460 255.720 ;
        RECT 1217.230 255.040 1217.550 255.300 ;
        RECT 1217.245 241.300 1217.535 241.345 ;
        RECT 1217.690 241.300 1218.010 241.360 ;
        RECT 1217.245 241.160 1218.010 241.300 ;
        RECT 1217.245 241.115 1217.535 241.160 ;
        RECT 1217.690 241.100 1218.010 241.160 ;
        RECT 1217.245 138.280 1217.535 138.325 ;
        RECT 1217.690 138.280 1218.010 138.340 ;
        RECT 1217.245 138.140 1218.010 138.280 ;
        RECT 1217.245 138.095 1217.535 138.140 ;
        RECT 1217.690 138.080 1218.010 138.140 ;
        RECT 1217.245 137.600 1217.535 137.645 ;
        RECT 1217.690 137.600 1218.010 137.660 ;
        RECT 1217.245 137.460 1218.010 137.600 ;
        RECT 1217.245 137.415 1217.535 137.460 ;
        RECT 1217.690 137.400 1218.010 137.460 ;
        RECT 1217.230 110.400 1217.550 110.460 ;
        RECT 1217.035 110.260 1217.550 110.400 ;
        RECT 1217.230 110.200 1217.550 110.260 ;
        RECT 1217.230 62.460 1217.550 62.520 ;
        RECT 1216.860 62.320 1217.550 62.460 ;
        RECT 1216.860 62.180 1217.000 62.320 ;
        RECT 1217.230 62.260 1217.550 62.320 ;
        RECT 1216.770 61.920 1217.090 62.180 ;
        RECT 662.930 37.980 663.250 38.040 ;
        RECT 1216.770 37.980 1217.090 38.040 ;
        RECT 662.930 37.840 1217.090 37.980 ;
        RECT 662.930 37.780 663.250 37.840 ;
        RECT 1216.770 37.780 1217.090 37.840 ;
      LAYER via ;
        RECT 1216.800 1593.960 1217.060 1594.220 ;
        RECT 1217.720 1593.960 1217.980 1594.220 ;
        RECT 1216.800 1545.680 1217.060 1545.940 ;
        RECT 1217.720 1545.680 1217.980 1545.940 ;
        RECT 1217.260 1448.780 1217.520 1449.040 ;
        RECT 1217.720 1400.840 1217.980 1401.100 ;
        RECT 1217.720 1393.360 1217.980 1393.620 ;
        RECT 1217.720 1283.540 1217.980 1283.800 ;
        RECT 1217.720 1276.060 1217.980 1276.320 ;
        RECT 1217.720 1200.920 1217.980 1201.180 ;
        RECT 1217.720 1186.640 1217.980 1186.900 ;
        RECT 1217.260 1097.220 1217.520 1097.480 ;
        RECT 1217.260 1096.540 1217.520 1096.800 ;
        RECT 1217.720 1014.260 1217.980 1014.520 ;
        RECT 1216.800 958.840 1217.060 959.100 ;
        RECT 1217.260 931.300 1217.520 931.560 ;
        RECT 1217.720 910.220 1217.980 910.480 ;
        RECT 1217.260 871.800 1217.520 872.060 ;
        RECT 1217.260 835.080 1217.520 835.340 ;
        RECT 1217.720 834.400 1217.980 834.660 ;
        RECT 1217.720 786.800 1217.980 787.060 ;
        RECT 1217.260 766.400 1217.520 766.660 ;
        RECT 1217.260 738.520 1217.520 738.780 ;
        RECT 1217.260 737.840 1217.520 738.100 ;
        RECT 1217.720 710.300 1217.980 710.560 ;
        RECT 1217.260 620.880 1217.520 621.140 ;
        RECT 1217.260 594.360 1217.520 594.620 ;
        RECT 1217.720 544.720 1217.980 544.980 ;
        RECT 1217.720 506.980 1217.980 507.240 ;
        RECT 1217.720 506.300 1217.980 506.560 ;
        RECT 1217.720 434.560 1217.980 434.820 ;
        RECT 1217.720 386.280 1217.980 386.540 ;
        RECT 1217.260 255.720 1217.520 255.980 ;
        RECT 1217.260 255.040 1217.520 255.300 ;
        RECT 1217.720 241.100 1217.980 241.360 ;
        RECT 1217.720 138.080 1217.980 138.340 ;
        RECT 1217.720 137.400 1217.980 137.660 ;
        RECT 1217.260 110.200 1217.520 110.460 ;
        RECT 1217.260 62.260 1217.520 62.520 ;
        RECT 1216.800 61.920 1217.060 62.180 ;
        RECT 662.960 37.780 663.220 38.040 ;
        RECT 1216.800 37.780 1217.060 38.040 ;
      LAYER met2 ;
        RECT 1217.620 1700.340 1217.900 1704.000 ;
        RECT 1217.620 1700.000 1217.920 1700.340 ;
        RECT 1217.780 1594.250 1217.920 1700.000 ;
        RECT 1216.800 1593.930 1217.060 1594.250 ;
        RECT 1217.720 1593.930 1217.980 1594.250 ;
        RECT 1216.860 1545.970 1217.000 1593.930 ;
        RECT 1216.800 1545.650 1217.060 1545.970 ;
        RECT 1217.720 1545.650 1217.980 1545.970 ;
        RECT 1217.780 1463.090 1217.920 1545.650 ;
        RECT 1217.320 1462.950 1217.920 1463.090 ;
        RECT 1217.320 1449.070 1217.460 1462.950 ;
        RECT 1217.260 1448.750 1217.520 1449.070 ;
        RECT 1217.720 1400.810 1217.980 1401.130 ;
        RECT 1217.780 1393.650 1217.920 1400.810 ;
        RECT 1217.720 1393.330 1217.980 1393.650 ;
        RECT 1217.720 1283.510 1217.980 1283.830 ;
        RECT 1217.780 1276.350 1217.920 1283.510 ;
        RECT 1217.720 1276.030 1217.980 1276.350 ;
        RECT 1217.720 1200.890 1217.980 1201.210 ;
        RECT 1217.780 1186.930 1217.920 1200.890 ;
        RECT 1217.720 1186.610 1217.980 1186.930 ;
        RECT 1217.260 1097.190 1217.520 1097.510 ;
        RECT 1217.320 1096.830 1217.460 1097.190 ;
        RECT 1217.260 1096.510 1217.520 1096.830 ;
        RECT 1217.720 1014.230 1217.980 1014.550 ;
        RECT 1217.780 983.010 1217.920 1014.230 ;
        RECT 1216.860 982.870 1217.920 983.010 ;
        RECT 1216.860 959.130 1217.000 982.870 ;
        RECT 1216.800 958.810 1217.060 959.130 ;
        RECT 1217.260 931.270 1217.520 931.590 ;
        RECT 1217.320 910.930 1217.460 931.270 ;
        RECT 1217.320 910.790 1217.920 910.930 ;
        RECT 1217.780 910.510 1217.920 910.790 ;
        RECT 1217.720 910.190 1217.980 910.510 ;
        RECT 1217.260 871.770 1217.520 872.090 ;
        RECT 1217.320 835.370 1217.460 871.770 ;
        RECT 1217.260 835.050 1217.520 835.370 ;
        RECT 1217.720 834.370 1217.980 834.690 ;
        RECT 1217.780 787.090 1217.920 834.370 ;
        RECT 1217.720 786.770 1217.980 787.090 ;
        RECT 1217.260 766.370 1217.520 766.690 ;
        RECT 1217.320 738.810 1217.460 766.370 ;
        RECT 1217.260 738.490 1217.520 738.810 ;
        RECT 1217.260 737.810 1217.520 738.130 ;
        RECT 1217.320 717.810 1217.460 737.810 ;
        RECT 1217.320 717.670 1217.920 717.810 ;
        RECT 1217.780 710.590 1217.920 717.670 ;
        RECT 1217.720 710.270 1217.980 710.590 ;
        RECT 1217.260 620.850 1217.520 621.170 ;
        RECT 1217.320 594.650 1217.460 620.850 ;
        RECT 1217.260 594.330 1217.520 594.650 ;
        RECT 1217.720 544.690 1217.980 545.010 ;
        RECT 1217.780 507.270 1217.920 544.690 ;
        RECT 1217.720 506.950 1217.980 507.270 ;
        RECT 1217.720 506.270 1217.980 506.590 ;
        RECT 1217.780 434.850 1217.920 506.270 ;
        RECT 1217.720 434.530 1217.980 434.850 ;
        RECT 1217.720 386.250 1217.980 386.570 ;
        RECT 1217.780 303.690 1217.920 386.250 ;
        RECT 1217.320 303.550 1217.920 303.690 ;
        RECT 1217.320 256.010 1217.460 303.550 ;
        RECT 1217.260 255.690 1217.520 256.010 ;
        RECT 1217.260 255.010 1217.520 255.330 ;
        RECT 1217.320 241.810 1217.460 255.010 ;
        RECT 1217.320 241.670 1217.920 241.810 ;
        RECT 1217.780 241.390 1217.920 241.670 ;
        RECT 1217.720 241.070 1217.980 241.390 ;
        RECT 1217.720 138.050 1217.980 138.370 ;
        RECT 1217.780 137.690 1217.920 138.050 ;
        RECT 1217.720 137.370 1217.980 137.690 ;
        RECT 1217.260 110.170 1217.520 110.490 ;
        RECT 1217.320 62.550 1217.460 110.170 ;
        RECT 1217.260 62.230 1217.520 62.550 ;
        RECT 1216.800 61.890 1217.060 62.210 ;
        RECT 1216.860 38.070 1217.000 61.890 ;
        RECT 662.960 37.750 663.220 38.070 ;
        RECT 1216.800 37.750 1217.060 38.070 ;
        RECT 663.020 2.400 663.160 37.750 ;
        RECT 662.810 -4.800 663.370 2.400 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1001.950 41.380 1002.270 41.440 ;
        RECT 1252.650 41.380 1252.970 41.440 ;
        RECT 1001.950 41.240 1252.970 41.380 ;
        RECT 1001.950 41.180 1002.270 41.240 ;
        RECT 1252.650 41.180 1252.970 41.240 ;
      LAYER via ;
        RECT 1001.980 41.180 1002.240 41.440 ;
        RECT 1252.680 41.180 1252.940 41.440 ;
      LAYER met2 ;
        RECT 1252.580 1700.340 1252.860 1704.000 ;
        RECT 1252.580 1700.000 1252.880 1700.340 ;
        RECT 1252.740 41.470 1252.880 1700.000 ;
        RECT 1001.980 41.150 1002.240 41.470 ;
        RECT 1252.680 41.150 1252.940 41.470 ;
        RECT 1002.040 2.400 1002.180 41.150 ;
        RECT 1001.830 -4.800 1002.390 2.400 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1019.430 37.640 1019.750 37.700 ;
        RECT 1254.490 37.640 1254.810 37.700 ;
        RECT 1019.430 37.500 1254.810 37.640 ;
        RECT 1019.430 37.440 1019.750 37.500 ;
        RECT 1254.490 37.440 1254.810 37.500 ;
      LAYER via ;
        RECT 1019.460 37.440 1019.720 37.700 ;
        RECT 1254.520 37.440 1254.780 37.700 ;
      LAYER met2 ;
        RECT 1254.420 1700.340 1254.700 1704.000 ;
        RECT 1254.420 1700.000 1254.720 1700.340 ;
        RECT 1254.580 37.730 1254.720 1700.000 ;
        RECT 1019.460 37.410 1019.720 37.730 ;
        RECT 1254.520 37.410 1254.780 37.730 ;
        RECT 1019.520 2.400 1019.660 37.410 ;
        RECT 1019.310 -4.800 1019.870 2.400 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1227.885 1674.925 1228.055 1678.835 ;
      LAYER mcon ;
        RECT 1227.885 1678.665 1228.055 1678.835 ;
      LAYER met1 ;
        RECT 1227.810 1686.980 1228.130 1687.040 ;
        RECT 1256.330 1686.980 1256.650 1687.040 ;
        RECT 1227.810 1686.840 1256.650 1686.980 ;
        RECT 1227.810 1686.780 1228.130 1686.840 ;
        RECT 1256.330 1686.780 1256.650 1686.840 ;
        RECT 1227.810 1678.820 1228.130 1678.880 ;
        RECT 1227.615 1678.680 1228.130 1678.820 ;
        RECT 1227.810 1678.620 1228.130 1678.680 ;
        RECT 1041.510 1675.080 1041.830 1675.140 ;
        RECT 1227.825 1675.080 1228.115 1675.125 ;
        RECT 1041.510 1674.940 1228.115 1675.080 ;
        RECT 1041.510 1674.880 1041.830 1674.940 ;
        RECT 1227.825 1674.895 1228.115 1674.940 ;
        RECT 1037.370 2.960 1037.690 3.020 ;
        RECT 1041.510 2.960 1041.830 3.020 ;
        RECT 1037.370 2.820 1041.830 2.960 ;
        RECT 1037.370 2.760 1037.690 2.820 ;
        RECT 1041.510 2.760 1041.830 2.820 ;
      LAYER via ;
        RECT 1227.840 1686.780 1228.100 1687.040 ;
        RECT 1256.360 1686.780 1256.620 1687.040 ;
        RECT 1227.840 1678.620 1228.100 1678.880 ;
        RECT 1041.540 1674.880 1041.800 1675.140 ;
        RECT 1037.400 2.760 1037.660 3.020 ;
        RECT 1041.540 2.760 1041.800 3.020 ;
      LAYER met2 ;
        RECT 1256.260 1700.340 1256.540 1704.000 ;
        RECT 1256.260 1700.000 1256.560 1700.340 ;
        RECT 1256.420 1687.070 1256.560 1700.000 ;
        RECT 1227.840 1686.750 1228.100 1687.070 ;
        RECT 1256.360 1686.750 1256.620 1687.070 ;
        RECT 1227.900 1678.910 1228.040 1686.750 ;
        RECT 1227.840 1678.590 1228.100 1678.910 ;
        RECT 1041.540 1674.850 1041.800 1675.170 ;
        RECT 1041.600 3.050 1041.740 1674.850 ;
        RECT 1037.400 2.730 1037.660 3.050 ;
        RECT 1041.540 2.730 1041.800 3.050 ;
        RECT 1037.460 2.400 1037.600 2.730 ;
        RECT 1037.250 -4.800 1037.810 2.400 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1258.170 1678.480 1258.490 1678.540 ;
        RECT 1260.470 1678.480 1260.790 1678.540 ;
        RECT 1258.170 1678.340 1260.790 1678.480 ;
        RECT 1258.170 1678.280 1258.490 1678.340 ;
        RECT 1260.470 1678.280 1260.790 1678.340 ;
        RECT 1260.470 1631.900 1260.790 1631.960 ;
        RECT 1261.390 1631.900 1261.710 1631.960 ;
        RECT 1260.470 1631.760 1261.710 1631.900 ;
        RECT 1260.470 1631.700 1260.790 1631.760 ;
        RECT 1261.390 1631.700 1261.710 1631.760 ;
        RECT 1054.850 1605.380 1055.170 1605.440 ;
        RECT 1261.390 1605.380 1261.710 1605.440 ;
        RECT 1054.850 1605.240 1261.710 1605.380 ;
        RECT 1054.850 1605.180 1055.170 1605.240 ;
        RECT 1261.390 1605.180 1261.710 1605.240 ;
      LAYER via ;
        RECT 1258.200 1678.280 1258.460 1678.540 ;
        RECT 1260.500 1678.280 1260.760 1678.540 ;
        RECT 1260.500 1631.700 1260.760 1631.960 ;
        RECT 1261.420 1631.700 1261.680 1631.960 ;
        RECT 1054.880 1605.180 1055.140 1605.440 ;
        RECT 1261.420 1605.180 1261.680 1605.440 ;
      LAYER met2 ;
        RECT 1258.100 1700.340 1258.380 1704.000 ;
        RECT 1258.100 1700.000 1258.400 1700.340 ;
        RECT 1258.260 1678.570 1258.400 1700.000 ;
        RECT 1258.200 1678.250 1258.460 1678.570 ;
        RECT 1260.500 1678.250 1260.760 1678.570 ;
        RECT 1260.560 1631.990 1260.700 1678.250 ;
        RECT 1260.500 1631.670 1260.760 1631.990 ;
        RECT 1261.420 1631.670 1261.680 1631.990 ;
        RECT 1261.480 1605.470 1261.620 1631.670 ;
        RECT 1054.880 1605.150 1055.140 1605.470 ;
        RECT 1261.420 1605.150 1261.680 1605.470 ;
        RECT 1054.940 17.410 1055.080 1605.150 ;
        RECT 1054.940 17.270 1055.540 17.410 ;
        RECT 1055.400 2.400 1055.540 17.270 ;
        RECT 1055.190 -4.800 1055.750 2.400 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1076.010 1598.240 1076.330 1598.300 ;
        RECT 1258.170 1598.240 1258.490 1598.300 ;
        RECT 1076.010 1598.100 1258.490 1598.240 ;
        RECT 1076.010 1598.040 1076.330 1598.100 ;
        RECT 1258.170 1598.040 1258.490 1598.100 ;
      LAYER via ;
        RECT 1076.040 1598.040 1076.300 1598.300 ;
        RECT 1258.200 1598.040 1258.460 1598.300 ;
      LAYER met2 ;
        RECT 1259.940 1700.340 1260.220 1704.000 ;
        RECT 1259.940 1700.000 1260.240 1700.340 ;
        RECT 1260.100 1678.765 1260.240 1700.000 ;
        RECT 1260.030 1678.395 1260.310 1678.765 ;
        RECT 1258.190 1677.035 1258.470 1677.405 ;
        RECT 1258.260 1598.330 1258.400 1677.035 ;
        RECT 1076.040 1598.010 1076.300 1598.330 ;
        RECT 1258.200 1598.010 1258.460 1598.330 ;
        RECT 1076.100 18.090 1076.240 1598.010 ;
        RECT 1073.340 17.950 1076.240 18.090 ;
        RECT 1073.340 2.400 1073.480 17.950 ;
        RECT 1073.130 -4.800 1073.690 2.400 ;
      LAYER via2 ;
        RECT 1260.030 1678.440 1260.310 1678.720 ;
        RECT 1258.190 1677.080 1258.470 1677.360 ;
      LAYER met3 ;
        RECT 1260.005 1678.730 1260.335 1678.745 ;
        RECT 1259.790 1678.415 1260.335 1678.730 ;
        RECT 1258.165 1677.370 1258.495 1677.385 ;
        RECT 1259.790 1677.370 1260.090 1678.415 ;
        RECT 1258.165 1677.070 1260.090 1677.370 ;
        RECT 1258.165 1677.055 1258.495 1677.070 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1096.250 610.540 1096.570 610.600 ;
        RECT 1260.930 610.540 1261.250 610.600 ;
        RECT 1096.250 610.400 1261.250 610.540 ;
        RECT 1096.250 610.340 1096.570 610.400 ;
        RECT 1260.930 610.340 1261.250 610.400 ;
      LAYER via ;
        RECT 1096.280 610.340 1096.540 610.600 ;
        RECT 1260.960 610.340 1261.220 610.600 ;
      LAYER met2 ;
        RECT 1261.780 1700.340 1262.060 1704.000 ;
        RECT 1261.780 1700.000 1262.080 1700.340 ;
        RECT 1261.940 1677.970 1262.080 1700.000 ;
        RECT 1261.020 1677.830 1262.080 1677.970 ;
        RECT 1261.020 610.630 1261.160 1677.830 ;
        RECT 1096.280 610.310 1096.540 610.630 ;
        RECT 1260.960 610.310 1261.220 610.630 ;
        RECT 1096.340 18.090 1096.480 610.310 ;
        RECT 1090.820 17.950 1096.480 18.090 ;
        RECT 1090.820 2.400 1090.960 17.950 ;
        RECT 1090.610 -4.800 1091.170 2.400 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1110.510 1640.060 1110.830 1640.120 ;
        RECT 1263.690 1640.060 1264.010 1640.120 ;
        RECT 1110.510 1639.920 1264.010 1640.060 ;
        RECT 1110.510 1639.860 1110.830 1639.920 ;
        RECT 1263.690 1639.860 1264.010 1639.920 ;
      LAYER via ;
        RECT 1110.540 1639.860 1110.800 1640.120 ;
        RECT 1263.720 1639.860 1263.980 1640.120 ;
      LAYER met2 ;
        RECT 1263.620 1700.340 1263.900 1704.000 ;
        RECT 1263.620 1700.000 1263.920 1700.340 ;
        RECT 1263.780 1640.150 1263.920 1700.000 ;
        RECT 1110.540 1639.830 1110.800 1640.150 ;
        RECT 1263.720 1639.830 1263.980 1640.150 ;
        RECT 1110.600 16.730 1110.740 1639.830 ;
        RECT 1108.760 16.590 1110.740 16.730 ;
        RECT 1108.760 2.400 1108.900 16.590 ;
        RECT 1108.550 -4.800 1109.110 2.400 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1131.210 1633.260 1131.530 1633.320 ;
        RECT 1265.530 1633.260 1265.850 1633.320 ;
        RECT 1131.210 1633.120 1265.850 1633.260 ;
        RECT 1131.210 1633.060 1131.530 1633.120 ;
        RECT 1265.530 1633.060 1265.850 1633.120 ;
      LAYER via ;
        RECT 1131.240 1633.060 1131.500 1633.320 ;
        RECT 1265.560 1633.060 1265.820 1633.320 ;
      LAYER met2 ;
        RECT 1265.460 1700.340 1265.740 1704.000 ;
        RECT 1265.460 1700.000 1265.760 1700.340 ;
        RECT 1265.620 1633.350 1265.760 1700.000 ;
        RECT 1131.240 1633.030 1131.500 1633.350 ;
        RECT 1265.560 1633.030 1265.820 1633.350 ;
        RECT 1131.300 16.730 1131.440 1633.030 ;
        RECT 1126.700 16.590 1131.440 16.730 ;
        RECT 1126.700 2.400 1126.840 16.590 ;
        RECT 1126.490 -4.800 1127.050 2.400 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1259.550 1683.920 1259.870 1683.980 ;
        RECT 1267.370 1683.920 1267.690 1683.980 ;
        RECT 1259.550 1683.780 1267.690 1683.920 ;
        RECT 1259.550 1683.720 1259.870 1683.780 ;
        RECT 1267.370 1683.720 1267.690 1683.780 ;
        RECT 1144.550 58.720 1144.870 58.780 ;
        RECT 1260.010 58.720 1260.330 58.780 ;
        RECT 1144.550 58.580 1260.330 58.720 ;
        RECT 1144.550 58.520 1144.870 58.580 ;
        RECT 1260.010 58.520 1260.330 58.580 ;
      LAYER via ;
        RECT 1259.580 1683.720 1259.840 1683.980 ;
        RECT 1267.400 1683.720 1267.660 1683.980 ;
        RECT 1144.580 58.520 1144.840 58.780 ;
        RECT 1260.040 58.520 1260.300 58.780 ;
      LAYER met2 ;
        RECT 1267.300 1700.340 1267.580 1704.000 ;
        RECT 1267.300 1700.000 1267.600 1700.340 ;
        RECT 1267.460 1684.010 1267.600 1700.000 ;
        RECT 1259.580 1683.690 1259.840 1684.010 ;
        RECT 1267.400 1683.690 1267.660 1684.010 ;
        RECT 1259.640 1677.970 1259.780 1683.690 ;
        RECT 1259.640 1677.830 1260.240 1677.970 ;
        RECT 1260.100 58.810 1260.240 1677.830 ;
        RECT 1144.580 58.490 1144.840 58.810 ;
        RECT 1260.040 58.490 1260.300 58.810 ;
        RECT 1144.640 2.400 1144.780 58.490 ;
        RECT 1144.430 -4.800 1144.990 2.400 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1264.610 1678.140 1264.930 1678.200 ;
        RECT 1269.210 1678.140 1269.530 1678.200 ;
        RECT 1264.610 1678.000 1269.530 1678.140 ;
        RECT 1264.610 1677.940 1264.930 1678.000 ;
        RECT 1269.210 1677.940 1269.530 1678.000 ;
        RECT 1165.710 51.920 1166.030 51.980 ;
        RECT 1264.610 51.920 1264.930 51.980 ;
        RECT 1165.710 51.780 1264.930 51.920 ;
        RECT 1165.710 51.720 1166.030 51.780 ;
        RECT 1264.610 51.720 1264.930 51.780 ;
        RECT 1162.490 17.580 1162.810 17.640 ;
        RECT 1165.710 17.580 1166.030 17.640 ;
        RECT 1162.490 17.440 1166.030 17.580 ;
        RECT 1162.490 17.380 1162.810 17.440 ;
        RECT 1165.710 17.380 1166.030 17.440 ;
      LAYER via ;
        RECT 1264.640 1677.940 1264.900 1678.200 ;
        RECT 1269.240 1677.940 1269.500 1678.200 ;
        RECT 1165.740 51.720 1166.000 51.980 ;
        RECT 1264.640 51.720 1264.900 51.980 ;
        RECT 1162.520 17.380 1162.780 17.640 ;
        RECT 1165.740 17.380 1166.000 17.640 ;
      LAYER met2 ;
        RECT 1269.140 1700.340 1269.420 1704.000 ;
        RECT 1269.140 1700.000 1269.440 1700.340 ;
        RECT 1269.300 1678.230 1269.440 1700.000 ;
        RECT 1264.640 1677.910 1264.900 1678.230 ;
        RECT 1269.240 1677.910 1269.500 1678.230 ;
        RECT 1264.700 52.010 1264.840 1677.910 ;
        RECT 1165.740 51.690 1166.000 52.010 ;
        RECT 1264.640 51.690 1264.900 52.010 ;
        RECT 1165.800 17.670 1165.940 51.690 ;
        RECT 1162.520 17.350 1162.780 17.670 ;
        RECT 1165.740 17.350 1166.000 17.670 ;
        RECT 1162.580 2.400 1162.720 17.350 ;
        RECT 1162.370 -4.800 1162.930 2.400 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 682.710 1605.040 683.030 1605.100 ;
        RECT 1219.530 1605.040 1219.850 1605.100 ;
        RECT 682.710 1604.900 1219.850 1605.040 ;
        RECT 682.710 1604.840 683.030 1604.900 ;
        RECT 1219.530 1604.840 1219.850 1604.900 ;
      LAYER via ;
        RECT 682.740 1604.840 683.000 1605.100 ;
        RECT 1219.560 1604.840 1219.820 1605.100 ;
      LAYER met2 ;
        RECT 1219.460 1700.340 1219.740 1704.000 ;
        RECT 1219.460 1700.000 1219.760 1700.340 ;
        RECT 1219.620 1605.130 1219.760 1700.000 ;
        RECT 682.740 1604.810 683.000 1605.130 ;
        RECT 1219.560 1604.810 1219.820 1605.130 ;
        RECT 682.800 24.210 682.940 1604.810 ;
        RECT 680.500 24.070 682.940 24.210 ;
        RECT 680.500 2.400 680.640 24.070 ;
        RECT 680.290 -4.800 680.850 2.400 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1265.990 1689.700 1266.310 1689.760 ;
        RECT 1271.050 1689.700 1271.370 1689.760 ;
        RECT 1265.990 1689.560 1271.370 1689.700 ;
        RECT 1265.990 1689.500 1266.310 1689.560 ;
        RECT 1271.050 1689.500 1271.370 1689.560 ;
        RECT 1179.970 52.260 1180.290 52.320 ;
        RECT 1265.990 52.260 1266.310 52.320 ;
        RECT 1179.970 52.120 1266.310 52.260 ;
        RECT 1179.970 52.060 1180.290 52.120 ;
        RECT 1265.990 52.060 1266.310 52.120 ;
      LAYER via ;
        RECT 1266.020 1689.500 1266.280 1689.760 ;
        RECT 1271.080 1689.500 1271.340 1689.760 ;
        RECT 1180.000 52.060 1180.260 52.320 ;
        RECT 1266.020 52.060 1266.280 52.320 ;
      LAYER met2 ;
        RECT 1270.980 1700.340 1271.260 1704.000 ;
        RECT 1270.980 1700.000 1271.280 1700.340 ;
        RECT 1271.140 1689.790 1271.280 1700.000 ;
        RECT 1266.020 1689.470 1266.280 1689.790 ;
        RECT 1271.080 1689.470 1271.340 1689.790 ;
        RECT 1266.080 52.350 1266.220 1689.470 ;
        RECT 1180.000 52.030 1180.260 52.350 ;
        RECT 1266.020 52.030 1266.280 52.350 ;
        RECT 1180.060 2.400 1180.200 52.030 ;
        RECT 1179.850 -4.800 1180.410 2.400 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1269.745 1290.385 1269.915 1304.495 ;
        RECT 1270.205 1151.325 1270.375 1193.655 ;
        RECT 1270.205 662.405 1270.375 710.515 ;
        RECT 1269.745 559.045 1269.915 613.955 ;
        RECT 1269.285 455.345 1269.455 476.255 ;
        RECT 1269.745 379.185 1269.915 400.775 ;
        RECT 1269.745 83.045 1269.915 90.355 ;
      LAYER mcon ;
        RECT 1269.745 1304.325 1269.915 1304.495 ;
        RECT 1270.205 1193.485 1270.375 1193.655 ;
        RECT 1270.205 710.345 1270.375 710.515 ;
        RECT 1269.745 613.785 1269.915 613.955 ;
        RECT 1269.285 476.085 1269.455 476.255 ;
        RECT 1269.745 400.605 1269.915 400.775 ;
        RECT 1269.745 90.185 1269.915 90.355 ;
      LAYER met1 ;
        RECT 1270.130 1594.160 1270.450 1594.220 ;
        RECT 1270.590 1594.160 1270.910 1594.220 ;
        RECT 1270.130 1594.020 1270.910 1594.160 ;
        RECT 1270.130 1593.960 1270.450 1594.020 ;
        RECT 1270.590 1593.960 1270.910 1594.020 ;
        RECT 1270.130 1491.280 1270.450 1491.540 ;
        RECT 1270.220 1490.860 1270.360 1491.280 ;
        RECT 1270.130 1490.600 1270.450 1490.860 ;
        RECT 1269.210 1435.380 1269.530 1435.440 ;
        RECT 1270.130 1435.380 1270.450 1435.440 ;
        RECT 1269.210 1435.240 1270.450 1435.380 ;
        RECT 1269.210 1435.180 1269.530 1435.240 ;
        RECT 1270.130 1435.180 1270.450 1435.240 ;
        RECT 1269.685 1304.480 1269.975 1304.525 ;
        RECT 1270.130 1304.480 1270.450 1304.540 ;
        RECT 1269.685 1304.340 1270.450 1304.480 ;
        RECT 1269.685 1304.295 1269.975 1304.340 ;
        RECT 1270.130 1304.280 1270.450 1304.340 ;
        RECT 1269.670 1290.540 1269.990 1290.600 ;
        RECT 1269.475 1290.400 1269.990 1290.540 ;
        RECT 1269.670 1290.340 1269.990 1290.400 ;
        RECT 1270.130 1193.640 1270.450 1193.700 ;
        RECT 1269.935 1193.500 1270.450 1193.640 ;
        RECT 1270.130 1193.440 1270.450 1193.500 ;
        RECT 1270.130 1151.480 1270.450 1151.540 ;
        RECT 1269.935 1151.340 1270.450 1151.480 ;
        RECT 1270.130 1151.280 1270.450 1151.340 ;
        RECT 1269.670 869.420 1269.990 869.680 ;
        RECT 1269.760 869.280 1269.900 869.420 ;
        RECT 1270.590 869.280 1270.910 869.340 ;
        RECT 1269.760 869.140 1270.910 869.280 ;
        RECT 1270.590 869.080 1270.910 869.140 ;
        RECT 1269.670 759.120 1269.990 759.180 ;
        RECT 1270.590 759.120 1270.910 759.180 ;
        RECT 1269.670 758.980 1270.910 759.120 ;
        RECT 1269.670 758.920 1269.990 758.980 ;
        RECT 1270.590 758.920 1270.910 758.980 ;
        RECT 1270.145 710.500 1270.435 710.545 ;
        RECT 1270.590 710.500 1270.910 710.560 ;
        RECT 1270.145 710.360 1270.910 710.500 ;
        RECT 1270.145 710.315 1270.435 710.360 ;
        RECT 1270.590 710.300 1270.910 710.360 ;
        RECT 1270.130 662.560 1270.450 662.620 ;
        RECT 1269.935 662.420 1270.450 662.560 ;
        RECT 1270.130 662.360 1270.450 662.420 ;
        RECT 1269.670 621.080 1269.990 621.140 ;
        RECT 1270.130 621.080 1270.450 621.140 ;
        RECT 1269.670 620.940 1270.450 621.080 ;
        RECT 1269.670 620.880 1269.990 620.940 ;
        RECT 1270.130 620.880 1270.450 620.940 ;
        RECT 1269.670 613.940 1269.990 614.000 ;
        RECT 1269.475 613.800 1269.990 613.940 ;
        RECT 1269.670 613.740 1269.990 613.800 ;
        RECT 1269.685 559.200 1269.975 559.245 ;
        RECT 1270.590 559.200 1270.910 559.260 ;
        RECT 1269.685 559.060 1270.910 559.200 ;
        RECT 1269.685 559.015 1269.975 559.060 ;
        RECT 1270.590 559.000 1270.910 559.060 ;
        RECT 1269.670 518.060 1269.990 518.120 ;
        RECT 1270.590 518.060 1270.910 518.120 ;
        RECT 1269.670 517.920 1270.910 518.060 ;
        RECT 1269.670 517.860 1269.990 517.920 ;
        RECT 1270.590 517.860 1270.910 517.920 ;
        RECT 1269.210 476.240 1269.530 476.300 ;
        RECT 1269.015 476.100 1269.530 476.240 ;
        RECT 1269.210 476.040 1269.530 476.100 ;
        RECT 1269.210 455.500 1269.530 455.560 ;
        RECT 1269.015 455.360 1269.530 455.500 ;
        RECT 1269.210 455.300 1269.530 455.360 ;
        RECT 1269.210 427.960 1269.530 428.020 ;
        RECT 1269.670 427.960 1269.990 428.020 ;
        RECT 1269.210 427.820 1269.990 427.960 ;
        RECT 1269.210 427.760 1269.530 427.820 ;
        RECT 1269.670 427.760 1269.990 427.820 ;
        RECT 1269.670 400.760 1269.990 400.820 ;
        RECT 1269.475 400.620 1269.990 400.760 ;
        RECT 1269.670 400.560 1269.990 400.620 ;
        RECT 1269.670 379.340 1269.990 379.400 ;
        RECT 1269.475 379.200 1269.990 379.340 ;
        RECT 1269.670 379.140 1269.990 379.200 ;
        RECT 1269.670 217.500 1269.990 217.560 ;
        RECT 1270.590 217.500 1270.910 217.560 ;
        RECT 1269.670 217.360 1270.910 217.500 ;
        RECT 1269.670 217.300 1269.990 217.360 ;
        RECT 1270.590 217.300 1270.910 217.360 ;
        RECT 1270.590 145.420 1270.910 145.480 ;
        RECT 1269.760 145.280 1270.910 145.420 ;
        RECT 1269.760 144.800 1269.900 145.280 ;
        RECT 1270.590 145.220 1270.910 145.280 ;
        RECT 1269.670 144.540 1269.990 144.800 ;
        RECT 1269.670 90.340 1269.990 90.400 ;
        RECT 1269.475 90.200 1269.990 90.340 ;
        RECT 1269.670 90.140 1269.990 90.200 ;
        RECT 1269.670 83.200 1269.990 83.260 ;
        RECT 1269.475 83.060 1269.990 83.200 ;
        RECT 1269.670 83.000 1269.990 83.060 ;
        RECT 1269.670 17.580 1269.990 17.640 ;
        RECT 1255.040 17.440 1269.990 17.580 ;
        RECT 1197.910 17.240 1198.230 17.300 ;
        RECT 1255.040 17.240 1255.180 17.440 ;
        RECT 1269.670 17.380 1269.990 17.440 ;
        RECT 1197.910 17.100 1255.180 17.240 ;
        RECT 1197.910 17.040 1198.230 17.100 ;
      LAYER via ;
        RECT 1270.160 1593.960 1270.420 1594.220 ;
        RECT 1270.620 1593.960 1270.880 1594.220 ;
        RECT 1270.160 1491.280 1270.420 1491.540 ;
        RECT 1270.160 1490.600 1270.420 1490.860 ;
        RECT 1269.240 1435.180 1269.500 1435.440 ;
        RECT 1270.160 1435.180 1270.420 1435.440 ;
        RECT 1270.160 1304.280 1270.420 1304.540 ;
        RECT 1269.700 1290.340 1269.960 1290.600 ;
        RECT 1270.160 1193.440 1270.420 1193.700 ;
        RECT 1270.160 1151.280 1270.420 1151.540 ;
        RECT 1269.700 869.420 1269.960 869.680 ;
        RECT 1270.620 869.080 1270.880 869.340 ;
        RECT 1269.700 758.920 1269.960 759.180 ;
        RECT 1270.620 758.920 1270.880 759.180 ;
        RECT 1270.620 710.300 1270.880 710.560 ;
        RECT 1270.160 662.360 1270.420 662.620 ;
        RECT 1269.700 620.880 1269.960 621.140 ;
        RECT 1270.160 620.880 1270.420 621.140 ;
        RECT 1269.700 613.740 1269.960 614.000 ;
        RECT 1270.620 559.000 1270.880 559.260 ;
        RECT 1269.700 517.860 1269.960 518.120 ;
        RECT 1270.620 517.860 1270.880 518.120 ;
        RECT 1269.240 476.040 1269.500 476.300 ;
        RECT 1269.240 455.300 1269.500 455.560 ;
        RECT 1269.240 427.760 1269.500 428.020 ;
        RECT 1269.700 427.760 1269.960 428.020 ;
        RECT 1269.700 400.560 1269.960 400.820 ;
        RECT 1269.700 379.140 1269.960 379.400 ;
        RECT 1269.700 217.300 1269.960 217.560 ;
        RECT 1270.620 217.300 1270.880 217.560 ;
        RECT 1270.620 145.220 1270.880 145.480 ;
        RECT 1269.700 144.540 1269.960 144.800 ;
        RECT 1269.700 90.140 1269.960 90.400 ;
        RECT 1269.700 83.000 1269.960 83.260 ;
        RECT 1197.940 17.040 1198.200 17.300 ;
        RECT 1269.700 17.380 1269.960 17.640 ;
      LAYER met2 ;
        RECT 1272.820 1700.340 1273.100 1704.000 ;
        RECT 1272.820 1700.000 1273.120 1700.340 ;
        RECT 1272.980 1677.405 1273.120 1700.000 ;
        RECT 1270.610 1677.035 1270.890 1677.405 ;
        RECT 1272.910 1677.035 1273.190 1677.405 ;
        RECT 1270.680 1594.250 1270.820 1677.035 ;
        RECT 1270.160 1593.930 1270.420 1594.250 ;
        RECT 1270.620 1593.930 1270.880 1594.250 ;
        RECT 1270.220 1491.570 1270.360 1593.930 ;
        RECT 1270.160 1491.250 1270.420 1491.570 ;
        RECT 1270.160 1490.570 1270.420 1490.890 ;
        RECT 1270.220 1483.605 1270.360 1490.570 ;
        RECT 1269.230 1483.235 1269.510 1483.605 ;
        RECT 1270.150 1483.235 1270.430 1483.605 ;
        RECT 1269.300 1435.470 1269.440 1483.235 ;
        RECT 1269.240 1435.150 1269.500 1435.470 ;
        RECT 1270.160 1435.150 1270.420 1435.470 ;
        RECT 1270.220 1304.570 1270.360 1435.150 ;
        RECT 1270.160 1304.250 1270.420 1304.570 ;
        RECT 1269.700 1290.310 1269.960 1290.630 ;
        RECT 1269.760 1193.810 1269.900 1290.310 ;
        RECT 1269.760 1193.730 1270.360 1193.810 ;
        RECT 1269.760 1193.670 1270.420 1193.730 ;
        RECT 1270.160 1193.410 1270.420 1193.670 ;
        RECT 1270.160 1151.250 1270.420 1151.570 ;
        RECT 1270.220 1128.530 1270.360 1151.250 ;
        RECT 1269.760 1128.390 1270.360 1128.530 ;
        RECT 1269.760 1007.605 1269.900 1128.390 ;
        RECT 1269.690 1007.235 1269.970 1007.605 ;
        RECT 1270.610 1007.235 1270.890 1007.605 ;
        RECT 1270.680 989.810 1270.820 1007.235 ;
        RECT 1270.220 989.670 1270.820 989.810 ;
        RECT 1270.220 932.010 1270.360 989.670 ;
        RECT 1270.220 931.870 1270.820 932.010 ;
        RECT 1270.680 931.330 1270.820 931.870 ;
        RECT 1269.760 931.190 1270.820 931.330 ;
        RECT 1269.760 869.710 1269.900 931.190 ;
        RECT 1269.700 869.390 1269.960 869.710 ;
        RECT 1270.620 869.050 1270.880 869.370 ;
        RECT 1270.680 759.210 1270.820 869.050 ;
        RECT 1269.700 758.890 1269.960 759.210 ;
        RECT 1270.620 758.890 1270.880 759.210 ;
        RECT 1269.760 724.725 1269.900 758.890 ;
        RECT 1269.690 724.355 1269.970 724.725 ;
        RECT 1270.610 724.355 1270.890 724.725 ;
        RECT 1270.680 710.590 1270.820 724.355 ;
        RECT 1270.620 710.270 1270.880 710.590 ;
        RECT 1270.160 662.330 1270.420 662.650 ;
        RECT 1270.220 621.170 1270.360 662.330 ;
        RECT 1269.700 620.850 1269.960 621.170 ;
        RECT 1270.160 620.850 1270.420 621.170 ;
        RECT 1269.760 614.030 1269.900 620.850 ;
        RECT 1269.700 613.710 1269.960 614.030 ;
        RECT 1270.620 558.970 1270.880 559.290 ;
        RECT 1270.680 518.150 1270.820 558.970 ;
        RECT 1269.700 517.830 1269.960 518.150 ;
        RECT 1270.620 517.830 1270.880 518.150 ;
        RECT 1269.760 503.610 1269.900 517.830 ;
        RECT 1269.300 503.470 1269.900 503.610 ;
        RECT 1269.300 476.330 1269.440 503.470 ;
        RECT 1269.240 476.010 1269.500 476.330 ;
        RECT 1269.240 455.270 1269.500 455.590 ;
        RECT 1269.300 428.050 1269.440 455.270 ;
        RECT 1269.240 427.730 1269.500 428.050 ;
        RECT 1269.700 427.730 1269.960 428.050 ;
        RECT 1269.760 400.850 1269.900 427.730 ;
        RECT 1269.700 400.530 1269.960 400.850 ;
        RECT 1269.700 379.110 1269.960 379.430 ;
        RECT 1269.760 217.590 1269.900 379.110 ;
        RECT 1269.700 217.270 1269.960 217.590 ;
        RECT 1270.620 217.270 1270.880 217.590 ;
        RECT 1270.680 145.510 1270.820 217.270 ;
        RECT 1270.620 145.190 1270.880 145.510 ;
        RECT 1269.700 144.510 1269.960 144.830 ;
        RECT 1269.760 90.430 1269.900 144.510 ;
        RECT 1269.700 90.110 1269.960 90.430 ;
        RECT 1269.700 82.970 1269.960 83.290 ;
        RECT 1269.760 17.670 1269.900 82.970 ;
        RECT 1269.700 17.350 1269.960 17.670 ;
        RECT 1197.940 17.010 1198.200 17.330 ;
        RECT 1198.000 2.400 1198.140 17.010 ;
        RECT 1197.790 -4.800 1198.350 2.400 ;
      LAYER via2 ;
        RECT 1270.610 1677.080 1270.890 1677.360 ;
        RECT 1272.910 1677.080 1273.190 1677.360 ;
        RECT 1269.230 1483.280 1269.510 1483.560 ;
        RECT 1270.150 1483.280 1270.430 1483.560 ;
        RECT 1269.690 1007.280 1269.970 1007.560 ;
        RECT 1270.610 1007.280 1270.890 1007.560 ;
        RECT 1269.690 724.400 1269.970 724.680 ;
        RECT 1270.610 724.400 1270.890 724.680 ;
      LAYER met3 ;
        RECT 1270.585 1677.370 1270.915 1677.385 ;
        RECT 1272.885 1677.370 1273.215 1677.385 ;
        RECT 1270.585 1677.070 1273.215 1677.370 ;
        RECT 1270.585 1677.055 1270.915 1677.070 ;
        RECT 1272.885 1677.055 1273.215 1677.070 ;
        RECT 1269.205 1483.570 1269.535 1483.585 ;
        RECT 1270.125 1483.570 1270.455 1483.585 ;
        RECT 1269.205 1483.270 1270.455 1483.570 ;
        RECT 1269.205 1483.255 1269.535 1483.270 ;
        RECT 1270.125 1483.255 1270.455 1483.270 ;
        RECT 1269.665 1007.570 1269.995 1007.585 ;
        RECT 1270.585 1007.570 1270.915 1007.585 ;
        RECT 1269.665 1007.270 1270.915 1007.570 ;
        RECT 1269.665 1007.255 1269.995 1007.270 ;
        RECT 1270.585 1007.255 1270.915 1007.270 ;
        RECT 1269.665 724.690 1269.995 724.705 ;
        RECT 1270.585 724.690 1270.915 724.705 ;
        RECT 1269.665 724.390 1270.915 724.690 ;
        RECT 1269.665 724.375 1269.995 724.390 ;
        RECT 1270.585 724.375 1270.915 724.390 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1244.905 17.425 1245.075 19.635 ;
      LAYER mcon ;
        RECT 1244.905 19.465 1245.075 19.635 ;
      LAYER met1 ;
        RECT 1244.845 19.620 1245.135 19.665 ;
        RECT 1274.730 19.620 1275.050 19.680 ;
        RECT 1244.845 19.480 1275.050 19.620 ;
        RECT 1244.845 19.435 1245.135 19.480 ;
        RECT 1274.730 19.420 1275.050 19.480 ;
        RECT 1215.850 17.580 1216.170 17.640 ;
        RECT 1244.845 17.580 1245.135 17.625 ;
        RECT 1215.850 17.440 1245.135 17.580 ;
        RECT 1215.850 17.380 1216.170 17.440 ;
        RECT 1244.845 17.395 1245.135 17.440 ;
      LAYER via ;
        RECT 1274.760 19.420 1275.020 19.680 ;
        RECT 1215.880 17.380 1216.140 17.640 ;
      LAYER met2 ;
        RECT 1274.660 1700.340 1274.940 1704.000 ;
        RECT 1274.660 1700.000 1274.960 1700.340 ;
        RECT 1274.820 19.710 1274.960 1700.000 ;
        RECT 1274.760 19.390 1275.020 19.710 ;
        RECT 1215.880 17.350 1216.140 17.670 ;
        RECT 1215.940 2.400 1216.080 17.350 ;
        RECT 1215.730 -4.800 1216.290 2.400 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1233.790 19.280 1234.110 19.340 ;
        RECT 1276.570 19.280 1276.890 19.340 ;
        RECT 1233.790 19.140 1276.890 19.280 ;
        RECT 1233.790 19.080 1234.110 19.140 ;
        RECT 1276.570 19.080 1276.890 19.140 ;
      LAYER via ;
        RECT 1233.820 19.080 1234.080 19.340 ;
        RECT 1276.600 19.080 1276.860 19.340 ;
      LAYER met2 ;
        RECT 1276.500 1700.340 1276.780 1704.000 ;
        RECT 1276.500 1700.000 1276.800 1700.340 ;
        RECT 1276.660 19.370 1276.800 1700.000 ;
        RECT 1233.820 19.050 1234.080 19.370 ;
        RECT 1276.600 19.050 1276.860 19.370 ;
        RECT 1233.880 2.400 1234.020 19.050 ;
        RECT 1233.670 -4.800 1234.230 2.400 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1278.410 1676.780 1278.730 1676.840 ;
        RECT 1280.250 1676.780 1280.570 1676.840 ;
        RECT 1278.410 1676.640 1280.570 1676.780 ;
        RECT 1278.410 1676.580 1278.730 1676.640 ;
        RECT 1280.250 1676.580 1280.570 1676.640 ;
        RECT 1251.730 14.520 1252.050 14.580 ;
        RECT 1280.250 14.520 1280.570 14.580 ;
        RECT 1251.730 14.380 1280.570 14.520 ;
        RECT 1251.730 14.320 1252.050 14.380 ;
        RECT 1280.250 14.320 1280.570 14.380 ;
      LAYER via ;
        RECT 1278.440 1676.580 1278.700 1676.840 ;
        RECT 1280.280 1676.580 1280.540 1676.840 ;
        RECT 1251.760 14.320 1252.020 14.580 ;
        RECT 1280.280 14.320 1280.540 14.580 ;
      LAYER met2 ;
        RECT 1278.340 1700.340 1278.620 1704.000 ;
        RECT 1278.340 1700.000 1278.640 1700.340 ;
        RECT 1278.500 1676.870 1278.640 1700.000 ;
        RECT 1278.440 1676.550 1278.700 1676.870 ;
        RECT 1280.280 1676.550 1280.540 1676.870 ;
        RECT 1280.340 14.610 1280.480 1676.550 ;
        RECT 1251.760 14.290 1252.020 14.610 ;
        RECT 1280.280 14.290 1280.540 14.610 ;
        RECT 1251.820 2.400 1251.960 14.290 ;
        RECT 1251.610 -4.800 1252.170 2.400 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1280.250 1677.800 1280.570 1677.860 ;
        RECT 1278.040 1677.660 1280.570 1677.800 ;
        RECT 1278.040 1676.100 1278.180 1677.660 ;
        RECT 1280.250 1677.600 1280.570 1677.660 ;
        RECT 1278.410 1676.100 1278.730 1676.160 ;
        RECT 1278.040 1675.960 1278.730 1676.100 ;
        RECT 1278.410 1675.900 1278.730 1675.960 ;
        RECT 1269.210 17.240 1269.530 17.300 ;
        RECT 1278.410 17.240 1278.730 17.300 ;
        RECT 1269.210 17.100 1278.730 17.240 ;
        RECT 1269.210 17.040 1269.530 17.100 ;
        RECT 1278.410 17.040 1278.730 17.100 ;
      LAYER via ;
        RECT 1280.280 1677.600 1280.540 1677.860 ;
        RECT 1278.440 1675.900 1278.700 1676.160 ;
        RECT 1269.240 17.040 1269.500 17.300 ;
        RECT 1278.440 17.040 1278.700 17.300 ;
      LAYER met2 ;
        RECT 1280.180 1700.340 1280.460 1704.000 ;
        RECT 1280.180 1700.000 1280.480 1700.340 ;
        RECT 1280.340 1677.890 1280.480 1700.000 ;
        RECT 1280.280 1677.570 1280.540 1677.890 ;
        RECT 1278.440 1675.870 1278.700 1676.190 ;
        RECT 1278.500 17.330 1278.640 1675.870 ;
        RECT 1269.240 17.010 1269.500 17.330 ;
        RECT 1278.440 17.010 1278.700 17.330 ;
        RECT 1269.300 2.400 1269.440 17.010 ;
        RECT 1269.090 -4.800 1269.650 2.400 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1282.165 1658.605 1282.335 1676.455 ;
        RECT 1282.625 848.725 1282.795 869.975 ;
        RECT 1282.165 697.085 1282.335 745.195 ;
        RECT 1282.625 565.845 1282.795 613.955 ;
        RECT 1283.085 131.325 1283.255 179.435 ;
      LAYER mcon ;
        RECT 1282.165 1676.285 1282.335 1676.455 ;
        RECT 1282.625 869.805 1282.795 869.975 ;
        RECT 1282.165 745.025 1282.335 745.195 ;
        RECT 1282.625 613.785 1282.795 613.955 ;
        RECT 1283.085 179.265 1283.255 179.435 ;
      LAYER met1 ;
        RECT 1282.090 1676.440 1282.410 1676.500 ;
        RECT 1281.895 1676.300 1282.410 1676.440 ;
        RECT 1282.090 1676.240 1282.410 1676.300 ;
        RECT 1282.105 1658.760 1282.395 1658.805 ;
        RECT 1283.010 1658.760 1283.330 1658.820 ;
        RECT 1282.105 1658.620 1283.330 1658.760 ;
        RECT 1282.105 1658.575 1282.395 1658.620 ;
        RECT 1283.010 1658.560 1283.330 1658.620 ;
        RECT 1282.090 1580.220 1282.410 1580.280 ;
        RECT 1283.010 1580.220 1283.330 1580.280 ;
        RECT 1282.090 1580.080 1283.330 1580.220 ;
        RECT 1282.090 1580.020 1282.410 1580.080 ;
        RECT 1283.010 1580.020 1283.330 1580.080 ;
        RECT 1282.090 1531.940 1282.410 1532.000 ;
        RECT 1283.470 1531.940 1283.790 1532.000 ;
        RECT 1282.090 1531.800 1283.790 1531.940 ;
        RECT 1282.090 1531.740 1282.410 1531.800 ;
        RECT 1283.470 1531.740 1283.790 1531.800 ;
        RECT 1282.550 1510.520 1282.870 1510.580 ;
        RECT 1283.470 1510.520 1283.790 1510.580 ;
        RECT 1282.550 1510.380 1283.790 1510.520 ;
        RECT 1282.550 1510.320 1282.870 1510.380 ;
        RECT 1283.470 1510.320 1283.790 1510.380 ;
        RECT 1282.550 1449.120 1282.870 1449.380 ;
        RECT 1282.640 1448.640 1282.780 1449.120 ;
        RECT 1283.010 1448.640 1283.330 1448.700 ;
        RECT 1282.640 1448.500 1283.330 1448.640 ;
        RECT 1283.010 1448.440 1283.330 1448.500 ;
        RECT 1282.550 1111.020 1282.870 1111.080 ;
        RECT 1283.010 1111.020 1283.330 1111.080 ;
        RECT 1282.550 1110.880 1283.330 1111.020 ;
        RECT 1282.550 1110.820 1282.870 1110.880 ;
        RECT 1283.010 1110.820 1283.330 1110.880 ;
        RECT 1282.565 869.960 1282.855 870.005 ;
        RECT 1283.010 869.960 1283.330 870.020 ;
        RECT 1282.565 869.820 1283.330 869.960 ;
        RECT 1282.565 869.775 1282.855 869.820 ;
        RECT 1283.010 869.760 1283.330 869.820 ;
        RECT 1282.550 848.880 1282.870 848.940 ;
        RECT 1282.355 848.740 1282.870 848.880 ;
        RECT 1282.550 848.680 1282.870 848.740 ;
        RECT 1283.010 759.120 1283.330 759.180 ;
        RECT 1284.390 759.120 1284.710 759.180 ;
        RECT 1283.010 758.980 1284.710 759.120 ;
        RECT 1283.010 758.920 1283.330 758.980 ;
        RECT 1284.390 758.920 1284.710 758.980 ;
        RECT 1282.105 745.180 1282.395 745.225 ;
        RECT 1283.930 745.180 1284.250 745.240 ;
        RECT 1282.105 745.040 1284.250 745.180 ;
        RECT 1282.105 744.995 1282.395 745.040 ;
        RECT 1283.930 744.980 1284.250 745.040 ;
        RECT 1282.090 697.240 1282.410 697.300 ;
        RECT 1281.895 697.100 1282.410 697.240 ;
        RECT 1282.090 697.040 1282.410 697.100 ;
        RECT 1282.550 613.940 1282.870 614.000 ;
        RECT 1282.355 613.800 1282.870 613.940 ;
        RECT 1282.550 613.740 1282.870 613.800 ;
        RECT 1282.565 566.000 1282.855 566.045 ;
        RECT 1283.010 566.000 1283.330 566.060 ;
        RECT 1282.565 565.860 1283.330 566.000 ;
        RECT 1282.565 565.815 1282.855 565.860 ;
        RECT 1283.010 565.800 1283.330 565.860 ;
        RECT 1282.550 427.960 1282.870 428.020 ;
        RECT 1283.470 427.960 1283.790 428.020 ;
        RECT 1282.550 427.820 1283.790 427.960 ;
        RECT 1282.550 427.760 1282.870 427.820 ;
        RECT 1283.470 427.760 1283.790 427.820 ;
        RECT 1282.550 400.220 1282.870 400.480 ;
        RECT 1282.640 399.740 1282.780 400.220 ;
        RECT 1283.010 399.740 1283.330 399.800 ;
        RECT 1282.640 399.600 1283.330 399.740 ;
        RECT 1283.010 399.540 1283.330 399.600 ;
        RECT 1282.550 331.400 1282.870 331.460 ;
        RECT 1283.010 331.400 1283.330 331.460 ;
        RECT 1282.550 331.260 1283.330 331.400 ;
        RECT 1282.550 331.200 1282.870 331.260 ;
        RECT 1283.010 331.200 1283.330 331.260 ;
        RECT 1282.550 283.120 1282.870 283.180 ;
        RECT 1283.010 283.120 1283.330 283.180 ;
        RECT 1282.550 282.980 1283.330 283.120 ;
        RECT 1282.550 282.920 1282.870 282.980 ;
        RECT 1283.010 282.920 1283.330 282.980 ;
        RECT 1283.010 186.220 1283.330 186.280 ;
        RECT 1283.470 186.220 1283.790 186.280 ;
        RECT 1283.010 186.080 1283.790 186.220 ;
        RECT 1283.010 186.020 1283.330 186.080 ;
        RECT 1283.470 186.020 1283.790 186.080 ;
        RECT 1283.025 179.420 1283.315 179.465 ;
        RECT 1283.470 179.420 1283.790 179.480 ;
        RECT 1283.025 179.280 1283.790 179.420 ;
        RECT 1283.025 179.235 1283.315 179.280 ;
        RECT 1283.470 179.220 1283.790 179.280 ;
        RECT 1283.010 131.480 1283.330 131.540 ;
        RECT 1282.815 131.340 1283.330 131.480 ;
        RECT 1283.010 131.280 1283.330 131.340 ;
        RECT 1282.550 83.540 1282.870 83.600 ;
        RECT 1282.550 83.400 1283.240 83.540 ;
        RECT 1282.550 83.340 1282.870 83.400 ;
        RECT 1283.100 83.260 1283.240 83.400 ;
        RECT 1283.010 83.000 1283.330 83.260 ;
        RECT 1282.550 41.380 1282.870 41.440 ;
        RECT 1287.150 41.380 1287.470 41.440 ;
        RECT 1282.550 41.240 1287.470 41.380 ;
        RECT 1282.550 41.180 1282.870 41.240 ;
        RECT 1287.150 41.180 1287.470 41.240 ;
      LAYER via ;
        RECT 1282.120 1676.240 1282.380 1676.500 ;
        RECT 1283.040 1658.560 1283.300 1658.820 ;
        RECT 1282.120 1580.020 1282.380 1580.280 ;
        RECT 1283.040 1580.020 1283.300 1580.280 ;
        RECT 1282.120 1531.740 1282.380 1532.000 ;
        RECT 1283.500 1531.740 1283.760 1532.000 ;
        RECT 1282.580 1510.320 1282.840 1510.580 ;
        RECT 1283.500 1510.320 1283.760 1510.580 ;
        RECT 1282.580 1449.120 1282.840 1449.380 ;
        RECT 1283.040 1448.440 1283.300 1448.700 ;
        RECT 1282.580 1110.820 1282.840 1111.080 ;
        RECT 1283.040 1110.820 1283.300 1111.080 ;
        RECT 1283.040 869.760 1283.300 870.020 ;
        RECT 1282.580 848.680 1282.840 848.940 ;
        RECT 1283.040 758.920 1283.300 759.180 ;
        RECT 1284.420 758.920 1284.680 759.180 ;
        RECT 1283.960 744.980 1284.220 745.240 ;
        RECT 1282.120 697.040 1282.380 697.300 ;
        RECT 1282.580 613.740 1282.840 614.000 ;
        RECT 1283.040 565.800 1283.300 566.060 ;
        RECT 1282.580 427.760 1282.840 428.020 ;
        RECT 1283.500 427.760 1283.760 428.020 ;
        RECT 1282.580 400.220 1282.840 400.480 ;
        RECT 1283.040 399.540 1283.300 399.800 ;
        RECT 1282.580 331.200 1282.840 331.460 ;
        RECT 1283.040 331.200 1283.300 331.460 ;
        RECT 1282.580 282.920 1282.840 283.180 ;
        RECT 1283.040 282.920 1283.300 283.180 ;
        RECT 1283.040 186.020 1283.300 186.280 ;
        RECT 1283.500 186.020 1283.760 186.280 ;
        RECT 1283.500 179.220 1283.760 179.480 ;
        RECT 1283.040 131.280 1283.300 131.540 ;
        RECT 1282.580 83.340 1282.840 83.600 ;
        RECT 1283.040 83.000 1283.300 83.260 ;
        RECT 1282.580 41.180 1282.840 41.440 ;
        RECT 1287.180 41.180 1287.440 41.440 ;
      LAYER met2 ;
        RECT 1282.020 1700.340 1282.300 1704.000 ;
        RECT 1282.020 1700.000 1282.320 1700.340 ;
        RECT 1282.180 1676.530 1282.320 1700.000 ;
        RECT 1282.120 1676.210 1282.380 1676.530 ;
        RECT 1283.040 1658.530 1283.300 1658.850 ;
        RECT 1283.100 1628.445 1283.240 1658.530 ;
        RECT 1282.110 1628.075 1282.390 1628.445 ;
        RECT 1283.030 1628.075 1283.310 1628.445 ;
        RECT 1282.180 1580.310 1282.320 1628.075 ;
        RECT 1282.120 1580.165 1282.380 1580.310 ;
        RECT 1283.040 1580.165 1283.300 1580.310 ;
        RECT 1282.110 1579.795 1282.390 1580.165 ;
        RECT 1283.030 1579.795 1283.310 1580.165 ;
        RECT 1282.180 1532.030 1282.320 1579.795 ;
        RECT 1282.120 1531.710 1282.380 1532.030 ;
        RECT 1283.500 1531.710 1283.760 1532.030 ;
        RECT 1283.560 1510.610 1283.700 1531.710 ;
        RECT 1282.580 1510.290 1282.840 1510.610 ;
        RECT 1283.500 1510.290 1283.760 1510.610 ;
        RECT 1282.640 1449.410 1282.780 1510.290 ;
        RECT 1282.580 1449.090 1282.840 1449.410 ;
        RECT 1283.040 1448.410 1283.300 1448.730 ;
        RECT 1283.100 1221.690 1283.240 1448.410 ;
        RECT 1282.640 1221.550 1283.240 1221.690 ;
        RECT 1282.640 1221.010 1282.780 1221.550 ;
        RECT 1282.640 1220.870 1283.240 1221.010 ;
        RECT 1283.100 1111.110 1283.240 1220.870 ;
        RECT 1282.580 1110.790 1282.840 1111.110 ;
        RECT 1283.040 1110.790 1283.300 1111.110 ;
        RECT 1282.640 1086.370 1282.780 1110.790 ;
        RECT 1282.640 1086.230 1283.240 1086.370 ;
        RECT 1283.100 932.010 1283.240 1086.230 ;
        RECT 1282.640 931.870 1283.240 932.010 ;
        RECT 1282.640 931.330 1282.780 931.870 ;
        RECT 1282.640 931.190 1283.240 931.330 ;
        RECT 1283.100 870.050 1283.240 931.190 ;
        RECT 1283.040 869.730 1283.300 870.050 ;
        RECT 1282.580 848.650 1282.840 848.970 ;
        RECT 1282.640 832.050 1282.780 848.650 ;
        RECT 1282.640 831.910 1283.240 832.050 ;
        RECT 1283.100 759.210 1283.240 831.910 ;
        RECT 1283.040 758.890 1283.300 759.210 ;
        RECT 1284.420 758.890 1284.680 759.210 ;
        RECT 1284.480 752.490 1284.620 758.890 ;
        RECT 1284.020 752.350 1284.620 752.490 ;
        RECT 1284.020 745.270 1284.160 752.350 ;
        RECT 1283.960 744.950 1284.220 745.270 ;
        RECT 1282.120 697.010 1282.380 697.330 ;
        RECT 1282.180 662.165 1282.320 697.010 ;
        RECT 1282.110 661.795 1282.390 662.165 ;
        RECT 1283.030 661.795 1283.310 662.165 ;
        RECT 1283.100 637.570 1283.240 661.795 ;
        RECT 1282.640 637.430 1283.240 637.570 ;
        RECT 1282.640 614.030 1282.780 637.430 ;
        RECT 1282.580 613.710 1282.840 614.030 ;
        RECT 1283.040 565.770 1283.300 566.090 ;
        RECT 1283.100 524.010 1283.240 565.770 ;
        RECT 1283.100 523.870 1283.700 524.010 ;
        RECT 1283.560 428.050 1283.700 523.870 ;
        RECT 1282.580 427.730 1282.840 428.050 ;
        RECT 1283.500 427.730 1283.760 428.050 ;
        RECT 1282.640 400.510 1282.780 427.730 ;
        RECT 1282.580 400.190 1282.840 400.510 ;
        RECT 1283.040 399.510 1283.300 399.830 ;
        RECT 1283.100 331.490 1283.240 399.510 ;
        RECT 1282.580 331.170 1282.840 331.490 ;
        RECT 1283.040 331.170 1283.300 331.490 ;
        RECT 1282.640 283.210 1282.780 331.170 ;
        RECT 1282.580 282.890 1282.840 283.210 ;
        RECT 1283.040 282.890 1283.300 283.210 ;
        RECT 1283.100 186.310 1283.240 282.890 ;
        RECT 1283.040 185.990 1283.300 186.310 ;
        RECT 1283.500 185.990 1283.760 186.310 ;
        RECT 1283.560 179.510 1283.700 185.990 ;
        RECT 1283.500 179.190 1283.760 179.510 ;
        RECT 1283.040 131.250 1283.300 131.570 ;
        RECT 1283.100 130.970 1283.240 131.250 ;
        RECT 1282.640 130.830 1283.240 130.970 ;
        RECT 1282.640 83.630 1282.780 130.830 ;
        RECT 1282.580 83.310 1282.840 83.630 ;
        RECT 1283.040 82.970 1283.300 83.290 ;
        RECT 1283.100 48.690 1283.240 82.970 ;
        RECT 1283.100 48.550 1283.700 48.690 ;
        RECT 1283.560 47.330 1283.700 48.550 ;
        RECT 1282.640 47.190 1283.700 47.330 ;
        RECT 1282.640 41.470 1282.780 47.190 ;
        RECT 1282.580 41.150 1282.840 41.470 ;
        RECT 1287.180 41.150 1287.440 41.470 ;
        RECT 1287.240 2.400 1287.380 41.150 ;
        RECT 1287.030 -4.800 1287.590 2.400 ;
      LAYER via2 ;
        RECT 1282.110 1628.120 1282.390 1628.400 ;
        RECT 1283.030 1628.120 1283.310 1628.400 ;
        RECT 1282.110 1579.840 1282.390 1580.120 ;
        RECT 1283.030 1579.840 1283.310 1580.120 ;
        RECT 1282.110 661.840 1282.390 662.120 ;
        RECT 1283.030 661.840 1283.310 662.120 ;
      LAYER met3 ;
        RECT 1282.085 1628.410 1282.415 1628.425 ;
        RECT 1283.005 1628.410 1283.335 1628.425 ;
        RECT 1282.085 1628.110 1283.335 1628.410 ;
        RECT 1282.085 1628.095 1282.415 1628.110 ;
        RECT 1283.005 1628.095 1283.335 1628.110 ;
        RECT 1282.085 1580.130 1282.415 1580.145 ;
        RECT 1283.005 1580.130 1283.335 1580.145 ;
        RECT 1282.085 1579.830 1283.335 1580.130 ;
        RECT 1282.085 1579.815 1282.415 1579.830 ;
        RECT 1283.005 1579.815 1283.335 1579.830 ;
        RECT 1282.085 662.130 1282.415 662.145 ;
        RECT 1283.005 662.130 1283.335 662.145 ;
        RECT 1282.085 661.830 1283.335 662.130 ;
        RECT 1282.085 661.815 1282.415 661.830 ;
        RECT 1283.005 661.815 1283.335 661.830 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1283.930 1677.460 1284.250 1677.520 ;
        RECT 1288.990 1677.460 1289.310 1677.520 ;
        RECT 1283.930 1677.320 1289.310 1677.460 ;
        RECT 1283.930 1677.260 1284.250 1677.320 ;
        RECT 1288.990 1677.260 1289.310 1677.320 ;
        RECT 1288.990 19.960 1289.310 20.020 ;
        RECT 1305.090 19.960 1305.410 20.020 ;
        RECT 1288.990 19.820 1305.410 19.960 ;
        RECT 1288.990 19.760 1289.310 19.820 ;
        RECT 1305.090 19.760 1305.410 19.820 ;
      LAYER via ;
        RECT 1283.960 1677.260 1284.220 1677.520 ;
        RECT 1289.020 1677.260 1289.280 1677.520 ;
        RECT 1289.020 19.760 1289.280 20.020 ;
        RECT 1305.120 19.760 1305.380 20.020 ;
      LAYER met2 ;
        RECT 1283.860 1700.340 1284.140 1704.000 ;
        RECT 1283.860 1700.000 1284.160 1700.340 ;
        RECT 1284.020 1677.550 1284.160 1700.000 ;
        RECT 1283.960 1677.230 1284.220 1677.550 ;
        RECT 1289.020 1677.230 1289.280 1677.550 ;
        RECT 1289.080 20.050 1289.220 1677.230 ;
        RECT 1289.020 19.730 1289.280 20.050 ;
        RECT 1305.120 19.730 1305.380 20.050 ;
        RECT 1305.180 2.400 1305.320 19.730 ;
        RECT 1304.970 -4.800 1305.530 2.400 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1285.770 1689.360 1286.090 1689.420 ;
        RECT 1317.050 1689.360 1317.370 1689.420 ;
        RECT 1285.770 1689.220 1317.370 1689.360 ;
        RECT 1285.770 1689.160 1286.090 1689.220 ;
        RECT 1317.050 1689.160 1317.370 1689.220 ;
        RECT 1314.290 1666.580 1314.610 1666.640 ;
        RECT 1317.050 1666.580 1317.370 1666.640 ;
        RECT 1314.290 1666.440 1317.370 1666.580 ;
        RECT 1314.290 1666.380 1314.610 1666.440 ;
        RECT 1317.050 1666.380 1317.370 1666.440 ;
        RECT 1314.290 20.640 1314.610 20.700 ;
        RECT 1323.030 20.640 1323.350 20.700 ;
        RECT 1314.290 20.500 1323.350 20.640 ;
        RECT 1314.290 20.440 1314.610 20.500 ;
        RECT 1323.030 20.440 1323.350 20.500 ;
      LAYER via ;
        RECT 1285.800 1689.160 1286.060 1689.420 ;
        RECT 1317.080 1689.160 1317.340 1689.420 ;
        RECT 1314.320 1666.380 1314.580 1666.640 ;
        RECT 1317.080 1666.380 1317.340 1666.640 ;
        RECT 1314.320 20.440 1314.580 20.700 ;
        RECT 1323.060 20.440 1323.320 20.700 ;
      LAYER met2 ;
        RECT 1285.700 1700.340 1285.980 1704.000 ;
        RECT 1285.700 1700.000 1286.000 1700.340 ;
        RECT 1285.860 1689.450 1286.000 1700.000 ;
        RECT 1285.800 1689.130 1286.060 1689.450 ;
        RECT 1317.080 1689.130 1317.340 1689.450 ;
        RECT 1317.140 1666.670 1317.280 1689.130 ;
        RECT 1314.320 1666.350 1314.580 1666.670 ;
        RECT 1317.080 1666.350 1317.340 1666.670 ;
        RECT 1314.380 20.730 1314.520 1666.350 ;
        RECT 1314.320 20.410 1314.580 20.730 ;
        RECT 1323.060 20.410 1323.320 20.730 ;
        RECT 1323.120 2.400 1323.260 20.410 ;
        RECT 1322.910 -4.800 1323.470 2.400 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1287.610 1688.680 1287.930 1688.740 ;
        RECT 1311.070 1688.680 1311.390 1688.740 ;
        RECT 1287.610 1688.540 1311.390 1688.680 ;
        RECT 1287.610 1688.480 1287.930 1688.540 ;
        RECT 1311.070 1688.480 1311.390 1688.540 ;
        RECT 1311.070 1683.920 1311.390 1683.980 ;
        RECT 1311.070 1683.780 1312.220 1683.920 ;
        RECT 1311.070 1683.720 1311.390 1683.780 ;
        RECT 1312.080 1683.240 1312.220 1683.780 ;
        RECT 1314.290 1683.240 1314.610 1683.300 ;
        RECT 1312.080 1683.100 1314.610 1683.240 ;
        RECT 1314.290 1683.040 1314.610 1683.100 ;
        RECT 1314.750 34.580 1315.070 34.640 ;
        RECT 1340.510 34.580 1340.830 34.640 ;
        RECT 1314.750 34.440 1340.830 34.580 ;
        RECT 1314.750 34.380 1315.070 34.440 ;
        RECT 1340.510 34.380 1340.830 34.440 ;
      LAYER via ;
        RECT 1287.640 1688.480 1287.900 1688.740 ;
        RECT 1311.100 1688.480 1311.360 1688.740 ;
        RECT 1311.100 1683.720 1311.360 1683.980 ;
        RECT 1314.320 1683.040 1314.580 1683.300 ;
        RECT 1314.780 34.380 1315.040 34.640 ;
        RECT 1340.540 34.380 1340.800 34.640 ;
      LAYER met2 ;
        RECT 1287.540 1700.340 1287.820 1704.000 ;
        RECT 1287.540 1700.000 1287.840 1700.340 ;
        RECT 1287.700 1688.770 1287.840 1700.000 ;
        RECT 1287.640 1688.450 1287.900 1688.770 ;
        RECT 1311.100 1688.450 1311.360 1688.770 ;
        RECT 1311.160 1684.010 1311.300 1688.450 ;
        RECT 1311.100 1683.690 1311.360 1684.010 ;
        RECT 1314.320 1683.010 1314.580 1683.330 ;
        RECT 1314.380 1667.090 1314.520 1683.010 ;
        RECT 1314.380 1666.950 1314.980 1667.090 ;
        RECT 1314.840 34.670 1314.980 1666.950 ;
        RECT 1314.780 34.350 1315.040 34.670 ;
        RECT 1340.540 34.350 1340.800 34.670 ;
        RECT 1340.600 2.400 1340.740 34.350 ;
        RECT 1340.390 -4.800 1340.950 2.400 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 703.410 1590.760 703.730 1590.820 ;
        RECT 1222.750 1590.760 1223.070 1590.820 ;
        RECT 703.410 1590.620 1223.070 1590.760 ;
        RECT 703.410 1590.560 703.730 1590.620 ;
        RECT 1222.750 1590.560 1223.070 1590.620 ;
      LAYER via ;
        RECT 703.440 1590.560 703.700 1590.820 ;
        RECT 1222.780 1590.560 1223.040 1590.820 ;
      LAYER met2 ;
        RECT 1221.300 1700.410 1221.580 1704.000 ;
        RECT 1221.300 1700.270 1222.060 1700.410 ;
        RECT 1221.300 1700.000 1221.580 1700.270 ;
        RECT 1221.920 1677.970 1222.060 1700.270 ;
        RECT 1221.920 1677.830 1222.980 1677.970 ;
        RECT 1222.840 1590.850 1222.980 1677.830 ;
        RECT 703.440 1590.530 703.700 1590.850 ;
        RECT 1222.780 1590.530 1223.040 1590.850 ;
        RECT 703.500 24.210 703.640 1590.530 ;
        RECT 698.440 24.070 703.640 24.210 ;
        RECT 698.440 2.400 698.580 24.070 ;
        RECT 698.230 -4.800 698.790 2.400 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1285.770 1684.600 1286.090 1684.660 ;
        RECT 1289.450 1684.600 1289.770 1684.660 ;
        RECT 1285.770 1684.460 1289.770 1684.600 ;
        RECT 1285.770 1684.400 1286.090 1684.460 ;
        RECT 1289.450 1684.400 1289.770 1684.460 ;
        RECT 1285.770 1583.620 1286.090 1583.680 ;
        RECT 1352.470 1583.620 1352.790 1583.680 ;
        RECT 1285.770 1583.480 1352.790 1583.620 ;
        RECT 1285.770 1583.420 1286.090 1583.480 ;
        RECT 1352.470 1583.420 1352.790 1583.480 ;
        RECT 1352.470 37.980 1352.790 38.040 ;
        RECT 1358.450 37.980 1358.770 38.040 ;
        RECT 1352.470 37.840 1358.770 37.980 ;
        RECT 1352.470 37.780 1352.790 37.840 ;
        RECT 1358.450 37.780 1358.770 37.840 ;
      LAYER via ;
        RECT 1285.800 1684.400 1286.060 1684.660 ;
        RECT 1289.480 1684.400 1289.740 1684.660 ;
        RECT 1285.800 1583.420 1286.060 1583.680 ;
        RECT 1352.500 1583.420 1352.760 1583.680 ;
        RECT 1352.500 37.780 1352.760 38.040 ;
        RECT 1358.480 37.780 1358.740 38.040 ;
      LAYER met2 ;
        RECT 1289.380 1700.340 1289.660 1704.000 ;
        RECT 1289.380 1700.000 1289.680 1700.340 ;
        RECT 1289.540 1684.690 1289.680 1700.000 ;
        RECT 1285.800 1684.370 1286.060 1684.690 ;
        RECT 1289.480 1684.370 1289.740 1684.690 ;
        RECT 1285.860 1583.710 1286.000 1684.370 ;
        RECT 1285.800 1583.390 1286.060 1583.710 ;
        RECT 1352.500 1583.390 1352.760 1583.710 ;
        RECT 1352.560 38.070 1352.700 1583.390 ;
        RECT 1352.500 37.750 1352.760 38.070 ;
        RECT 1358.480 37.750 1358.740 38.070 ;
        RECT 1358.540 2.400 1358.680 37.750 ;
        RECT 1358.330 -4.800 1358.890 2.400 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1314.825 1683.765 1314.995 1688.015 ;
        RECT 1318.505 1683.765 1318.675 1684.615 ;
        RECT 1355.305 1655.885 1355.475 1685.975 ;
      LAYER mcon ;
        RECT 1314.825 1687.845 1314.995 1688.015 ;
        RECT 1355.305 1685.805 1355.475 1685.975 ;
        RECT 1318.505 1684.445 1318.675 1684.615 ;
      LAYER met1 ;
        RECT 1291.290 1688.000 1291.610 1688.060 ;
        RECT 1314.765 1688.000 1315.055 1688.045 ;
        RECT 1291.290 1687.860 1315.055 1688.000 ;
        RECT 1291.290 1687.800 1291.610 1687.860 ;
        RECT 1314.765 1687.815 1315.055 1687.860 ;
        RECT 1355.245 1685.960 1355.535 1686.005 ;
        RECT 1318.980 1685.820 1355.535 1685.960 ;
        RECT 1318.445 1684.600 1318.735 1684.645 ;
        RECT 1318.980 1684.600 1319.120 1685.820 ;
        RECT 1355.245 1685.775 1355.535 1685.820 ;
        RECT 1318.445 1684.460 1319.120 1684.600 ;
        RECT 1318.445 1684.415 1318.735 1684.460 ;
        RECT 1314.765 1683.920 1315.055 1683.965 ;
        RECT 1318.445 1683.920 1318.735 1683.965 ;
        RECT 1314.765 1683.780 1318.735 1683.920 ;
        RECT 1314.765 1683.735 1315.055 1683.780 ;
        RECT 1318.445 1683.735 1318.735 1683.780 ;
        RECT 1355.245 1656.040 1355.535 1656.085 ;
        RECT 1362.590 1656.040 1362.910 1656.100 ;
        RECT 1355.245 1655.900 1362.910 1656.040 ;
        RECT 1355.245 1655.855 1355.535 1655.900 ;
        RECT 1362.590 1655.840 1362.910 1655.900 ;
        RECT 1362.590 1632.040 1362.910 1632.300 ;
        RECT 1362.680 1631.280 1362.820 1632.040 ;
        RECT 1362.590 1631.020 1362.910 1631.280 ;
        RECT 1362.590 20.980 1362.910 21.040 ;
        RECT 1376.390 20.980 1376.710 21.040 ;
        RECT 1362.590 20.840 1376.710 20.980 ;
        RECT 1362.590 20.780 1362.910 20.840 ;
        RECT 1376.390 20.780 1376.710 20.840 ;
      LAYER via ;
        RECT 1291.320 1687.800 1291.580 1688.060 ;
        RECT 1362.620 1655.840 1362.880 1656.100 ;
        RECT 1362.620 1632.040 1362.880 1632.300 ;
        RECT 1362.620 1631.020 1362.880 1631.280 ;
        RECT 1362.620 20.780 1362.880 21.040 ;
        RECT 1376.420 20.780 1376.680 21.040 ;
      LAYER met2 ;
        RECT 1291.220 1700.340 1291.500 1704.000 ;
        RECT 1291.220 1700.000 1291.520 1700.340 ;
        RECT 1291.380 1688.090 1291.520 1700.000 ;
        RECT 1291.320 1687.770 1291.580 1688.090 ;
        RECT 1362.620 1655.810 1362.880 1656.130 ;
        RECT 1362.680 1632.330 1362.820 1655.810 ;
        RECT 1362.620 1632.010 1362.880 1632.330 ;
        RECT 1362.620 1630.990 1362.880 1631.310 ;
        RECT 1362.680 21.070 1362.820 1630.990 ;
        RECT 1362.620 20.750 1362.880 21.070 ;
        RECT 1376.420 20.750 1376.680 21.070 ;
        RECT 1376.480 2.400 1376.620 20.750 ;
        RECT 1376.270 -4.800 1376.830 2.400 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1293.130 1685.620 1293.450 1685.680 ;
        RECT 1304.630 1685.620 1304.950 1685.680 ;
        RECT 1293.130 1685.480 1304.950 1685.620 ;
        RECT 1293.130 1685.420 1293.450 1685.480 ;
        RECT 1304.630 1685.420 1304.950 1685.480 ;
        RECT 1304.630 1683.920 1304.950 1683.980 ;
        RECT 1304.630 1683.780 1306.240 1683.920 ;
        RECT 1304.630 1683.720 1304.950 1683.780 ;
        RECT 1306.100 1683.580 1306.240 1683.780 ;
        RECT 1307.850 1683.580 1308.170 1683.640 ;
        RECT 1306.100 1683.440 1308.170 1683.580 ;
        RECT 1307.850 1683.380 1308.170 1683.440 ;
        RECT 1307.850 1597.220 1308.170 1597.280 ;
        RECT 1393.870 1597.220 1394.190 1597.280 ;
        RECT 1307.850 1597.080 1394.190 1597.220 ;
        RECT 1307.850 1597.020 1308.170 1597.080 ;
        RECT 1393.870 1597.020 1394.190 1597.080 ;
      LAYER via ;
        RECT 1293.160 1685.420 1293.420 1685.680 ;
        RECT 1304.660 1685.420 1304.920 1685.680 ;
        RECT 1304.660 1683.720 1304.920 1683.980 ;
        RECT 1307.880 1683.380 1308.140 1683.640 ;
        RECT 1307.880 1597.020 1308.140 1597.280 ;
        RECT 1393.900 1597.020 1394.160 1597.280 ;
      LAYER met2 ;
        RECT 1293.060 1700.340 1293.340 1704.000 ;
        RECT 1293.060 1700.000 1293.360 1700.340 ;
        RECT 1293.220 1685.710 1293.360 1700.000 ;
        RECT 1293.160 1685.390 1293.420 1685.710 ;
        RECT 1304.660 1685.390 1304.920 1685.710 ;
        RECT 1304.720 1684.010 1304.860 1685.390 ;
        RECT 1304.660 1683.690 1304.920 1684.010 ;
        RECT 1307.880 1683.350 1308.140 1683.670 ;
        RECT 1307.940 1597.310 1308.080 1683.350 ;
        RECT 1307.880 1596.990 1308.140 1597.310 ;
        RECT 1393.900 1596.990 1394.160 1597.310 ;
        RECT 1393.960 3.130 1394.100 1596.990 ;
        RECT 1393.960 2.990 1394.560 3.130 ;
        RECT 1394.420 2.400 1394.560 2.990 ;
        RECT 1394.210 -4.800 1394.770 2.400 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1294.970 1590.420 1295.290 1590.480 ;
        RECT 1407.670 1590.420 1407.990 1590.480 ;
        RECT 1294.970 1590.280 1407.990 1590.420 ;
        RECT 1294.970 1590.220 1295.290 1590.280 ;
        RECT 1407.670 1590.220 1407.990 1590.280 ;
        RECT 1407.670 2.960 1407.990 3.020 ;
        RECT 1412.270 2.960 1412.590 3.020 ;
        RECT 1407.670 2.820 1412.590 2.960 ;
        RECT 1407.670 2.760 1407.990 2.820 ;
        RECT 1412.270 2.760 1412.590 2.820 ;
      LAYER via ;
        RECT 1295.000 1590.220 1295.260 1590.480 ;
        RECT 1407.700 1590.220 1407.960 1590.480 ;
        RECT 1407.700 2.760 1407.960 3.020 ;
        RECT 1412.300 2.760 1412.560 3.020 ;
      LAYER met2 ;
        RECT 1294.900 1700.340 1295.180 1704.000 ;
        RECT 1294.900 1700.000 1295.200 1700.340 ;
        RECT 1295.060 1590.510 1295.200 1700.000 ;
        RECT 1295.000 1590.190 1295.260 1590.510 ;
        RECT 1407.700 1590.190 1407.960 1590.510 ;
        RECT 1407.760 3.050 1407.900 1590.190 ;
        RECT 1407.700 2.730 1407.960 3.050 ;
        RECT 1412.300 2.730 1412.560 3.050 ;
        RECT 1412.360 2.400 1412.500 2.730 ;
        RECT 1412.150 -4.800 1412.710 2.400 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1296.810 1617.960 1297.130 1618.020 ;
        RECT 1428.370 1617.960 1428.690 1618.020 ;
        RECT 1296.810 1617.820 1428.690 1617.960 ;
        RECT 1296.810 1617.760 1297.130 1617.820 ;
        RECT 1428.370 1617.760 1428.690 1617.820 ;
        RECT 1428.370 2.960 1428.690 3.020 ;
        RECT 1429.750 2.960 1430.070 3.020 ;
        RECT 1428.370 2.820 1430.070 2.960 ;
        RECT 1428.370 2.760 1428.690 2.820 ;
        RECT 1429.750 2.760 1430.070 2.820 ;
      LAYER via ;
        RECT 1296.840 1617.760 1297.100 1618.020 ;
        RECT 1428.400 1617.760 1428.660 1618.020 ;
        RECT 1428.400 2.760 1428.660 3.020 ;
        RECT 1429.780 2.760 1430.040 3.020 ;
      LAYER met2 ;
        RECT 1296.740 1700.340 1297.020 1704.000 ;
        RECT 1296.740 1700.000 1297.040 1700.340 ;
        RECT 1296.900 1618.050 1297.040 1700.000 ;
        RECT 1296.840 1617.730 1297.100 1618.050 ;
        RECT 1428.400 1617.730 1428.660 1618.050 ;
        RECT 1428.460 3.050 1428.600 1617.730 ;
        RECT 1428.400 2.730 1428.660 3.050 ;
        RECT 1429.780 2.730 1430.040 3.050 ;
        RECT 1429.840 2.400 1429.980 2.730 ;
        RECT 1429.630 -4.800 1430.190 2.400 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1352.560 1652.840 1421.700 1652.980 ;
        RECT 1298.650 1652.300 1298.970 1652.360 ;
        RECT 1352.560 1652.300 1352.700 1652.840 ;
        RECT 1421.560 1652.640 1421.700 1652.840 ;
        RECT 1442.170 1652.640 1442.490 1652.700 ;
        RECT 1421.560 1652.500 1442.490 1652.640 ;
        RECT 1442.170 1652.440 1442.490 1652.500 ;
        RECT 1298.650 1652.160 1352.700 1652.300 ;
        RECT 1298.650 1652.100 1298.970 1652.160 ;
        RECT 1442.170 2.960 1442.490 3.020 ;
        RECT 1447.690 2.960 1448.010 3.020 ;
        RECT 1442.170 2.820 1448.010 2.960 ;
        RECT 1442.170 2.760 1442.490 2.820 ;
        RECT 1447.690 2.760 1448.010 2.820 ;
      LAYER via ;
        RECT 1298.680 1652.100 1298.940 1652.360 ;
        RECT 1442.200 1652.440 1442.460 1652.700 ;
        RECT 1442.200 2.760 1442.460 3.020 ;
        RECT 1447.720 2.760 1447.980 3.020 ;
      LAYER met2 ;
        RECT 1298.580 1700.340 1298.860 1704.000 ;
        RECT 1298.580 1700.000 1298.880 1700.340 ;
        RECT 1298.740 1652.390 1298.880 1700.000 ;
        RECT 1442.200 1652.410 1442.460 1652.730 ;
        RECT 1298.680 1652.070 1298.940 1652.390 ;
        RECT 1442.260 3.050 1442.400 1652.410 ;
        RECT 1442.200 2.730 1442.460 3.050 ;
        RECT 1447.720 2.730 1447.980 3.050 ;
        RECT 1447.780 2.400 1447.920 2.730 ;
        RECT 1447.570 -4.800 1448.130 2.400 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1300.490 1685.280 1300.810 1685.340 ;
        RECT 1302.790 1685.280 1303.110 1685.340 ;
        RECT 1300.490 1685.140 1303.110 1685.280 ;
        RECT 1300.490 1685.080 1300.810 1685.140 ;
        RECT 1302.790 1685.080 1303.110 1685.140 ;
        RECT 1302.790 1668.620 1303.110 1668.680 ;
        RECT 1462.870 1668.620 1463.190 1668.680 ;
        RECT 1302.790 1668.480 1463.190 1668.620 ;
        RECT 1302.790 1668.420 1303.110 1668.480 ;
        RECT 1462.870 1668.420 1463.190 1668.480 ;
        RECT 1462.870 2.960 1463.190 3.020 ;
        RECT 1465.630 2.960 1465.950 3.020 ;
        RECT 1462.870 2.820 1465.950 2.960 ;
        RECT 1462.870 2.760 1463.190 2.820 ;
        RECT 1465.630 2.760 1465.950 2.820 ;
      LAYER via ;
        RECT 1300.520 1685.080 1300.780 1685.340 ;
        RECT 1302.820 1685.080 1303.080 1685.340 ;
        RECT 1302.820 1668.420 1303.080 1668.680 ;
        RECT 1462.900 1668.420 1463.160 1668.680 ;
        RECT 1462.900 2.760 1463.160 3.020 ;
        RECT 1465.660 2.760 1465.920 3.020 ;
      LAYER met2 ;
        RECT 1300.420 1700.340 1300.700 1704.000 ;
        RECT 1300.420 1700.000 1300.720 1700.340 ;
        RECT 1300.580 1685.370 1300.720 1700.000 ;
        RECT 1300.520 1685.050 1300.780 1685.370 ;
        RECT 1302.820 1685.050 1303.080 1685.370 ;
        RECT 1302.880 1668.710 1303.020 1685.050 ;
        RECT 1302.820 1668.390 1303.080 1668.710 ;
        RECT 1462.900 1668.390 1463.160 1668.710 ;
        RECT 1462.960 3.050 1463.100 1668.390 ;
        RECT 1462.900 2.730 1463.160 3.050 ;
        RECT 1465.660 2.730 1465.920 3.050 ;
        RECT 1465.720 2.400 1465.860 2.730 ;
        RECT 1465.510 -4.800 1466.070 2.400 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1303.325 1683.765 1303.495 1685.975 ;
      LAYER mcon ;
        RECT 1303.325 1685.805 1303.495 1685.975 ;
      LAYER met1 ;
        RECT 1302.330 1685.960 1302.650 1686.020 ;
        RECT 1303.265 1685.960 1303.555 1686.005 ;
        RECT 1302.330 1685.820 1303.555 1685.960 ;
        RECT 1302.330 1685.760 1302.650 1685.820 ;
        RECT 1303.265 1685.775 1303.555 1685.820 ;
        RECT 1303.250 1683.920 1303.570 1683.980 ;
        RECT 1303.055 1683.780 1303.570 1683.920 ;
        RECT 1303.250 1683.720 1303.570 1683.780 ;
        RECT 1303.250 1661.820 1303.570 1661.880 ;
        RECT 1484.030 1661.820 1484.350 1661.880 ;
        RECT 1303.250 1661.680 1484.350 1661.820 ;
        RECT 1303.250 1661.620 1303.570 1661.680 ;
        RECT 1484.030 1661.620 1484.350 1661.680 ;
      LAYER via ;
        RECT 1302.360 1685.760 1302.620 1686.020 ;
        RECT 1303.280 1683.720 1303.540 1683.980 ;
        RECT 1303.280 1661.620 1303.540 1661.880 ;
        RECT 1484.060 1661.620 1484.320 1661.880 ;
      LAYER met2 ;
        RECT 1302.260 1700.340 1302.540 1704.000 ;
        RECT 1302.260 1700.000 1302.560 1700.340 ;
        RECT 1302.420 1686.050 1302.560 1700.000 ;
        RECT 1302.360 1685.730 1302.620 1686.050 ;
        RECT 1303.280 1683.690 1303.540 1684.010 ;
        RECT 1303.340 1661.910 1303.480 1683.690 ;
        RECT 1303.280 1661.590 1303.540 1661.910 ;
        RECT 1484.060 1661.590 1484.320 1661.910 ;
        RECT 1484.120 7.210 1484.260 1661.590 ;
        RECT 1483.660 7.070 1484.260 7.210 ;
        RECT 1483.660 2.400 1483.800 7.070 ;
        RECT 1483.450 -4.800 1484.010 2.400 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1304.170 1685.280 1304.490 1685.340 ;
        RECT 1309.230 1685.280 1309.550 1685.340 ;
        RECT 1304.170 1685.140 1309.550 1685.280 ;
        RECT 1304.170 1685.080 1304.490 1685.140 ;
        RECT 1309.230 1685.080 1309.550 1685.140 ;
        RECT 1309.230 1640.400 1309.550 1640.460 ;
        RECT 1497.370 1640.400 1497.690 1640.460 ;
        RECT 1309.230 1640.260 1497.690 1640.400 ;
        RECT 1309.230 1640.200 1309.550 1640.260 ;
        RECT 1497.370 1640.200 1497.690 1640.260 ;
        RECT 1497.370 2.960 1497.690 3.020 ;
        RECT 1501.510 2.960 1501.830 3.020 ;
        RECT 1497.370 2.820 1501.830 2.960 ;
        RECT 1497.370 2.760 1497.690 2.820 ;
        RECT 1501.510 2.760 1501.830 2.820 ;
      LAYER via ;
        RECT 1304.200 1685.080 1304.460 1685.340 ;
        RECT 1309.260 1685.080 1309.520 1685.340 ;
        RECT 1309.260 1640.200 1309.520 1640.460 ;
        RECT 1497.400 1640.200 1497.660 1640.460 ;
        RECT 1497.400 2.760 1497.660 3.020 ;
        RECT 1501.540 2.760 1501.800 3.020 ;
      LAYER met2 ;
        RECT 1304.100 1700.340 1304.380 1704.000 ;
        RECT 1304.100 1700.000 1304.400 1700.340 ;
        RECT 1304.260 1685.370 1304.400 1700.000 ;
        RECT 1304.200 1685.050 1304.460 1685.370 ;
        RECT 1309.260 1685.050 1309.520 1685.370 ;
        RECT 1309.320 1640.490 1309.460 1685.050 ;
        RECT 1309.260 1640.170 1309.520 1640.490 ;
        RECT 1497.400 1640.170 1497.660 1640.490 ;
        RECT 1497.460 3.050 1497.600 1640.170 ;
        RECT 1497.400 2.730 1497.660 3.050 ;
        RECT 1501.540 2.730 1501.800 3.050 ;
        RECT 1501.600 2.400 1501.740 2.730 ;
        RECT 1501.390 -4.800 1501.950 2.400 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1306.010 1684.600 1306.330 1684.660 ;
        RECT 1310.150 1684.600 1310.470 1684.660 ;
        RECT 1306.010 1684.460 1310.470 1684.600 ;
        RECT 1306.010 1684.400 1306.330 1684.460 ;
        RECT 1310.150 1684.400 1310.470 1684.460 ;
        RECT 1310.150 1647.540 1310.470 1647.600 ;
        RECT 1518.070 1647.540 1518.390 1647.600 ;
        RECT 1310.150 1647.400 1518.390 1647.540 ;
        RECT 1310.150 1647.340 1310.470 1647.400 ;
        RECT 1518.070 1647.340 1518.390 1647.400 ;
        RECT 1518.070 2.960 1518.390 3.020 ;
        RECT 1518.990 2.960 1519.310 3.020 ;
        RECT 1518.070 2.820 1519.310 2.960 ;
        RECT 1518.070 2.760 1518.390 2.820 ;
        RECT 1518.990 2.760 1519.310 2.820 ;
      LAYER via ;
        RECT 1306.040 1684.400 1306.300 1684.660 ;
        RECT 1310.180 1684.400 1310.440 1684.660 ;
        RECT 1310.180 1647.340 1310.440 1647.600 ;
        RECT 1518.100 1647.340 1518.360 1647.600 ;
        RECT 1518.100 2.760 1518.360 3.020 ;
        RECT 1519.020 2.760 1519.280 3.020 ;
      LAYER met2 ;
        RECT 1305.940 1700.340 1306.220 1704.000 ;
        RECT 1305.940 1700.000 1306.240 1700.340 ;
        RECT 1306.100 1684.690 1306.240 1700.000 ;
        RECT 1306.040 1684.370 1306.300 1684.690 ;
        RECT 1310.180 1684.370 1310.440 1684.690 ;
        RECT 1310.240 1647.630 1310.380 1684.370 ;
        RECT 1310.180 1647.310 1310.440 1647.630 ;
        RECT 1518.100 1647.310 1518.360 1647.630 ;
        RECT 1518.160 3.050 1518.300 1647.310 ;
        RECT 1518.100 2.730 1518.360 3.050 ;
        RECT 1519.020 2.730 1519.280 3.050 ;
        RECT 1519.080 2.400 1519.220 2.730 ;
        RECT 1518.870 -4.800 1519.430 2.400 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1223.210 1679.500 1223.530 1679.560 ;
        RECT 1225.510 1679.500 1225.830 1679.560 ;
        RECT 1223.210 1679.360 1225.830 1679.500 ;
        RECT 1223.210 1679.300 1223.530 1679.360 ;
        RECT 1225.510 1679.300 1225.830 1679.360 ;
        RECT 717.210 1583.960 717.530 1584.020 ;
        RECT 1225.510 1583.960 1225.830 1584.020 ;
        RECT 717.210 1583.820 1225.830 1583.960 ;
        RECT 717.210 1583.760 717.530 1583.820 ;
        RECT 1225.510 1583.760 1225.830 1583.820 ;
      LAYER via ;
        RECT 1223.240 1679.300 1223.500 1679.560 ;
        RECT 1225.540 1679.300 1225.800 1679.560 ;
        RECT 717.240 1583.760 717.500 1584.020 ;
        RECT 1225.540 1583.760 1225.800 1584.020 ;
      LAYER met2 ;
        RECT 1223.140 1700.340 1223.420 1704.000 ;
        RECT 1223.140 1700.000 1223.440 1700.340 ;
        RECT 1223.300 1679.590 1223.440 1700.000 ;
        RECT 1223.240 1679.270 1223.500 1679.590 ;
        RECT 1225.540 1679.270 1225.800 1679.590 ;
        RECT 1225.600 1584.050 1225.740 1679.270 ;
        RECT 717.240 1583.730 717.500 1584.050 ;
        RECT 1225.540 1583.730 1225.800 1584.050 ;
        RECT 717.300 16.730 717.440 1583.730 ;
        RECT 716.380 16.590 717.440 16.730 ;
        RECT 716.380 2.400 716.520 16.590 ;
        RECT 716.170 -4.800 716.730 2.400 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1304.170 1684.260 1304.490 1684.320 ;
        RECT 1307.850 1684.260 1308.170 1684.320 ;
        RECT 1304.170 1684.120 1308.170 1684.260 ;
        RECT 1304.170 1684.060 1304.490 1684.120 ;
        RECT 1307.850 1684.060 1308.170 1684.120 ;
        RECT 1304.170 1612.520 1304.490 1612.580 ;
        RECT 1531.870 1612.520 1532.190 1612.580 ;
        RECT 1304.170 1612.380 1532.190 1612.520 ;
        RECT 1304.170 1612.320 1304.490 1612.380 ;
        RECT 1531.870 1612.320 1532.190 1612.380 ;
      LAYER via ;
        RECT 1304.200 1684.060 1304.460 1684.320 ;
        RECT 1307.880 1684.060 1308.140 1684.320 ;
        RECT 1304.200 1612.320 1304.460 1612.580 ;
        RECT 1531.900 1612.320 1532.160 1612.580 ;
      LAYER met2 ;
        RECT 1307.780 1700.340 1308.060 1704.000 ;
        RECT 1307.780 1700.000 1308.080 1700.340 ;
        RECT 1307.940 1684.350 1308.080 1700.000 ;
        RECT 1304.200 1684.030 1304.460 1684.350 ;
        RECT 1307.880 1684.030 1308.140 1684.350 ;
        RECT 1304.260 1612.610 1304.400 1684.030 ;
        RECT 1304.200 1612.290 1304.460 1612.610 ;
        RECT 1531.900 1612.290 1532.160 1612.610 ;
        RECT 1531.960 17.410 1532.100 1612.290 ;
        RECT 1531.960 17.270 1537.160 17.410 ;
        RECT 1537.020 2.400 1537.160 17.270 ;
        RECT 1536.810 -4.800 1537.370 2.400 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1305.090 1684.940 1305.410 1685.000 ;
        RECT 1309.690 1684.940 1310.010 1685.000 ;
        RECT 1305.090 1684.800 1310.010 1684.940 ;
        RECT 1305.090 1684.740 1305.410 1684.800 ;
        RECT 1309.690 1684.740 1310.010 1684.800 ;
        RECT 1305.090 1549.960 1305.410 1550.020 ;
        RECT 1552.570 1549.960 1552.890 1550.020 ;
        RECT 1305.090 1549.820 1552.890 1549.960 ;
        RECT 1305.090 1549.760 1305.410 1549.820 ;
        RECT 1552.570 1549.760 1552.890 1549.820 ;
      LAYER via ;
        RECT 1305.120 1684.740 1305.380 1685.000 ;
        RECT 1309.720 1684.740 1309.980 1685.000 ;
        RECT 1305.120 1549.760 1305.380 1550.020 ;
        RECT 1552.600 1549.760 1552.860 1550.020 ;
      LAYER met2 ;
        RECT 1309.620 1700.340 1309.900 1704.000 ;
        RECT 1309.620 1700.000 1309.920 1700.340 ;
        RECT 1309.780 1685.030 1309.920 1700.000 ;
        RECT 1305.120 1684.710 1305.380 1685.030 ;
        RECT 1309.720 1684.710 1309.980 1685.030 ;
        RECT 1305.180 1550.050 1305.320 1684.710 ;
        RECT 1305.120 1549.730 1305.380 1550.050 ;
        RECT 1552.600 1549.730 1552.860 1550.050 ;
        RECT 1552.660 17.410 1552.800 1549.730 ;
        RECT 1552.660 17.270 1555.100 17.410 ;
        RECT 1554.960 2.400 1555.100 17.270 ;
        RECT 1554.750 -4.800 1555.310 2.400 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1389.805 1688.185 1389.975 1689.375 ;
        RECT 1404.065 1683.765 1404.235 1688.355 ;
      LAYER mcon ;
        RECT 1389.805 1689.205 1389.975 1689.375 ;
        RECT 1404.065 1688.185 1404.235 1688.355 ;
      LAYER met1 ;
        RECT 1389.745 1689.360 1390.035 1689.405 ;
        RECT 1376.480 1689.220 1390.035 1689.360 ;
        RECT 1311.530 1688.680 1311.850 1688.740 ;
        RECT 1376.480 1688.680 1376.620 1689.220 ;
        RECT 1389.745 1689.175 1390.035 1689.220 ;
        RECT 1311.530 1688.540 1376.620 1688.680 ;
        RECT 1311.530 1688.480 1311.850 1688.540 ;
        RECT 1389.745 1688.340 1390.035 1688.385 ;
        RECT 1404.005 1688.340 1404.295 1688.385 ;
        RECT 1389.745 1688.200 1404.295 1688.340 ;
        RECT 1389.745 1688.155 1390.035 1688.200 ;
        RECT 1404.005 1688.155 1404.295 1688.200 ;
        RECT 1403.990 1683.920 1404.310 1683.980 ;
        RECT 1403.795 1683.780 1404.310 1683.920 ;
        RECT 1403.990 1683.720 1404.310 1683.780 ;
        RECT 1403.990 37.980 1404.310 38.040 ;
        RECT 1572.810 37.980 1573.130 38.040 ;
        RECT 1403.990 37.840 1573.130 37.980 ;
        RECT 1403.990 37.780 1404.310 37.840 ;
        RECT 1572.810 37.780 1573.130 37.840 ;
      LAYER via ;
        RECT 1311.560 1688.480 1311.820 1688.740 ;
        RECT 1404.020 1683.720 1404.280 1683.980 ;
        RECT 1404.020 37.780 1404.280 38.040 ;
        RECT 1572.840 37.780 1573.100 38.040 ;
      LAYER met2 ;
        RECT 1311.460 1700.340 1311.740 1704.000 ;
        RECT 1311.460 1700.000 1311.760 1700.340 ;
        RECT 1311.620 1688.770 1311.760 1700.000 ;
        RECT 1311.560 1688.450 1311.820 1688.770 ;
        RECT 1404.020 1683.690 1404.280 1684.010 ;
        RECT 1404.080 1682.730 1404.220 1683.690 ;
        RECT 1403.620 1682.590 1404.220 1682.730 ;
        RECT 1403.620 1632.410 1403.760 1682.590 ;
        RECT 1403.620 1632.270 1404.220 1632.410 ;
        RECT 1404.080 38.070 1404.220 1632.270 ;
        RECT 1404.020 37.750 1404.280 38.070 ;
        RECT 1572.840 37.750 1573.100 38.070 ;
        RECT 1572.900 2.400 1573.040 37.750 ;
        RECT 1572.690 -4.800 1573.250 2.400 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1312.910 1598.580 1313.230 1598.640 ;
        RECT 1587.070 1598.580 1587.390 1598.640 ;
        RECT 1312.910 1598.440 1587.390 1598.580 ;
        RECT 1312.910 1598.380 1313.230 1598.440 ;
        RECT 1587.070 1598.380 1587.390 1598.440 ;
      LAYER via ;
        RECT 1312.940 1598.380 1313.200 1598.640 ;
        RECT 1587.100 1598.380 1587.360 1598.640 ;
      LAYER met2 ;
        RECT 1313.300 1700.410 1313.580 1704.000 ;
        RECT 1313.000 1700.270 1313.580 1700.410 ;
        RECT 1313.000 1598.670 1313.140 1700.270 ;
        RECT 1313.300 1700.000 1313.580 1700.270 ;
        RECT 1312.940 1598.350 1313.200 1598.670 ;
        RECT 1587.100 1598.350 1587.360 1598.670 ;
        RECT 1587.160 17.410 1587.300 1598.350 ;
        RECT 1587.160 17.270 1590.520 17.410 ;
        RECT 1590.380 2.400 1590.520 17.270 ;
        RECT 1590.170 -4.800 1590.730 2.400 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1311.990 1684.940 1312.310 1685.000 ;
        RECT 1315.210 1684.940 1315.530 1685.000 ;
        RECT 1311.990 1684.800 1315.530 1684.940 ;
        RECT 1311.990 1684.740 1312.310 1684.800 ;
        RECT 1315.210 1684.740 1315.530 1684.800 ;
        RECT 1311.990 1591.440 1312.310 1591.500 ;
        RECT 1607.770 1591.440 1608.090 1591.500 ;
        RECT 1311.990 1591.300 1608.090 1591.440 ;
        RECT 1311.990 1591.240 1312.310 1591.300 ;
        RECT 1607.770 1591.240 1608.090 1591.300 ;
      LAYER via ;
        RECT 1312.020 1684.740 1312.280 1685.000 ;
        RECT 1315.240 1684.740 1315.500 1685.000 ;
        RECT 1312.020 1591.240 1312.280 1591.500 ;
        RECT 1607.800 1591.240 1608.060 1591.500 ;
      LAYER met2 ;
        RECT 1315.140 1700.340 1315.420 1704.000 ;
        RECT 1315.140 1700.000 1315.440 1700.340 ;
        RECT 1315.300 1685.030 1315.440 1700.000 ;
        RECT 1312.020 1684.710 1312.280 1685.030 ;
        RECT 1315.240 1684.710 1315.500 1685.030 ;
        RECT 1312.080 1591.530 1312.220 1684.710 ;
        RECT 1312.020 1591.210 1312.280 1591.530 ;
        RECT 1607.800 1591.210 1608.060 1591.530 ;
        RECT 1607.860 17.410 1608.000 1591.210 ;
        RECT 1607.860 17.270 1608.460 17.410 ;
        RECT 1608.320 2.400 1608.460 17.270 ;
        RECT 1608.110 -4.800 1608.670 2.400 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1316.590 1466.660 1316.910 1466.720 ;
        RECT 1621.570 1466.660 1621.890 1466.720 ;
        RECT 1316.590 1466.520 1621.890 1466.660 ;
        RECT 1316.590 1466.460 1316.910 1466.520 ;
        RECT 1621.570 1466.460 1621.890 1466.520 ;
      LAYER via ;
        RECT 1316.620 1466.460 1316.880 1466.720 ;
        RECT 1621.600 1466.460 1621.860 1466.720 ;
      LAYER met2 ;
        RECT 1316.980 1700.410 1317.260 1704.000 ;
        RECT 1316.680 1700.270 1317.260 1700.410 ;
        RECT 1316.680 1466.750 1316.820 1700.270 ;
        RECT 1316.980 1700.000 1317.260 1700.270 ;
        RECT 1316.620 1466.430 1316.880 1466.750 ;
        RECT 1621.600 1466.430 1621.860 1466.750 ;
        RECT 1621.660 17.410 1621.800 1466.430 ;
        RECT 1621.660 17.270 1626.400 17.410 ;
        RECT 1626.260 2.400 1626.400 17.270 ;
        RECT 1626.050 -4.800 1626.610 2.400 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1318.430 1654.340 1318.750 1654.400 ;
        RECT 1642.270 1654.340 1642.590 1654.400 ;
        RECT 1318.430 1654.200 1642.590 1654.340 ;
        RECT 1318.430 1654.140 1318.750 1654.200 ;
        RECT 1642.270 1654.140 1642.590 1654.200 ;
      LAYER via ;
        RECT 1318.460 1654.140 1318.720 1654.400 ;
        RECT 1642.300 1654.140 1642.560 1654.400 ;
      LAYER met2 ;
        RECT 1318.820 1700.340 1319.100 1704.000 ;
        RECT 1318.820 1700.000 1319.120 1700.340 ;
        RECT 1318.980 1684.600 1319.120 1700.000 ;
        RECT 1318.520 1684.460 1319.120 1684.600 ;
        RECT 1318.520 1654.430 1318.660 1684.460 ;
        RECT 1318.460 1654.110 1318.720 1654.430 ;
        RECT 1642.300 1654.110 1642.560 1654.430 ;
        RECT 1642.360 17.410 1642.500 1654.110 ;
        RECT 1642.360 17.270 1644.340 17.410 ;
        RECT 1644.200 2.400 1644.340 17.270 ;
        RECT 1643.990 -4.800 1644.550 2.400 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1318.890 1683.920 1319.210 1683.980 ;
        RECT 1320.730 1683.920 1321.050 1683.980 ;
        RECT 1318.890 1683.780 1321.050 1683.920 ;
        RECT 1318.890 1683.720 1319.210 1683.780 ;
        RECT 1320.730 1683.720 1321.050 1683.780 ;
        RECT 1318.890 1626.120 1319.210 1626.180 ;
        RECT 1656.530 1626.120 1656.850 1626.180 ;
        RECT 1318.890 1625.980 1656.850 1626.120 ;
        RECT 1318.890 1625.920 1319.210 1625.980 ;
        RECT 1656.530 1625.920 1656.850 1625.980 ;
      LAYER via ;
        RECT 1318.920 1683.720 1319.180 1683.980 ;
        RECT 1320.760 1683.720 1321.020 1683.980 ;
        RECT 1318.920 1625.920 1319.180 1626.180 ;
        RECT 1656.560 1625.920 1656.820 1626.180 ;
      LAYER met2 ;
        RECT 1320.660 1700.340 1320.940 1704.000 ;
        RECT 1320.660 1700.000 1320.960 1700.340 ;
        RECT 1320.820 1684.010 1320.960 1700.000 ;
        RECT 1318.920 1683.690 1319.180 1684.010 ;
        RECT 1320.760 1683.690 1321.020 1684.010 ;
        RECT 1318.980 1626.210 1319.120 1683.690 ;
        RECT 1318.920 1625.890 1319.180 1626.210 ;
        RECT 1656.560 1625.890 1656.820 1626.210 ;
        RECT 1656.620 17.410 1656.760 1625.890 ;
        RECT 1656.620 17.270 1662.280 17.410 ;
        RECT 1662.140 2.400 1662.280 17.270 ;
        RECT 1661.930 -4.800 1662.490 2.400 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1322.570 1612.180 1322.890 1612.240 ;
        RECT 1676.770 1612.180 1677.090 1612.240 ;
        RECT 1322.570 1612.040 1677.090 1612.180 ;
        RECT 1322.570 1611.980 1322.890 1612.040 ;
        RECT 1676.770 1611.980 1677.090 1612.040 ;
      LAYER via ;
        RECT 1322.600 1611.980 1322.860 1612.240 ;
        RECT 1676.800 1611.980 1677.060 1612.240 ;
      LAYER met2 ;
        RECT 1322.500 1700.340 1322.780 1704.000 ;
        RECT 1322.500 1700.000 1322.800 1700.340 ;
        RECT 1322.660 1612.270 1322.800 1700.000 ;
        RECT 1322.600 1611.950 1322.860 1612.270 ;
        RECT 1676.800 1611.950 1677.060 1612.270 ;
        RECT 1676.860 17.410 1677.000 1611.950 ;
        RECT 1676.860 17.270 1679.760 17.410 ;
        RECT 1679.620 2.400 1679.760 17.270 ;
        RECT 1679.410 -4.800 1679.970 2.400 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1319.810 1684.260 1320.130 1684.320 ;
        RECT 1324.410 1684.260 1324.730 1684.320 ;
        RECT 1319.810 1684.120 1324.730 1684.260 ;
        RECT 1319.810 1684.060 1320.130 1684.120 ;
        RECT 1324.410 1684.060 1324.730 1684.120 ;
        RECT 1319.810 1542.820 1320.130 1542.880 ;
        RECT 1697.470 1542.820 1697.790 1542.880 ;
        RECT 1319.810 1542.680 1697.790 1542.820 ;
        RECT 1319.810 1542.620 1320.130 1542.680 ;
        RECT 1697.470 1542.620 1697.790 1542.680 ;
      LAYER via ;
        RECT 1319.840 1684.060 1320.100 1684.320 ;
        RECT 1324.440 1684.060 1324.700 1684.320 ;
        RECT 1319.840 1542.620 1320.100 1542.880 ;
        RECT 1697.500 1542.620 1697.760 1542.880 ;
      LAYER met2 ;
        RECT 1324.340 1700.340 1324.620 1704.000 ;
        RECT 1324.340 1700.000 1324.640 1700.340 ;
        RECT 1324.500 1684.350 1324.640 1700.000 ;
        RECT 1319.840 1684.030 1320.100 1684.350 ;
        RECT 1324.440 1684.030 1324.700 1684.350 ;
        RECT 1319.900 1542.910 1320.040 1684.030 ;
        RECT 1319.840 1542.590 1320.100 1542.910 ;
        RECT 1697.500 1542.590 1697.760 1542.910 ;
        RECT 1697.560 2.400 1697.700 1542.590 ;
        RECT 1697.350 -4.800 1697.910 2.400 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1225.050 1678.140 1225.370 1678.200 ;
        RECT 1227.810 1678.140 1228.130 1678.200 ;
        RECT 1225.050 1678.000 1228.130 1678.140 ;
        RECT 1225.050 1677.940 1225.370 1678.000 ;
        RECT 1227.810 1677.940 1228.130 1678.000 ;
        RECT 737.910 1576.820 738.230 1576.880 ;
        RECT 1227.810 1576.820 1228.130 1576.880 ;
        RECT 737.910 1576.680 1228.130 1576.820 ;
        RECT 737.910 1576.620 738.230 1576.680 ;
        RECT 1227.810 1576.620 1228.130 1576.680 ;
      LAYER via ;
        RECT 1225.080 1677.940 1225.340 1678.200 ;
        RECT 1227.840 1677.940 1228.100 1678.200 ;
        RECT 737.940 1576.620 738.200 1576.880 ;
        RECT 1227.840 1576.620 1228.100 1576.880 ;
      LAYER met2 ;
        RECT 1224.980 1700.340 1225.260 1704.000 ;
        RECT 1224.980 1700.000 1225.280 1700.340 ;
        RECT 1225.140 1678.230 1225.280 1700.000 ;
        RECT 1225.080 1677.910 1225.340 1678.230 ;
        RECT 1227.840 1677.910 1228.100 1678.230 ;
        RECT 1227.900 1576.910 1228.040 1677.910 ;
        RECT 737.940 1576.590 738.200 1576.910 ;
        RECT 1227.840 1576.590 1228.100 1576.910 ;
        RECT 738.000 16.730 738.140 1576.590 ;
        RECT 734.320 16.590 738.140 16.730 ;
        RECT 734.320 2.400 734.460 16.590 ;
        RECT 734.110 -4.800 734.670 2.400 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1330.465 1683.765 1330.635 1686.315 ;
      LAYER mcon ;
        RECT 1330.465 1686.145 1330.635 1686.315 ;
      LAYER met1 ;
        RECT 1326.250 1686.300 1326.570 1686.360 ;
        RECT 1330.405 1686.300 1330.695 1686.345 ;
        RECT 1326.250 1686.160 1330.695 1686.300 ;
        RECT 1326.250 1686.100 1326.570 1686.160 ;
        RECT 1330.405 1686.115 1330.695 1686.160 ;
        RECT 1330.390 1683.920 1330.710 1683.980 ;
        RECT 1330.195 1683.780 1330.710 1683.920 ;
        RECT 1330.390 1683.720 1330.710 1683.780 ;
        RECT 1330.390 1667.600 1330.710 1667.660 ;
        RECT 1711.270 1667.600 1711.590 1667.660 ;
        RECT 1330.390 1667.460 1711.590 1667.600 ;
        RECT 1330.390 1667.400 1330.710 1667.460 ;
        RECT 1711.270 1667.400 1711.590 1667.460 ;
      LAYER via ;
        RECT 1326.280 1686.100 1326.540 1686.360 ;
        RECT 1330.420 1683.720 1330.680 1683.980 ;
        RECT 1330.420 1667.400 1330.680 1667.660 ;
        RECT 1711.300 1667.400 1711.560 1667.660 ;
      LAYER met2 ;
        RECT 1326.180 1700.340 1326.460 1704.000 ;
        RECT 1326.180 1700.000 1326.480 1700.340 ;
        RECT 1326.340 1686.390 1326.480 1700.000 ;
        RECT 1326.280 1686.070 1326.540 1686.390 ;
        RECT 1330.420 1683.690 1330.680 1684.010 ;
        RECT 1330.480 1667.690 1330.620 1683.690 ;
        RECT 1330.420 1667.370 1330.680 1667.690 ;
        RECT 1711.300 1667.370 1711.560 1667.690 ;
        RECT 1711.360 17.410 1711.500 1667.370 ;
        RECT 1711.360 17.270 1715.640 17.410 ;
        RECT 1715.500 2.400 1715.640 17.270 ;
        RECT 1715.290 -4.800 1715.850 2.400 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1376.465 1687.165 1376.635 1688.355 ;
        RECT 1389.345 1687.165 1389.515 1688.355 ;
      LAYER mcon ;
        RECT 1376.465 1688.185 1376.635 1688.355 ;
        RECT 1389.345 1688.185 1389.515 1688.355 ;
      LAYER met1 ;
        RECT 1376.405 1688.340 1376.695 1688.385 ;
        RECT 1389.285 1688.340 1389.575 1688.385 ;
        RECT 1376.405 1688.200 1389.575 1688.340 ;
        RECT 1376.405 1688.155 1376.695 1688.200 ;
        RECT 1389.285 1688.155 1389.575 1688.200 ;
        RECT 1328.090 1687.320 1328.410 1687.380 ;
        RECT 1376.405 1687.320 1376.695 1687.365 ;
        RECT 1328.090 1687.180 1376.695 1687.320 ;
        RECT 1328.090 1687.120 1328.410 1687.180 ;
        RECT 1376.405 1687.135 1376.695 1687.180 ;
        RECT 1389.285 1687.320 1389.575 1687.365 ;
        RECT 1731.970 1687.320 1732.290 1687.380 ;
        RECT 1389.285 1687.180 1732.290 1687.320 ;
        RECT 1389.285 1687.135 1389.575 1687.180 ;
        RECT 1731.970 1687.120 1732.290 1687.180 ;
      LAYER via ;
        RECT 1328.120 1687.120 1328.380 1687.380 ;
        RECT 1732.000 1687.120 1732.260 1687.380 ;
      LAYER met2 ;
        RECT 1328.020 1700.340 1328.300 1704.000 ;
        RECT 1328.020 1700.000 1328.320 1700.340 ;
        RECT 1328.180 1687.410 1328.320 1700.000 ;
        RECT 1328.120 1687.090 1328.380 1687.410 ;
        RECT 1732.000 1687.090 1732.260 1687.410 ;
        RECT 1732.060 17.410 1732.200 1687.090 ;
        RECT 1732.060 17.270 1733.580 17.410 ;
        RECT 1733.440 2.400 1733.580 17.270 ;
        RECT 1733.230 -4.800 1733.790 2.400 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1325.790 1685.280 1326.110 1685.340 ;
        RECT 1329.930 1685.280 1330.250 1685.340 ;
        RECT 1325.790 1685.140 1330.250 1685.280 ;
        RECT 1325.790 1685.080 1326.110 1685.140 ;
        RECT 1329.930 1685.080 1330.250 1685.140 ;
        RECT 1325.790 1619.320 1326.110 1619.380 ;
        RECT 1745.770 1619.320 1746.090 1619.380 ;
        RECT 1325.790 1619.180 1746.090 1619.320 ;
        RECT 1325.790 1619.120 1326.110 1619.180 ;
        RECT 1745.770 1619.120 1746.090 1619.180 ;
      LAYER via ;
        RECT 1325.820 1685.080 1326.080 1685.340 ;
        RECT 1329.960 1685.080 1330.220 1685.340 ;
        RECT 1325.820 1619.120 1326.080 1619.380 ;
        RECT 1745.800 1619.120 1746.060 1619.380 ;
      LAYER met2 ;
        RECT 1329.860 1700.340 1330.140 1704.000 ;
        RECT 1329.860 1700.000 1330.160 1700.340 ;
        RECT 1330.020 1685.370 1330.160 1700.000 ;
        RECT 1325.820 1685.050 1326.080 1685.370 ;
        RECT 1329.960 1685.050 1330.220 1685.370 ;
        RECT 1325.880 1619.410 1326.020 1685.050 ;
        RECT 1325.820 1619.090 1326.080 1619.410 ;
        RECT 1745.800 1619.090 1746.060 1619.410 ;
        RECT 1745.860 17.410 1746.000 1619.090 ;
        RECT 1745.860 17.270 1751.520 17.410 ;
        RECT 1751.380 2.400 1751.520 17.270 ;
        RECT 1751.170 -4.800 1751.730 2.400 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1331.770 1689.020 1332.090 1689.080 ;
        RECT 1334.990 1689.020 1335.310 1689.080 ;
        RECT 1331.770 1688.880 1335.310 1689.020 ;
        RECT 1331.770 1688.820 1332.090 1688.880 ;
        RECT 1334.990 1688.820 1335.310 1688.880 ;
        RECT 1334.990 1681.540 1335.310 1681.600 ;
        RECT 1766.470 1681.540 1766.790 1681.600 ;
        RECT 1334.990 1681.400 1766.790 1681.540 ;
        RECT 1334.990 1681.340 1335.310 1681.400 ;
        RECT 1766.470 1681.340 1766.790 1681.400 ;
      LAYER via ;
        RECT 1331.800 1688.820 1332.060 1689.080 ;
        RECT 1335.020 1688.820 1335.280 1689.080 ;
        RECT 1335.020 1681.340 1335.280 1681.600 ;
        RECT 1766.500 1681.340 1766.760 1681.600 ;
      LAYER met2 ;
        RECT 1331.700 1700.340 1331.980 1704.000 ;
        RECT 1331.700 1700.000 1332.000 1700.340 ;
        RECT 1331.860 1689.110 1332.000 1700.000 ;
        RECT 1331.800 1688.790 1332.060 1689.110 ;
        RECT 1335.020 1688.790 1335.280 1689.110 ;
        RECT 1335.080 1681.630 1335.220 1688.790 ;
        RECT 1335.020 1681.310 1335.280 1681.630 ;
        RECT 1766.500 1681.310 1766.760 1681.630 ;
        RECT 1766.560 6.530 1766.700 1681.310 ;
        RECT 1766.560 6.390 1769.000 6.530 ;
        RECT 1768.860 2.400 1769.000 6.390 ;
        RECT 1768.650 -4.800 1769.210 2.400 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1333.610 1685.280 1333.930 1685.340 ;
        RECT 1333.610 1685.140 1338.900 1685.280 ;
        RECT 1333.610 1685.080 1333.930 1685.140 ;
        RECT 1338.760 1684.600 1338.900 1685.140 ;
        RECT 1338.300 1684.460 1338.900 1684.600 ;
        RECT 1338.300 1684.320 1338.440 1684.460 ;
        RECT 1338.210 1684.060 1338.530 1684.320 ;
        RECT 1338.210 1660.800 1338.530 1660.860 ;
        RECT 1780.270 1660.800 1780.590 1660.860 ;
        RECT 1338.210 1660.660 1780.590 1660.800 ;
        RECT 1338.210 1660.600 1338.530 1660.660 ;
        RECT 1780.270 1660.600 1780.590 1660.660 ;
        RECT 1780.270 20.980 1780.590 21.040 ;
        RECT 1786.710 20.980 1787.030 21.040 ;
        RECT 1780.270 20.840 1787.030 20.980 ;
        RECT 1780.270 20.780 1780.590 20.840 ;
        RECT 1786.710 20.780 1787.030 20.840 ;
      LAYER via ;
        RECT 1333.640 1685.080 1333.900 1685.340 ;
        RECT 1338.240 1684.060 1338.500 1684.320 ;
        RECT 1338.240 1660.600 1338.500 1660.860 ;
        RECT 1780.300 1660.600 1780.560 1660.860 ;
        RECT 1780.300 20.780 1780.560 21.040 ;
        RECT 1786.740 20.780 1787.000 21.040 ;
      LAYER met2 ;
        RECT 1333.540 1700.340 1333.820 1704.000 ;
        RECT 1333.540 1700.000 1333.840 1700.340 ;
        RECT 1333.700 1685.370 1333.840 1700.000 ;
        RECT 1333.640 1685.050 1333.900 1685.370 ;
        RECT 1338.240 1684.030 1338.500 1684.350 ;
        RECT 1338.300 1660.890 1338.440 1684.030 ;
        RECT 1338.240 1660.570 1338.500 1660.890 ;
        RECT 1780.300 1660.570 1780.560 1660.890 ;
        RECT 1780.360 21.070 1780.500 1660.570 ;
        RECT 1780.300 20.750 1780.560 21.070 ;
        RECT 1786.740 20.750 1787.000 21.070 ;
        RECT 1786.800 2.400 1786.940 20.750 ;
        RECT 1786.590 -4.800 1787.150 2.400 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1333.150 1683.920 1333.470 1683.980 ;
        RECT 1335.450 1683.920 1335.770 1683.980 ;
        RECT 1333.150 1683.780 1335.770 1683.920 ;
        RECT 1333.150 1683.720 1333.470 1683.780 ;
        RECT 1335.450 1683.720 1335.770 1683.780 ;
        RECT 1333.150 1633.260 1333.470 1633.320 ;
        RECT 1800.970 1633.260 1801.290 1633.320 ;
        RECT 1333.150 1633.120 1801.290 1633.260 ;
        RECT 1333.150 1633.060 1333.470 1633.120 ;
        RECT 1800.970 1633.060 1801.290 1633.120 ;
      LAYER via ;
        RECT 1333.180 1683.720 1333.440 1683.980 ;
        RECT 1335.480 1683.720 1335.740 1683.980 ;
        RECT 1333.180 1633.060 1333.440 1633.320 ;
        RECT 1801.000 1633.060 1801.260 1633.320 ;
      LAYER met2 ;
        RECT 1335.380 1700.340 1335.660 1704.000 ;
        RECT 1335.380 1700.000 1335.680 1700.340 ;
        RECT 1335.540 1684.010 1335.680 1700.000 ;
        RECT 1333.180 1683.690 1333.440 1684.010 ;
        RECT 1335.480 1683.690 1335.740 1684.010 ;
        RECT 1333.240 1633.350 1333.380 1683.690 ;
        RECT 1333.180 1633.030 1333.440 1633.350 ;
        RECT 1801.000 1633.030 1801.260 1633.350 ;
        RECT 1801.060 17.410 1801.200 1633.030 ;
        RECT 1801.060 17.270 1804.880 17.410 ;
        RECT 1804.740 2.400 1804.880 17.270 ;
        RECT 1804.530 -4.800 1805.090 2.400 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1335.910 1683.920 1336.230 1683.980 ;
        RECT 1337.290 1683.920 1337.610 1683.980 ;
        RECT 1335.910 1683.780 1337.610 1683.920 ;
        RECT 1335.910 1683.720 1336.230 1683.780 ;
        RECT 1337.290 1683.720 1337.610 1683.780 ;
        RECT 1335.910 1584.640 1336.230 1584.700 ;
        RECT 1821.670 1584.640 1821.990 1584.700 ;
        RECT 1335.910 1584.500 1821.990 1584.640 ;
        RECT 1335.910 1584.440 1336.230 1584.500 ;
        RECT 1821.670 1584.440 1821.990 1584.500 ;
      LAYER via ;
        RECT 1335.940 1683.720 1336.200 1683.980 ;
        RECT 1337.320 1683.720 1337.580 1683.980 ;
        RECT 1335.940 1584.440 1336.200 1584.700 ;
        RECT 1821.700 1584.440 1821.960 1584.700 ;
      LAYER met2 ;
        RECT 1337.220 1700.340 1337.500 1704.000 ;
        RECT 1337.220 1700.000 1337.520 1700.340 ;
        RECT 1337.380 1684.010 1337.520 1700.000 ;
        RECT 1335.940 1683.690 1336.200 1684.010 ;
        RECT 1337.320 1683.690 1337.580 1684.010 ;
        RECT 1336.000 1584.730 1336.140 1683.690 ;
        RECT 1335.940 1584.410 1336.200 1584.730 ;
        RECT 1821.700 1584.410 1821.960 1584.730 ;
        RECT 1821.760 17.410 1821.900 1584.410 ;
        RECT 1821.760 17.270 1822.820 17.410 ;
        RECT 1822.680 2.400 1822.820 17.270 ;
        RECT 1822.470 -4.800 1823.030 2.400 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1339.130 1646.860 1339.450 1646.920 ;
        RECT 1835.470 1646.860 1835.790 1646.920 ;
        RECT 1339.130 1646.720 1835.790 1646.860 ;
        RECT 1339.130 1646.660 1339.450 1646.720 ;
        RECT 1835.470 1646.660 1835.790 1646.720 ;
      LAYER via ;
        RECT 1339.160 1646.660 1339.420 1646.920 ;
        RECT 1835.500 1646.660 1835.760 1646.920 ;
      LAYER met2 ;
        RECT 1339.060 1700.340 1339.340 1704.000 ;
        RECT 1339.060 1700.000 1339.360 1700.340 ;
        RECT 1339.220 1646.950 1339.360 1700.000 ;
        RECT 1339.160 1646.630 1339.420 1646.950 ;
        RECT 1835.500 1646.630 1835.760 1646.950 ;
        RECT 1835.560 17.410 1835.700 1646.630 ;
        RECT 1835.560 17.270 1840.300 17.410 ;
        RECT 1840.160 2.400 1840.300 17.270 ;
        RECT 1839.950 -4.800 1840.510 2.400 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1340.970 1598.240 1341.290 1598.300 ;
        RECT 1856.170 1598.240 1856.490 1598.300 ;
        RECT 1340.970 1598.100 1856.490 1598.240 ;
        RECT 1340.970 1598.040 1341.290 1598.100 ;
        RECT 1856.170 1598.040 1856.490 1598.100 ;
      LAYER via ;
        RECT 1341.000 1598.040 1341.260 1598.300 ;
        RECT 1856.200 1598.040 1856.460 1598.300 ;
      LAYER met2 ;
        RECT 1340.900 1700.340 1341.180 1704.000 ;
        RECT 1340.900 1700.000 1341.200 1700.340 ;
        RECT 1341.060 1598.330 1341.200 1700.000 ;
        RECT 1341.000 1598.010 1341.260 1598.330 ;
        RECT 1856.200 1598.010 1856.460 1598.330 ;
        RECT 1856.260 17.410 1856.400 1598.010 ;
        RECT 1856.260 17.270 1858.240 17.410 ;
        RECT 1858.100 2.400 1858.240 17.270 ;
        RECT 1857.890 -4.800 1858.450 2.400 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1341.430 1683.920 1341.750 1683.980 ;
        RECT 1342.810 1683.920 1343.130 1683.980 ;
        RECT 1341.430 1683.780 1343.130 1683.920 ;
        RECT 1341.430 1683.720 1341.750 1683.780 ;
        RECT 1342.810 1683.720 1343.130 1683.780 ;
        RECT 1341.430 1577.500 1341.750 1577.560 ;
        RECT 1869.970 1577.500 1870.290 1577.560 ;
        RECT 1341.430 1577.360 1870.290 1577.500 ;
        RECT 1341.430 1577.300 1341.750 1577.360 ;
        RECT 1869.970 1577.300 1870.290 1577.360 ;
        RECT 1869.970 20.980 1870.290 21.040 ;
        RECT 1875.950 20.980 1876.270 21.040 ;
        RECT 1869.970 20.840 1876.270 20.980 ;
        RECT 1869.970 20.780 1870.290 20.840 ;
        RECT 1875.950 20.780 1876.270 20.840 ;
      LAYER via ;
        RECT 1341.460 1683.720 1341.720 1683.980 ;
        RECT 1342.840 1683.720 1343.100 1683.980 ;
        RECT 1341.460 1577.300 1341.720 1577.560 ;
        RECT 1870.000 1577.300 1870.260 1577.560 ;
        RECT 1870.000 20.780 1870.260 21.040 ;
        RECT 1875.980 20.780 1876.240 21.040 ;
      LAYER met2 ;
        RECT 1342.740 1700.340 1343.020 1704.000 ;
        RECT 1342.740 1700.000 1343.040 1700.340 ;
        RECT 1342.900 1684.010 1343.040 1700.000 ;
        RECT 1341.460 1683.690 1341.720 1684.010 ;
        RECT 1342.840 1683.690 1343.100 1684.010 ;
        RECT 1341.520 1577.590 1341.660 1683.690 ;
        RECT 1341.460 1577.270 1341.720 1577.590 ;
        RECT 1870.000 1577.270 1870.260 1577.590 ;
        RECT 1870.060 21.070 1870.200 1577.270 ;
        RECT 1870.000 20.750 1870.260 21.070 ;
        RECT 1875.980 20.750 1876.240 21.070 ;
        RECT 1876.040 2.400 1876.180 20.750 ;
        RECT 1875.830 -4.800 1876.390 2.400 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 758.150 79.460 758.470 79.520 ;
        RECT 1225.970 79.460 1226.290 79.520 ;
        RECT 758.150 79.320 1226.290 79.460 ;
        RECT 758.150 79.260 758.470 79.320 ;
        RECT 1225.970 79.260 1226.290 79.320 ;
        RECT 752.170 20.980 752.490 21.040 ;
        RECT 758.150 20.980 758.470 21.040 ;
        RECT 752.170 20.840 758.470 20.980 ;
        RECT 752.170 20.780 752.490 20.840 ;
        RECT 758.150 20.780 758.470 20.840 ;
      LAYER via ;
        RECT 758.180 79.260 758.440 79.520 ;
        RECT 1226.000 79.260 1226.260 79.520 ;
        RECT 752.200 20.780 752.460 21.040 ;
        RECT 758.180 20.780 758.440 21.040 ;
      LAYER met2 ;
        RECT 1226.820 1700.340 1227.100 1704.000 ;
        RECT 1226.820 1700.000 1227.120 1700.340 ;
        RECT 1226.980 1666.410 1227.120 1700.000 ;
        RECT 1226.060 1666.270 1227.120 1666.410 ;
        RECT 1226.060 79.550 1226.200 1666.270 ;
        RECT 758.180 79.230 758.440 79.550 ;
        RECT 1226.000 79.230 1226.260 79.550 ;
        RECT 758.240 21.070 758.380 79.230 ;
        RECT 752.200 20.750 752.460 21.070 ;
        RECT 758.180 20.750 758.440 21.070 ;
        RECT 752.260 2.400 752.400 20.750 ;
        RECT 752.050 -4.800 752.610 2.400 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1343.270 1683.920 1343.590 1683.980 ;
        RECT 1344.650 1683.920 1344.970 1683.980 ;
        RECT 1343.270 1683.780 1344.970 1683.920 ;
        RECT 1343.270 1683.720 1343.590 1683.780 ;
        RECT 1344.650 1683.720 1344.970 1683.780 ;
        RECT 1343.270 1549.620 1343.590 1549.680 ;
        RECT 1890.670 1549.620 1890.990 1549.680 ;
        RECT 1343.270 1549.480 1890.990 1549.620 ;
        RECT 1343.270 1549.420 1343.590 1549.480 ;
        RECT 1890.670 1549.420 1890.990 1549.480 ;
      LAYER via ;
        RECT 1343.300 1683.720 1343.560 1683.980 ;
        RECT 1344.680 1683.720 1344.940 1683.980 ;
        RECT 1343.300 1549.420 1343.560 1549.680 ;
        RECT 1890.700 1549.420 1890.960 1549.680 ;
      LAYER met2 ;
        RECT 1344.580 1700.340 1344.860 1704.000 ;
        RECT 1344.580 1700.000 1344.880 1700.340 ;
        RECT 1344.740 1684.010 1344.880 1700.000 ;
        RECT 1343.300 1683.690 1343.560 1684.010 ;
        RECT 1344.680 1683.690 1344.940 1684.010 ;
        RECT 1343.360 1549.710 1343.500 1683.690 ;
        RECT 1343.300 1549.390 1343.560 1549.710 ;
        RECT 1890.700 1549.390 1890.960 1549.710 ;
        RECT 1890.760 17.410 1890.900 1549.390 ;
        RECT 1890.760 17.270 1894.120 17.410 ;
        RECT 1893.980 2.400 1894.120 17.270 ;
        RECT 1893.770 -4.800 1894.330 2.400 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1346.030 1654.000 1346.350 1654.060 ;
        RECT 1911.370 1654.000 1911.690 1654.060 ;
        RECT 1346.030 1653.860 1911.690 1654.000 ;
        RECT 1346.030 1653.800 1346.350 1653.860 ;
        RECT 1911.370 1653.800 1911.690 1653.860 ;
      LAYER via ;
        RECT 1346.060 1653.800 1346.320 1654.060 ;
        RECT 1911.400 1653.800 1911.660 1654.060 ;
      LAYER met2 ;
        RECT 1346.420 1700.340 1346.700 1704.000 ;
        RECT 1346.420 1700.000 1346.720 1700.340 ;
        RECT 1346.580 1684.770 1346.720 1700.000 ;
        RECT 1346.120 1684.630 1346.720 1684.770 ;
        RECT 1346.120 1654.090 1346.260 1684.630 ;
        RECT 1346.060 1653.770 1346.320 1654.090 ;
        RECT 1911.400 1653.770 1911.660 1654.090 ;
        RECT 1911.460 17.410 1911.600 1653.770 ;
        RECT 1911.460 17.270 1912.060 17.410 ;
        RECT 1911.920 2.400 1912.060 17.270 ;
        RECT 1911.710 -4.800 1912.270 2.400 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1348.330 1611.840 1348.650 1611.900 ;
        RECT 1925.170 1611.840 1925.490 1611.900 ;
        RECT 1348.330 1611.700 1925.490 1611.840 ;
        RECT 1348.330 1611.640 1348.650 1611.700 ;
        RECT 1925.170 1611.640 1925.490 1611.700 ;
      LAYER via ;
        RECT 1348.360 1611.640 1348.620 1611.900 ;
        RECT 1925.200 1611.640 1925.460 1611.900 ;
      LAYER met2 ;
        RECT 1348.260 1700.340 1348.540 1704.000 ;
        RECT 1348.260 1700.000 1348.560 1700.340 ;
        RECT 1348.420 1611.930 1348.560 1700.000 ;
        RECT 1348.360 1611.610 1348.620 1611.930 ;
        RECT 1925.200 1611.610 1925.460 1611.930 ;
        RECT 1925.260 17.410 1925.400 1611.610 ;
        RECT 1925.260 17.270 1929.540 17.410 ;
        RECT 1929.400 2.400 1929.540 17.270 ;
        RECT 1929.190 -4.800 1929.750 2.400 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1349.250 1570.700 1349.570 1570.760 ;
        RECT 1945.870 1570.700 1946.190 1570.760 ;
        RECT 1349.250 1570.560 1946.190 1570.700 ;
        RECT 1349.250 1570.500 1349.570 1570.560 ;
        RECT 1945.870 1570.500 1946.190 1570.560 ;
      LAYER via ;
        RECT 1349.280 1570.500 1349.540 1570.760 ;
        RECT 1945.900 1570.500 1946.160 1570.760 ;
      LAYER met2 ;
        RECT 1350.100 1700.410 1350.380 1704.000 ;
        RECT 1349.800 1700.270 1350.380 1700.410 ;
        RECT 1349.800 1677.970 1349.940 1700.270 ;
        RECT 1350.100 1700.000 1350.380 1700.270 ;
        RECT 1349.340 1677.830 1349.940 1677.970 ;
        RECT 1349.340 1570.790 1349.480 1677.830 ;
        RECT 1349.280 1570.470 1349.540 1570.790 ;
        RECT 1945.900 1570.470 1946.160 1570.790 ;
        RECT 1945.960 17.410 1946.100 1570.470 ;
        RECT 1945.960 17.270 1947.480 17.410 ;
        RECT 1947.340 2.400 1947.480 17.270 ;
        RECT 1947.130 -4.800 1947.690 2.400 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1347.870 1676.780 1348.190 1676.840 ;
        RECT 1351.550 1676.780 1351.870 1676.840 ;
        RECT 1347.870 1676.640 1351.870 1676.780 ;
        RECT 1347.870 1676.580 1348.190 1676.640 ;
        RECT 1351.550 1676.580 1351.870 1676.640 ;
        RECT 1347.870 14.180 1348.190 14.240 ;
        RECT 1965.190 14.180 1965.510 14.240 ;
        RECT 1347.870 14.040 1952.540 14.180 ;
        RECT 1347.870 13.980 1348.190 14.040 ;
        RECT 1952.400 13.840 1952.540 14.040 ;
        RECT 1959.760 14.040 1965.510 14.180 ;
        RECT 1959.760 13.840 1959.900 14.040 ;
        RECT 1965.190 13.980 1965.510 14.040 ;
        RECT 1952.400 13.700 1959.900 13.840 ;
      LAYER via ;
        RECT 1347.900 1676.580 1348.160 1676.840 ;
        RECT 1351.580 1676.580 1351.840 1676.840 ;
        RECT 1347.900 13.980 1348.160 14.240 ;
        RECT 1965.220 13.980 1965.480 14.240 ;
      LAYER met2 ;
        RECT 1351.940 1700.410 1352.220 1704.000 ;
        RECT 1351.640 1700.270 1352.220 1700.410 ;
        RECT 1351.640 1676.870 1351.780 1700.270 ;
        RECT 1351.940 1700.000 1352.220 1700.270 ;
        RECT 1347.900 1676.550 1348.160 1676.870 ;
        RECT 1351.580 1676.550 1351.840 1676.870 ;
        RECT 1347.960 14.270 1348.100 1676.550 ;
        RECT 1347.900 13.950 1348.160 14.270 ;
        RECT 1965.220 13.950 1965.480 14.270 ;
        RECT 1965.280 2.400 1965.420 13.950 ;
        RECT 1965.070 -4.800 1965.630 2.400 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1354.845 1055.785 1355.015 1103.895 ;
        RECT 1354.845 910.945 1355.015 959.055 ;
        RECT 1353.925 855.525 1354.095 903.975 ;
      LAYER mcon ;
        RECT 1354.845 1103.725 1355.015 1103.895 ;
        RECT 1354.845 958.885 1355.015 959.055 ;
        RECT 1353.925 903.805 1354.095 903.975 ;
      LAYER met1 ;
        RECT 1354.310 1345.620 1354.630 1345.680 ;
        RECT 1354.770 1345.620 1355.090 1345.680 ;
        RECT 1354.310 1345.480 1355.090 1345.620 ;
        RECT 1354.310 1345.420 1354.630 1345.480 ;
        RECT 1354.770 1345.420 1355.090 1345.480 ;
        RECT 1353.850 1297.340 1354.170 1297.400 ;
        RECT 1354.770 1297.340 1355.090 1297.400 ;
        RECT 1353.850 1297.200 1355.090 1297.340 ;
        RECT 1353.850 1297.140 1354.170 1297.200 ;
        RECT 1354.770 1297.140 1355.090 1297.200 ;
        RECT 1353.850 1200.780 1354.170 1200.840 ;
        RECT 1354.770 1200.780 1355.090 1200.840 ;
        RECT 1353.850 1200.640 1355.090 1200.780 ;
        RECT 1353.850 1200.580 1354.170 1200.640 ;
        RECT 1354.770 1200.580 1355.090 1200.640 ;
        RECT 1354.770 1103.880 1355.090 1103.940 ;
        RECT 1354.575 1103.740 1355.090 1103.880 ;
        RECT 1354.770 1103.680 1355.090 1103.740 ;
        RECT 1354.770 1055.940 1355.090 1056.000 ;
        RECT 1354.575 1055.800 1355.090 1055.940 ;
        RECT 1354.770 1055.740 1355.090 1055.800 ;
        RECT 1354.770 959.040 1355.090 959.100 ;
        RECT 1354.575 958.900 1355.090 959.040 ;
        RECT 1354.770 958.840 1355.090 958.900 ;
        RECT 1354.770 911.100 1355.090 911.160 ;
        RECT 1354.575 910.960 1355.090 911.100 ;
        RECT 1354.770 910.900 1355.090 910.960 ;
        RECT 1353.865 903.960 1354.155 904.005 ;
        RECT 1354.770 903.960 1355.090 904.020 ;
        RECT 1353.865 903.820 1355.090 903.960 ;
        RECT 1353.865 903.775 1354.155 903.820 ;
        RECT 1354.770 903.760 1355.090 903.820 ;
        RECT 1353.850 855.680 1354.170 855.740 ;
        RECT 1353.655 855.540 1354.170 855.680 ;
        RECT 1353.850 855.480 1354.170 855.540 ;
        RECT 1354.770 593.340 1355.090 593.600 ;
        RECT 1354.860 592.920 1355.000 593.340 ;
        RECT 1354.770 592.660 1355.090 592.920 ;
        RECT 1354.770 14.520 1355.090 14.580 ;
        RECT 1983.130 14.520 1983.450 14.580 ;
        RECT 1354.770 14.380 1983.450 14.520 ;
        RECT 1354.770 14.320 1355.090 14.380 ;
        RECT 1983.130 14.320 1983.450 14.380 ;
      LAYER via ;
        RECT 1354.340 1345.420 1354.600 1345.680 ;
        RECT 1354.800 1345.420 1355.060 1345.680 ;
        RECT 1353.880 1297.140 1354.140 1297.400 ;
        RECT 1354.800 1297.140 1355.060 1297.400 ;
        RECT 1353.880 1200.580 1354.140 1200.840 ;
        RECT 1354.800 1200.580 1355.060 1200.840 ;
        RECT 1354.800 1103.680 1355.060 1103.940 ;
        RECT 1354.800 1055.740 1355.060 1056.000 ;
        RECT 1354.800 958.840 1355.060 959.100 ;
        RECT 1354.800 910.900 1355.060 911.160 ;
        RECT 1354.800 903.760 1355.060 904.020 ;
        RECT 1353.880 855.480 1354.140 855.740 ;
        RECT 1354.800 593.340 1355.060 593.600 ;
        RECT 1354.800 592.660 1355.060 592.920 ;
        RECT 1354.800 14.320 1355.060 14.580 ;
        RECT 1983.160 14.320 1983.420 14.580 ;
      LAYER met2 ;
        RECT 1353.780 1701.090 1354.060 1704.000 ;
        RECT 1353.480 1700.950 1354.060 1701.090 ;
        RECT 1353.480 1685.565 1353.620 1700.950 ;
        RECT 1353.780 1700.000 1354.060 1700.950 ;
        RECT 1353.410 1685.195 1353.690 1685.565 ;
        RECT 1353.870 1683.665 1354.150 1684.035 ;
        RECT 1353.940 1611.330 1354.080 1683.665 ;
        RECT 1353.940 1611.190 1355.000 1611.330 ;
        RECT 1354.860 1393.730 1355.000 1611.190 ;
        RECT 1354.400 1393.590 1355.000 1393.730 ;
        RECT 1354.400 1345.710 1354.540 1393.590 ;
        RECT 1353.870 1345.195 1354.150 1345.565 ;
        RECT 1354.340 1345.390 1354.600 1345.710 ;
        RECT 1354.800 1345.565 1355.060 1345.710 ;
        RECT 1354.790 1345.195 1355.070 1345.565 ;
        RECT 1353.940 1297.430 1354.080 1345.195 ;
        RECT 1353.880 1297.110 1354.140 1297.430 ;
        RECT 1354.800 1297.110 1355.060 1297.430 ;
        RECT 1354.860 1249.005 1355.000 1297.110 ;
        RECT 1353.870 1248.635 1354.150 1249.005 ;
        RECT 1354.790 1248.635 1355.070 1249.005 ;
        RECT 1353.940 1200.870 1354.080 1248.635 ;
        RECT 1353.880 1200.550 1354.140 1200.870 ;
        RECT 1354.800 1200.550 1355.060 1200.870 ;
        RECT 1354.860 1103.970 1355.000 1200.550 ;
        RECT 1354.800 1103.650 1355.060 1103.970 ;
        RECT 1354.800 1055.710 1355.060 1056.030 ;
        RECT 1354.860 959.130 1355.000 1055.710 ;
        RECT 1354.800 958.810 1355.060 959.130 ;
        RECT 1354.800 910.870 1355.060 911.190 ;
        RECT 1354.860 904.050 1355.000 910.870 ;
        RECT 1354.800 903.730 1355.060 904.050 ;
        RECT 1353.880 855.450 1354.140 855.770 ;
        RECT 1353.940 814.485 1354.080 855.450 ;
        RECT 1353.870 814.115 1354.150 814.485 ;
        RECT 1353.870 812.755 1354.150 813.125 ;
        RECT 1353.940 766.205 1354.080 812.755 ;
        RECT 1353.870 765.835 1354.150 766.205 ;
        RECT 1354.790 765.835 1355.070 766.205 ;
        RECT 1354.860 593.630 1355.000 765.835 ;
        RECT 1354.800 593.310 1355.060 593.630 ;
        RECT 1354.800 592.630 1355.060 592.950 ;
        RECT 1354.860 14.610 1355.000 592.630 ;
        RECT 1354.800 14.290 1355.060 14.610 ;
        RECT 1983.160 14.290 1983.420 14.610 ;
        RECT 1983.220 2.400 1983.360 14.290 ;
        RECT 1983.010 -4.800 1983.570 2.400 ;
      LAYER via2 ;
        RECT 1353.410 1685.240 1353.690 1685.520 ;
        RECT 1353.870 1683.710 1354.150 1683.990 ;
        RECT 1353.870 1345.240 1354.150 1345.520 ;
        RECT 1354.790 1345.240 1355.070 1345.520 ;
        RECT 1353.870 1248.680 1354.150 1248.960 ;
        RECT 1354.790 1248.680 1355.070 1248.960 ;
        RECT 1353.870 814.160 1354.150 814.440 ;
        RECT 1353.870 812.800 1354.150 813.080 ;
        RECT 1353.870 765.880 1354.150 766.160 ;
        RECT 1354.790 765.880 1355.070 766.160 ;
      LAYER met3 ;
        RECT 1353.385 1685.530 1353.715 1685.545 ;
        RECT 1353.385 1685.230 1354.850 1685.530 ;
        RECT 1353.385 1685.215 1353.715 1685.230 ;
        RECT 1353.845 1684.000 1354.175 1684.015 ;
        RECT 1354.550 1684.000 1354.850 1685.230 ;
        RECT 1353.845 1683.700 1354.850 1684.000 ;
        RECT 1353.845 1683.685 1354.175 1683.700 ;
        RECT 1353.845 1345.530 1354.175 1345.545 ;
        RECT 1354.765 1345.530 1355.095 1345.545 ;
        RECT 1353.845 1345.230 1355.095 1345.530 ;
        RECT 1353.845 1345.215 1354.175 1345.230 ;
        RECT 1354.765 1345.215 1355.095 1345.230 ;
        RECT 1353.845 1248.970 1354.175 1248.985 ;
        RECT 1354.765 1248.970 1355.095 1248.985 ;
        RECT 1353.845 1248.670 1355.095 1248.970 ;
        RECT 1353.845 1248.655 1354.175 1248.670 ;
        RECT 1354.765 1248.655 1355.095 1248.670 ;
        RECT 1353.845 814.450 1354.175 814.465 ;
        RECT 1353.845 814.150 1354.850 814.450 ;
        RECT 1353.845 814.135 1354.175 814.150 ;
        RECT 1353.845 813.090 1354.175 813.105 ;
        RECT 1354.550 813.090 1354.850 814.150 ;
        RECT 1353.845 812.790 1354.850 813.090 ;
        RECT 1353.845 812.775 1354.175 812.790 ;
        RECT 1353.845 766.170 1354.175 766.185 ;
        RECT 1354.765 766.170 1355.095 766.185 ;
        RECT 1353.845 765.870 1355.095 766.170 ;
        RECT 1353.845 765.855 1354.175 765.870 ;
        RECT 1354.765 765.855 1355.095 765.870 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1353.465 1683.765 1353.635 1687.675 ;
      LAYER mcon ;
        RECT 1353.465 1687.505 1353.635 1687.675 ;
      LAYER met1 ;
        RECT 1353.405 1687.660 1353.695 1687.705 ;
        RECT 1355.690 1687.660 1356.010 1687.720 ;
        RECT 1353.405 1687.520 1356.010 1687.660 ;
        RECT 1353.405 1687.475 1353.695 1687.520 ;
        RECT 1355.690 1687.460 1356.010 1687.520 ;
        RECT 1353.390 1683.920 1353.710 1683.980 ;
        RECT 1353.195 1683.780 1353.710 1683.920 ;
        RECT 1353.390 1683.720 1353.710 1683.780 ;
        RECT 1353.390 14.860 1353.710 14.920 ;
        RECT 2001.070 14.860 2001.390 14.920 ;
        RECT 1353.390 14.720 2001.390 14.860 ;
        RECT 1353.390 14.660 1353.710 14.720 ;
        RECT 2001.070 14.660 2001.390 14.720 ;
      LAYER via ;
        RECT 1355.720 1687.460 1355.980 1687.720 ;
        RECT 1353.420 1683.720 1353.680 1683.980 ;
        RECT 1353.420 14.660 1353.680 14.920 ;
        RECT 2001.100 14.660 2001.360 14.920 ;
      LAYER met2 ;
        RECT 1355.620 1700.340 1355.900 1704.000 ;
        RECT 1355.620 1700.000 1355.920 1700.340 ;
        RECT 1355.780 1687.750 1355.920 1700.000 ;
        RECT 1355.720 1687.430 1355.980 1687.750 ;
        RECT 1353.420 1683.690 1353.680 1684.010 ;
        RECT 1353.480 14.950 1353.620 1683.690 ;
        RECT 1353.420 14.630 1353.680 14.950 ;
        RECT 2001.100 14.630 2001.360 14.950 ;
        RECT 2001.160 2.400 2001.300 14.630 ;
        RECT 2000.950 -4.800 2001.510 2.400 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1355.230 1683.920 1355.550 1683.980 ;
        RECT 1357.530 1683.920 1357.850 1683.980 ;
        RECT 1355.230 1683.780 1357.850 1683.920 ;
        RECT 1355.230 1683.720 1355.550 1683.780 ;
        RECT 1357.530 1683.720 1357.850 1683.780 ;
        RECT 1355.230 15.200 1355.550 15.260 ;
        RECT 2018.550 15.200 2018.870 15.260 ;
        RECT 1355.230 15.060 2018.870 15.200 ;
        RECT 1355.230 15.000 1355.550 15.060 ;
        RECT 2018.550 15.000 2018.870 15.060 ;
      LAYER via ;
        RECT 1355.260 1683.720 1355.520 1683.980 ;
        RECT 1357.560 1683.720 1357.820 1683.980 ;
        RECT 1355.260 15.000 1355.520 15.260 ;
        RECT 2018.580 15.000 2018.840 15.260 ;
      LAYER met2 ;
        RECT 1357.460 1700.340 1357.740 1704.000 ;
        RECT 1357.460 1700.000 1357.760 1700.340 ;
        RECT 1357.620 1684.010 1357.760 1700.000 ;
        RECT 1355.260 1683.690 1355.520 1684.010 ;
        RECT 1357.560 1683.690 1357.820 1684.010 ;
        RECT 1355.320 15.290 1355.460 1683.690 ;
        RECT 1355.260 14.970 1355.520 15.290 ;
        RECT 2018.580 14.970 2018.840 15.290 ;
        RECT 2018.640 2.400 2018.780 14.970 ;
        RECT 2018.430 -4.800 2018.990 2.400 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1359.370 1684.260 1359.690 1684.320 ;
        RECT 1360.750 1684.260 1361.070 1684.320 ;
        RECT 1359.370 1684.120 1361.070 1684.260 ;
        RECT 1359.370 1684.060 1359.690 1684.120 ;
        RECT 1360.750 1684.060 1361.070 1684.120 ;
        RECT 1361.210 15.540 1361.530 15.600 ;
        RECT 2036.490 15.540 2036.810 15.600 ;
        RECT 1361.210 15.400 2036.810 15.540 ;
        RECT 1361.210 15.340 1361.530 15.400 ;
        RECT 2036.490 15.340 2036.810 15.400 ;
      LAYER via ;
        RECT 1359.400 1684.060 1359.660 1684.320 ;
        RECT 1360.780 1684.060 1361.040 1684.320 ;
        RECT 1361.240 15.340 1361.500 15.600 ;
        RECT 2036.520 15.340 2036.780 15.600 ;
      LAYER met2 ;
        RECT 1359.300 1700.340 1359.580 1704.000 ;
        RECT 1359.300 1700.000 1359.600 1700.340 ;
        RECT 1359.460 1684.350 1359.600 1700.000 ;
        RECT 1359.400 1684.030 1359.660 1684.350 ;
        RECT 1360.780 1684.030 1361.040 1684.350 ;
        RECT 1360.840 1677.970 1360.980 1684.030 ;
        RECT 1360.840 1677.830 1361.440 1677.970 ;
        RECT 1361.300 15.630 1361.440 1677.830 ;
        RECT 1361.240 15.310 1361.500 15.630 ;
        RECT 2036.520 15.310 2036.780 15.630 ;
        RECT 2036.580 2.400 2036.720 15.310 ;
        RECT 2036.370 -4.800 2036.930 2.400 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1359.830 1683.920 1360.150 1683.980 ;
        RECT 1361.210 1683.920 1361.530 1683.980 ;
        RECT 1359.830 1683.780 1361.530 1683.920 ;
        RECT 1359.830 1683.720 1360.150 1683.780 ;
        RECT 1361.210 1683.720 1361.530 1683.780 ;
        RECT 1359.830 15.880 1360.150 15.940 ;
        RECT 2054.430 15.880 2054.750 15.940 ;
        RECT 1359.830 15.740 2054.750 15.880 ;
        RECT 1359.830 15.680 1360.150 15.740 ;
        RECT 2054.430 15.680 2054.750 15.740 ;
      LAYER via ;
        RECT 1359.860 1683.720 1360.120 1683.980 ;
        RECT 1361.240 1683.720 1361.500 1683.980 ;
        RECT 1359.860 15.680 1360.120 15.940 ;
        RECT 2054.460 15.680 2054.720 15.940 ;
      LAYER met2 ;
        RECT 1361.140 1700.340 1361.420 1704.000 ;
        RECT 1361.140 1700.000 1361.440 1700.340 ;
        RECT 1361.300 1684.010 1361.440 1700.000 ;
        RECT 1359.860 1683.690 1360.120 1684.010 ;
        RECT 1361.240 1683.690 1361.500 1684.010 ;
        RECT 1359.920 15.970 1360.060 1683.690 ;
        RECT 1359.860 15.650 1360.120 15.970 ;
        RECT 2054.460 15.650 2054.720 15.970 ;
        RECT 2054.520 2.400 2054.660 15.650 ;
        RECT 2054.310 -4.800 2054.870 2.400 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1228.730 1678.280 1229.050 1678.540 ;
        RECT 1228.820 1677.800 1228.960 1678.280 ;
        RECT 1228.820 1677.660 1232.180 1677.800 ;
        RECT 1232.040 1677.520 1232.180 1677.660 ;
        RECT 1231.950 1677.260 1232.270 1677.520 ;
        RECT 772.410 1597.900 772.730 1597.960 ;
        RECT 1231.950 1597.900 1232.270 1597.960 ;
        RECT 772.410 1597.760 1232.270 1597.900 ;
        RECT 772.410 1597.700 772.730 1597.760 ;
        RECT 1231.950 1597.700 1232.270 1597.760 ;
      LAYER via ;
        RECT 1228.760 1678.280 1229.020 1678.540 ;
        RECT 1231.980 1677.260 1232.240 1677.520 ;
        RECT 772.440 1597.700 772.700 1597.960 ;
        RECT 1231.980 1597.700 1232.240 1597.960 ;
      LAYER met2 ;
        RECT 1228.660 1700.340 1228.940 1704.000 ;
        RECT 1228.660 1700.000 1228.960 1700.340 ;
        RECT 1228.820 1678.570 1228.960 1700.000 ;
        RECT 1228.760 1678.250 1229.020 1678.570 ;
        RECT 1231.980 1677.230 1232.240 1677.550 ;
        RECT 1232.040 1597.990 1232.180 1677.230 ;
        RECT 772.440 1597.670 772.700 1597.990 ;
        RECT 1231.980 1597.670 1232.240 1597.990 ;
        RECT 772.500 18.090 772.640 1597.670 ;
        RECT 769.740 17.950 772.640 18.090 ;
        RECT 769.740 2.400 769.880 17.950 ;
        RECT 769.530 -4.800 770.090 2.400 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1362.205 559.045 1362.375 607.155 ;
        RECT 1361.745 510.765 1361.915 558.535 ;
        RECT 1361.745 372.725 1361.915 486.455 ;
      LAYER mcon ;
        RECT 1362.205 606.985 1362.375 607.155 ;
        RECT 1361.745 558.365 1361.915 558.535 ;
        RECT 1361.745 486.285 1361.915 486.455 ;
      LAYER met1 ;
        RECT 1362.130 1587.360 1362.450 1587.420 ;
        RECT 1363.050 1587.360 1363.370 1587.420 ;
        RECT 1362.130 1587.220 1363.370 1587.360 ;
        RECT 1362.130 1587.160 1362.450 1587.220 ;
        RECT 1363.050 1587.160 1363.370 1587.220 ;
        RECT 1362.130 1366.700 1362.450 1366.760 ;
        RECT 1361.760 1366.560 1362.450 1366.700 ;
        RECT 1361.760 1366.080 1361.900 1366.560 ;
        RECT 1362.130 1366.500 1362.450 1366.560 ;
        RECT 1361.670 1365.820 1361.990 1366.080 ;
        RECT 1361.670 1207.580 1361.990 1207.640 ;
        RECT 1362.130 1207.580 1362.450 1207.640 ;
        RECT 1361.670 1207.440 1362.450 1207.580 ;
        RECT 1361.670 1207.380 1361.990 1207.440 ;
        RECT 1362.130 1207.380 1362.450 1207.440 ;
        RECT 1362.130 1077.020 1362.450 1077.080 ;
        RECT 1361.760 1076.880 1362.450 1077.020 ;
        RECT 1361.760 1076.400 1361.900 1076.880 ;
        RECT 1362.130 1076.820 1362.450 1076.880 ;
        RECT 1361.670 1076.140 1361.990 1076.400 ;
        RECT 1361.670 627.880 1361.990 627.940 ;
        RECT 1362.130 627.880 1362.450 627.940 ;
        RECT 1361.670 627.740 1362.450 627.880 ;
        RECT 1361.670 627.680 1361.990 627.740 ;
        RECT 1362.130 627.680 1362.450 627.740 ;
        RECT 1362.130 620.740 1362.450 620.800 ;
        RECT 1363.050 620.740 1363.370 620.800 ;
        RECT 1362.130 620.600 1363.370 620.740 ;
        RECT 1362.130 620.540 1362.450 620.600 ;
        RECT 1363.050 620.540 1363.370 620.600 ;
        RECT 1362.145 607.140 1362.435 607.185 ;
        RECT 1363.050 607.140 1363.370 607.200 ;
        RECT 1362.145 607.000 1363.370 607.140 ;
        RECT 1362.145 606.955 1362.435 607.000 ;
        RECT 1363.050 606.940 1363.370 607.000 ;
        RECT 1362.130 559.200 1362.450 559.260 ;
        RECT 1361.935 559.060 1362.450 559.200 ;
        RECT 1362.130 559.000 1362.450 559.060 ;
        RECT 1361.685 558.520 1361.975 558.565 ;
        RECT 1362.130 558.520 1362.450 558.580 ;
        RECT 1361.685 558.380 1362.450 558.520 ;
        RECT 1361.685 558.335 1361.975 558.380 ;
        RECT 1362.130 558.320 1362.450 558.380 ;
        RECT 1361.670 510.920 1361.990 510.980 ;
        RECT 1361.475 510.780 1361.990 510.920 ;
        RECT 1361.670 510.720 1361.990 510.780 ;
        RECT 1361.685 486.440 1361.975 486.485 ;
        RECT 1362.130 486.440 1362.450 486.500 ;
        RECT 1361.685 486.300 1362.450 486.440 ;
        RECT 1361.685 486.255 1361.975 486.300 ;
        RECT 1362.130 486.240 1362.450 486.300 ;
        RECT 1361.670 372.880 1361.990 372.940 ;
        RECT 1361.475 372.740 1361.990 372.880 ;
        RECT 1361.670 372.680 1361.990 372.740 ;
        RECT 1362.130 324.260 1362.450 324.320 ;
        RECT 1361.760 324.120 1362.450 324.260 ;
        RECT 1361.760 323.980 1361.900 324.120 ;
        RECT 1362.130 324.060 1362.450 324.120 ;
        RECT 1361.670 323.720 1361.990 323.980 ;
        RECT 1361.670 16.220 1361.990 16.280 ;
        RECT 2072.370 16.220 2072.690 16.280 ;
        RECT 1361.670 16.080 2072.690 16.220 ;
        RECT 1361.670 16.020 1361.990 16.080 ;
        RECT 2072.370 16.020 2072.690 16.080 ;
      LAYER via ;
        RECT 1362.160 1587.160 1362.420 1587.420 ;
        RECT 1363.080 1587.160 1363.340 1587.420 ;
        RECT 1362.160 1366.500 1362.420 1366.760 ;
        RECT 1361.700 1365.820 1361.960 1366.080 ;
        RECT 1361.700 1207.380 1361.960 1207.640 ;
        RECT 1362.160 1207.380 1362.420 1207.640 ;
        RECT 1362.160 1076.820 1362.420 1077.080 ;
        RECT 1361.700 1076.140 1361.960 1076.400 ;
        RECT 1361.700 627.680 1361.960 627.940 ;
        RECT 1362.160 627.680 1362.420 627.940 ;
        RECT 1362.160 620.540 1362.420 620.800 ;
        RECT 1363.080 620.540 1363.340 620.800 ;
        RECT 1363.080 606.940 1363.340 607.200 ;
        RECT 1362.160 559.000 1362.420 559.260 ;
        RECT 1362.160 558.320 1362.420 558.580 ;
        RECT 1361.700 510.720 1361.960 510.980 ;
        RECT 1362.160 486.240 1362.420 486.500 ;
        RECT 1361.700 372.680 1361.960 372.940 ;
        RECT 1362.160 324.060 1362.420 324.320 ;
        RECT 1361.700 323.720 1361.960 323.980 ;
        RECT 1361.700 16.020 1361.960 16.280 ;
        RECT 2072.400 16.020 2072.660 16.280 ;
      LAYER met2 ;
        RECT 1362.980 1700.340 1363.260 1704.000 ;
        RECT 1362.980 1700.000 1363.280 1700.340 ;
        RECT 1363.140 1587.450 1363.280 1700.000 ;
        RECT 1362.160 1587.130 1362.420 1587.450 ;
        RECT 1363.080 1587.130 1363.340 1587.450 ;
        RECT 1362.220 1366.790 1362.360 1587.130 ;
        RECT 1362.160 1366.470 1362.420 1366.790 ;
        RECT 1361.700 1365.790 1361.960 1366.110 ;
        RECT 1361.760 1207.670 1361.900 1365.790 ;
        RECT 1361.700 1207.350 1361.960 1207.670 ;
        RECT 1362.160 1207.350 1362.420 1207.670 ;
        RECT 1362.220 1077.110 1362.360 1207.350 ;
        RECT 1362.160 1076.790 1362.420 1077.110 ;
        RECT 1361.700 1076.110 1361.960 1076.430 ;
        RECT 1361.760 869.565 1361.900 1076.110 ;
        RECT 1360.770 869.195 1361.050 869.565 ;
        RECT 1361.690 869.195 1361.970 869.565 ;
        RECT 1360.840 821.285 1360.980 869.195 ;
        RECT 1360.770 820.915 1361.050 821.285 ;
        RECT 1361.690 820.915 1361.970 821.285 ;
        RECT 1361.760 786.490 1361.900 820.915 ;
        RECT 1361.760 786.350 1362.360 786.490 ;
        RECT 1362.220 651.850 1362.360 786.350 ;
        RECT 1361.760 651.710 1362.360 651.850 ;
        RECT 1361.760 627.970 1361.900 651.710 ;
        RECT 1361.700 627.650 1361.960 627.970 ;
        RECT 1362.160 627.650 1362.420 627.970 ;
        RECT 1362.220 620.830 1362.360 627.650 ;
        RECT 1362.160 620.510 1362.420 620.830 ;
        RECT 1363.080 620.510 1363.340 620.830 ;
        RECT 1363.140 607.230 1363.280 620.510 ;
        RECT 1363.080 606.910 1363.340 607.230 ;
        RECT 1362.160 558.970 1362.420 559.290 ;
        RECT 1362.220 558.610 1362.360 558.970 ;
        RECT 1362.160 558.290 1362.420 558.610 ;
        RECT 1361.700 510.690 1361.960 511.010 ;
        RECT 1361.760 510.410 1361.900 510.690 ;
        RECT 1361.760 510.270 1362.360 510.410 ;
        RECT 1362.220 486.530 1362.360 510.270 ;
        RECT 1362.160 486.210 1362.420 486.530 ;
        RECT 1361.700 372.650 1361.960 372.970 ;
        RECT 1361.760 372.485 1361.900 372.650 ;
        RECT 1360.770 372.115 1361.050 372.485 ;
        RECT 1361.690 372.115 1361.970 372.485 ;
        RECT 1360.840 324.885 1360.980 372.115 ;
        RECT 1360.770 324.515 1361.050 324.885 ;
        RECT 1362.150 324.515 1362.430 324.885 ;
        RECT 1362.220 324.350 1362.360 324.515 ;
        RECT 1362.160 324.030 1362.420 324.350 ;
        RECT 1361.700 323.690 1361.960 324.010 ;
        RECT 1361.760 16.310 1361.900 323.690 ;
        RECT 1361.700 15.990 1361.960 16.310 ;
        RECT 2072.400 15.990 2072.660 16.310 ;
        RECT 2072.460 2.400 2072.600 15.990 ;
        RECT 2072.250 -4.800 2072.810 2.400 ;
      LAYER via2 ;
        RECT 1360.770 869.240 1361.050 869.520 ;
        RECT 1361.690 869.240 1361.970 869.520 ;
        RECT 1360.770 820.960 1361.050 821.240 ;
        RECT 1361.690 820.960 1361.970 821.240 ;
        RECT 1360.770 372.160 1361.050 372.440 ;
        RECT 1361.690 372.160 1361.970 372.440 ;
        RECT 1360.770 324.560 1361.050 324.840 ;
        RECT 1362.150 324.560 1362.430 324.840 ;
      LAYER met3 ;
        RECT 1360.745 869.530 1361.075 869.545 ;
        RECT 1361.665 869.530 1361.995 869.545 ;
        RECT 1360.745 869.230 1361.995 869.530 ;
        RECT 1360.745 869.215 1361.075 869.230 ;
        RECT 1361.665 869.215 1361.995 869.230 ;
        RECT 1360.745 821.250 1361.075 821.265 ;
        RECT 1361.665 821.250 1361.995 821.265 ;
        RECT 1360.745 820.950 1361.995 821.250 ;
        RECT 1360.745 820.935 1361.075 820.950 ;
        RECT 1361.665 820.935 1361.995 820.950 ;
        RECT 1360.745 372.450 1361.075 372.465 ;
        RECT 1361.665 372.450 1361.995 372.465 ;
        RECT 1360.745 372.150 1361.995 372.450 ;
        RECT 1360.745 372.135 1361.075 372.150 ;
        RECT 1361.665 372.135 1361.995 372.150 ;
        RECT 1360.745 324.850 1361.075 324.865 ;
        RECT 1362.125 324.850 1362.455 324.865 ;
        RECT 1360.745 324.550 1362.455 324.850 ;
        RECT 1360.745 324.535 1361.075 324.550 ;
        RECT 1362.125 324.535 1362.455 324.550 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1364.890 16.560 1365.210 16.620 ;
        RECT 2089.850 16.560 2090.170 16.620 ;
        RECT 1364.890 16.420 2090.170 16.560 ;
        RECT 1364.890 16.360 1365.210 16.420 ;
        RECT 2089.850 16.360 2090.170 16.420 ;
      LAYER via ;
        RECT 1364.920 16.360 1365.180 16.620 ;
        RECT 2089.880 16.360 2090.140 16.620 ;
      LAYER met2 ;
        RECT 1364.820 1700.340 1365.100 1704.000 ;
        RECT 1364.820 1700.000 1365.120 1700.340 ;
        RECT 1364.980 16.650 1365.120 1700.000 ;
        RECT 1364.920 16.330 1365.180 16.650 ;
        RECT 2089.880 16.330 2090.140 16.650 ;
        RECT 2089.940 2.400 2090.080 16.330 ;
        RECT 2089.730 -4.800 2090.290 2.400 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1366.730 1685.280 1367.050 1685.340 ;
        RECT 1371.790 1685.280 1372.110 1685.340 ;
        RECT 1366.730 1685.140 1372.110 1685.280 ;
        RECT 1366.730 1685.080 1367.050 1685.140 ;
        RECT 1371.790 1685.080 1372.110 1685.140 ;
        RECT 1369.030 1631.900 1369.350 1631.960 ;
        RECT 1371.790 1631.900 1372.110 1631.960 ;
        RECT 1369.030 1631.760 1372.110 1631.900 ;
        RECT 1369.030 1631.700 1369.350 1631.760 ;
        RECT 1371.790 1631.700 1372.110 1631.760 ;
        RECT 1369.030 16.900 1369.350 16.960 ;
        RECT 2107.790 16.900 2108.110 16.960 ;
        RECT 1369.030 16.760 2108.110 16.900 ;
        RECT 1369.030 16.700 1369.350 16.760 ;
        RECT 2107.790 16.700 2108.110 16.760 ;
      LAYER via ;
        RECT 1366.760 1685.080 1367.020 1685.340 ;
        RECT 1371.820 1685.080 1372.080 1685.340 ;
        RECT 1369.060 1631.700 1369.320 1631.960 ;
        RECT 1371.820 1631.700 1372.080 1631.960 ;
        RECT 1369.060 16.700 1369.320 16.960 ;
        RECT 2107.820 16.700 2108.080 16.960 ;
      LAYER met2 ;
        RECT 1366.660 1700.340 1366.940 1704.000 ;
        RECT 1366.660 1700.000 1366.960 1700.340 ;
        RECT 1366.820 1685.370 1366.960 1700.000 ;
        RECT 1366.760 1685.050 1367.020 1685.370 ;
        RECT 1371.820 1685.050 1372.080 1685.370 ;
        RECT 1371.880 1631.990 1372.020 1685.050 ;
        RECT 1369.060 1631.670 1369.320 1631.990 ;
        RECT 1371.820 1631.670 1372.080 1631.990 ;
        RECT 1369.120 16.990 1369.260 1631.670 ;
        RECT 1369.060 16.670 1369.320 16.990 ;
        RECT 2107.820 16.670 2108.080 16.990 ;
        RECT 2107.880 2.400 2108.020 16.670 ;
        RECT 2107.670 -4.800 2108.230 2.400 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1369.490 20.640 1369.810 20.700 ;
        RECT 2125.270 20.640 2125.590 20.700 ;
        RECT 1369.490 20.500 2125.590 20.640 ;
        RECT 1369.490 20.440 1369.810 20.500 ;
        RECT 2125.270 20.440 2125.590 20.500 ;
      LAYER via ;
        RECT 1369.520 20.440 1369.780 20.700 ;
        RECT 2125.300 20.440 2125.560 20.700 ;
      LAYER met2 ;
        RECT 1368.500 1700.340 1368.780 1704.000 ;
        RECT 1368.500 1700.000 1368.800 1700.340 ;
        RECT 1368.660 1635.810 1368.800 1700.000 ;
        RECT 1368.660 1635.670 1369.720 1635.810 ;
        RECT 1369.580 20.730 1369.720 1635.670 ;
        RECT 1369.520 20.410 1369.780 20.730 ;
        RECT 2125.300 20.410 2125.560 20.730 ;
        RECT 2125.360 14.010 2125.500 20.410 ;
        RECT 2125.360 13.870 2125.960 14.010 ;
        RECT 2125.820 2.400 2125.960 13.870 ;
        RECT 2125.610 -4.800 2126.170 2.400 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1366.270 1684.600 1366.590 1684.660 ;
        RECT 1370.410 1684.600 1370.730 1684.660 ;
        RECT 1366.270 1684.460 1370.730 1684.600 ;
        RECT 1366.270 1684.400 1366.590 1684.460 ;
        RECT 1370.410 1684.400 1370.730 1684.460 ;
        RECT 1366.270 1631.900 1366.590 1631.960 ;
        RECT 1368.570 1631.900 1368.890 1631.960 ;
        RECT 1366.270 1631.760 1368.890 1631.900 ;
        RECT 1366.270 1631.700 1366.590 1631.760 ;
        RECT 1368.570 1631.700 1368.890 1631.760 ;
        RECT 1368.570 20.300 1368.890 20.360 ;
        RECT 2143.670 20.300 2143.990 20.360 ;
        RECT 1368.570 20.160 2143.990 20.300 ;
        RECT 1368.570 20.100 1368.890 20.160 ;
        RECT 2143.670 20.100 2143.990 20.160 ;
      LAYER via ;
        RECT 1366.300 1684.400 1366.560 1684.660 ;
        RECT 1370.440 1684.400 1370.700 1684.660 ;
        RECT 1366.300 1631.700 1366.560 1631.960 ;
        RECT 1368.600 1631.700 1368.860 1631.960 ;
        RECT 1368.600 20.100 1368.860 20.360 ;
        RECT 2143.700 20.100 2143.960 20.360 ;
      LAYER met2 ;
        RECT 1370.340 1700.340 1370.620 1704.000 ;
        RECT 1370.340 1700.000 1370.640 1700.340 ;
        RECT 1370.500 1684.690 1370.640 1700.000 ;
        RECT 1366.300 1684.370 1366.560 1684.690 ;
        RECT 1370.440 1684.370 1370.700 1684.690 ;
        RECT 1366.360 1631.990 1366.500 1684.370 ;
        RECT 1366.300 1631.670 1366.560 1631.990 ;
        RECT 1368.600 1631.670 1368.860 1631.990 ;
        RECT 1368.660 20.390 1368.800 1631.670 ;
        RECT 1368.600 20.070 1368.860 20.390 ;
        RECT 2143.700 20.070 2143.960 20.390 ;
        RECT 2143.760 2.400 2143.900 20.070 ;
        RECT 2143.550 -4.800 2144.110 2.400 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1367.190 1684.940 1367.510 1685.000 ;
        RECT 1372.250 1684.940 1372.570 1685.000 ;
        RECT 1367.190 1684.800 1372.570 1684.940 ;
        RECT 1367.190 1684.740 1367.510 1684.800 ;
        RECT 1372.250 1684.740 1372.570 1684.800 ;
        RECT 1367.190 19.960 1367.510 20.020 ;
        RECT 2161.610 19.960 2161.930 20.020 ;
        RECT 1367.190 19.820 2161.930 19.960 ;
        RECT 1367.190 19.760 1367.510 19.820 ;
        RECT 2161.610 19.760 2161.930 19.820 ;
      LAYER via ;
        RECT 1367.220 1684.740 1367.480 1685.000 ;
        RECT 1372.280 1684.740 1372.540 1685.000 ;
        RECT 1367.220 19.760 1367.480 20.020 ;
        RECT 2161.640 19.760 2161.900 20.020 ;
      LAYER met2 ;
        RECT 1372.180 1700.340 1372.460 1704.000 ;
        RECT 1372.180 1700.000 1372.480 1700.340 ;
        RECT 1372.340 1685.030 1372.480 1700.000 ;
        RECT 1367.220 1684.710 1367.480 1685.030 ;
        RECT 1372.280 1684.710 1372.540 1685.030 ;
        RECT 1367.280 20.050 1367.420 1684.710 ;
        RECT 1367.220 19.730 1367.480 20.050 ;
        RECT 2161.640 19.730 2161.900 20.050 ;
        RECT 2161.700 2.400 2161.840 19.730 ;
        RECT 2161.490 -4.800 2162.050 2.400 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1374.165 1655.545 1374.335 1685.635 ;
      LAYER mcon ;
        RECT 1374.165 1685.465 1374.335 1685.635 ;
      LAYER met1 ;
        RECT 1374.090 1685.620 1374.410 1685.680 ;
        RECT 1373.895 1685.480 1374.410 1685.620 ;
        RECT 1374.090 1685.420 1374.410 1685.480 ;
        RECT 1374.105 1655.700 1374.395 1655.745 ;
        RECT 1378.690 1655.700 1379.010 1655.760 ;
        RECT 1374.105 1655.560 1379.010 1655.700 ;
        RECT 1374.105 1655.515 1374.395 1655.560 ;
        RECT 1378.690 1655.500 1379.010 1655.560 ;
        RECT 1378.690 19.620 1379.010 19.680 ;
        RECT 2179.090 19.620 2179.410 19.680 ;
        RECT 1378.690 19.480 2179.410 19.620 ;
        RECT 1378.690 19.420 1379.010 19.480 ;
        RECT 2179.090 19.420 2179.410 19.480 ;
      LAYER via ;
        RECT 1374.120 1685.420 1374.380 1685.680 ;
        RECT 1378.720 1655.500 1378.980 1655.760 ;
        RECT 1378.720 19.420 1378.980 19.680 ;
        RECT 2179.120 19.420 2179.380 19.680 ;
      LAYER met2 ;
        RECT 1374.020 1700.340 1374.300 1704.000 ;
        RECT 1374.020 1700.000 1374.320 1700.340 ;
        RECT 1374.180 1685.710 1374.320 1700.000 ;
        RECT 1374.120 1685.390 1374.380 1685.710 ;
        RECT 1378.720 1655.470 1378.980 1655.790 ;
        RECT 1378.780 19.710 1378.920 1655.470 ;
        RECT 1378.720 19.390 1378.980 19.710 ;
        RECT 2179.120 19.390 2179.380 19.710 ;
        RECT 2179.180 2.400 2179.320 19.390 ;
        RECT 2178.970 -4.800 2179.530 2.400 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 2166.745 19.125 2166.915 19.975 ;
      LAYER mcon ;
        RECT 2166.745 19.805 2166.915 19.975 ;
      LAYER met1 ;
        RECT 2166.685 19.960 2166.975 20.005 ;
        RECT 2197.030 19.960 2197.350 20.020 ;
        RECT 2166.685 19.820 2197.350 19.960 ;
        RECT 2166.685 19.775 2166.975 19.820 ;
        RECT 2197.030 19.760 2197.350 19.820 ;
        RECT 1375.470 19.280 1375.790 19.340 ;
        RECT 2166.685 19.280 2166.975 19.325 ;
        RECT 1375.470 19.140 2166.975 19.280 ;
        RECT 1375.470 19.080 1375.790 19.140 ;
        RECT 2166.685 19.095 2166.975 19.140 ;
      LAYER via ;
        RECT 2197.060 19.760 2197.320 20.020 ;
        RECT 1375.500 19.080 1375.760 19.340 ;
      LAYER met2 ;
        RECT 1375.400 1700.340 1375.680 1704.000 ;
        RECT 1375.400 1700.000 1375.700 1700.340 ;
        RECT 1375.560 19.370 1375.700 1700.000 ;
        RECT 2197.060 19.730 2197.320 20.050 ;
        RECT 1375.500 19.050 1375.760 19.370 ;
        RECT 2197.120 2.400 2197.260 19.730 ;
        RECT 2196.910 -4.800 2197.470 2.400 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1374.550 1684.260 1374.870 1684.320 ;
        RECT 1377.310 1684.260 1377.630 1684.320 ;
        RECT 1374.550 1684.120 1377.630 1684.260 ;
        RECT 1374.550 1684.060 1374.870 1684.120 ;
        RECT 1377.310 1684.060 1377.630 1684.120 ;
        RECT 1375.010 18.940 1375.330 19.000 ;
        RECT 2214.970 18.940 2215.290 19.000 ;
        RECT 1375.010 18.800 2215.290 18.940 ;
        RECT 1375.010 18.740 1375.330 18.800 ;
        RECT 2214.970 18.740 2215.290 18.800 ;
      LAYER via ;
        RECT 1374.580 1684.060 1374.840 1684.320 ;
        RECT 1377.340 1684.060 1377.600 1684.320 ;
        RECT 1375.040 18.740 1375.300 19.000 ;
        RECT 2215.000 18.740 2215.260 19.000 ;
      LAYER met2 ;
        RECT 1377.240 1700.340 1377.520 1704.000 ;
        RECT 1377.240 1700.000 1377.540 1700.340 ;
        RECT 1377.400 1684.350 1377.540 1700.000 ;
        RECT 1374.580 1684.030 1374.840 1684.350 ;
        RECT 1377.340 1684.030 1377.600 1684.350 ;
        RECT 1374.640 1677.970 1374.780 1684.030 ;
        RECT 1374.640 1677.830 1375.240 1677.970 ;
        RECT 1375.100 19.030 1375.240 1677.830 ;
        RECT 1375.040 18.710 1375.300 19.030 ;
        RECT 2215.000 18.710 2215.260 19.030 ;
        RECT 2215.060 2.400 2215.200 18.710 ;
        RECT 2214.850 -4.800 2215.410 2.400 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1376.465 1242.105 1376.635 1249.075 ;
        RECT 1376.465 1027.905 1376.635 1048.815 ;
        RECT 1376.465 952.425 1376.635 953.275 ;
        RECT 1376.005 855.525 1376.175 903.975 ;
        RECT 1376.005 807.245 1376.175 855.015 ;
        RECT 1376.925 620.925 1377.095 669.375 ;
        RECT 1376.465 421.005 1376.635 469.115 ;
        RECT 1376.465 255.085 1376.635 282.795 ;
        RECT 1374.625 83.045 1374.795 131.155 ;
        RECT 1376.925 18.445 1377.095 41.395 ;
      LAYER mcon ;
        RECT 1376.465 1248.905 1376.635 1249.075 ;
        RECT 1376.465 1048.645 1376.635 1048.815 ;
        RECT 1376.465 953.105 1376.635 953.275 ;
        RECT 1376.005 903.805 1376.175 903.975 ;
        RECT 1376.005 854.845 1376.175 855.015 ;
        RECT 1376.925 669.205 1377.095 669.375 ;
        RECT 1376.465 468.945 1376.635 469.115 ;
        RECT 1376.465 282.625 1376.635 282.795 ;
        RECT 1374.625 130.985 1374.795 131.155 ;
        RECT 1376.925 41.225 1377.095 41.395 ;
      LAYER met1 ;
        RECT 1375.930 1525.140 1376.250 1525.200 ;
        RECT 1376.390 1525.140 1376.710 1525.200 ;
        RECT 1375.930 1525.000 1376.710 1525.140 ;
        RECT 1375.930 1524.940 1376.250 1525.000 ;
        RECT 1376.390 1524.940 1376.710 1525.000 ;
        RECT 1376.390 1511.340 1376.710 1511.600 ;
        RECT 1376.480 1510.520 1376.620 1511.340 ;
        RECT 1376.850 1510.520 1377.170 1510.580 ;
        RECT 1376.480 1510.380 1377.170 1510.520 ;
        RECT 1376.850 1510.320 1377.170 1510.380 ;
        RECT 1376.850 1463.260 1377.170 1463.320 ;
        RECT 1376.480 1463.120 1377.170 1463.260 ;
        RECT 1376.480 1462.640 1376.620 1463.120 ;
        RECT 1376.850 1463.060 1377.170 1463.120 ;
        RECT 1376.390 1462.380 1376.710 1462.640 ;
        RECT 1376.850 1414.640 1377.170 1414.700 ;
        RECT 1376.480 1414.500 1377.170 1414.640 ;
        RECT 1376.480 1414.360 1376.620 1414.500 ;
        RECT 1376.850 1414.440 1377.170 1414.500 ;
        RECT 1376.390 1414.100 1376.710 1414.360 ;
        RECT 1376.850 1304.820 1377.170 1304.880 ;
        RECT 1376.480 1304.680 1377.170 1304.820 ;
        RECT 1376.480 1303.860 1376.620 1304.680 ;
        RECT 1376.850 1304.620 1377.170 1304.680 ;
        RECT 1376.390 1303.600 1376.710 1303.860 ;
        RECT 1376.390 1249.060 1376.710 1249.120 ;
        RECT 1376.195 1248.920 1376.710 1249.060 ;
        RECT 1376.390 1248.860 1376.710 1248.920 ;
        RECT 1376.390 1242.260 1376.710 1242.320 ;
        RECT 1376.195 1242.120 1376.710 1242.260 ;
        RECT 1376.390 1242.060 1376.710 1242.120 ;
        RECT 1376.390 1200.780 1376.710 1200.840 ;
        RECT 1376.850 1200.780 1377.170 1200.840 ;
        RECT 1376.390 1200.640 1377.170 1200.780 ;
        RECT 1376.390 1200.580 1376.710 1200.640 ;
        RECT 1376.850 1200.580 1377.170 1200.640 ;
        RECT 1376.850 1193.640 1377.170 1193.700 ;
        RECT 1377.770 1193.640 1378.090 1193.700 ;
        RECT 1376.850 1193.500 1378.090 1193.640 ;
        RECT 1376.850 1193.440 1377.170 1193.500 ;
        RECT 1377.770 1193.440 1378.090 1193.500 ;
        RECT 1376.390 1048.800 1376.710 1048.860 ;
        RECT 1376.195 1048.660 1376.710 1048.800 ;
        RECT 1376.390 1048.600 1376.710 1048.660 ;
        RECT 1376.390 1028.060 1376.710 1028.120 ;
        RECT 1376.195 1027.920 1376.710 1028.060 ;
        RECT 1376.390 1027.860 1376.710 1027.920 ;
        RECT 1376.405 953.260 1376.695 953.305 ;
        RECT 1376.850 953.260 1377.170 953.320 ;
        RECT 1376.405 953.120 1377.170 953.260 ;
        RECT 1376.405 953.075 1376.695 953.120 ;
        RECT 1376.850 953.060 1377.170 953.120 ;
        RECT 1376.390 952.580 1376.710 952.640 ;
        RECT 1376.195 952.440 1376.710 952.580 ;
        RECT 1376.390 952.380 1376.710 952.440 ;
        RECT 1376.390 931.640 1376.710 931.900 ;
        RECT 1376.480 931.160 1376.620 931.640 ;
        RECT 1376.850 931.160 1377.170 931.220 ;
        RECT 1376.480 931.020 1377.170 931.160 ;
        RECT 1376.850 930.960 1377.170 931.020 ;
        RECT 1375.945 903.960 1376.235 904.005 ;
        RECT 1376.850 903.960 1377.170 904.020 ;
        RECT 1375.945 903.820 1377.170 903.960 ;
        RECT 1375.945 903.775 1376.235 903.820 ;
        RECT 1376.850 903.760 1377.170 903.820 ;
        RECT 1375.930 855.680 1376.250 855.740 ;
        RECT 1375.735 855.540 1376.250 855.680 ;
        RECT 1375.930 855.480 1376.250 855.540 ;
        RECT 1375.930 855.000 1376.250 855.060 ;
        RECT 1375.735 854.860 1376.250 855.000 ;
        RECT 1375.930 854.800 1376.250 854.860 ;
        RECT 1375.945 807.400 1376.235 807.445 ;
        RECT 1376.850 807.400 1377.170 807.460 ;
        RECT 1375.945 807.260 1377.170 807.400 ;
        RECT 1375.945 807.215 1376.235 807.260 ;
        RECT 1376.850 807.200 1377.170 807.260 ;
        RECT 1376.850 710.840 1377.170 710.900 ;
        RECT 1377.310 710.840 1377.630 710.900 ;
        RECT 1376.850 710.700 1377.630 710.840 ;
        RECT 1376.850 710.640 1377.170 710.700 ;
        RECT 1377.310 710.640 1377.630 710.700 ;
        RECT 1377.310 676.500 1377.630 676.560 ;
        RECT 1376.940 676.360 1377.630 676.500 ;
        RECT 1376.940 676.220 1377.080 676.360 ;
        RECT 1377.310 676.300 1377.630 676.360 ;
        RECT 1376.850 675.960 1377.170 676.220 ;
        RECT 1376.850 669.360 1377.170 669.420 ;
        RECT 1376.655 669.220 1377.170 669.360 ;
        RECT 1376.850 669.160 1377.170 669.220 ;
        RECT 1376.850 621.080 1377.170 621.140 ;
        RECT 1376.655 620.940 1377.170 621.080 ;
        RECT 1376.850 620.880 1377.170 620.940 ;
        RECT 1376.390 469.100 1376.710 469.160 ;
        RECT 1376.195 468.960 1376.710 469.100 ;
        RECT 1376.390 468.900 1376.710 468.960 ;
        RECT 1376.390 421.160 1376.710 421.220 ;
        RECT 1376.195 421.020 1376.710 421.160 ;
        RECT 1376.390 420.960 1376.710 421.020 ;
        RECT 1376.390 282.780 1376.710 282.840 ;
        RECT 1376.195 282.640 1376.710 282.780 ;
        RECT 1376.390 282.580 1376.710 282.640 ;
        RECT 1376.390 255.240 1376.710 255.300 ;
        RECT 1376.195 255.100 1376.710 255.240 ;
        RECT 1376.390 255.040 1376.710 255.100 ;
        RECT 1374.550 137.940 1374.870 138.000 ;
        RECT 1376.850 137.940 1377.170 138.000 ;
        RECT 1374.550 137.800 1377.170 137.940 ;
        RECT 1374.550 137.740 1374.870 137.800 ;
        RECT 1376.850 137.740 1377.170 137.800 ;
        RECT 1374.550 131.140 1374.870 131.200 ;
        RECT 1374.355 131.000 1374.870 131.140 ;
        RECT 1374.550 130.940 1374.870 131.000 ;
        RECT 1374.550 83.200 1374.870 83.260 ;
        RECT 1374.355 83.060 1374.870 83.200 ;
        RECT 1374.550 83.000 1374.870 83.060 ;
        RECT 1374.550 47.840 1374.870 47.900 ;
        RECT 1376.850 47.840 1377.170 47.900 ;
        RECT 1374.550 47.700 1377.170 47.840 ;
        RECT 1374.550 47.640 1374.870 47.700 ;
        RECT 1376.850 47.640 1377.170 47.700 ;
        RECT 1376.850 41.380 1377.170 41.440 ;
        RECT 1376.655 41.240 1377.170 41.380 ;
        RECT 1376.850 41.180 1377.170 41.240 ;
        RECT 1376.865 18.600 1377.155 18.645 ;
        RECT 2232.910 18.600 2233.230 18.660 ;
        RECT 1376.865 18.460 2233.230 18.600 ;
        RECT 1376.865 18.415 1377.155 18.460 ;
        RECT 2232.910 18.400 2233.230 18.460 ;
      LAYER via ;
        RECT 1375.960 1524.940 1376.220 1525.200 ;
        RECT 1376.420 1524.940 1376.680 1525.200 ;
        RECT 1376.420 1511.340 1376.680 1511.600 ;
        RECT 1376.880 1510.320 1377.140 1510.580 ;
        RECT 1376.880 1463.060 1377.140 1463.320 ;
        RECT 1376.420 1462.380 1376.680 1462.640 ;
        RECT 1376.880 1414.440 1377.140 1414.700 ;
        RECT 1376.420 1414.100 1376.680 1414.360 ;
        RECT 1376.880 1304.620 1377.140 1304.880 ;
        RECT 1376.420 1303.600 1376.680 1303.860 ;
        RECT 1376.420 1248.860 1376.680 1249.120 ;
        RECT 1376.420 1242.060 1376.680 1242.320 ;
        RECT 1376.420 1200.580 1376.680 1200.840 ;
        RECT 1376.880 1200.580 1377.140 1200.840 ;
        RECT 1376.880 1193.440 1377.140 1193.700 ;
        RECT 1377.800 1193.440 1378.060 1193.700 ;
        RECT 1376.420 1048.600 1376.680 1048.860 ;
        RECT 1376.420 1027.860 1376.680 1028.120 ;
        RECT 1376.880 953.060 1377.140 953.320 ;
        RECT 1376.420 952.380 1376.680 952.640 ;
        RECT 1376.420 931.640 1376.680 931.900 ;
        RECT 1376.880 930.960 1377.140 931.220 ;
        RECT 1376.880 903.760 1377.140 904.020 ;
        RECT 1375.960 855.480 1376.220 855.740 ;
        RECT 1375.960 854.800 1376.220 855.060 ;
        RECT 1376.880 807.200 1377.140 807.460 ;
        RECT 1376.880 710.640 1377.140 710.900 ;
        RECT 1377.340 710.640 1377.600 710.900 ;
        RECT 1377.340 676.300 1377.600 676.560 ;
        RECT 1376.880 675.960 1377.140 676.220 ;
        RECT 1376.880 669.160 1377.140 669.420 ;
        RECT 1376.880 620.880 1377.140 621.140 ;
        RECT 1376.420 468.900 1376.680 469.160 ;
        RECT 1376.420 420.960 1376.680 421.220 ;
        RECT 1376.420 282.580 1376.680 282.840 ;
        RECT 1376.420 255.040 1376.680 255.300 ;
        RECT 1374.580 137.740 1374.840 138.000 ;
        RECT 1376.880 137.740 1377.140 138.000 ;
        RECT 1374.580 130.940 1374.840 131.200 ;
        RECT 1374.580 83.000 1374.840 83.260 ;
        RECT 1374.580 47.640 1374.840 47.900 ;
        RECT 1376.880 47.640 1377.140 47.900 ;
        RECT 1376.880 41.180 1377.140 41.440 ;
        RECT 2232.940 18.400 2233.200 18.660 ;
      LAYER met2 ;
        RECT 1379.080 1700.340 1379.360 1704.000 ;
        RECT 1379.080 1700.000 1379.380 1700.340 ;
        RECT 1379.240 1629.125 1379.380 1700.000 ;
        RECT 1379.170 1628.755 1379.450 1629.125 ;
        RECT 1376.410 1573.675 1376.690 1574.045 ;
        RECT 1376.480 1573.250 1376.620 1573.675 ;
        RECT 1376.020 1573.110 1376.620 1573.250 ;
        RECT 1376.020 1525.230 1376.160 1573.110 ;
        RECT 1375.960 1524.910 1376.220 1525.230 ;
        RECT 1376.420 1524.910 1376.680 1525.230 ;
        RECT 1376.480 1511.630 1376.620 1524.910 ;
        RECT 1376.420 1511.310 1376.680 1511.630 ;
        RECT 1376.880 1510.290 1377.140 1510.610 ;
        RECT 1376.940 1463.350 1377.080 1510.290 ;
        RECT 1376.880 1463.030 1377.140 1463.350 ;
        RECT 1376.420 1462.350 1376.680 1462.670 ;
        RECT 1376.480 1435.210 1376.620 1462.350 ;
        RECT 1376.480 1435.070 1377.080 1435.210 ;
        RECT 1376.940 1414.730 1377.080 1435.070 ;
        RECT 1376.880 1414.410 1377.140 1414.730 ;
        RECT 1376.420 1414.070 1376.680 1414.390 ;
        RECT 1376.480 1369.250 1376.620 1414.070 ;
        RECT 1376.480 1369.110 1377.080 1369.250 ;
        RECT 1376.940 1304.910 1377.080 1369.110 ;
        RECT 1376.880 1304.590 1377.140 1304.910 ;
        RECT 1376.420 1303.570 1376.680 1303.890 ;
        RECT 1376.480 1249.150 1376.620 1303.570 ;
        RECT 1376.420 1248.830 1376.680 1249.150 ;
        RECT 1376.420 1242.030 1376.680 1242.350 ;
        RECT 1376.480 1200.870 1376.620 1242.030 ;
        RECT 1376.420 1200.550 1376.680 1200.870 ;
        RECT 1376.880 1200.550 1377.140 1200.870 ;
        RECT 1376.940 1193.730 1377.080 1200.550 ;
        RECT 1376.880 1193.410 1377.140 1193.730 ;
        RECT 1377.800 1193.410 1378.060 1193.730 ;
        RECT 1377.860 1145.645 1378.000 1193.410 ;
        RECT 1376.870 1145.275 1377.150 1145.645 ;
        RECT 1377.790 1145.275 1378.070 1145.645 ;
        RECT 1376.940 1128.530 1377.080 1145.275 ;
        RECT 1376.480 1128.390 1377.080 1128.530 ;
        RECT 1376.480 1048.890 1376.620 1128.390 ;
        RECT 1376.420 1048.570 1376.680 1048.890 ;
        RECT 1376.420 1027.830 1376.680 1028.150 ;
        RECT 1376.480 1000.690 1376.620 1027.830 ;
        RECT 1376.480 1000.550 1377.080 1000.690 ;
        RECT 1376.940 953.350 1377.080 1000.550 ;
        RECT 1376.880 953.030 1377.140 953.350 ;
        RECT 1376.420 952.350 1376.680 952.670 ;
        RECT 1376.480 931.930 1376.620 952.350 ;
        RECT 1376.420 931.610 1376.680 931.930 ;
        RECT 1376.880 930.930 1377.140 931.250 ;
        RECT 1376.940 904.050 1377.080 930.930 ;
        RECT 1376.880 903.730 1377.140 904.050 ;
        RECT 1375.960 855.450 1376.220 855.770 ;
        RECT 1376.020 855.090 1376.160 855.450 ;
        RECT 1375.960 854.770 1376.220 855.090 ;
        RECT 1376.880 807.170 1377.140 807.490 ;
        RECT 1376.940 710.930 1377.080 807.170 ;
        RECT 1376.880 710.610 1377.140 710.930 ;
        RECT 1377.340 710.610 1377.600 710.930 ;
        RECT 1377.400 676.590 1377.540 710.610 ;
        RECT 1377.340 676.270 1377.600 676.590 ;
        RECT 1376.880 675.930 1377.140 676.250 ;
        RECT 1376.940 669.450 1377.080 675.930 ;
        RECT 1376.880 669.130 1377.140 669.450 ;
        RECT 1376.880 620.850 1377.140 621.170 ;
        RECT 1376.940 596.770 1377.080 620.850 ;
        RECT 1376.480 596.630 1377.080 596.770 ;
        RECT 1376.480 469.190 1376.620 596.630 ;
        RECT 1376.420 468.870 1376.680 469.190 ;
        RECT 1376.420 420.930 1376.680 421.250 ;
        RECT 1376.480 282.870 1376.620 420.930 ;
        RECT 1376.420 282.550 1376.680 282.870 ;
        RECT 1376.420 255.010 1376.680 255.330 ;
        RECT 1376.480 186.050 1376.620 255.010 ;
        RECT 1376.480 185.910 1377.080 186.050 ;
        RECT 1376.940 138.030 1377.080 185.910 ;
        RECT 1374.580 137.710 1374.840 138.030 ;
        RECT 1376.880 137.710 1377.140 138.030 ;
        RECT 1374.640 131.230 1374.780 137.710 ;
        RECT 1374.580 130.910 1374.840 131.230 ;
        RECT 1374.580 82.970 1374.840 83.290 ;
        RECT 1374.640 47.930 1374.780 82.970 ;
        RECT 1374.580 47.610 1374.840 47.930 ;
        RECT 1376.880 47.610 1377.140 47.930 ;
        RECT 1376.940 41.470 1377.080 47.610 ;
        RECT 1376.880 41.150 1377.140 41.470 ;
        RECT 2232.940 18.370 2233.200 18.690 ;
        RECT 2233.000 2.400 2233.140 18.370 ;
        RECT 2232.790 -4.800 2233.350 2.400 ;
      LAYER via2 ;
        RECT 1379.170 1628.800 1379.450 1629.080 ;
        RECT 1376.410 1573.720 1376.690 1574.000 ;
        RECT 1376.870 1145.320 1377.150 1145.600 ;
        RECT 1377.790 1145.320 1378.070 1145.600 ;
      LAYER met3 ;
        RECT 1379.145 1629.090 1379.475 1629.105 ;
        RECT 1376.630 1628.790 1379.475 1629.090 ;
        RECT 1376.630 1628.420 1376.930 1628.790 ;
        RECT 1379.145 1628.775 1379.475 1628.790 ;
        RECT 1376.590 1628.100 1376.970 1628.420 ;
        RECT 1376.590 1574.690 1376.970 1574.700 ;
        RECT 1376.400 1574.380 1376.970 1574.690 ;
        RECT 1376.400 1574.025 1376.700 1574.380 ;
        RECT 1376.385 1573.695 1376.715 1574.025 ;
        RECT 1376.845 1145.610 1377.175 1145.625 ;
        RECT 1377.765 1145.610 1378.095 1145.625 ;
        RECT 1376.845 1145.310 1378.095 1145.610 ;
        RECT 1376.845 1145.295 1377.175 1145.310 ;
        RECT 1377.765 1145.295 1378.095 1145.310 ;
      LAYER via3 ;
        RECT 1376.620 1628.100 1376.940 1628.420 ;
        RECT 1376.620 1574.380 1376.940 1574.700 ;
      LAYER met4 ;
        RECT 1376.615 1628.095 1376.945 1628.425 ;
        RECT 1376.630 1574.705 1376.930 1628.095 ;
        RECT 1376.615 1574.375 1376.945 1574.705 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 793.110 1570.020 793.430 1570.080 ;
        RECT 1230.570 1570.020 1230.890 1570.080 ;
        RECT 793.110 1569.880 1230.890 1570.020 ;
        RECT 793.110 1569.820 793.430 1569.880 ;
        RECT 1230.570 1569.820 1230.890 1569.880 ;
      LAYER via ;
        RECT 793.140 1569.820 793.400 1570.080 ;
        RECT 1230.600 1569.820 1230.860 1570.080 ;
      LAYER met2 ;
        RECT 1230.500 1700.340 1230.780 1704.000 ;
        RECT 1230.500 1700.000 1230.800 1700.340 ;
        RECT 1230.660 1570.110 1230.800 1700.000 ;
        RECT 793.140 1569.790 793.400 1570.110 ;
        RECT 1230.600 1569.790 1230.860 1570.110 ;
        RECT 793.200 18.090 793.340 1569.790 ;
        RECT 787.680 17.950 793.340 18.090 ;
        RECT 787.680 2.400 787.820 17.950 ;
        RECT 787.470 -4.800 788.030 2.400 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1380.990 1672.700 1381.310 1672.760 ;
        RECT 1385.590 1672.700 1385.910 1672.760 ;
        RECT 1380.990 1672.560 1385.910 1672.700 ;
        RECT 1380.990 1672.500 1381.310 1672.560 ;
        RECT 1385.590 1672.500 1385.910 1672.560 ;
        RECT 1385.590 18.260 1385.910 18.320 ;
        RECT 2250.850 18.260 2251.170 18.320 ;
        RECT 1385.590 18.120 2251.170 18.260 ;
        RECT 1385.590 18.060 1385.910 18.120 ;
        RECT 2250.850 18.060 2251.170 18.120 ;
      LAYER via ;
        RECT 1381.020 1672.500 1381.280 1672.760 ;
        RECT 1385.620 1672.500 1385.880 1672.760 ;
        RECT 1385.620 18.060 1385.880 18.320 ;
        RECT 2250.880 18.060 2251.140 18.320 ;
      LAYER met2 ;
        RECT 1380.920 1700.340 1381.200 1704.000 ;
        RECT 1380.920 1700.000 1381.220 1700.340 ;
        RECT 1381.080 1672.790 1381.220 1700.000 ;
        RECT 1381.020 1672.470 1381.280 1672.790 ;
        RECT 1385.620 1672.470 1385.880 1672.790 ;
        RECT 1385.680 18.350 1385.820 1672.470 ;
        RECT 1385.620 18.030 1385.880 18.350 ;
        RECT 2250.880 18.030 2251.140 18.350 ;
        RECT 2250.940 2.400 2251.080 18.030 ;
        RECT 2250.730 -4.800 2251.290 2.400 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1382.445 676.345 1382.615 724.455 ;
        RECT 1382.445 537.965 1382.615 596.955 ;
        RECT 1382.445 48.365 1382.615 96.475 ;
      LAYER mcon ;
        RECT 1382.445 724.285 1382.615 724.455 ;
        RECT 1382.445 596.785 1382.615 596.955 ;
        RECT 1382.445 96.305 1382.615 96.475 ;
      LAYER met1 ;
        RECT 1382.370 724.440 1382.690 724.500 ;
        RECT 1382.175 724.300 1382.690 724.440 ;
        RECT 1382.370 724.240 1382.690 724.300 ;
        RECT 1382.370 676.500 1382.690 676.560 ;
        RECT 1382.370 676.360 1382.885 676.500 ;
        RECT 1382.370 676.300 1382.690 676.360 ;
        RECT 1382.385 596.940 1382.675 596.985 ;
        RECT 1382.830 596.940 1383.150 597.000 ;
        RECT 1382.385 596.800 1383.150 596.940 ;
        RECT 1382.385 596.755 1382.675 596.800 ;
        RECT 1382.830 596.740 1383.150 596.800 ;
        RECT 1382.370 538.120 1382.690 538.180 ;
        RECT 1382.175 537.980 1382.690 538.120 ;
        RECT 1382.370 537.920 1382.690 537.980 ;
        RECT 1382.370 96.460 1382.690 96.520 ;
        RECT 1382.175 96.320 1382.690 96.460 ;
        RECT 1382.370 96.260 1382.690 96.320 ;
        RECT 1382.370 48.520 1382.690 48.580 ;
        RECT 1382.175 48.380 1382.690 48.520 ;
        RECT 1382.370 48.320 1382.690 48.380 ;
        RECT 1382.830 17.920 1383.150 17.980 ;
        RECT 2268.330 17.920 2268.650 17.980 ;
        RECT 1382.830 17.780 2268.650 17.920 ;
        RECT 1382.830 17.720 1383.150 17.780 ;
        RECT 2268.330 17.720 2268.650 17.780 ;
      LAYER via ;
        RECT 1382.400 724.240 1382.660 724.500 ;
        RECT 1382.400 676.300 1382.660 676.560 ;
        RECT 1382.860 596.740 1383.120 597.000 ;
        RECT 1382.400 537.920 1382.660 538.180 ;
        RECT 1382.400 96.260 1382.660 96.520 ;
        RECT 1382.400 48.320 1382.660 48.580 ;
        RECT 1382.860 17.720 1383.120 17.980 ;
        RECT 2268.360 17.720 2268.620 17.980 ;
      LAYER met2 ;
        RECT 1382.760 1700.340 1383.040 1704.000 ;
        RECT 1382.760 1700.000 1383.060 1700.340 ;
        RECT 1382.920 1650.260 1383.060 1700.000 ;
        RECT 1382.460 1650.120 1383.060 1650.260 ;
        RECT 1382.460 724.530 1382.600 1650.120 ;
        RECT 1382.400 724.210 1382.660 724.530 ;
        RECT 1382.400 676.270 1382.660 676.590 ;
        RECT 1382.460 628.050 1382.600 676.270 ;
        RECT 1382.460 627.910 1383.060 628.050 ;
        RECT 1382.920 597.030 1383.060 627.910 ;
        RECT 1382.860 596.710 1383.120 597.030 ;
        RECT 1382.400 537.890 1382.660 538.210 ;
        RECT 1382.460 96.550 1382.600 537.890 ;
        RECT 1382.400 96.230 1382.660 96.550 ;
        RECT 1382.400 48.290 1382.660 48.610 ;
        RECT 1382.460 39.850 1382.600 48.290 ;
        RECT 1382.460 39.710 1383.060 39.850 ;
        RECT 1382.920 18.010 1383.060 39.710 ;
        RECT 1382.860 17.690 1383.120 18.010 ;
        RECT 2268.360 17.690 2268.620 18.010 ;
        RECT 2268.420 2.400 2268.560 17.690 ;
        RECT 2268.210 -4.800 2268.770 2.400 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1381.985 1646.365 1382.155 1684.615 ;
      LAYER mcon ;
        RECT 1381.985 1684.445 1382.155 1684.615 ;
      LAYER met1 ;
        RECT 1381.925 1684.600 1382.215 1684.645 ;
        RECT 1384.670 1684.600 1384.990 1684.660 ;
        RECT 1381.925 1684.460 1384.990 1684.600 ;
        RECT 1381.925 1684.415 1382.215 1684.460 ;
        RECT 1384.670 1684.400 1384.990 1684.460 ;
        RECT 1381.910 1646.520 1382.230 1646.580 ;
        RECT 1381.715 1646.380 1382.230 1646.520 ;
        RECT 1381.910 1646.320 1382.230 1646.380 ;
        RECT 1381.910 17.580 1382.230 17.640 ;
        RECT 2286.270 17.580 2286.590 17.640 ;
        RECT 1381.910 17.440 2286.590 17.580 ;
        RECT 1381.910 17.380 1382.230 17.440 ;
        RECT 2286.270 17.380 2286.590 17.440 ;
      LAYER via ;
        RECT 1384.700 1684.400 1384.960 1684.660 ;
        RECT 1381.940 1646.320 1382.200 1646.580 ;
        RECT 1381.940 17.380 1382.200 17.640 ;
        RECT 2286.300 17.380 2286.560 17.640 ;
      LAYER met2 ;
        RECT 1384.600 1700.340 1384.880 1704.000 ;
        RECT 1384.600 1700.000 1384.900 1700.340 ;
        RECT 1384.760 1684.690 1384.900 1700.000 ;
        RECT 1384.700 1684.370 1384.960 1684.690 ;
        RECT 1381.940 1646.290 1382.200 1646.610 ;
        RECT 1382.000 17.670 1382.140 1646.290 ;
        RECT 1381.940 17.350 1382.200 17.670 ;
        RECT 2286.300 17.350 2286.560 17.670 ;
        RECT 2286.360 2.400 2286.500 17.350 ;
        RECT 2286.150 -4.800 2286.710 2.400 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1386.510 1684.260 1386.830 1684.320 ;
        RECT 1383.840 1684.120 1386.830 1684.260 ;
        RECT 1380.530 1683.580 1380.850 1683.640 ;
        RECT 1383.840 1683.580 1383.980 1684.120 ;
        RECT 1386.510 1684.060 1386.830 1684.120 ;
        RECT 1380.530 1683.440 1383.980 1683.580 ;
        RECT 1380.530 1683.380 1380.850 1683.440 ;
        RECT 1380.530 17.240 1380.850 17.300 ;
        RECT 2304.210 17.240 2304.530 17.300 ;
        RECT 1380.530 17.100 2304.530 17.240 ;
        RECT 1380.530 17.040 1380.850 17.100 ;
        RECT 2304.210 17.040 2304.530 17.100 ;
      LAYER via ;
        RECT 1380.560 1683.380 1380.820 1683.640 ;
        RECT 1386.540 1684.060 1386.800 1684.320 ;
        RECT 1380.560 17.040 1380.820 17.300 ;
        RECT 2304.240 17.040 2304.500 17.300 ;
      LAYER met2 ;
        RECT 1386.440 1700.340 1386.720 1704.000 ;
        RECT 1386.440 1700.000 1386.740 1700.340 ;
        RECT 1386.600 1684.350 1386.740 1700.000 ;
        RECT 1386.540 1684.030 1386.800 1684.350 ;
        RECT 1380.560 1683.350 1380.820 1683.670 ;
        RECT 1380.620 17.330 1380.760 1683.350 ;
        RECT 1380.560 17.010 1380.820 17.330 ;
        RECT 2304.240 17.010 2304.500 17.330 ;
        RECT 2304.300 2.400 2304.440 17.010 ;
        RECT 2304.090 -4.800 2304.650 2.400 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1388.350 1677.600 1388.670 1677.860 ;
        RECT 1388.440 1676.840 1388.580 1677.600 ;
        RECT 1388.350 1676.580 1388.670 1676.840 ;
      LAYER via ;
        RECT 1388.380 1677.600 1388.640 1677.860 ;
        RECT 1388.380 1676.580 1388.640 1676.840 ;
      LAYER met2 ;
        RECT 1388.280 1700.340 1388.560 1704.000 ;
        RECT 1388.280 1700.000 1388.580 1700.340 ;
        RECT 1388.440 1677.890 1388.580 1700.000 ;
        RECT 1388.380 1677.570 1388.640 1677.890 ;
        RECT 1388.380 1676.550 1388.640 1676.870 ;
        RECT 1388.440 41.210 1388.580 1676.550 ;
        RECT 1387.980 41.070 1388.580 41.210 ;
        RECT 1387.980 20.245 1388.120 41.070 ;
        RECT 1387.910 19.875 1388.190 20.245 ;
        RECT 2322.170 19.875 2322.450 20.245 ;
        RECT 2322.240 2.400 2322.380 19.875 ;
        RECT 2322.030 -4.800 2322.590 2.400 ;
      LAYER via2 ;
        RECT 1387.910 19.920 1388.190 20.200 ;
        RECT 2322.170 19.920 2322.450 20.200 ;
      LAYER met3 ;
        RECT 1387.885 20.210 1388.215 20.225 ;
        RECT 2322.145 20.210 2322.475 20.225 ;
        RECT 1387.885 19.910 2322.475 20.210 ;
        RECT 1387.885 19.895 1388.215 19.910 ;
        RECT 2322.145 19.895 2322.475 19.910 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1389.345 1386.945 1389.515 1447.975 ;
        RECT 1389.805 1104.065 1389.975 1125.995 ;
        RECT 1389.345 1048.985 1389.515 1097.095 ;
      LAYER mcon ;
        RECT 1389.345 1447.805 1389.515 1447.975 ;
        RECT 1389.805 1125.825 1389.975 1125.995 ;
        RECT 1389.345 1096.925 1389.515 1097.095 ;
      LAYER met1 ;
        RECT 1390.190 1665.900 1390.510 1665.960 ;
        RECT 1389.820 1665.760 1390.510 1665.900 ;
        RECT 1389.820 1665.620 1389.960 1665.760 ;
        RECT 1390.190 1665.700 1390.510 1665.760 ;
        RECT 1389.730 1665.360 1390.050 1665.620 ;
        RECT 1389.270 1587.360 1389.590 1587.420 ;
        RECT 1389.730 1587.360 1390.050 1587.420 ;
        RECT 1389.270 1587.220 1390.050 1587.360 ;
        RECT 1389.270 1587.160 1389.590 1587.220 ;
        RECT 1389.730 1587.160 1390.050 1587.220 ;
        RECT 1389.270 1524.800 1389.590 1524.860 ;
        RECT 1391.110 1524.800 1391.430 1524.860 ;
        RECT 1389.270 1524.660 1391.430 1524.800 ;
        RECT 1389.270 1524.600 1389.590 1524.660 ;
        RECT 1391.110 1524.600 1391.430 1524.660 ;
        RECT 1389.285 1447.960 1389.575 1448.005 ;
        RECT 1389.730 1447.960 1390.050 1448.020 ;
        RECT 1389.285 1447.820 1390.050 1447.960 ;
        RECT 1389.285 1447.775 1389.575 1447.820 ;
        RECT 1389.730 1447.760 1390.050 1447.820 ;
        RECT 1389.270 1387.100 1389.590 1387.160 ;
        RECT 1389.075 1386.960 1389.590 1387.100 ;
        RECT 1389.270 1386.900 1389.590 1386.960 ;
        RECT 1389.270 1272.860 1389.590 1272.920 ;
        RECT 1390.190 1272.860 1390.510 1272.920 ;
        RECT 1389.270 1272.720 1390.510 1272.860 ;
        RECT 1389.270 1272.660 1389.590 1272.720 ;
        RECT 1390.190 1272.660 1390.510 1272.720 ;
        RECT 1389.270 1241.920 1389.590 1241.980 ;
        RECT 1390.190 1241.920 1390.510 1241.980 ;
        RECT 1389.270 1241.780 1390.510 1241.920 ;
        RECT 1389.270 1241.720 1389.590 1241.780 ;
        RECT 1390.190 1241.720 1390.510 1241.780 ;
        RECT 1388.810 1193.640 1389.130 1193.700 ;
        RECT 1390.190 1193.640 1390.510 1193.700 ;
        RECT 1388.810 1193.500 1390.510 1193.640 ;
        RECT 1388.810 1193.440 1389.130 1193.500 ;
        RECT 1390.190 1193.440 1390.510 1193.500 ;
        RECT 1389.730 1125.980 1390.050 1126.040 ;
        RECT 1389.535 1125.840 1390.050 1125.980 ;
        RECT 1389.730 1125.780 1390.050 1125.840 ;
        RECT 1389.730 1104.220 1390.050 1104.280 ;
        RECT 1389.535 1104.080 1390.050 1104.220 ;
        RECT 1389.730 1104.020 1390.050 1104.080 ;
        RECT 1389.285 1097.080 1389.575 1097.125 ;
        RECT 1389.730 1097.080 1390.050 1097.140 ;
        RECT 1389.285 1096.940 1390.050 1097.080 ;
        RECT 1389.285 1096.895 1389.575 1096.940 ;
        RECT 1389.730 1096.880 1390.050 1096.940 ;
        RECT 1389.270 1049.140 1389.590 1049.200 ;
        RECT 1389.075 1049.000 1389.590 1049.140 ;
        RECT 1389.270 1048.940 1389.590 1049.000 ;
        RECT 1389.730 959.180 1390.050 959.440 ;
        RECT 1389.820 958.700 1389.960 959.180 ;
        RECT 1390.190 958.700 1390.510 958.760 ;
        RECT 1389.820 958.560 1390.510 958.700 ;
        RECT 1390.190 958.500 1390.510 958.560 ;
        RECT 1388.810 952.240 1389.130 952.300 ;
        RECT 1390.190 952.240 1390.510 952.300 ;
        RECT 1388.810 952.100 1390.510 952.240 ;
        RECT 1388.810 952.040 1389.130 952.100 ;
        RECT 1390.190 952.040 1390.510 952.100 ;
        RECT 1389.270 855.680 1389.590 855.740 ;
        RECT 1389.730 855.680 1390.050 855.740 ;
        RECT 1389.270 855.540 1390.050 855.680 ;
        RECT 1389.270 855.480 1389.590 855.540 ;
        RECT 1389.730 855.480 1390.050 855.540 ;
        RECT 1389.270 807.400 1389.590 807.460 ;
        RECT 1390.650 807.400 1390.970 807.460 ;
        RECT 1389.270 807.260 1390.970 807.400 ;
        RECT 1389.270 807.200 1389.590 807.260 ;
        RECT 1390.650 807.200 1390.970 807.260 ;
      LAYER via ;
        RECT 1390.220 1665.700 1390.480 1665.960 ;
        RECT 1389.760 1665.360 1390.020 1665.620 ;
        RECT 1389.300 1587.160 1389.560 1587.420 ;
        RECT 1389.760 1587.160 1390.020 1587.420 ;
        RECT 1389.300 1524.600 1389.560 1524.860 ;
        RECT 1391.140 1524.600 1391.400 1524.860 ;
        RECT 1389.760 1447.760 1390.020 1448.020 ;
        RECT 1389.300 1386.900 1389.560 1387.160 ;
        RECT 1389.300 1272.660 1389.560 1272.920 ;
        RECT 1390.220 1272.660 1390.480 1272.920 ;
        RECT 1389.300 1241.720 1389.560 1241.980 ;
        RECT 1390.220 1241.720 1390.480 1241.980 ;
        RECT 1388.840 1193.440 1389.100 1193.700 ;
        RECT 1390.220 1193.440 1390.480 1193.700 ;
        RECT 1389.760 1125.780 1390.020 1126.040 ;
        RECT 1389.760 1104.020 1390.020 1104.280 ;
        RECT 1389.760 1096.880 1390.020 1097.140 ;
        RECT 1389.300 1048.940 1389.560 1049.200 ;
        RECT 1389.760 959.180 1390.020 959.440 ;
        RECT 1390.220 958.500 1390.480 958.760 ;
        RECT 1388.840 952.040 1389.100 952.300 ;
        RECT 1390.220 952.040 1390.480 952.300 ;
        RECT 1389.300 855.480 1389.560 855.740 ;
        RECT 1389.760 855.480 1390.020 855.740 ;
        RECT 1389.300 807.200 1389.560 807.460 ;
        RECT 1390.680 807.200 1390.940 807.460 ;
      LAYER met2 ;
        RECT 1390.120 1700.340 1390.400 1704.000 ;
        RECT 1390.120 1700.000 1390.420 1700.340 ;
        RECT 1390.280 1665.990 1390.420 1700.000 ;
        RECT 1390.220 1665.670 1390.480 1665.990 ;
        RECT 1389.760 1665.330 1390.020 1665.650 ;
        RECT 1389.820 1587.450 1389.960 1665.330 ;
        RECT 1389.300 1587.130 1389.560 1587.450 ;
        RECT 1389.760 1587.130 1390.020 1587.450 ;
        RECT 1389.360 1524.890 1389.500 1587.130 ;
        RECT 1389.300 1524.570 1389.560 1524.890 ;
        RECT 1391.140 1524.570 1391.400 1524.890 ;
        RECT 1391.200 1476.805 1391.340 1524.570 ;
        RECT 1389.750 1476.435 1390.030 1476.805 ;
        RECT 1391.130 1476.435 1391.410 1476.805 ;
        RECT 1389.820 1448.050 1389.960 1476.435 ;
        RECT 1389.760 1447.730 1390.020 1448.050 ;
        RECT 1389.300 1386.870 1389.560 1387.190 ;
        RECT 1389.360 1272.950 1389.500 1386.870 ;
        RECT 1389.300 1272.630 1389.560 1272.950 ;
        RECT 1390.220 1272.630 1390.480 1272.950 ;
        RECT 1390.280 1242.010 1390.420 1272.630 ;
        RECT 1389.300 1241.690 1389.560 1242.010 ;
        RECT 1390.220 1241.690 1390.480 1242.010 ;
        RECT 1389.360 1193.925 1389.500 1241.690 ;
        RECT 1388.840 1193.410 1389.100 1193.730 ;
        RECT 1389.290 1193.555 1389.570 1193.925 ;
        RECT 1390.210 1193.555 1390.490 1193.925 ;
        RECT 1390.220 1193.410 1390.480 1193.555 ;
        RECT 1388.900 1145.645 1389.040 1193.410 ;
        RECT 1388.830 1145.275 1389.110 1145.645 ;
        RECT 1389.750 1145.275 1390.030 1145.645 ;
        RECT 1389.820 1126.070 1389.960 1145.275 ;
        RECT 1389.760 1125.750 1390.020 1126.070 ;
        RECT 1389.760 1103.990 1390.020 1104.310 ;
        RECT 1389.820 1097.170 1389.960 1103.990 ;
        RECT 1389.760 1096.850 1390.020 1097.170 ;
        RECT 1389.300 1048.910 1389.560 1049.230 ;
        RECT 1389.360 1027.890 1389.500 1048.910 ;
        RECT 1389.360 1027.750 1389.960 1027.890 ;
        RECT 1389.820 959.470 1389.960 1027.750 ;
        RECT 1389.760 959.150 1390.020 959.470 ;
        RECT 1390.220 958.470 1390.480 958.790 ;
        RECT 1390.280 952.330 1390.420 958.470 ;
        RECT 1388.840 952.010 1389.100 952.330 ;
        RECT 1390.220 952.010 1390.480 952.330 ;
        RECT 1388.900 904.245 1389.040 952.010 ;
        RECT 1388.830 903.875 1389.110 904.245 ;
        RECT 1389.750 903.875 1390.030 904.245 ;
        RECT 1389.820 855.770 1389.960 903.875 ;
        RECT 1389.300 855.450 1389.560 855.770 ;
        RECT 1389.760 855.450 1390.020 855.770 ;
        RECT 1389.360 807.490 1389.500 855.450 ;
        RECT 1389.300 807.170 1389.560 807.490 ;
        RECT 1390.680 807.170 1390.940 807.490 ;
        RECT 1390.740 766.090 1390.880 807.170 ;
        RECT 1390.280 765.950 1390.880 766.090 ;
        RECT 1390.280 724.440 1390.420 765.950 ;
        RECT 1389.360 724.300 1390.420 724.440 ;
        RECT 1389.360 641.650 1389.500 724.300 ;
        RECT 1389.360 641.510 1390.420 641.650 ;
        RECT 1390.280 603.570 1390.420 641.510 ;
        RECT 1389.820 603.430 1390.420 603.570 ;
        RECT 1389.820 545.770 1389.960 603.430 ;
        RECT 1389.360 545.630 1389.960 545.770 ;
        RECT 1389.360 545.090 1389.500 545.630 ;
        RECT 1389.360 544.950 1390.420 545.090 ;
        RECT 1390.280 507.010 1390.420 544.950 ;
        RECT 1389.360 506.870 1390.420 507.010 ;
        RECT 1389.360 496.130 1389.500 506.870 ;
        RECT 1389.360 495.990 1389.960 496.130 ;
        RECT 1389.820 448.530 1389.960 495.990 ;
        RECT 1388.900 448.390 1389.960 448.530 ;
        RECT 1388.900 313.890 1389.040 448.390 ;
        RECT 1388.900 313.750 1389.960 313.890 ;
        RECT 1389.820 134.370 1389.960 313.750 ;
        RECT 1389.820 134.230 1390.420 134.370 ;
        RECT 1390.280 62.290 1390.420 134.230 ;
        RECT 1389.360 62.150 1390.420 62.290 ;
        RECT 1389.360 19.565 1389.500 62.150 ;
        RECT 1389.290 19.195 1389.570 19.565 ;
        RECT 2339.650 19.195 2339.930 19.565 ;
        RECT 2339.720 2.400 2339.860 19.195 ;
        RECT 2339.510 -4.800 2340.070 2.400 ;
      LAYER via2 ;
        RECT 1389.750 1476.480 1390.030 1476.760 ;
        RECT 1391.130 1476.480 1391.410 1476.760 ;
        RECT 1389.290 1193.600 1389.570 1193.880 ;
        RECT 1390.210 1193.600 1390.490 1193.880 ;
        RECT 1388.830 1145.320 1389.110 1145.600 ;
        RECT 1389.750 1145.320 1390.030 1145.600 ;
        RECT 1388.830 903.920 1389.110 904.200 ;
        RECT 1389.750 903.920 1390.030 904.200 ;
        RECT 1389.290 19.240 1389.570 19.520 ;
        RECT 2339.650 19.240 2339.930 19.520 ;
      LAYER met3 ;
        RECT 1389.725 1476.770 1390.055 1476.785 ;
        RECT 1391.105 1476.770 1391.435 1476.785 ;
        RECT 1389.725 1476.470 1391.435 1476.770 ;
        RECT 1389.725 1476.455 1390.055 1476.470 ;
        RECT 1391.105 1476.455 1391.435 1476.470 ;
        RECT 1389.265 1193.890 1389.595 1193.905 ;
        RECT 1390.185 1193.890 1390.515 1193.905 ;
        RECT 1389.265 1193.590 1390.515 1193.890 ;
        RECT 1389.265 1193.575 1389.595 1193.590 ;
        RECT 1390.185 1193.575 1390.515 1193.590 ;
        RECT 1388.805 1145.610 1389.135 1145.625 ;
        RECT 1389.725 1145.610 1390.055 1145.625 ;
        RECT 1388.805 1145.310 1390.055 1145.610 ;
        RECT 1388.805 1145.295 1389.135 1145.310 ;
        RECT 1389.725 1145.295 1390.055 1145.310 ;
        RECT 1388.805 904.210 1389.135 904.225 ;
        RECT 1389.725 904.210 1390.055 904.225 ;
        RECT 1388.805 903.910 1390.055 904.210 ;
        RECT 1388.805 903.895 1389.135 903.910 ;
        RECT 1389.725 903.895 1390.055 903.910 ;
        RECT 1389.265 19.530 1389.595 19.545 ;
        RECT 2339.625 19.530 2339.955 19.545 ;
        RECT 1389.265 19.230 2339.955 19.530 ;
        RECT 1389.265 19.215 1389.595 19.230 ;
        RECT 2339.625 19.215 2339.955 19.230 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1390.725 641.325 1390.895 676.175 ;
        RECT 1391.645 524.365 1391.815 572.475 ;
        RECT 1390.265 186.405 1390.435 234.515 ;
        RECT 1391.185 48.365 1391.355 137.615 ;
      LAYER mcon ;
        RECT 1390.725 676.005 1390.895 676.175 ;
        RECT 1391.645 572.305 1391.815 572.475 ;
        RECT 1390.265 234.345 1390.435 234.515 ;
        RECT 1391.185 137.445 1391.355 137.615 ;
      LAYER met1 ;
        RECT 1390.190 1665.220 1390.510 1665.280 ;
        RECT 1392.030 1665.220 1392.350 1665.280 ;
        RECT 1390.190 1665.080 1392.350 1665.220 ;
        RECT 1390.190 1665.020 1390.510 1665.080 ;
        RECT 1392.030 1665.020 1392.350 1665.080 ;
        RECT 1390.190 1539.080 1390.510 1539.140 ;
        RECT 1390.650 1539.080 1390.970 1539.140 ;
        RECT 1390.190 1538.940 1390.970 1539.080 ;
        RECT 1390.190 1538.880 1390.510 1538.940 ;
        RECT 1390.650 1538.880 1390.970 1538.940 ;
        RECT 1390.650 1483.660 1390.970 1483.720 ;
        RECT 1391.570 1483.660 1391.890 1483.720 ;
        RECT 1390.650 1483.520 1391.890 1483.660 ;
        RECT 1390.650 1483.460 1390.970 1483.520 ;
        RECT 1391.570 1483.460 1391.890 1483.520 ;
        RECT 1391.110 1207.580 1391.430 1207.640 ;
        RECT 1391.570 1207.580 1391.890 1207.640 ;
        RECT 1391.110 1207.440 1391.890 1207.580 ;
        RECT 1391.110 1207.380 1391.430 1207.440 ;
        RECT 1391.570 1207.380 1391.890 1207.440 ;
        RECT 1391.110 931.500 1391.430 931.560 ;
        RECT 1392.030 931.500 1392.350 931.560 ;
        RECT 1391.110 931.360 1392.350 931.500 ;
        RECT 1391.110 931.300 1391.430 931.360 ;
        RECT 1392.030 931.300 1392.350 931.360 ;
        RECT 1390.650 738.380 1390.970 738.440 ;
        RECT 1391.570 738.380 1391.890 738.440 ;
        RECT 1390.650 738.240 1391.890 738.380 ;
        RECT 1390.650 738.180 1390.970 738.240 ;
        RECT 1391.570 738.180 1391.890 738.240 ;
        RECT 1390.650 676.160 1390.970 676.220 ;
        RECT 1390.455 676.020 1390.970 676.160 ;
        RECT 1390.650 675.960 1390.970 676.020 ;
        RECT 1390.665 641.480 1390.955 641.525 ;
        RECT 1391.110 641.480 1391.430 641.540 ;
        RECT 1390.665 641.340 1391.430 641.480 ;
        RECT 1390.665 641.295 1390.955 641.340 ;
        RECT 1391.110 641.280 1391.430 641.340 ;
        RECT 1391.110 572.800 1391.430 572.860 ;
        RECT 1391.110 572.660 1392.260 572.800 ;
        RECT 1391.110 572.600 1391.430 572.660 ;
        RECT 1391.585 572.460 1391.875 572.505 ;
        RECT 1392.120 572.460 1392.260 572.660 ;
        RECT 1391.585 572.320 1392.260 572.460 ;
        RECT 1391.585 572.275 1391.875 572.320 ;
        RECT 1391.570 524.520 1391.890 524.580 ;
        RECT 1391.375 524.380 1391.890 524.520 ;
        RECT 1391.570 524.320 1391.890 524.380 ;
        RECT 1390.190 338.200 1390.510 338.260 ;
        RECT 1390.650 338.200 1390.970 338.260 ;
        RECT 1390.190 338.060 1390.970 338.200 ;
        RECT 1390.190 338.000 1390.510 338.060 ;
        RECT 1390.650 338.000 1390.970 338.060 ;
        RECT 1390.190 255.240 1390.510 255.300 ;
        RECT 1391.110 255.240 1391.430 255.300 ;
        RECT 1390.190 255.100 1391.430 255.240 ;
        RECT 1390.190 255.040 1390.510 255.100 ;
        RECT 1391.110 255.040 1391.430 255.100 ;
        RECT 1390.205 234.500 1390.495 234.545 ;
        RECT 1391.110 234.500 1391.430 234.560 ;
        RECT 1390.205 234.360 1391.430 234.500 ;
        RECT 1390.205 234.315 1390.495 234.360 ;
        RECT 1391.110 234.300 1391.430 234.360 ;
        RECT 1390.190 186.560 1390.510 186.620 ;
        RECT 1389.995 186.420 1390.510 186.560 ;
        RECT 1390.190 186.360 1390.510 186.420 ;
        RECT 1390.190 137.600 1390.510 137.660 ;
        RECT 1391.125 137.600 1391.415 137.645 ;
        RECT 1390.190 137.460 1391.415 137.600 ;
        RECT 1390.190 137.400 1390.510 137.460 ;
        RECT 1391.125 137.415 1391.415 137.460 ;
        RECT 1391.110 48.520 1391.430 48.580 ;
        RECT 1390.915 48.380 1391.430 48.520 ;
        RECT 1391.110 48.320 1391.430 48.380 ;
      LAYER via ;
        RECT 1390.220 1665.020 1390.480 1665.280 ;
        RECT 1392.060 1665.020 1392.320 1665.280 ;
        RECT 1390.220 1538.880 1390.480 1539.140 ;
        RECT 1390.680 1538.880 1390.940 1539.140 ;
        RECT 1390.680 1483.460 1390.940 1483.720 ;
        RECT 1391.600 1483.460 1391.860 1483.720 ;
        RECT 1391.140 1207.380 1391.400 1207.640 ;
        RECT 1391.600 1207.380 1391.860 1207.640 ;
        RECT 1391.140 931.300 1391.400 931.560 ;
        RECT 1392.060 931.300 1392.320 931.560 ;
        RECT 1390.680 738.180 1390.940 738.440 ;
        RECT 1391.600 738.180 1391.860 738.440 ;
        RECT 1390.680 675.960 1390.940 676.220 ;
        RECT 1391.140 641.280 1391.400 641.540 ;
        RECT 1391.140 572.600 1391.400 572.860 ;
        RECT 1391.600 524.320 1391.860 524.580 ;
        RECT 1390.220 338.000 1390.480 338.260 ;
        RECT 1390.680 338.000 1390.940 338.260 ;
        RECT 1390.220 255.040 1390.480 255.300 ;
        RECT 1391.140 255.040 1391.400 255.300 ;
        RECT 1391.140 234.300 1391.400 234.560 ;
        RECT 1390.220 186.360 1390.480 186.620 ;
        RECT 1390.220 137.400 1390.480 137.660 ;
        RECT 1391.140 48.320 1391.400 48.580 ;
      LAYER met2 ;
        RECT 1391.960 1700.340 1392.240 1704.000 ;
        RECT 1391.960 1700.000 1392.260 1700.340 ;
        RECT 1392.120 1665.310 1392.260 1700.000 ;
        RECT 1390.220 1664.990 1390.480 1665.310 ;
        RECT 1392.060 1664.990 1392.320 1665.310 ;
        RECT 1390.280 1618.130 1390.420 1664.990 ;
        RECT 1390.280 1617.990 1390.880 1618.130 ;
        RECT 1390.740 1539.170 1390.880 1617.990 ;
        RECT 1390.220 1538.850 1390.480 1539.170 ;
        RECT 1390.680 1538.850 1390.940 1539.170 ;
        RECT 1390.280 1531.885 1390.420 1538.850 ;
        RECT 1390.210 1531.515 1390.490 1531.885 ;
        RECT 1391.590 1531.515 1391.870 1531.885 ;
        RECT 1391.660 1483.750 1391.800 1531.515 ;
        RECT 1390.680 1483.430 1390.940 1483.750 ;
        RECT 1391.600 1483.430 1391.860 1483.750 ;
        RECT 1390.210 1386.930 1390.490 1387.045 ;
        RECT 1390.740 1386.930 1390.880 1483.430 ;
        RECT 1390.210 1386.790 1390.880 1386.930 ;
        RECT 1390.210 1386.675 1390.490 1386.790 ;
        RECT 1391.590 1385.995 1391.870 1386.365 ;
        RECT 1391.660 1207.670 1391.800 1385.995 ;
        RECT 1391.140 1207.350 1391.400 1207.670 ;
        RECT 1391.600 1207.350 1391.860 1207.670 ;
        RECT 1391.200 1028.570 1391.340 1207.350 ;
        RECT 1390.280 1028.430 1391.340 1028.570 ;
        RECT 1390.280 1014.405 1390.420 1028.430 ;
        RECT 1390.210 1014.035 1390.490 1014.405 ;
        RECT 1391.130 1014.035 1391.410 1014.405 ;
        RECT 1391.200 931.590 1391.340 1014.035 ;
        RECT 1391.140 931.270 1391.400 931.590 ;
        RECT 1392.060 931.270 1392.320 931.590 ;
        RECT 1392.120 893.930 1392.260 931.270 ;
        RECT 1391.660 893.790 1392.260 893.930 ;
        RECT 1391.660 738.470 1391.800 893.790 ;
        RECT 1390.680 738.150 1390.940 738.470 ;
        RECT 1391.600 738.150 1391.860 738.470 ;
        RECT 1390.740 714.410 1390.880 738.150 ;
        RECT 1390.280 714.270 1390.880 714.410 ;
        RECT 1390.280 689.930 1390.420 714.270 ;
        RECT 1390.280 689.790 1390.880 689.930 ;
        RECT 1390.740 676.250 1390.880 689.790 ;
        RECT 1390.680 675.930 1390.940 676.250 ;
        RECT 1391.140 641.250 1391.400 641.570 ;
        RECT 1391.200 572.890 1391.340 641.250 ;
        RECT 1391.140 572.570 1391.400 572.890 ;
        RECT 1391.600 524.290 1391.860 524.610 ;
        RECT 1391.660 483.325 1391.800 524.290 ;
        RECT 1390.670 482.955 1390.950 483.325 ;
        RECT 1391.590 482.955 1391.870 483.325 ;
        RECT 1390.740 400.930 1390.880 482.955 ;
        RECT 1390.280 400.790 1390.880 400.930 ;
        RECT 1390.280 400.250 1390.420 400.790 ;
        RECT 1390.280 400.110 1390.880 400.250 ;
        RECT 1390.740 338.290 1390.880 400.110 ;
        RECT 1390.220 337.970 1390.480 338.290 ;
        RECT 1390.680 337.970 1390.940 338.290 ;
        RECT 1390.280 255.330 1390.420 337.970 ;
        RECT 1390.220 255.010 1390.480 255.330 ;
        RECT 1391.140 255.010 1391.400 255.330 ;
        RECT 1391.200 234.590 1391.340 255.010 ;
        RECT 1391.140 234.270 1391.400 234.590 ;
        RECT 1390.220 186.330 1390.480 186.650 ;
        RECT 1390.280 137.690 1390.420 186.330 ;
        RECT 1390.220 137.370 1390.480 137.690 ;
        RECT 1391.140 48.290 1391.400 48.610 ;
        RECT 1391.200 18.885 1391.340 48.290 ;
        RECT 1391.130 18.515 1391.410 18.885 ;
        RECT 2357.590 18.515 2357.870 18.885 ;
        RECT 2357.660 2.400 2357.800 18.515 ;
        RECT 2357.450 -4.800 2358.010 2.400 ;
      LAYER via2 ;
        RECT 1390.210 1531.560 1390.490 1531.840 ;
        RECT 1391.590 1531.560 1391.870 1531.840 ;
        RECT 1390.210 1386.720 1390.490 1387.000 ;
        RECT 1391.590 1386.040 1391.870 1386.320 ;
        RECT 1390.210 1014.080 1390.490 1014.360 ;
        RECT 1391.130 1014.080 1391.410 1014.360 ;
        RECT 1390.670 483.000 1390.950 483.280 ;
        RECT 1391.590 483.000 1391.870 483.280 ;
        RECT 1391.130 18.560 1391.410 18.840 ;
        RECT 2357.590 18.560 2357.870 18.840 ;
      LAYER met3 ;
        RECT 1390.185 1531.850 1390.515 1531.865 ;
        RECT 1391.565 1531.850 1391.895 1531.865 ;
        RECT 1390.185 1531.550 1391.895 1531.850 ;
        RECT 1390.185 1531.535 1390.515 1531.550 ;
        RECT 1391.565 1531.535 1391.895 1531.550 ;
        RECT 1390.185 1387.010 1390.515 1387.025 ;
        RECT 1389.510 1386.710 1390.515 1387.010 ;
        RECT 1389.510 1386.330 1389.810 1386.710 ;
        RECT 1390.185 1386.695 1390.515 1386.710 ;
        RECT 1391.565 1386.330 1391.895 1386.345 ;
        RECT 1389.510 1386.030 1391.895 1386.330 ;
        RECT 1391.565 1386.015 1391.895 1386.030 ;
        RECT 1390.185 1014.370 1390.515 1014.385 ;
        RECT 1391.105 1014.370 1391.435 1014.385 ;
        RECT 1390.185 1014.070 1391.435 1014.370 ;
        RECT 1390.185 1014.055 1390.515 1014.070 ;
        RECT 1391.105 1014.055 1391.435 1014.070 ;
        RECT 1390.645 483.290 1390.975 483.305 ;
        RECT 1391.565 483.290 1391.895 483.305 ;
        RECT 1390.645 482.990 1391.895 483.290 ;
        RECT 1390.645 482.975 1390.975 482.990 ;
        RECT 1391.565 482.975 1391.895 482.990 ;
        RECT 1391.105 18.850 1391.435 18.865 ;
        RECT 2357.565 18.850 2357.895 18.865 ;
        RECT 1391.105 18.550 2357.895 18.850 ;
        RECT 1391.105 18.535 1391.435 18.550 ;
        RECT 2357.565 18.535 2357.895 18.550 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1395.710 1650.260 1396.030 1650.320 ;
        RECT 1399.390 1650.260 1399.710 1650.320 ;
        RECT 1395.710 1650.120 1399.710 1650.260 ;
        RECT 1395.710 1650.060 1396.030 1650.120 ;
        RECT 1399.390 1650.060 1399.710 1650.120 ;
      LAYER via ;
        RECT 1395.740 1650.060 1396.000 1650.320 ;
        RECT 1399.420 1650.060 1399.680 1650.320 ;
      LAYER met2 ;
        RECT 1393.800 1700.410 1394.080 1704.000 ;
        RECT 1393.800 1700.270 1394.560 1700.410 ;
        RECT 1393.800 1700.000 1394.080 1700.270 ;
        RECT 1394.420 1677.290 1394.560 1700.270 ;
        RECT 1394.420 1677.150 1395.940 1677.290 ;
        RECT 1395.800 1650.350 1395.940 1677.150 ;
        RECT 1395.740 1650.030 1396.000 1650.350 ;
        RECT 1399.420 1650.030 1399.680 1650.350 ;
        RECT 1399.480 18.205 1399.620 1650.030 ;
        RECT 1399.410 17.835 1399.690 18.205 ;
        RECT 2375.530 17.835 2375.810 18.205 ;
        RECT 2375.600 2.400 2375.740 17.835 ;
        RECT 2375.390 -4.800 2375.950 2.400 ;
      LAYER via2 ;
        RECT 1399.410 17.880 1399.690 18.160 ;
        RECT 2375.530 17.880 2375.810 18.160 ;
      LAYER met3 ;
        RECT 1399.385 18.170 1399.715 18.185 ;
        RECT 2375.505 18.170 2375.835 18.185 ;
        RECT 1399.385 17.870 2375.835 18.170 ;
        RECT 1399.385 17.855 1399.715 17.870 ;
        RECT 2375.505 17.855 2375.835 17.870 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1395.710 1685.280 1396.030 1685.340 ;
        RECT 1400.310 1685.280 1400.630 1685.340 ;
        RECT 1395.710 1685.140 1400.630 1685.280 ;
        RECT 1395.710 1685.080 1396.030 1685.140 ;
        RECT 1400.310 1685.080 1400.630 1685.140 ;
      LAYER via ;
        RECT 1395.740 1685.080 1396.000 1685.340 ;
        RECT 1400.340 1685.080 1400.600 1685.340 ;
      LAYER met2 ;
        RECT 1395.640 1700.340 1395.920 1704.000 ;
        RECT 1395.640 1700.000 1395.940 1700.340 ;
        RECT 1395.800 1685.370 1395.940 1700.000 ;
        RECT 1395.740 1685.050 1396.000 1685.370 ;
        RECT 1400.340 1685.050 1400.600 1685.370 ;
        RECT 1400.400 39.850 1400.540 1685.050 ;
        RECT 1399.940 39.710 1400.540 39.850 ;
        RECT 1399.940 17.525 1400.080 39.710 ;
        RECT 1399.870 17.155 1400.150 17.525 ;
        RECT 2393.470 17.155 2393.750 17.525 ;
        RECT 2393.540 2.400 2393.680 17.155 ;
        RECT 2393.330 -4.800 2393.890 2.400 ;
      LAYER via2 ;
        RECT 1399.870 17.200 1400.150 17.480 ;
        RECT 2393.470 17.200 2393.750 17.480 ;
      LAYER met3 ;
        RECT 1399.845 17.490 1400.175 17.505 ;
        RECT 2393.445 17.490 2393.775 17.505 ;
        RECT 1399.845 17.190 2393.775 17.490 ;
        RECT 1399.845 17.175 1400.175 17.190 ;
        RECT 2393.445 17.175 2393.775 17.190 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1397.550 1683.920 1397.870 1683.980 ;
        RECT 1399.850 1683.920 1400.170 1683.980 ;
        RECT 1397.550 1683.780 1400.170 1683.920 ;
        RECT 1397.550 1683.720 1397.870 1683.780 ;
        RECT 1399.850 1683.720 1400.170 1683.780 ;
        RECT 1398.930 40.360 1399.250 40.420 ;
        RECT 1399.850 40.360 1400.170 40.420 ;
        RECT 1398.930 40.220 1400.170 40.360 ;
        RECT 1398.930 40.160 1399.250 40.220 ;
        RECT 1399.850 40.160 1400.170 40.220 ;
      LAYER via ;
        RECT 1397.580 1683.720 1397.840 1683.980 ;
        RECT 1399.880 1683.720 1400.140 1683.980 ;
        RECT 1398.960 40.160 1399.220 40.420 ;
        RECT 1399.880 40.160 1400.140 40.420 ;
      LAYER met2 ;
        RECT 1397.480 1700.340 1397.760 1704.000 ;
        RECT 1397.480 1700.000 1397.780 1700.340 ;
        RECT 1397.640 1684.010 1397.780 1700.000 ;
        RECT 1397.580 1683.690 1397.840 1684.010 ;
        RECT 1399.880 1683.690 1400.140 1684.010 ;
        RECT 1399.940 40.450 1400.080 1683.690 ;
        RECT 1398.960 40.130 1399.220 40.450 ;
        RECT 1399.880 40.130 1400.140 40.450 ;
        RECT 1399.020 16.845 1399.160 40.130 ;
        RECT 1398.950 16.475 1399.230 16.845 ;
        RECT 2411.410 16.475 2411.690 16.845 ;
        RECT 2411.480 2.400 2411.620 16.475 ;
        RECT 2411.270 -4.800 2411.830 2.400 ;
      LAYER via2 ;
        RECT 1398.950 16.520 1399.230 16.800 ;
        RECT 2411.410 16.520 2411.690 16.800 ;
      LAYER met3 ;
        RECT 1398.925 16.810 1399.255 16.825 ;
        RECT 2411.385 16.810 2411.715 16.825 ;
        RECT 1398.925 16.510 2411.715 16.810 ;
        RECT 1398.925 16.495 1399.255 16.510 ;
        RECT 2411.385 16.495 2411.715 16.510 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 806.910 1563.220 807.230 1563.280 ;
        RECT 1231.490 1563.220 1231.810 1563.280 ;
        RECT 806.910 1563.080 1231.810 1563.220 ;
        RECT 806.910 1563.020 807.230 1563.080 ;
        RECT 1231.490 1563.020 1231.810 1563.080 ;
      LAYER via ;
        RECT 806.940 1563.020 807.200 1563.280 ;
        RECT 1231.520 1563.020 1231.780 1563.280 ;
      LAYER met2 ;
        RECT 1232.340 1700.340 1232.620 1704.000 ;
        RECT 1232.340 1700.000 1232.640 1700.340 ;
        RECT 1232.500 1677.970 1232.640 1700.000 ;
        RECT 1231.580 1677.830 1232.640 1677.970 ;
        RECT 1231.580 1563.310 1231.720 1677.830 ;
        RECT 806.940 1562.990 807.200 1563.310 ;
        RECT 1231.520 1562.990 1231.780 1563.310 ;
        RECT 807.000 18.090 807.140 1562.990 ;
        RECT 805.620 17.950 807.140 18.090 ;
        RECT 805.620 2.400 805.760 17.950 ;
        RECT 805.410 -4.800 805.970 2.400 ;
    END
  END la_oen[9]
  PIN user_clock2
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2916.810 -4.800 2917.370 2.400 ;
    END
  END user_clock2
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1121.165 23.885 1121.335 25.075 ;
      LAYER mcon ;
        RECT 1121.165 24.905 1121.335 25.075 ;
      LAYER met1 ;
        RECT 1121.105 25.060 1121.395 25.105 ;
        RECT 1145.930 25.060 1146.250 25.120 ;
        RECT 1121.105 24.920 1146.250 25.060 ;
        RECT 1121.105 24.875 1121.395 24.920 ;
        RECT 1145.930 24.860 1146.250 24.920 ;
        RECT 2.830 24.040 3.150 24.100 ;
        RECT 1121.105 24.040 1121.395 24.085 ;
        RECT 2.830 23.900 1121.395 24.040 ;
        RECT 2.830 23.840 3.150 23.900 ;
        RECT 1121.105 23.855 1121.395 23.900 ;
      LAYER via ;
        RECT 1145.960 24.860 1146.220 25.120 ;
        RECT 2.860 23.840 3.120 24.100 ;
      LAYER met2 ;
        RECT 1150.000 1700.410 1150.280 1704.000 ;
        RECT 1146.020 1700.270 1150.280 1700.410 ;
        RECT 1146.020 25.150 1146.160 1700.270 ;
        RECT 1150.000 1700.000 1150.280 1700.270 ;
        RECT 1145.960 24.830 1146.220 25.150 ;
        RECT 2.860 23.810 3.120 24.130 ;
        RECT 2.920 2.400 3.060 23.810 ;
        RECT 2.710 -4.800 3.270 2.400 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 8.350 24.380 8.670 24.440 ;
        RECT 8.350 24.240 1121.780 24.380 ;
        RECT 8.350 24.180 8.670 24.240 ;
        RECT 1121.640 24.040 1121.780 24.240 ;
        RECT 1146.390 24.040 1146.710 24.100 ;
        RECT 1121.640 23.900 1146.710 24.040 ;
        RECT 1146.390 23.840 1146.710 23.900 ;
      LAYER via ;
        RECT 8.380 24.180 8.640 24.440 ;
        RECT 1146.420 23.840 1146.680 24.100 ;
      LAYER met2 ;
        RECT 1150.460 1700.340 1150.740 1704.000 ;
        RECT 1150.460 1700.000 1150.760 1700.340 ;
        RECT 1150.620 1678.650 1150.760 1700.000 ;
        RECT 1146.480 1678.510 1150.760 1678.650 ;
        RECT 8.380 24.150 8.640 24.470 ;
        RECT 8.440 2.400 8.580 24.150 ;
        RECT 1146.480 24.130 1146.620 1678.510 ;
        RECT 1146.420 23.810 1146.680 24.130 ;
        RECT 8.230 -4.800 8.790 2.400 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1150.990 1678.480 1151.310 1678.540 ;
        RECT 1146.940 1678.340 1151.310 1678.480 ;
        RECT 1146.940 1678.200 1147.080 1678.340 ;
        RECT 1150.990 1678.280 1151.310 1678.340 ;
        RECT 1146.850 1677.940 1147.170 1678.200 ;
        RECT 14.330 24.720 14.650 24.780 ;
        RECT 1146.850 24.720 1147.170 24.780 ;
        RECT 14.330 24.580 1147.170 24.720 ;
        RECT 14.330 24.520 14.650 24.580 ;
        RECT 1146.850 24.520 1147.170 24.580 ;
      LAYER via ;
        RECT 1151.020 1678.280 1151.280 1678.540 ;
        RECT 1146.880 1677.940 1147.140 1678.200 ;
        RECT 14.360 24.520 14.620 24.780 ;
        RECT 1146.880 24.520 1147.140 24.780 ;
      LAYER met2 ;
        RECT 1150.920 1700.340 1151.200 1704.000 ;
        RECT 1150.920 1700.000 1151.220 1700.340 ;
        RECT 1151.080 1678.570 1151.220 1700.000 ;
        RECT 1151.020 1678.250 1151.280 1678.570 ;
        RECT 1146.880 1677.910 1147.140 1678.230 ;
        RECT 1146.940 24.810 1147.080 1677.910 ;
        RECT 14.360 24.490 14.620 24.810 ;
        RECT 1146.880 24.490 1147.140 24.810 ;
        RECT 14.420 2.400 14.560 24.490 ;
        RECT 14.210 -4.800 14.770 2.400 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1120.705 22.865 1120.875 25.075 ;
      LAYER mcon ;
        RECT 1120.705 24.905 1120.875 25.075 ;
      LAYER met1 ;
        RECT 38.250 25.060 38.570 25.120 ;
        RECT 1120.645 25.060 1120.935 25.105 ;
        RECT 38.250 24.920 1120.935 25.060 ;
        RECT 38.250 24.860 38.570 24.920 ;
        RECT 1120.645 24.875 1120.935 24.920 ;
        RECT 1120.645 23.020 1120.935 23.065 ;
        RECT 1153.750 23.020 1154.070 23.080 ;
        RECT 1120.645 22.880 1154.070 23.020 ;
        RECT 1120.645 22.835 1120.935 22.880 ;
        RECT 1153.750 22.820 1154.070 22.880 ;
      LAYER via ;
        RECT 38.280 24.860 38.540 25.120 ;
        RECT 1153.780 22.820 1154.040 23.080 ;
      LAYER met2 ;
        RECT 1153.220 1700.410 1153.500 1704.000 ;
        RECT 1153.220 1700.270 1153.980 1700.410 ;
        RECT 1153.220 1700.000 1153.500 1700.270 ;
        RECT 38.280 24.830 38.540 25.150 ;
        RECT 38.340 2.400 38.480 24.830 ;
        RECT 1153.840 23.110 1153.980 1700.270 ;
        RECT 1153.780 22.790 1154.040 23.110 ;
        RECT 38.130 -4.800 38.690 2.400 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1159.730 1685.620 1160.050 1685.680 ;
        RECT 1174.450 1685.620 1174.770 1685.680 ;
        RECT 1159.730 1685.480 1174.770 1685.620 ;
        RECT 1159.730 1685.420 1160.050 1685.480 ;
        RECT 1174.450 1685.420 1174.770 1685.480 ;
        RECT 241.110 1659.780 241.430 1659.840 ;
        RECT 1159.730 1659.780 1160.050 1659.840 ;
        RECT 241.110 1659.640 1160.050 1659.780 ;
        RECT 241.110 1659.580 241.430 1659.640 ;
        RECT 1159.730 1659.580 1160.050 1659.640 ;
      LAYER via ;
        RECT 1159.760 1685.420 1160.020 1685.680 ;
        RECT 1174.480 1685.420 1174.740 1685.680 ;
        RECT 241.140 1659.580 241.400 1659.840 ;
        RECT 1159.760 1659.580 1160.020 1659.840 ;
      LAYER met2 ;
        RECT 1174.380 1700.340 1174.660 1704.000 ;
        RECT 1174.380 1700.000 1174.680 1700.340 ;
        RECT 1174.540 1685.710 1174.680 1700.000 ;
        RECT 1159.760 1685.390 1160.020 1685.710 ;
        RECT 1174.480 1685.390 1174.740 1685.710 ;
        RECT 1159.820 1659.870 1159.960 1685.390 ;
        RECT 241.140 1659.550 241.400 1659.870 ;
        RECT 1159.760 1659.550 1160.020 1659.870 ;
        RECT 241.200 17.410 241.340 1659.550 ;
        RECT 240.740 17.270 241.340 17.410 ;
        RECT 240.740 2.400 240.880 17.270 ;
        RECT 240.530 -4.800 241.090 2.400 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 289.945 1680.025 290.115 1680.875 ;
        RECT 313.865 1679.685 314.035 1680.875 ;
        RECT 338.245 1679.005 338.415 1679.855 ;
        RECT 386.085 1679.005 386.255 1679.855 ;
        RECT 386.545 1679.005 386.715 1679.855 ;
        RECT 408.165 1679.005 408.335 1679.855 ;
        RECT 434.845 1679.005 435.015 1679.855 ;
        RECT 482.685 1679.005 482.855 1679.855 ;
        RECT 483.145 1679.005 483.315 1679.855 ;
        RECT 531.445 1679.685 532.535 1679.855 ;
        RECT 531.445 1679.345 531.615 1679.685 ;
        RECT 579.745 1679.005 579.915 1679.855 ;
        RECT 645.525 1679.515 645.695 1680.195 ;
        RECT 882.885 1680.025 883.975 1680.195 ;
        RECT 645.065 1679.345 645.695 1679.515 ;
        RECT 662.545 1679.005 662.715 1679.855 ;
        RECT 710.385 1679.005 710.555 1679.855 ;
        RECT 717.745 1679.685 718.375 1679.855 ;
        RECT 883.805 1679.685 883.975 1680.025 ;
        RECT 718.205 1679.345 718.375 1679.685 ;
        RECT 897.145 1679.005 897.315 1679.855 ;
        RECT 944.985 1679.005 945.155 1679.855 ;
        RECT 945.445 1679.005 945.615 1679.855 ;
        RECT 980.405 1679.005 980.575 1679.855 ;
        RECT 993.745 1679.005 993.915 1679.855 ;
        RECT 1041.585 1679.005 1041.755 1679.855 ;
        RECT 1048.485 1679.685 1049.115 1679.855 ;
      LAYER mcon ;
        RECT 289.945 1680.705 290.115 1680.875 ;
        RECT 313.865 1680.705 314.035 1680.875 ;
        RECT 645.525 1680.025 645.695 1680.195 ;
        RECT 338.245 1679.685 338.415 1679.855 ;
        RECT 386.085 1679.685 386.255 1679.855 ;
        RECT 386.545 1679.685 386.715 1679.855 ;
        RECT 408.165 1679.685 408.335 1679.855 ;
        RECT 434.845 1679.685 435.015 1679.855 ;
        RECT 482.685 1679.685 482.855 1679.855 ;
        RECT 483.145 1679.685 483.315 1679.855 ;
        RECT 532.365 1679.685 532.535 1679.855 ;
        RECT 579.745 1679.685 579.915 1679.855 ;
        RECT 662.545 1679.685 662.715 1679.855 ;
        RECT 710.385 1679.685 710.555 1679.855 ;
        RECT 897.145 1679.685 897.315 1679.855 ;
        RECT 944.985 1679.685 945.155 1679.855 ;
        RECT 945.445 1679.685 945.615 1679.855 ;
        RECT 980.405 1679.685 980.575 1679.855 ;
        RECT 993.745 1679.685 993.915 1679.855 ;
        RECT 1041.585 1679.685 1041.755 1679.855 ;
        RECT 1048.945 1679.685 1049.115 1679.855 ;
      LAYER met1 ;
        RECT 1166.170 1683.920 1166.490 1683.980 ;
        RECT 1176.290 1683.920 1176.610 1683.980 ;
        RECT 1166.170 1683.780 1176.610 1683.920 ;
        RECT 1166.170 1683.720 1166.490 1683.780 ;
        RECT 1176.290 1683.720 1176.610 1683.780 ;
        RECT 289.885 1680.860 290.175 1680.905 ;
        RECT 313.805 1680.860 314.095 1680.905 ;
        RECT 289.885 1680.720 314.095 1680.860 ;
        RECT 289.885 1680.675 290.175 1680.720 ;
        RECT 313.805 1680.675 314.095 1680.720 ;
        RECT 261.810 1680.180 262.130 1680.240 ;
        RECT 289.885 1680.180 290.175 1680.225 ;
        RECT 645.465 1680.180 645.755 1680.225 ;
        RECT 765.510 1680.180 765.830 1680.240 ;
        RECT 882.825 1680.180 883.115 1680.225 ;
        RECT 261.810 1680.040 290.175 1680.180 ;
        RECT 261.810 1679.980 262.130 1680.040 ;
        RECT 289.885 1679.995 290.175 1680.040 ;
        RECT 386.100 1680.040 386.700 1680.180 ;
        RECT 386.100 1679.885 386.240 1680.040 ;
        RECT 386.560 1679.885 386.700 1680.040 ;
        RECT 482.700 1680.040 483.300 1680.180 ;
        RECT 482.700 1679.885 482.840 1680.040 ;
        RECT 483.160 1679.885 483.300 1680.040 ;
        RECT 546.180 1680.040 579.900 1680.180 ;
        RECT 313.805 1679.840 314.095 1679.885 ;
        RECT 338.185 1679.840 338.475 1679.885 ;
        RECT 313.805 1679.700 338.475 1679.840 ;
        RECT 313.805 1679.655 314.095 1679.700 ;
        RECT 338.185 1679.655 338.475 1679.700 ;
        RECT 386.025 1679.655 386.315 1679.885 ;
        RECT 386.485 1679.655 386.775 1679.885 ;
        RECT 408.105 1679.840 408.395 1679.885 ;
        RECT 434.785 1679.840 435.075 1679.885 ;
        RECT 408.105 1679.700 435.075 1679.840 ;
        RECT 408.105 1679.655 408.395 1679.700 ;
        RECT 434.785 1679.655 435.075 1679.700 ;
        RECT 482.625 1679.655 482.915 1679.885 ;
        RECT 483.085 1679.655 483.375 1679.885 ;
        RECT 532.305 1679.840 532.595 1679.885 ;
        RECT 546.180 1679.840 546.320 1680.040 ;
        RECT 579.760 1679.885 579.900 1680.040 ;
        RECT 645.465 1680.040 662.700 1680.180 ;
        RECT 645.465 1679.995 645.755 1680.040 ;
        RECT 662.560 1679.885 662.700 1680.040 ;
        RECT 765.510 1680.040 766.200 1680.180 ;
        RECT 765.510 1679.980 765.830 1680.040 ;
        RECT 531.000 1679.700 531.600 1679.840 ;
        RECT 338.185 1679.160 338.475 1679.205 ;
        RECT 386.025 1679.160 386.315 1679.205 ;
        RECT 338.185 1679.020 386.315 1679.160 ;
        RECT 338.185 1678.975 338.475 1679.020 ;
        RECT 386.025 1678.975 386.315 1679.020 ;
        RECT 386.485 1679.160 386.775 1679.205 ;
        RECT 408.105 1679.160 408.395 1679.205 ;
        RECT 386.485 1679.020 408.395 1679.160 ;
        RECT 386.485 1678.975 386.775 1679.020 ;
        RECT 408.105 1678.975 408.395 1679.020 ;
        RECT 434.785 1679.160 435.075 1679.205 ;
        RECT 482.625 1679.160 482.915 1679.205 ;
        RECT 434.785 1679.020 482.915 1679.160 ;
        RECT 434.785 1678.975 435.075 1679.020 ;
        RECT 482.625 1678.975 482.915 1679.020 ;
        RECT 483.085 1679.160 483.375 1679.205 ;
        RECT 531.000 1679.160 531.140 1679.700 ;
        RECT 531.460 1679.545 531.600 1679.700 ;
        RECT 532.305 1679.700 546.320 1679.840 ;
        RECT 532.305 1679.655 532.595 1679.700 ;
        RECT 579.685 1679.655 579.975 1679.885 ;
        RECT 662.485 1679.655 662.775 1679.885 ;
        RECT 710.325 1679.840 710.615 1679.885 ;
        RECT 717.685 1679.840 717.975 1679.885 ;
        RECT 710.325 1679.700 717.975 1679.840 ;
        RECT 766.060 1679.840 766.200 1680.040 ;
        RECT 766.520 1680.040 883.115 1680.180 ;
        RECT 766.520 1679.840 766.660 1680.040 ;
        RECT 882.825 1679.995 883.115 1680.040 ;
        RECT 945.000 1680.040 945.600 1680.180 ;
        RECT 945.000 1679.885 945.140 1680.040 ;
        RECT 945.460 1679.885 945.600 1680.040 ;
        RECT 766.060 1679.700 766.660 1679.840 ;
        RECT 883.745 1679.840 884.035 1679.885 ;
        RECT 897.085 1679.840 897.375 1679.885 ;
        RECT 883.745 1679.700 897.375 1679.840 ;
        RECT 710.325 1679.655 710.615 1679.700 ;
        RECT 717.685 1679.655 717.975 1679.700 ;
        RECT 883.745 1679.655 884.035 1679.700 ;
        RECT 897.085 1679.655 897.375 1679.700 ;
        RECT 944.925 1679.655 945.215 1679.885 ;
        RECT 945.385 1679.655 945.675 1679.885 ;
        RECT 980.345 1679.840 980.635 1679.885 ;
        RECT 993.685 1679.840 993.975 1679.885 ;
        RECT 980.345 1679.700 993.975 1679.840 ;
        RECT 980.345 1679.655 980.635 1679.700 ;
        RECT 993.685 1679.655 993.975 1679.700 ;
        RECT 1041.525 1679.840 1041.815 1679.885 ;
        RECT 1048.425 1679.840 1048.715 1679.885 ;
        RECT 1041.525 1679.700 1048.715 1679.840 ;
        RECT 1041.525 1679.655 1041.815 1679.700 ;
        RECT 1048.425 1679.655 1048.715 1679.700 ;
        RECT 1048.885 1679.840 1049.175 1679.885 ;
        RECT 1048.885 1679.700 1090.040 1679.840 ;
        RECT 1048.885 1679.655 1049.175 1679.700 ;
        RECT 531.385 1679.315 531.675 1679.545 ;
        RECT 645.005 1679.500 645.295 1679.545 ;
        RECT 595.860 1679.360 645.295 1679.500 ;
        RECT 483.085 1679.020 531.140 1679.160 ;
        RECT 579.685 1679.160 579.975 1679.205 ;
        RECT 595.860 1679.160 596.000 1679.360 ;
        RECT 645.005 1679.315 645.295 1679.360 ;
        RECT 718.145 1679.500 718.435 1679.545 ;
        RECT 765.510 1679.500 765.830 1679.560 ;
        RECT 718.145 1679.360 765.830 1679.500 ;
        RECT 1089.900 1679.500 1090.040 1679.700 ;
        RECT 1166.170 1679.500 1166.490 1679.560 ;
        RECT 1089.900 1679.360 1166.490 1679.500 ;
        RECT 718.145 1679.315 718.435 1679.360 ;
        RECT 765.510 1679.300 765.830 1679.360 ;
        RECT 1166.170 1679.300 1166.490 1679.360 ;
        RECT 579.685 1679.020 596.000 1679.160 ;
        RECT 662.485 1679.160 662.775 1679.205 ;
        RECT 710.325 1679.160 710.615 1679.205 ;
        RECT 662.485 1679.020 710.615 1679.160 ;
        RECT 483.085 1678.975 483.375 1679.020 ;
        RECT 579.685 1678.975 579.975 1679.020 ;
        RECT 662.485 1678.975 662.775 1679.020 ;
        RECT 710.325 1678.975 710.615 1679.020 ;
        RECT 897.085 1679.160 897.375 1679.205 ;
        RECT 944.925 1679.160 945.215 1679.205 ;
        RECT 897.085 1679.020 945.215 1679.160 ;
        RECT 897.085 1678.975 897.375 1679.020 ;
        RECT 944.925 1678.975 945.215 1679.020 ;
        RECT 945.385 1679.160 945.675 1679.205 ;
        RECT 980.345 1679.160 980.635 1679.205 ;
        RECT 945.385 1679.020 980.635 1679.160 ;
        RECT 945.385 1678.975 945.675 1679.020 ;
        RECT 980.345 1678.975 980.635 1679.020 ;
        RECT 993.685 1679.160 993.975 1679.205 ;
        RECT 1041.525 1679.160 1041.815 1679.205 ;
        RECT 993.685 1679.020 1041.815 1679.160 ;
        RECT 993.685 1678.975 993.975 1679.020 ;
        RECT 1041.525 1678.975 1041.815 1679.020 ;
        RECT 258.130 17.920 258.450 17.980 ;
        RECT 261.810 17.920 262.130 17.980 ;
        RECT 258.130 17.780 262.130 17.920 ;
        RECT 258.130 17.720 258.450 17.780 ;
        RECT 261.810 17.720 262.130 17.780 ;
      LAYER via ;
        RECT 1166.200 1683.720 1166.460 1683.980 ;
        RECT 1176.320 1683.720 1176.580 1683.980 ;
        RECT 261.840 1679.980 262.100 1680.240 ;
        RECT 765.540 1679.980 765.800 1680.240 ;
        RECT 765.540 1679.300 765.800 1679.560 ;
        RECT 1166.200 1679.300 1166.460 1679.560 ;
        RECT 258.160 17.720 258.420 17.980 ;
        RECT 261.840 17.720 262.100 17.980 ;
      LAYER met2 ;
        RECT 1176.220 1700.340 1176.500 1704.000 ;
        RECT 1176.220 1700.000 1176.520 1700.340 ;
        RECT 1176.380 1684.010 1176.520 1700.000 ;
        RECT 1166.200 1683.690 1166.460 1684.010 ;
        RECT 1176.320 1683.690 1176.580 1684.010 ;
        RECT 261.840 1679.950 262.100 1680.270 ;
        RECT 765.540 1679.950 765.800 1680.270 ;
        RECT 261.900 18.010 262.040 1679.950 ;
        RECT 765.600 1679.590 765.740 1679.950 ;
        RECT 1166.260 1679.590 1166.400 1683.690 ;
        RECT 765.540 1679.270 765.800 1679.590 ;
        RECT 1166.200 1679.270 1166.460 1679.590 ;
        RECT 258.160 17.690 258.420 18.010 ;
        RECT 261.840 17.690 262.100 18.010 ;
        RECT 258.220 2.400 258.360 17.690 ;
        RECT 258.010 -4.800 258.570 2.400 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 282.510 1673.040 282.830 1673.100 ;
        RECT 1178.130 1673.040 1178.450 1673.100 ;
        RECT 282.510 1672.900 1178.450 1673.040 ;
        RECT 282.510 1672.840 282.830 1672.900 ;
        RECT 1178.130 1672.840 1178.450 1672.900 ;
        RECT 276.070 16.900 276.390 16.960 ;
        RECT 282.510 16.900 282.830 16.960 ;
        RECT 276.070 16.760 282.830 16.900 ;
        RECT 276.070 16.700 276.390 16.760 ;
        RECT 282.510 16.700 282.830 16.760 ;
      LAYER via ;
        RECT 282.540 1672.840 282.800 1673.100 ;
        RECT 1178.160 1672.840 1178.420 1673.100 ;
        RECT 276.100 16.700 276.360 16.960 ;
        RECT 282.540 16.700 282.800 16.960 ;
      LAYER met2 ;
        RECT 1178.060 1700.340 1178.340 1704.000 ;
        RECT 1178.060 1700.000 1178.360 1700.340 ;
        RECT 1178.220 1673.130 1178.360 1700.000 ;
        RECT 282.540 1672.810 282.800 1673.130 ;
        RECT 1178.160 1672.810 1178.420 1673.130 ;
        RECT 282.600 16.990 282.740 1672.810 ;
        RECT 276.100 16.670 276.360 16.990 ;
        RECT 282.540 16.670 282.800 16.990 ;
        RECT 276.160 2.400 276.300 16.670 ;
        RECT 275.950 -4.800 276.510 2.400 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1179.970 1677.460 1180.290 1677.520 ;
        RECT 1182.270 1677.460 1182.590 1677.520 ;
        RECT 1179.970 1677.320 1182.590 1677.460 ;
        RECT 1179.970 1677.260 1180.290 1677.320 ;
        RECT 1182.270 1677.260 1182.590 1677.320 ;
        RECT 294.010 45.120 294.330 45.180 ;
        RECT 1182.270 45.120 1182.590 45.180 ;
        RECT 294.010 44.980 1182.590 45.120 ;
        RECT 294.010 44.920 294.330 44.980 ;
        RECT 1182.270 44.920 1182.590 44.980 ;
      LAYER via ;
        RECT 1180.000 1677.260 1180.260 1677.520 ;
        RECT 1182.300 1677.260 1182.560 1677.520 ;
        RECT 294.040 44.920 294.300 45.180 ;
        RECT 1182.300 44.920 1182.560 45.180 ;
      LAYER met2 ;
        RECT 1179.900 1700.340 1180.180 1704.000 ;
        RECT 1179.900 1700.000 1180.200 1700.340 ;
        RECT 1180.060 1677.550 1180.200 1700.000 ;
        RECT 1180.000 1677.230 1180.260 1677.550 ;
        RECT 1182.300 1677.230 1182.560 1677.550 ;
        RECT 1182.360 45.210 1182.500 1677.230 ;
        RECT 294.040 44.890 294.300 45.210 ;
        RECT 1182.300 44.890 1182.560 45.210 ;
        RECT 294.100 2.400 294.240 44.890 ;
        RECT 293.890 -4.800 294.450 2.400 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1181.810 1678.480 1182.130 1678.540 ;
        RECT 1183.190 1678.480 1183.510 1678.540 ;
        RECT 1181.810 1678.340 1183.510 1678.480 ;
        RECT 1181.810 1678.280 1182.130 1678.340 ;
        RECT 1183.190 1678.280 1183.510 1678.340 ;
        RECT 311.950 45.460 312.270 45.520 ;
        RECT 1183.190 45.460 1183.510 45.520 ;
        RECT 311.950 45.320 1183.510 45.460 ;
        RECT 311.950 45.260 312.270 45.320 ;
        RECT 1183.190 45.260 1183.510 45.320 ;
      LAYER via ;
        RECT 1181.840 1678.280 1182.100 1678.540 ;
        RECT 1183.220 1678.280 1183.480 1678.540 ;
        RECT 311.980 45.260 312.240 45.520 ;
        RECT 1183.220 45.260 1183.480 45.520 ;
      LAYER met2 ;
        RECT 1181.740 1700.340 1182.020 1704.000 ;
        RECT 1181.740 1700.000 1182.040 1700.340 ;
        RECT 1181.900 1678.570 1182.040 1700.000 ;
        RECT 1181.840 1678.250 1182.100 1678.570 ;
        RECT 1183.220 1678.250 1183.480 1678.570 ;
        RECT 1183.280 45.550 1183.420 1678.250 ;
        RECT 311.980 45.230 312.240 45.550 ;
        RECT 1183.220 45.230 1183.480 45.550 ;
        RECT 312.040 2.400 312.180 45.230 ;
        RECT 311.830 -4.800 312.390 2.400 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 329.890 45.800 330.210 45.860 ;
        RECT 1181.810 45.800 1182.130 45.860 ;
        RECT 329.890 45.660 1182.130 45.800 ;
        RECT 329.890 45.600 330.210 45.660 ;
        RECT 1181.810 45.600 1182.130 45.660 ;
      LAYER via ;
        RECT 329.920 45.600 330.180 45.860 ;
        RECT 1181.840 45.600 1182.100 45.860 ;
      LAYER met2 ;
        RECT 1183.580 1700.410 1183.860 1704.000 ;
        RECT 1183.280 1700.270 1183.860 1700.410 ;
        RECT 1183.280 1679.330 1183.420 1700.270 ;
        RECT 1183.580 1700.000 1183.860 1700.270 ;
        RECT 1182.820 1679.190 1183.420 1679.330 ;
        RECT 1182.820 1677.970 1182.960 1679.190 ;
        RECT 1181.900 1677.830 1182.960 1677.970 ;
        RECT 1181.900 45.890 1182.040 1677.830 ;
        RECT 329.920 45.570 330.180 45.890 ;
        RECT 1181.840 45.570 1182.100 45.890 ;
        RECT 329.980 2.400 330.120 45.570 ;
        RECT 329.770 -4.800 330.330 2.400 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 347.370 46.140 347.690 46.200 ;
        RECT 1185.490 46.140 1185.810 46.200 ;
        RECT 347.370 46.000 1185.810 46.140 ;
        RECT 347.370 45.940 347.690 46.000 ;
        RECT 1185.490 45.940 1185.810 46.000 ;
      LAYER via ;
        RECT 347.400 45.940 347.660 46.200 ;
        RECT 1185.520 45.940 1185.780 46.200 ;
      LAYER met2 ;
        RECT 1185.420 1700.340 1185.700 1704.000 ;
        RECT 1185.420 1700.000 1185.720 1700.340 ;
        RECT 1185.580 46.230 1185.720 1700.000 ;
        RECT 347.400 45.910 347.660 46.230 ;
        RECT 1185.520 45.910 1185.780 46.230 ;
        RECT 347.460 2.400 347.600 45.910 ;
        RECT 347.250 -4.800 347.810 2.400 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1187.865 1587.205 1188.035 1635.315 ;
        RECT 1187.865 1442.025 1188.035 1490.475 ;
        RECT 1187.865 1220.685 1188.035 1241.935 ;
        RECT 1187.405 1138.745 1187.575 1159.995 ;
        RECT 1188.325 1072.785 1188.495 1096.755 ;
        RECT 1187.865 834.785 1188.035 862.495 ;
        RECT 1187.865 737.885 1188.035 765.935 ;
        RECT 1187.865 669.885 1188.035 717.315 ;
        RECT 1187.865 427.805 1188.035 475.915 ;
        RECT 1187.865 365.925 1188.035 414.035 ;
        RECT 1187.865 179.605 1188.035 227.715 ;
        RECT 1187.865 46.325 1188.035 82.875 ;
      LAYER mcon ;
        RECT 1187.865 1635.145 1188.035 1635.315 ;
        RECT 1187.865 1490.305 1188.035 1490.475 ;
        RECT 1187.865 1241.765 1188.035 1241.935 ;
        RECT 1187.405 1159.825 1187.575 1159.995 ;
        RECT 1188.325 1096.585 1188.495 1096.755 ;
        RECT 1187.865 862.325 1188.035 862.495 ;
        RECT 1187.865 765.765 1188.035 765.935 ;
        RECT 1187.865 717.145 1188.035 717.315 ;
        RECT 1187.865 475.745 1188.035 475.915 ;
        RECT 1187.865 413.865 1188.035 414.035 ;
        RECT 1187.865 227.545 1188.035 227.715 ;
        RECT 1187.865 82.705 1188.035 82.875 ;
      LAYER met1 ;
        RECT 1187.805 1635.300 1188.095 1635.345 ;
        RECT 1188.250 1635.300 1188.570 1635.360 ;
        RECT 1187.805 1635.160 1188.570 1635.300 ;
        RECT 1187.805 1635.115 1188.095 1635.160 ;
        RECT 1188.250 1635.100 1188.570 1635.160 ;
        RECT 1187.790 1587.360 1188.110 1587.420 ;
        RECT 1187.595 1587.220 1188.110 1587.360 ;
        RECT 1187.790 1587.160 1188.110 1587.220 ;
        RECT 1187.790 1545.340 1188.110 1545.600 ;
        RECT 1187.880 1545.200 1188.020 1545.340 ;
        RECT 1188.250 1545.200 1188.570 1545.260 ;
        RECT 1187.880 1545.060 1188.570 1545.200 ;
        RECT 1188.250 1545.000 1188.570 1545.060 ;
        RECT 1187.805 1490.460 1188.095 1490.505 ;
        RECT 1188.250 1490.460 1188.570 1490.520 ;
        RECT 1187.805 1490.320 1188.570 1490.460 ;
        RECT 1187.805 1490.275 1188.095 1490.320 ;
        RECT 1188.250 1490.260 1188.570 1490.320 ;
        RECT 1187.790 1442.180 1188.110 1442.240 ;
        RECT 1187.595 1442.040 1188.110 1442.180 ;
        RECT 1187.790 1441.980 1188.110 1442.040 ;
        RECT 1188.250 1297.820 1188.570 1298.080 ;
        RECT 1188.340 1297.400 1188.480 1297.820 ;
        RECT 1188.250 1297.140 1188.570 1297.400 ;
        RECT 1188.250 1270.140 1188.570 1270.200 ;
        RECT 1187.880 1270.000 1188.570 1270.140 ;
        RECT 1187.880 1269.520 1188.020 1270.000 ;
        RECT 1188.250 1269.940 1188.570 1270.000 ;
        RECT 1187.790 1269.260 1188.110 1269.520 ;
        RECT 1187.790 1241.920 1188.110 1241.980 ;
        RECT 1187.595 1241.780 1188.110 1241.920 ;
        RECT 1187.790 1241.720 1188.110 1241.780 ;
        RECT 1187.805 1220.840 1188.095 1220.885 ;
        RECT 1188.250 1220.840 1188.570 1220.900 ;
        RECT 1187.805 1220.700 1188.570 1220.840 ;
        RECT 1187.805 1220.655 1188.095 1220.700 ;
        RECT 1188.250 1220.640 1188.570 1220.700 ;
        RECT 1187.345 1159.980 1187.635 1160.025 ;
        RECT 1188.250 1159.980 1188.570 1160.040 ;
        RECT 1187.345 1159.840 1188.570 1159.980 ;
        RECT 1187.345 1159.795 1187.635 1159.840 ;
        RECT 1188.250 1159.780 1188.570 1159.840 ;
        RECT 1187.330 1138.900 1187.650 1138.960 ;
        RECT 1187.135 1138.760 1187.650 1138.900 ;
        RECT 1187.330 1138.700 1187.650 1138.760 ;
        RECT 1188.250 1096.740 1188.570 1096.800 ;
        RECT 1188.055 1096.600 1188.570 1096.740 ;
        RECT 1188.250 1096.540 1188.570 1096.600 ;
        RECT 1188.250 1072.940 1188.570 1073.000 ;
        RECT 1188.055 1072.800 1188.570 1072.940 ;
        RECT 1188.250 1072.740 1188.570 1072.800 ;
        RECT 1187.790 1007.320 1188.110 1007.380 ;
        RECT 1188.250 1007.320 1188.570 1007.380 ;
        RECT 1187.790 1007.180 1188.570 1007.320 ;
        RECT 1187.790 1007.120 1188.110 1007.180 ;
        RECT 1188.250 1007.120 1188.570 1007.180 ;
        RECT 1187.790 931.640 1188.110 931.900 ;
        RECT 1187.880 931.160 1188.020 931.640 ;
        RECT 1188.250 931.160 1188.570 931.220 ;
        RECT 1187.880 931.020 1188.570 931.160 ;
        RECT 1188.250 930.960 1188.570 931.020 ;
        RECT 1187.790 869.960 1188.110 870.020 ;
        RECT 1188.250 869.960 1188.570 870.020 ;
        RECT 1187.790 869.820 1188.570 869.960 ;
        RECT 1187.790 869.760 1188.110 869.820 ;
        RECT 1188.250 869.760 1188.570 869.820 ;
        RECT 1187.790 862.480 1188.110 862.540 ;
        RECT 1187.595 862.340 1188.110 862.480 ;
        RECT 1187.790 862.280 1188.110 862.340 ;
        RECT 1187.790 834.940 1188.110 835.000 ;
        RECT 1187.595 834.800 1188.110 834.940 ;
        RECT 1187.790 834.740 1188.110 834.800 ;
        RECT 1187.790 814.200 1188.110 814.260 ;
        RECT 1188.250 814.200 1188.570 814.260 ;
        RECT 1187.790 814.060 1188.570 814.200 ;
        RECT 1187.790 814.000 1188.110 814.060 ;
        RECT 1188.250 814.000 1188.570 814.060 ;
        RECT 1187.790 765.920 1188.110 765.980 ;
        RECT 1187.595 765.780 1188.110 765.920 ;
        RECT 1187.790 765.720 1188.110 765.780 ;
        RECT 1187.790 738.040 1188.110 738.100 ;
        RECT 1187.595 737.900 1188.110 738.040 ;
        RECT 1187.790 737.840 1188.110 737.900 ;
        RECT 1187.805 717.300 1188.095 717.345 ;
        RECT 1188.250 717.300 1188.570 717.360 ;
        RECT 1187.805 717.160 1188.570 717.300 ;
        RECT 1187.805 717.115 1188.095 717.160 ;
        RECT 1188.250 717.100 1188.570 717.160 ;
        RECT 1187.790 670.040 1188.110 670.100 ;
        RECT 1187.595 669.900 1188.110 670.040 ;
        RECT 1187.790 669.840 1188.110 669.900 ;
        RECT 1187.790 566.000 1188.110 566.060 ;
        RECT 1188.250 566.000 1188.570 566.060 ;
        RECT 1187.790 565.860 1188.570 566.000 ;
        RECT 1187.790 565.800 1188.110 565.860 ;
        RECT 1188.250 565.800 1188.570 565.860 ;
        RECT 1188.250 496.980 1188.570 497.040 ;
        RECT 1187.880 496.840 1188.570 496.980 ;
        RECT 1187.880 496.700 1188.020 496.840 ;
        RECT 1188.250 496.780 1188.570 496.840 ;
        RECT 1187.790 496.440 1188.110 496.700 ;
        RECT 1187.790 475.900 1188.110 475.960 ;
        RECT 1187.595 475.760 1188.110 475.900 ;
        RECT 1187.790 475.700 1188.110 475.760 ;
        RECT 1187.805 427.960 1188.095 428.005 ;
        RECT 1188.250 427.960 1188.570 428.020 ;
        RECT 1187.805 427.820 1188.570 427.960 ;
        RECT 1187.805 427.775 1188.095 427.820 ;
        RECT 1188.250 427.760 1188.570 427.820 ;
        RECT 1187.805 414.020 1188.095 414.065 ;
        RECT 1188.250 414.020 1188.570 414.080 ;
        RECT 1187.805 413.880 1188.570 414.020 ;
        RECT 1187.805 413.835 1188.095 413.880 ;
        RECT 1188.250 413.820 1188.570 413.880 ;
        RECT 1187.790 366.080 1188.110 366.140 ;
        RECT 1187.595 365.940 1188.110 366.080 ;
        RECT 1187.790 365.880 1188.110 365.940 ;
        RECT 1187.790 331.740 1188.110 331.800 ;
        RECT 1187.420 331.600 1188.110 331.740 ;
        RECT 1187.420 331.120 1187.560 331.600 ;
        RECT 1187.790 331.540 1188.110 331.600 ;
        RECT 1187.330 330.860 1187.650 331.120 ;
        RECT 1187.330 234.840 1187.650 234.900 ;
        RECT 1187.790 234.840 1188.110 234.900 ;
        RECT 1187.330 234.700 1188.110 234.840 ;
        RECT 1187.330 234.640 1187.650 234.700 ;
        RECT 1187.790 234.640 1188.110 234.700 ;
        RECT 1187.790 227.700 1188.110 227.760 ;
        RECT 1187.595 227.560 1188.110 227.700 ;
        RECT 1187.790 227.500 1188.110 227.560 ;
        RECT 1187.805 179.760 1188.095 179.805 ;
        RECT 1188.250 179.760 1188.570 179.820 ;
        RECT 1187.805 179.620 1188.570 179.760 ;
        RECT 1187.805 179.575 1188.095 179.620 ;
        RECT 1188.250 179.560 1188.570 179.620 ;
        RECT 1187.790 96.800 1188.110 96.860 ;
        RECT 1188.250 96.800 1188.570 96.860 ;
        RECT 1187.790 96.660 1188.570 96.800 ;
        RECT 1187.790 96.600 1188.110 96.660 ;
        RECT 1188.250 96.600 1188.570 96.660 ;
        RECT 1187.790 82.860 1188.110 82.920 ;
        RECT 1187.595 82.720 1188.110 82.860 ;
        RECT 1187.790 82.660 1188.110 82.720 ;
        RECT 365.310 46.480 365.630 46.540 ;
        RECT 1187.805 46.480 1188.095 46.525 ;
        RECT 365.310 46.340 1188.095 46.480 ;
        RECT 365.310 46.280 365.630 46.340 ;
        RECT 1187.805 46.295 1188.095 46.340 ;
      LAYER via ;
        RECT 1188.280 1635.100 1188.540 1635.360 ;
        RECT 1187.820 1587.160 1188.080 1587.420 ;
        RECT 1187.820 1545.340 1188.080 1545.600 ;
        RECT 1188.280 1545.000 1188.540 1545.260 ;
        RECT 1188.280 1490.260 1188.540 1490.520 ;
        RECT 1187.820 1441.980 1188.080 1442.240 ;
        RECT 1188.280 1297.820 1188.540 1298.080 ;
        RECT 1188.280 1297.140 1188.540 1297.400 ;
        RECT 1188.280 1269.940 1188.540 1270.200 ;
        RECT 1187.820 1269.260 1188.080 1269.520 ;
        RECT 1187.820 1241.720 1188.080 1241.980 ;
        RECT 1188.280 1220.640 1188.540 1220.900 ;
        RECT 1188.280 1159.780 1188.540 1160.040 ;
        RECT 1187.360 1138.700 1187.620 1138.960 ;
        RECT 1188.280 1096.540 1188.540 1096.800 ;
        RECT 1188.280 1072.740 1188.540 1073.000 ;
        RECT 1187.820 1007.120 1188.080 1007.380 ;
        RECT 1188.280 1007.120 1188.540 1007.380 ;
        RECT 1187.820 931.640 1188.080 931.900 ;
        RECT 1188.280 930.960 1188.540 931.220 ;
        RECT 1187.820 869.760 1188.080 870.020 ;
        RECT 1188.280 869.760 1188.540 870.020 ;
        RECT 1187.820 862.280 1188.080 862.540 ;
        RECT 1187.820 834.740 1188.080 835.000 ;
        RECT 1187.820 814.000 1188.080 814.260 ;
        RECT 1188.280 814.000 1188.540 814.260 ;
        RECT 1187.820 765.720 1188.080 765.980 ;
        RECT 1187.820 737.840 1188.080 738.100 ;
        RECT 1188.280 717.100 1188.540 717.360 ;
        RECT 1187.820 669.840 1188.080 670.100 ;
        RECT 1187.820 565.800 1188.080 566.060 ;
        RECT 1188.280 565.800 1188.540 566.060 ;
        RECT 1188.280 496.780 1188.540 497.040 ;
        RECT 1187.820 496.440 1188.080 496.700 ;
        RECT 1187.820 475.700 1188.080 475.960 ;
        RECT 1188.280 427.760 1188.540 428.020 ;
        RECT 1188.280 413.820 1188.540 414.080 ;
        RECT 1187.820 365.880 1188.080 366.140 ;
        RECT 1187.820 331.540 1188.080 331.800 ;
        RECT 1187.360 330.860 1187.620 331.120 ;
        RECT 1187.360 234.640 1187.620 234.900 ;
        RECT 1187.820 234.640 1188.080 234.900 ;
        RECT 1187.820 227.500 1188.080 227.760 ;
        RECT 1188.280 179.560 1188.540 179.820 ;
        RECT 1187.820 96.600 1188.080 96.860 ;
        RECT 1188.280 96.600 1188.540 96.860 ;
        RECT 1187.820 82.660 1188.080 82.920 ;
        RECT 365.340 46.280 365.600 46.540 ;
      LAYER met2 ;
        RECT 1187.260 1700.340 1187.540 1704.000 ;
        RECT 1187.260 1700.000 1187.560 1700.340 ;
        RECT 1187.420 1665.050 1187.560 1700.000 ;
        RECT 1187.420 1664.910 1188.480 1665.050 ;
        RECT 1188.340 1635.390 1188.480 1664.910 ;
        RECT 1188.280 1635.070 1188.540 1635.390 ;
        RECT 1187.820 1587.130 1188.080 1587.450 ;
        RECT 1187.880 1545.630 1188.020 1587.130 ;
        RECT 1187.820 1545.310 1188.080 1545.630 ;
        RECT 1188.280 1544.970 1188.540 1545.290 ;
        RECT 1188.340 1490.550 1188.480 1544.970 ;
        RECT 1188.280 1490.230 1188.540 1490.550 ;
        RECT 1187.820 1441.950 1188.080 1442.270 ;
        RECT 1187.880 1414.130 1188.020 1441.950 ;
        RECT 1187.880 1413.990 1188.480 1414.130 ;
        RECT 1188.340 1393.845 1188.480 1413.990 ;
        RECT 1188.270 1393.475 1188.550 1393.845 ;
        RECT 1188.270 1321.395 1188.550 1321.765 ;
        RECT 1188.340 1298.110 1188.480 1321.395 ;
        RECT 1188.280 1297.790 1188.540 1298.110 ;
        RECT 1188.280 1297.110 1188.540 1297.430 ;
        RECT 1188.340 1270.230 1188.480 1297.110 ;
        RECT 1188.280 1269.910 1188.540 1270.230 ;
        RECT 1187.820 1269.230 1188.080 1269.550 ;
        RECT 1187.880 1242.010 1188.020 1269.230 ;
        RECT 1187.820 1241.690 1188.080 1242.010 ;
        RECT 1188.280 1220.610 1188.540 1220.930 ;
        RECT 1188.340 1160.070 1188.480 1220.610 ;
        RECT 1188.280 1159.750 1188.540 1160.070 ;
        RECT 1187.360 1138.670 1187.620 1138.990 ;
        RECT 1187.420 1097.365 1187.560 1138.670 ;
        RECT 1187.350 1096.995 1187.630 1097.365 ;
        RECT 1188.270 1096.995 1188.550 1097.365 ;
        RECT 1188.340 1096.830 1188.480 1096.995 ;
        RECT 1188.280 1096.510 1188.540 1096.830 ;
        RECT 1188.280 1072.710 1188.540 1073.030 ;
        RECT 1188.340 1007.410 1188.480 1072.710 ;
        RECT 1187.820 1007.090 1188.080 1007.410 ;
        RECT 1188.280 1007.090 1188.540 1007.410 ;
        RECT 1187.880 931.930 1188.020 1007.090 ;
        RECT 1187.820 931.610 1188.080 931.930 ;
        RECT 1188.280 930.930 1188.540 931.250 ;
        RECT 1188.340 870.050 1188.480 930.930 ;
        RECT 1187.820 869.730 1188.080 870.050 ;
        RECT 1188.280 869.730 1188.540 870.050 ;
        RECT 1187.880 862.570 1188.020 869.730 ;
        RECT 1187.820 862.250 1188.080 862.570 ;
        RECT 1187.820 834.710 1188.080 835.030 ;
        RECT 1187.880 814.370 1188.020 834.710 ;
        RECT 1187.880 814.290 1188.480 814.370 ;
        RECT 1187.820 814.230 1188.540 814.290 ;
        RECT 1187.820 813.970 1188.080 814.230 ;
        RECT 1188.280 813.970 1188.540 814.230 ;
        RECT 1187.880 766.885 1188.020 813.970 ;
        RECT 1187.810 766.515 1188.090 766.885 ;
        RECT 1187.810 765.835 1188.090 766.205 ;
        RECT 1187.820 765.690 1188.080 765.835 ;
        RECT 1187.820 737.810 1188.080 738.130 ;
        RECT 1187.880 717.810 1188.020 737.810 ;
        RECT 1187.880 717.670 1188.480 717.810 ;
        RECT 1188.340 717.390 1188.480 717.670 ;
        RECT 1188.280 717.070 1188.540 717.390 ;
        RECT 1187.820 669.810 1188.080 670.130 ;
        RECT 1187.880 622.045 1188.020 669.810 ;
        RECT 1187.810 621.675 1188.090 622.045 ;
        RECT 1188.270 620.995 1188.550 621.365 ;
        RECT 1188.340 566.090 1188.480 620.995 ;
        RECT 1187.820 565.770 1188.080 566.090 ;
        RECT 1188.280 565.770 1188.540 566.090 ;
        RECT 1187.880 565.490 1188.020 565.770 ;
        RECT 1187.880 565.350 1188.480 565.490 ;
        RECT 1188.340 497.070 1188.480 565.350 ;
        RECT 1188.280 496.750 1188.540 497.070 ;
        RECT 1187.820 496.410 1188.080 496.730 ;
        RECT 1187.880 475.990 1188.020 496.410 ;
        RECT 1187.820 475.670 1188.080 475.990 ;
        RECT 1188.280 427.730 1188.540 428.050 ;
        RECT 1188.340 414.110 1188.480 427.730 ;
        RECT 1188.280 413.790 1188.540 414.110 ;
        RECT 1187.820 365.850 1188.080 366.170 ;
        RECT 1187.880 331.830 1188.020 365.850 ;
        RECT 1187.820 331.510 1188.080 331.830 ;
        RECT 1187.360 330.830 1187.620 331.150 ;
        RECT 1187.420 324.090 1187.560 330.830 ;
        RECT 1187.420 323.950 1188.480 324.090 ;
        RECT 1188.340 282.610 1188.480 323.950 ;
        RECT 1187.420 282.470 1188.480 282.610 ;
        RECT 1187.420 234.930 1187.560 282.470 ;
        RECT 1187.360 234.610 1187.620 234.930 ;
        RECT 1187.820 234.610 1188.080 234.930 ;
        RECT 1187.880 227.790 1188.020 234.610 ;
        RECT 1187.820 227.470 1188.080 227.790 ;
        RECT 1188.280 179.530 1188.540 179.850 ;
        RECT 1188.340 96.890 1188.480 179.530 ;
        RECT 1187.820 96.570 1188.080 96.890 ;
        RECT 1188.280 96.570 1188.540 96.890 ;
        RECT 1187.880 82.950 1188.020 96.570 ;
        RECT 1187.820 82.630 1188.080 82.950 ;
        RECT 365.340 46.250 365.600 46.570 ;
        RECT 365.400 2.400 365.540 46.250 ;
        RECT 365.190 -4.800 365.750 2.400 ;
      LAYER via2 ;
        RECT 1188.270 1393.520 1188.550 1393.800 ;
        RECT 1188.270 1321.440 1188.550 1321.720 ;
        RECT 1187.350 1097.040 1187.630 1097.320 ;
        RECT 1188.270 1097.040 1188.550 1097.320 ;
        RECT 1187.810 766.560 1188.090 766.840 ;
        RECT 1187.810 765.880 1188.090 766.160 ;
        RECT 1187.810 621.720 1188.090 622.000 ;
        RECT 1188.270 621.040 1188.550 621.320 ;
      LAYER met3 ;
        RECT 1188.245 1393.810 1188.575 1393.825 ;
        RECT 1188.910 1393.810 1189.290 1393.820 ;
        RECT 1188.245 1393.510 1189.290 1393.810 ;
        RECT 1188.245 1393.495 1188.575 1393.510 ;
        RECT 1188.910 1393.500 1189.290 1393.510 ;
        RECT 1188.245 1321.730 1188.575 1321.745 ;
        RECT 1188.910 1321.730 1189.290 1321.740 ;
        RECT 1188.245 1321.430 1189.290 1321.730 ;
        RECT 1188.245 1321.415 1188.575 1321.430 ;
        RECT 1188.910 1321.420 1189.290 1321.430 ;
        RECT 1187.325 1097.330 1187.655 1097.345 ;
        RECT 1188.245 1097.330 1188.575 1097.345 ;
        RECT 1187.325 1097.030 1188.575 1097.330 ;
        RECT 1187.325 1097.015 1187.655 1097.030 ;
        RECT 1188.245 1097.015 1188.575 1097.030 ;
        RECT 1187.785 766.850 1188.115 766.865 ;
        RECT 1187.785 766.535 1188.330 766.850 ;
        RECT 1188.030 766.185 1188.330 766.535 ;
        RECT 1187.785 765.870 1188.330 766.185 ;
        RECT 1187.785 765.855 1188.115 765.870 ;
        RECT 1187.785 622.010 1188.115 622.025 ;
        RECT 1187.785 621.695 1188.330 622.010 ;
        RECT 1188.030 621.345 1188.330 621.695 ;
        RECT 1188.030 621.030 1188.575 621.345 ;
        RECT 1188.245 621.015 1188.575 621.030 ;
      LAYER via3 ;
        RECT 1188.940 1393.500 1189.260 1393.820 ;
        RECT 1188.940 1321.420 1189.260 1321.740 ;
      LAYER met4 ;
        RECT 1188.935 1393.495 1189.265 1393.825 ;
        RECT 1188.950 1321.745 1189.250 1393.495 ;
        RECT 1188.935 1321.415 1189.265 1321.745 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 383.250 46.820 383.570 46.880 ;
        RECT 1189.170 46.820 1189.490 46.880 ;
        RECT 383.250 46.680 1189.490 46.820 ;
        RECT 383.250 46.620 383.570 46.680 ;
        RECT 1189.170 46.620 1189.490 46.680 ;
      LAYER via ;
        RECT 383.280 46.620 383.540 46.880 ;
        RECT 1189.200 46.620 1189.460 46.880 ;
      LAYER met2 ;
        RECT 1189.100 1700.340 1189.380 1704.000 ;
        RECT 1189.100 1700.000 1189.400 1700.340 ;
        RECT 1189.260 46.910 1189.400 1700.000 ;
        RECT 383.280 46.590 383.540 46.910 ;
        RECT 1189.200 46.590 1189.460 46.910 ;
        RECT 383.340 2.400 383.480 46.590 ;
        RECT 383.130 -4.800 383.690 2.400 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1188.710 1678.140 1189.030 1678.200 ;
        RECT 1190.550 1678.140 1190.870 1678.200 ;
        RECT 1188.710 1678.000 1190.870 1678.140 ;
        RECT 1188.710 1677.940 1189.030 1678.000 ;
        RECT 1190.550 1677.940 1190.870 1678.000 ;
        RECT 401.190 47.160 401.510 47.220 ;
        RECT 1188.710 47.160 1189.030 47.220 ;
        RECT 401.190 47.020 1189.030 47.160 ;
        RECT 401.190 46.960 401.510 47.020 ;
        RECT 1188.710 46.960 1189.030 47.020 ;
      LAYER via ;
        RECT 1188.740 1677.940 1189.000 1678.200 ;
        RECT 1190.580 1677.940 1190.840 1678.200 ;
        RECT 401.220 46.960 401.480 47.220 ;
        RECT 1188.740 46.960 1189.000 47.220 ;
      LAYER met2 ;
        RECT 1190.940 1700.410 1191.220 1704.000 ;
        RECT 1190.640 1700.270 1191.220 1700.410 ;
        RECT 1190.640 1678.230 1190.780 1700.270 ;
        RECT 1190.940 1700.000 1191.220 1700.270 ;
        RECT 1188.740 1677.910 1189.000 1678.230 ;
        RECT 1190.580 1677.910 1190.840 1678.230 ;
        RECT 1188.800 47.250 1188.940 1677.910 ;
        RECT 401.220 46.930 401.480 47.250 ;
        RECT 1188.740 46.930 1189.000 47.250 ;
        RECT 401.280 2.400 401.420 46.930 ;
        RECT 401.070 -4.800 401.630 2.400 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1154.210 1028.400 1154.530 1028.460 ;
        RECT 1155.130 1028.400 1155.450 1028.460 ;
        RECT 1154.210 1028.260 1155.450 1028.400 ;
        RECT 1154.210 1028.200 1154.530 1028.260 ;
        RECT 1155.130 1028.200 1155.450 1028.260 ;
        RECT 1154.210 979.780 1154.530 979.840 ;
        RECT 1155.130 979.780 1155.450 979.840 ;
        RECT 1154.210 979.640 1155.450 979.780 ;
        RECT 1154.210 979.580 1154.530 979.640 ;
        RECT 1155.130 979.580 1155.450 979.640 ;
        RECT 1154.210 931.840 1154.530 931.900 ;
        RECT 1155.130 931.840 1155.450 931.900 ;
        RECT 1154.210 931.700 1155.450 931.840 ;
        RECT 1154.210 931.640 1154.530 931.700 ;
        RECT 1155.130 931.640 1155.450 931.700 ;
        RECT 1154.210 883.220 1154.530 883.280 ;
        RECT 1155.130 883.220 1155.450 883.280 ;
        RECT 1154.210 883.080 1155.450 883.220 ;
        RECT 1154.210 883.020 1154.530 883.080 ;
        RECT 1155.130 883.020 1155.450 883.080 ;
        RECT 1154.210 835.280 1154.530 835.340 ;
        RECT 1155.130 835.280 1155.450 835.340 ;
        RECT 1154.210 835.140 1155.450 835.280 ;
        RECT 1154.210 835.080 1154.530 835.140 ;
        RECT 1155.130 835.080 1155.450 835.140 ;
        RECT 1154.210 786.660 1154.530 786.720 ;
        RECT 1155.130 786.660 1155.450 786.720 ;
        RECT 1154.210 786.520 1155.450 786.660 ;
        RECT 1154.210 786.460 1154.530 786.520 ;
        RECT 1155.130 786.460 1155.450 786.520 ;
        RECT 1154.210 255.580 1154.530 255.640 ;
        RECT 1155.130 255.580 1155.450 255.640 ;
        RECT 1154.210 255.440 1155.450 255.580 ;
        RECT 1154.210 255.380 1154.530 255.440 ;
        RECT 1155.130 255.380 1155.450 255.440 ;
        RECT 1154.210 206.960 1154.530 207.020 ;
        RECT 1155.130 206.960 1155.450 207.020 ;
        RECT 1154.210 206.820 1155.450 206.960 ;
        RECT 1154.210 206.760 1154.530 206.820 ;
        RECT 1155.130 206.760 1155.450 206.820 ;
        RECT 1154.210 159.020 1154.530 159.080 ;
        RECT 1155.130 159.020 1155.450 159.080 ;
        RECT 1154.210 158.880 1155.450 159.020 ;
        RECT 1154.210 158.820 1154.530 158.880 ;
        RECT 1155.130 158.820 1155.450 158.880 ;
        RECT 1154.210 110.400 1154.530 110.460 ;
        RECT 1155.130 110.400 1155.450 110.460 ;
        RECT 1154.210 110.260 1155.450 110.400 ;
        RECT 1154.210 110.200 1154.530 110.260 ;
        RECT 1155.130 110.200 1155.450 110.260 ;
        RECT 1154.210 62.460 1154.530 62.520 ;
        RECT 1155.130 62.460 1155.450 62.520 ;
        RECT 1154.210 62.320 1155.450 62.460 ;
        RECT 1154.210 62.260 1154.530 62.320 ;
        RECT 1155.130 62.260 1155.450 62.320 ;
        RECT 62.170 30.840 62.490 30.900 ;
        RECT 1154.210 30.840 1154.530 30.900 ;
        RECT 62.170 30.700 1154.530 30.840 ;
        RECT 62.170 30.640 62.490 30.700 ;
        RECT 1154.210 30.640 1154.530 30.700 ;
      LAYER via ;
        RECT 1154.240 1028.200 1154.500 1028.460 ;
        RECT 1155.160 1028.200 1155.420 1028.460 ;
        RECT 1154.240 979.580 1154.500 979.840 ;
        RECT 1155.160 979.580 1155.420 979.840 ;
        RECT 1154.240 931.640 1154.500 931.900 ;
        RECT 1155.160 931.640 1155.420 931.900 ;
        RECT 1154.240 883.020 1154.500 883.280 ;
        RECT 1155.160 883.020 1155.420 883.280 ;
        RECT 1154.240 835.080 1154.500 835.340 ;
        RECT 1155.160 835.080 1155.420 835.340 ;
        RECT 1154.240 786.460 1154.500 786.720 ;
        RECT 1155.160 786.460 1155.420 786.720 ;
        RECT 1154.240 255.380 1154.500 255.640 ;
        RECT 1155.160 255.380 1155.420 255.640 ;
        RECT 1154.240 206.760 1154.500 207.020 ;
        RECT 1155.160 206.760 1155.420 207.020 ;
        RECT 1154.240 158.820 1154.500 159.080 ;
        RECT 1155.160 158.820 1155.420 159.080 ;
        RECT 1154.240 110.200 1154.500 110.460 ;
        RECT 1155.160 110.200 1155.420 110.460 ;
        RECT 1154.240 62.260 1154.500 62.520 ;
        RECT 1155.160 62.260 1155.420 62.520 ;
        RECT 62.200 30.640 62.460 30.900 ;
        RECT 1154.240 30.640 1154.500 30.900 ;
      LAYER met2 ;
        RECT 1155.980 1700.410 1156.260 1704.000 ;
        RECT 1155.680 1700.270 1156.260 1700.410 ;
        RECT 1155.680 1666.410 1155.820 1700.270 ;
        RECT 1155.980 1700.000 1156.260 1700.270 ;
        RECT 1155.220 1666.270 1155.820 1666.410 ;
        RECT 1155.220 1028.490 1155.360 1666.270 ;
        RECT 1154.240 1028.170 1154.500 1028.490 ;
        RECT 1155.160 1028.170 1155.420 1028.490 ;
        RECT 1154.300 979.870 1154.440 1028.170 ;
        RECT 1154.240 979.550 1154.500 979.870 ;
        RECT 1155.160 979.550 1155.420 979.870 ;
        RECT 1155.220 931.930 1155.360 979.550 ;
        RECT 1154.240 931.610 1154.500 931.930 ;
        RECT 1155.160 931.610 1155.420 931.930 ;
        RECT 1154.300 883.310 1154.440 931.610 ;
        RECT 1154.240 882.990 1154.500 883.310 ;
        RECT 1155.160 882.990 1155.420 883.310 ;
        RECT 1155.220 835.370 1155.360 882.990 ;
        RECT 1154.240 835.050 1154.500 835.370 ;
        RECT 1155.160 835.050 1155.420 835.370 ;
        RECT 1154.300 786.750 1154.440 835.050 ;
        RECT 1154.240 786.430 1154.500 786.750 ;
        RECT 1155.160 786.430 1155.420 786.750 ;
        RECT 1155.220 255.670 1155.360 786.430 ;
        RECT 1154.240 255.350 1154.500 255.670 ;
        RECT 1155.160 255.350 1155.420 255.670 ;
        RECT 1154.300 207.050 1154.440 255.350 ;
        RECT 1154.240 206.730 1154.500 207.050 ;
        RECT 1155.160 206.730 1155.420 207.050 ;
        RECT 1155.220 159.110 1155.360 206.730 ;
        RECT 1154.240 158.790 1154.500 159.110 ;
        RECT 1155.160 158.790 1155.420 159.110 ;
        RECT 1154.300 110.490 1154.440 158.790 ;
        RECT 1154.240 110.170 1154.500 110.490 ;
        RECT 1155.160 110.170 1155.420 110.490 ;
        RECT 1155.220 62.550 1155.360 110.170 ;
        RECT 1154.240 62.230 1154.500 62.550 ;
        RECT 1155.160 62.230 1155.420 62.550 ;
        RECT 1154.300 30.930 1154.440 62.230 ;
        RECT 62.200 30.610 62.460 30.930 ;
        RECT 1154.240 30.610 1154.500 30.930 ;
        RECT 62.260 2.400 62.400 30.610 ;
        RECT 62.050 -4.800 62.610 2.400 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 419.130 47.500 419.450 47.560 ;
        RECT 1192.850 47.500 1193.170 47.560 ;
        RECT 419.130 47.360 1193.170 47.500 ;
        RECT 419.130 47.300 419.450 47.360 ;
        RECT 1192.850 47.300 1193.170 47.360 ;
      LAYER via ;
        RECT 419.160 47.300 419.420 47.560 ;
        RECT 1192.880 47.300 1193.140 47.560 ;
      LAYER met2 ;
        RECT 1192.780 1700.340 1193.060 1704.000 ;
        RECT 1192.780 1700.000 1193.080 1700.340 ;
        RECT 1192.940 47.590 1193.080 1700.000 ;
        RECT 419.160 47.270 419.420 47.590 ;
        RECT 1192.880 47.270 1193.140 47.590 ;
        RECT 419.220 2.400 419.360 47.270 ;
        RECT 419.010 -4.800 419.570 2.400 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 436.610 47.840 436.930 47.900 ;
        RECT 1195.150 47.840 1195.470 47.900 ;
        RECT 436.610 47.700 1195.470 47.840 ;
        RECT 436.610 47.640 436.930 47.700 ;
        RECT 1195.150 47.640 1195.470 47.700 ;
      LAYER via ;
        RECT 436.640 47.640 436.900 47.900 ;
        RECT 1195.180 47.640 1195.440 47.900 ;
      LAYER met2 ;
        RECT 1194.620 1700.340 1194.900 1704.000 ;
        RECT 1194.620 1700.000 1194.920 1700.340 ;
        RECT 1194.780 1667.090 1194.920 1700.000 ;
        RECT 1194.780 1666.950 1195.380 1667.090 ;
        RECT 1195.240 47.930 1195.380 1666.950 ;
        RECT 436.640 47.610 436.900 47.930 ;
        RECT 1195.180 47.610 1195.440 47.930 ;
        RECT 436.700 2.400 436.840 47.610 ;
        RECT 436.490 -4.800 437.050 2.400 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 454.550 48.180 454.870 48.240 ;
        RECT 1196.530 48.180 1196.850 48.240 ;
        RECT 454.550 48.040 1196.850 48.180 ;
        RECT 454.550 47.980 454.870 48.040 ;
        RECT 1196.530 47.980 1196.850 48.040 ;
      LAYER via ;
        RECT 454.580 47.980 454.840 48.240 ;
        RECT 1196.560 47.980 1196.820 48.240 ;
      LAYER met2 ;
        RECT 1196.460 1700.340 1196.740 1704.000 ;
        RECT 1196.460 1700.000 1196.760 1700.340 ;
        RECT 1196.620 48.270 1196.760 1700.000 ;
        RECT 454.580 47.950 454.840 48.270 ;
        RECT 1196.560 47.950 1196.820 48.270 ;
        RECT 454.640 2.400 454.780 47.950 ;
        RECT 454.430 -4.800 454.990 2.400 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1196.070 1668.960 1196.390 1669.020 ;
        RECT 1197.910 1668.960 1198.230 1669.020 ;
        RECT 1196.070 1668.820 1198.230 1668.960 ;
        RECT 1196.070 1668.760 1196.390 1668.820 ;
        RECT 1197.910 1668.760 1198.230 1668.820 ;
        RECT 472.490 44.440 472.810 44.500 ;
        RECT 1196.070 44.440 1196.390 44.500 ;
        RECT 472.490 44.300 1196.390 44.440 ;
        RECT 472.490 44.240 472.810 44.300 ;
        RECT 1196.070 44.240 1196.390 44.300 ;
      LAYER via ;
        RECT 1196.100 1668.760 1196.360 1669.020 ;
        RECT 1197.940 1668.760 1198.200 1669.020 ;
        RECT 472.520 44.240 472.780 44.500 ;
        RECT 1196.100 44.240 1196.360 44.500 ;
      LAYER met2 ;
        RECT 1198.300 1700.410 1198.580 1704.000 ;
        RECT 1198.000 1700.270 1198.580 1700.410 ;
        RECT 1198.000 1669.050 1198.140 1700.270 ;
        RECT 1198.300 1700.000 1198.580 1700.270 ;
        RECT 1196.100 1668.730 1196.360 1669.050 ;
        RECT 1197.940 1668.730 1198.200 1669.050 ;
        RECT 1196.160 44.530 1196.300 1668.730 ;
        RECT 472.520 44.210 472.780 44.530 ;
        RECT 1196.100 44.210 1196.360 44.530 ;
        RECT 472.580 2.400 472.720 44.210 ;
        RECT 472.370 -4.800 472.930 2.400 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 490.430 44.100 490.750 44.160 ;
        RECT 1200.210 44.100 1200.530 44.160 ;
        RECT 490.430 43.960 1200.530 44.100 ;
        RECT 490.430 43.900 490.750 43.960 ;
        RECT 1200.210 43.900 1200.530 43.960 ;
      LAYER via ;
        RECT 490.460 43.900 490.720 44.160 ;
        RECT 1200.240 43.900 1200.500 44.160 ;
      LAYER met2 ;
        RECT 1200.140 1700.340 1200.420 1704.000 ;
        RECT 1200.140 1700.000 1200.440 1700.340 ;
        RECT 1200.300 44.190 1200.440 1700.000 ;
        RECT 490.460 43.870 490.720 44.190 ;
        RECT 1200.240 43.870 1200.500 44.190 ;
        RECT 490.520 2.400 490.660 43.870 ;
        RECT 490.310 -4.800 490.870 2.400 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1202.585 289.765 1202.755 337.875 ;
      LAYER mcon ;
        RECT 1202.585 337.705 1202.755 337.875 ;
      LAYER met1 ;
        RECT 1202.510 1656.180 1202.830 1656.440 ;
        RECT 1202.600 1655.760 1202.740 1656.180 ;
        RECT 1202.510 1655.500 1202.830 1655.760 ;
        RECT 1202.510 337.860 1202.830 337.920 ;
        RECT 1202.315 337.720 1202.830 337.860 ;
        RECT 1202.510 337.660 1202.830 337.720 ;
        RECT 1202.510 289.920 1202.830 289.980 ;
        RECT 1202.315 289.780 1202.830 289.920 ;
        RECT 1202.510 289.720 1202.830 289.780 ;
        RECT 507.910 43.760 508.230 43.820 ;
        RECT 1202.510 43.760 1202.830 43.820 ;
        RECT 507.910 43.620 1202.830 43.760 ;
        RECT 507.910 43.560 508.230 43.620 ;
        RECT 1202.510 43.560 1202.830 43.620 ;
      LAYER via ;
        RECT 1202.540 1656.180 1202.800 1656.440 ;
        RECT 1202.540 1655.500 1202.800 1655.760 ;
        RECT 1202.540 337.660 1202.800 337.920 ;
        RECT 1202.540 289.720 1202.800 289.980 ;
        RECT 507.940 43.560 508.200 43.820 ;
        RECT 1202.540 43.560 1202.800 43.820 ;
      LAYER met2 ;
        RECT 1201.980 1700.340 1202.260 1704.000 ;
        RECT 1201.980 1700.000 1202.280 1700.340 ;
        RECT 1202.140 1678.480 1202.280 1700.000 ;
        RECT 1202.140 1678.340 1202.740 1678.480 ;
        RECT 1202.600 1656.470 1202.740 1678.340 ;
        RECT 1202.540 1656.150 1202.800 1656.470 ;
        RECT 1202.540 1655.470 1202.800 1655.790 ;
        RECT 1202.600 337.950 1202.740 1655.470 ;
        RECT 1202.540 337.630 1202.800 337.950 ;
        RECT 1202.540 289.690 1202.800 290.010 ;
        RECT 1202.600 43.850 1202.740 289.690 ;
        RECT 507.940 43.530 508.200 43.850 ;
        RECT 1202.540 43.530 1202.800 43.850 ;
        RECT 508.000 2.400 508.140 43.530 ;
        RECT 507.790 -4.800 508.350 2.400 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1202.050 1677.800 1202.370 1677.860 ;
        RECT 1203.890 1677.800 1204.210 1677.860 ;
        RECT 1202.050 1677.660 1204.210 1677.800 ;
        RECT 1202.050 1677.600 1202.370 1677.660 ;
        RECT 1203.890 1677.600 1204.210 1677.660 ;
        RECT 525.850 43.420 526.170 43.480 ;
        RECT 1202.050 43.420 1202.370 43.480 ;
        RECT 525.850 43.280 1202.370 43.420 ;
        RECT 525.850 43.220 526.170 43.280 ;
        RECT 1202.050 43.220 1202.370 43.280 ;
      LAYER via ;
        RECT 1202.080 1677.600 1202.340 1677.860 ;
        RECT 1203.920 1677.600 1204.180 1677.860 ;
        RECT 525.880 43.220 526.140 43.480 ;
        RECT 1202.080 43.220 1202.340 43.480 ;
      LAYER met2 ;
        RECT 1203.820 1700.340 1204.100 1704.000 ;
        RECT 1203.820 1700.000 1204.120 1700.340 ;
        RECT 1203.980 1677.890 1204.120 1700.000 ;
        RECT 1202.080 1677.570 1202.340 1677.890 ;
        RECT 1203.920 1677.570 1204.180 1677.890 ;
        RECT 1202.140 43.510 1202.280 1677.570 ;
        RECT 525.880 43.190 526.140 43.510 ;
        RECT 1202.080 43.190 1202.340 43.510 ;
        RECT 525.940 2.400 526.080 43.190 ;
        RECT 525.730 -4.800 526.290 2.400 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1201.590 1678.480 1201.910 1678.540 ;
        RECT 1205.270 1678.480 1205.590 1678.540 ;
        RECT 1201.590 1678.340 1205.590 1678.480 ;
        RECT 1201.590 1678.280 1201.910 1678.340 ;
        RECT 1205.270 1678.280 1205.590 1678.340 ;
        RECT 543.790 43.080 544.110 43.140 ;
        RECT 1201.590 43.080 1201.910 43.140 ;
        RECT 543.790 42.940 1201.910 43.080 ;
        RECT 543.790 42.880 544.110 42.940 ;
        RECT 1201.590 42.880 1201.910 42.940 ;
      LAYER via ;
        RECT 1201.620 1678.280 1201.880 1678.540 ;
        RECT 1205.300 1678.280 1205.560 1678.540 ;
        RECT 543.820 42.880 544.080 43.140 ;
        RECT 1201.620 42.880 1201.880 43.140 ;
      LAYER met2 ;
        RECT 1205.660 1700.410 1205.940 1704.000 ;
        RECT 1205.360 1700.270 1205.940 1700.410 ;
        RECT 1205.360 1678.570 1205.500 1700.270 ;
        RECT 1205.660 1700.000 1205.940 1700.270 ;
        RECT 1201.620 1678.250 1201.880 1678.570 ;
        RECT 1205.300 1678.250 1205.560 1678.570 ;
        RECT 1201.680 43.170 1201.820 1678.250 ;
        RECT 543.820 42.850 544.080 43.170 ;
        RECT 1201.620 42.850 1201.880 43.170 ;
        RECT 543.880 2.400 544.020 42.850 ;
        RECT 543.670 -4.800 544.230 2.400 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1207.570 1678.140 1207.890 1678.200 ;
        RECT 1209.410 1678.140 1209.730 1678.200 ;
        RECT 1207.570 1678.000 1209.730 1678.140 ;
        RECT 1207.570 1677.940 1207.890 1678.000 ;
        RECT 1209.410 1677.940 1209.730 1678.000 ;
        RECT 561.730 42.740 562.050 42.800 ;
        RECT 1209.410 42.740 1209.730 42.800 ;
        RECT 561.730 42.600 1209.730 42.740 ;
        RECT 561.730 42.540 562.050 42.600 ;
        RECT 1209.410 42.540 1209.730 42.600 ;
      LAYER via ;
        RECT 1207.600 1677.940 1207.860 1678.200 ;
        RECT 1209.440 1677.940 1209.700 1678.200 ;
        RECT 561.760 42.540 562.020 42.800 ;
        RECT 1209.440 42.540 1209.700 42.800 ;
      LAYER met2 ;
        RECT 1207.500 1700.340 1207.780 1704.000 ;
        RECT 1207.500 1700.000 1207.800 1700.340 ;
        RECT 1207.660 1678.230 1207.800 1700.000 ;
        RECT 1207.600 1677.910 1207.860 1678.230 ;
        RECT 1209.440 1677.910 1209.700 1678.230 ;
        RECT 1209.500 42.830 1209.640 1677.910 ;
        RECT 561.760 42.510 562.020 42.830 ;
        RECT 1209.440 42.510 1209.700 42.830 ;
        RECT 561.820 2.400 561.960 42.510 ;
        RECT 561.610 -4.800 562.170 2.400 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 579.670 42.400 579.990 42.460 ;
        RECT 1208.950 42.400 1209.270 42.460 ;
        RECT 579.670 42.260 1209.270 42.400 ;
        RECT 579.670 42.200 579.990 42.260 ;
        RECT 1208.950 42.200 1209.270 42.260 ;
      LAYER via ;
        RECT 579.700 42.200 579.960 42.460 ;
        RECT 1208.980 42.200 1209.240 42.460 ;
      LAYER met2 ;
        RECT 1209.340 1700.410 1209.620 1704.000 ;
        RECT 1209.040 1700.270 1209.620 1700.410 ;
        RECT 1209.040 42.490 1209.180 1700.270 ;
        RECT 1209.340 1700.000 1209.620 1700.270 ;
        RECT 579.700 42.170 579.960 42.490 ;
        RECT 1208.980 42.170 1209.240 42.490 ;
        RECT 579.760 2.400 579.900 42.170 ;
        RECT 579.550 -4.800 580.110 2.400 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1158.350 1669.440 1158.670 1669.700 ;
        RECT 1158.440 1669.020 1158.580 1669.440 ;
        RECT 1158.350 1668.760 1158.670 1669.020 ;
        RECT 86.550 44.780 86.870 44.840 ;
        RECT 1158.350 44.780 1158.670 44.840 ;
        RECT 86.550 44.640 1158.670 44.780 ;
        RECT 86.550 44.580 86.870 44.640 ;
        RECT 1158.350 44.580 1158.670 44.640 ;
      LAYER via ;
        RECT 1158.380 1669.440 1158.640 1669.700 ;
        RECT 1158.380 1668.760 1158.640 1669.020 ;
        RECT 86.580 44.580 86.840 44.840 ;
        RECT 1158.380 44.580 1158.640 44.840 ;
      LAYER met2 ;
        RECT 1158.280 1700.340 1158.560 1704.000 ;
        RECT 1158.280 1700.000 1158.580 1700.340 ;
        RECT 1158.440 1669.730 1158.580 1700.000 ;
        RECT 1158.380 1669.410 1158.640 1669.730 ;
        RECT 1158.380 1668.730 1158.640 1669.050 ;
        RECT 1158.440 44.870 1158.580 1668.730 ;
        RECT 86.580 44.550 86.840 44.870 ;
        RECT 1158.380 44.550 1158.640 44.870 ;
        RECT 86.640 7.210 86.780 44.550 ;
        RECT 86.180 7.070 86.780 7.210 ;
        RECT 86.180 2.400 86.320 7.070 ;
        RECT 85.970 -4.800 86.530 2.400 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 597.150 42.060 597.470 42.120 ;
        RECT 1211.250 42.060 1211.570 42.120 ;
        RECT 597.150 41.920 1211.570 42.060 ;
        RECT 597.150 41.860 597.470 41.920 ;
        RECT 1211.250 41.860 1211.570 41.920 ;
      LAYER via ;
        RECT 597.180 41.860 597.440 42.120 ;
        RECT 1211.280 41.860 1211.540 42.120 ;
      LAYER met2 ;
        RECT 1211.180 1700.340 1211.460 1704.000 ;
        RECT 1211.180 1700.000 1211.480 1700.340 ;
        RECT 1211.340 42.150 1211.480 1700.000 ;
        RECT 597.180 41.830 597.440 42.150 ;
        RECT 1211.280 41.830 1211.540 42.150 ;
        RECT 597.240 2.400 597.380 41.830 ;
        RECT 597.030 -4.800 597.590 2.400 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 615.090 41.720 615.410 41.780 ;
        RECT 1213.090 41.720 1213.410 41.780 ;
        RECT 615.090 41.580 1213.410 41.720 ;
        RECT 615.090 41.520 615.410 41.580 ;
        RECT 1213.090 41.520 1213.410 41.580 ;
      LAYER via ;
        RECT 615.120 41.520 615.380 41.780 ;
        RECT 1213.120 41.520 1213.380 41.780 ;
      LAYER met2 ;
        RECT 1213.020 1700.340 1213.300 1704.000 ;
        RECT 1213.020 1700.000 1213.320 1700.340 ;
        RECT 1213.180 41.810 1213.320 1700.000 ;
        RECT 615.120 41.490 615.380 41.810 ;
        RECT 1213.120 41.490 1213.380 41.810 ;
        RECT 615.180 2.400 615.320 41.490 ;
        RECT 614.970 -4.800 615.530 2.400 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1160.650 1670.320 1160.970 1670.380 ;
        RECT 1160.280 1670.180 1160.970 1670.320 ;
        RECT 1160.280 1669.360 1160.420 1670.180 ;
        RECT 1160.650 1670.120 1160.970 1670.180 ;
        RECT 1160.190 1669.100 1160.510 1669.360 ;
        RECT 110.010 52.260 110.330 52.320 ;
        RECT 1160.190 52.260 1160.510 52.320 ;
        RECT 110.010 52.120 1160.510 52.260 ;
        RECT 110.010 52.060 110.330 52.120 ;
        RECT 1160.190 52.060 1160.510 52.120 ;
      LAYER via ;
        RECT 1160.680 1670.120 1160.940 1670.380 ;
        RECT 1160.220 1669.100 1160.480 1669.360 ;
        RECT 110.040 52.060 110.300 52.320 ;
        RECT 1160.220 52.060 1160.480 52.320 ;
      LAYER met2 ;
        RECT 1160.580 1700.340 1160.860 1704.000 ;
        RECT 1160.580 1700.000 1160.880 1700.340 ;
        RECT 1160.740 1670.410 1160.880 1700.000 ;
        RECT 1160.680 1670.090 1160.940 1670.410 ;
        RECT 1160.220 1669.070 1160.480 1669.390 ;
        RECT 1160.280 52.350 1160.420 1669.070 ;
        RECT 110.040 52.030 110.300 52.350 ;
        RECT 1160.220 52.030 1160.480 52.350 ;
        RECT 110.100 17.410 110.240 52.030 ;
        RECT 109.640 17.270 110.240 17.410 ;
        RECT 109.640 2.400 109.780 17.270 ;
        RECT 109.430 -4.800 109.990 2.400 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1160.190 1680.180 1160.510 1680.240 ;
        RECT 1163.410 1680.180 1163.730 1680.240 ;
        RECT 1160.190 1680.040 1163.730 1680.180 ;
        RECT 1160.190 1679.980 1160.510 1680.040 ;
        RECT 1163.410 1679.980 1163.730 1680.040 ;
        RECT 137.610 52.600 137.930 52.660 ;
        RECT 1160.650 52.600 1160.970 52.660 ;
        RECT 137.610 52.460 1160.970 52.600 ;
        RECT 137.610 52.400 137.930 52.460 ;
        RECT 1160.650 52.400 1160.970 52.460 ;
        RECT 133.470 17.580 133.790 17.640 ;
        RECT 137.610 17.580 137.930 17.640 ;
        RECT 133.470 17.440 137.930 17.580 ;
        RECT 133.470 17.380 133.790 17.440 ;
        RECT 137.610 17.380 137.930 17.440 ;
      LAYER via ;
        RECT 1160.220 1679.980 1160.480 1680.240 ;
        RECT 1163.440 1679.980 1163.700 1680.240 ;
        RECT 137.640 52.400 137.900 52.660 ;
        RECT 1160.680 52.400 1160.940 52.660 ;
        RECT 133.500 17.380 133.760 17.640 ;
        RECT 137.640 17.380 137.900 17.640 ;
      LAYER met2 ;
        RECT 1163.340 1700.340 1163.620 1704.000 ;
        RECT 1163.340 1700.000 1163.640 1700.340 ;
        RECT 1163.500 1680.270 1163.640 1700.000 ;
        RECT 1160.220 1679.950 1160.480 1680.270 ;
        RECT 1163.440 1679.950 1163.700 1680.270 ;
        RECT 1160.280 1669.810 1160.420 1679.950 ;
        RECT 1160.280 1669.670 1160.880 1669.810 ;
        RECT 1160.740 52.690 1160.880 1669.670 ;
        RECT 137.640 52.370 137.900 52.690 ;
        RECT 1160.680 52.370 1160.940 52.690 ;
        RECT 137.700 17.670 137.840 52.370 ;
        RECT 133.500 17.350 133.760 17.670 ;
        RECT 137.640 17.350 137.900 17.670 ;
        RECT 133.560 2.400 133.700 17.350 ;
        RECT 133.350 -4.800 133.910 2.400 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1161.110 1665.900 1161.430 1665.960 ;
        RECT 1165.250 1665.900 1165.570 1665.960 ;
        RECT 1161.110 1665.760 1165.570 1665.900 ;
        RECT 1161.110 1665.700 1161.430 1665.760 ;
        RECT 1165.250 1665.700 1165.570 1665.760 ;
        RECT 151.410 52.940 151.730 53.000 ;
        RECT 1161.110 52.940 1161.430 53.000 ;
        RECT 151.410 52.800 1161.430 52.940 ;
        RECT 151.410 52.740 151.730 52.800 ;
        RECT 1161.110 52.740 1161.430 52.800 ;
      LAYER via ;
        RECT 1161.140 1665.700 1161.400 1665.960 ;
        RECT 1165.280 1665.700 1165.540 1665.960 ;
        RECT 151.440 52.740 151.700 53.000 ;
        RECT 1161.140 52.740 1161.400 53.000 ;
      LAYER met2 ;
        RECT 1165.180 1700.340 1165.460 1704.000 ;
        RECT 1165.180 1700.000 1165.480 1700.340 ;
        RECT 1165.340 1665.990 1165.480 1700.000 ;
        RECT 1161.140 1665.670 1161.400 1665.990 ;
        RECT 1165.280 1665.670 1165.540 1665.990 ;
        RECT 1161.200 53.030 1161.340 1665.670 ;
        RECT 151.440 52.710 151.700 53.030 ;
        RECT 1161.140 52.710 1161.400 53.030 ;
        RECT 151.500 2.400 151.640 52.710 ;
        RECT 151.290 -4.800 151.850 2.400 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 172.110 1645.500 172.430 1645.560 ;
        RECT 1166.170 1645.500 1166.490 1645.560 ;
        RECT 172.110 1645.360 1166.490 1645.500 ;
        RECT 172.110 1645.300 172.430 1645.360 ;
        RECT 1166.170 1645.300 1166.490 1645.360 ;
        RECT 169.350 17.580 169.670 17.640 ;
        RECT 172.110 17.580 172.430 17.640 ;
        RECT 169.350 17.440 172.430 17.580 ;
        RECT 169.350 17.380 169.670 17.440 ;
        RECT 172.110 17.380 172.430 17.440 ;
      LAYER via ;
        RECT 172.140 1645.300 172.400 1645.560 ;
        RECT 1166.200 1645.300 1166.460 1645.560 ;
        RECT 169.380 17.380 169.640 17.640 ;
        RECT 172.140 17.380 172.400 17.640 ;
      LAYER met2 ;
        RECT 1167.020 1700.410 1167.300 1704.000 ;
        RECT 1166.720 1700.270 1167.300 1700.410 ;
        RECT 1166.720 1677.970 1166.860 1700.270 ;
        RECT 1167.020 1700.000 1167.300 1700.270 ;
        RECT 1166.260 1677.830 1166.860 1677.970 ;
        RECT 1166.260 1645.590 1166.400 1677.830 ;
        RECT 172.140 1645.270 172.400 1645.590 ;
        RECT 1166.200 1645.270 1166.460 1645.590 ;
        RECT 172.200 17.670 172.340 1645.270 ;
        RECT 169.380 17.350 169.640 17.670 ;
        RECT 172.140 17.350 172.400 17.670 ;
        RECT 169.440 2.400 169.580 17.350 ;
        RECT 169.230 -4.800 169.790 2.400 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1167.550 1679.160 1167.870 1679.220 ;
        RECT 1168.470 1679.160 1168.790 1679.220 ;
        RECT 1167.550 1679.020 1168.790 1679.160 ;
        RECT 1167.550 1678.960 1167.870 1679.020 ;
        RECT 1168.470 1678.960 1168.790 1679.020 ;
        RECT 192.810 1638.700 193.130 1638.760 ;
        RECT 1167.550 1638.700 1167.870 1638.760 ;
        RECT 192.810 1638.560 1167.870 1638.700 ;
        RECT 192.810 1638.500 193.130 1638.560 ;
        RECT 1167.550 1638.500 1167.870 1638.560 ;
        RECT 186.830 17.920 187.150 17.980 ;
        RECT 192.810 17.920 193.130 17.980 ;
        RECT 186.830 17.780 193.130 17.920 ;
        RECT 186.830 17.720 187.150 17.780 ;
        RECT 192.810 17.720 193.130 17.780 ;
      LAYER via ;
        RECT 1167.580 1678.960 1167.840 1679.220 ;
        RECT 1168.500 1678.960 1168.760 1679.220 ;
        RECT 192.840 1638.500 193.100 1638.760 ;
        RECT 1167.580 1638.500 1167.840 1638.760 ;
        RECT 186.860 17.720 187.120 17.980 ;
        RECT 192.840 17.720 193.100 17.980 ;
      LAYER met2 ;
        RECT 1168.860 1700.410 1169.140 1704.000 ;
        RECT 1168.560 1700.270 1169.140 1700.410 ;
        RECT 1168.560 1679.250 1168.700 1700.270 ;
        RECT 1168.860 1700.000 1169.140 1700.270 ;
        RECT 1167.580 1678.930 1167.840 1679.250 ;
        RECT 1168.500 1678.930 1168.760 1679.250 ;
        RECT 1167.640 1638.790 1167.780 1678.930 ;
        RECT 192.840 1638.470 193.100 1638.790 ;
        RECT 1167.580 1638.470 1167.840 1638.790 ;
        RECT 192.900 18.010 193.040 1638.470 ;
        RECT 186.860 17.690 187.120 18.010 ;
        RECT 192.840 17.690 193.100 18.010 ;
        RECT 186.920 2.400 187.060 17.690 ;
        RECT 186.710 -4.800 187.270 2.400 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1166.630 1677.460 1166.950 1677.520 ;
        RECT 1170.770 1677.460 1171.090 1677.520 ;
        RECT 1166.630 1677.320 1171.090 1677.460 ;
        RECT 1166.630 1677.260 1166.950 1677.320 ;
        RECT 1170.770 1677.260 1171.090 1677.320 ;
        RECT 210.290 1624.760 210.610 1624.820 ;
        RECT 1166.630 1624.760 1166.950 1624.820 ;
        RECT 210.290 1624.620 1166.950 1624.760 ;
        RECT 210.290 1624.560 210.610 1624.620 ;
        RECT 1166.630 1624.560 1166.950 1624.620 ;
        RECT 204.770 17.580 205.090 17.640 ;
        RECT 210.290 17.580 210.610 17.640 ;
        RECT 204.770 17.440 210.610 17.580 ;
        RECT 204.770 17.380 205.090 17.440 ;
        RECT 210.290 17.380 210.610 17.440 ;
      LAYER via ;
        RECT 1166.660 1677.260 1166.920 1677.520 ;
        RECT 1170.800 1677.260 1171.060 1677.520 ;
        RECT 210.320 1624.560 210.580 1624.820 ;
        RECT 1166.660 1624.560 1166.920 1624.820 ;
        RECT 204.800 17.380 205.060 17.640 ;
        RECT 210.320 17.380 210.580 17.640 ;
      LAYER met2 ;
        RECT 1170.700 1700.340 1170.980 1704.000 ;
        RECT 1170.700 1700.000 1171.000 1700.340 ;
        RECT 1170.860 1677.550 1171.000 1700.000 ;
        RECT 1166.660 1677.230 1166.920 1677.550 ;
        RECT 1170.800 1677.230 1171.060 1677.550 ;
        RECT 1166.720 1624.850 1166.860 1677.230 ;
        RECT 210.320 1624.530 210.580 1624.850 ;
        RECT 1166.660 1624.530 1166.920 1624.850 ;
        RECT 210.380 17.670 210.520 1624.530 ;
        RECT 204.800 17.350 205.060 17.670 ;
        RECT 210.320 17.350 210.580 17.670 ;
        RECT 204.860 2.400 205.000 17.350 ;
        RECT 204.650 -4.800 205.210 2.400 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 230.990 1617.960 231.310 1618.020 ;
        RECT 1172.610 1617.960 1172.930 1618.020 ;
        RECT 230.990 1617.820 1172.930 1617.960 ;
        RECT 230.990 1617.760 231.310 1617.820 ;
        RECT 1172.610 1617.760 1172.930 1617.820 ;
        RECT 222.710 18.600 223.030 18.660 ;
        RECT 230.990 18.600 231.310 18.660 ;
        RECT 222.710 18.460 231.310 18.600 ;
        RECT 222.710 18.400 223.030 18.460 ;
        RECT 230.990 18.400 231.310 18.460 ;
      LAYER via ;
        RECT 231.020 1617.760 231.280 1618.020 ;
        RECT 1172.640 1617.760 1172.900 1618.020 ;
        RECT 222.740 18.400 223.000 18.660 ;
        RECT 231.020 18.400 231.280 18.660 ;
      LAYER met2 ;
        RECT 1172.540 1700.340 1172.820 1704.000 ;
        RECT 1172.540 1700.000 1172.840 1700.340 ;
        RECT 1172.700 1618.050 1172.840 1700.000 ;
        RECT 231.020 1617.730 231.280 1618.050 ;
        RECT 1172.640 1617.730 1172.900 1618.050 ;
        RECT 231.080 18.690 231.220 1617.730 ;
        RECT 222.740 18.370 223.000 18.690 ;
        RECT 231.020 18.370 231.280 18.690 ;
        RECT 222.800 2.400 222.940 18.370 ;
        RECT 222.590 -4.800 223.150 2.400 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1147.845 1642.285 1148.015 1671.015 ;
        RECT 1147.385 1546.065 1147.555 1593.835 ;
        RECT 1147.385 1497.445 1147.555 1545.555 ;
        RECT 1147.845 1352.605 1148.015 1400.715 ;
        RECT 1147.845 1256.045 1148.015 1304.155 ;
        RECT 1147.845 386.665 1148.015 400.775 ;
        RECT 1147.845 338.045 1148.015 386.155 ;
        RECT 1147.845 241.485 1148.015 289.595 ;
        RECT 1147.845 144.925 1148.015 193.035 ;
      LAYER mcon ;
        RECT 1147.845 1670.845 1148.015 1671.015 ;
        RECT 1147.385 1593.665 1147.555 1593.835 ;
        RECT 1147.385 1545.385 1147.555 1545.555 ;
        RECT 1147.845 1400.545 1148.015 1400.715 ;
        RECT 1147.845 1303.985 1148.015 1304.155 ;
        RECT 1147.845 400.605 1148.015 400.775 ;
        RECT 1147.845 385.985 1148.015 386.155 ;
        RECT 1147.845 289.425 1148.015 289.595 ;
        RECT 1147.845 192.865 1148.015 193.035 ;
      LAYER met1 ;
        RECT 1147.785 1671.000 1148.075 1671.045 ;
        RECT 1151.450 1671.000 1151.770 1671.060 ;
        RECT 1147.785 1670.860 1151.770 1671.000 ;
        RECT 1147.785 1670.815 1148.075 1670.860 ;
        RECT 1151.450 1670.800 1151.770 1670.860 ;
        RECT 1147.770 1642.440 1148.090 1642.500 ;
        RECT 1147.575 1642.300 1148.090 1642.440 ;
        RECT 1147.770 1642.240 1148.090 1642.300 ;
        RECT 1147.325 1593.820 1147.615 1593.865 ;
        RECT 1147.770 1593.820 1148.090 1593.880 ;
        RECT 1147.325 1593.680 1148.090 1593.820 ;
        RECT 1147.325 1593.635 1147.615 1593.680 ;
        RECT 1147.770 1593.620 1148.090 1593.680 ;
        RECT 1147.310 1546.220 1147.630 1546.280 ;
        RECT 1147.115 1546.080 1147.630 1546.220 ;
        RECT 1147.310 1546.020 1147.630 1546.080 ;
        RECT 1147.310 1545.540 1147.630 1545.600 ;
        RECT 1147.115 1545.400 1147.630 1545.540 ;
        RECT 1147.310 1545.340 1147.630 1545.400 ;
        RECT 1147.325 1497.600 1147.615 1497.645 ;
        RECT 1147.770 1497.600 1148.090 1497.660 ;
        RECT 1147.325 1497.460 1148.090 1497.600 ;
        RECT 1147.325 1497.415 1147.615 1497.460 ;
        RECT 1147.770 1497.400 1148.090 1497.460 ;
        RECT 1147.770 1400.700 1148.090 1400.760 ;
        RECT 1147.575 1400.560 1148.090 1400.700 ;
        RECT 1147.770 1400.500 1148.090 1400.560 ;
        RECT 1147.785 1352.760 1148.075 1352.805 ;
        RECT 1148.230 1352.760 1148.550 1352.820 ;
        RECT 1147.785 1352.620 1148.550 1352.760 ;
        RECT 1147.785 1352.575 1148.075 1352.620 ;
        RECT 1148.230 1352.560 1148.550 1352.620 ;
        RECT 1147.770 1304.140 1148.090 1304.200 ;
        RECT 1147.575 1304.000 1148.090 1304.140 ;
        RECT 1147.770 1303.940 1148.090 1304.000 ;
        RECT 1147.785 1256.200 1148.075 1256.245 ;
        RECT 1148.230 1256.200 1148.550 1256.260 ;
        RECT 1147.785 1256.060 1148.550 1256.200 ;
        RECT 1147.785 1256.015 1148.075 1256.060 ;
        RECT 1148.230 1256.000 1148.550 1256.060 ;
        RECT 1148.230 1159.300 1148.550 1159.360 ;
        RECT 1149.150 1159.300 1149.470 1159.360 ;
        RECT 1148.230 1159.160 1149.470 1159.300 ;
        RECT 1148.230 1159.100 1148.550 1159.160 ;
        RECT 1149.150 1159.100 1149.470 1159.160 ;
        RECT 1148.230 1062.740 1148.550 1062.800 ;
        RECT 1149.150 1062.740 1149.470 1062.800 ;
        RECT 1148.230 1062.600 1149.470 1062.740 ;
        RECT 1148.230 1062.540 1148.550 1062.600 ;
        RECT 1149.150 1062.540 1149.470 1062.600 ;
        RECT 1148.230 966.180 1148.550 966.240 ;
        RECT 1149.150 966.180 1149.470 966.240 ;
        RECT 1148.230 966.040 1149.470 966.180 ;
        RECT 1148.230 965.980 1148.550 966.040 ;
        RECT 1149.150 965.980 1149.470 966.040 ;
        RECT 1148.230 869.620 1148.550 869.680 ;
        RECT 1149.150 869.620 1149.470 869.680 ;
        RECT 1148.230 869.480 1149.470 869.620 ;
        RECT 1148.230 869.420 1148.550 869.480 ;
        RECT 1149.150 869.420 1149.470 869.480 ;
        RECT 1147.770 821.000 1148.090 821.060 ;
        RECT 1149.150 821.000 1149.470 821.060 ;
        RECT 1147.770 820.860 1149.470 821.000 ;
        RECT 1147.770 820.800 1148.090 820.860 ;
        RECT 1149.150 820.800 1149.470 820.860 ;
        RECT 1147.770 689.900 1148.090 690.160 ;
        RECT 1147.310 689.760 1147.630 689.820 ;
        RECT 1147.860 689.760 1148.000 689.900 ;
        RECT 1147.310 689.620 1148.000 689.760 ;
        RECT 1147.310 689.560 1147.630 689.620 ;
        RECT 1147.770 593.340 1148.090 593.600 ;
        RECT 1147.310 593.200 1147.630 593.260 ;
        RECT 1147.860 593.200 1148.000 593.340 ;
        RECT 1147.310 593.060 1148.000 593.200 ;
        RECT 1147.310 593.000 1147.630 593.060 ;
        RECT 1147.770 496.780 1148.090 497.040 ;
        RECT 1147.310 496.640 1147.630 496.700 ;
        RECT 1147.860 496.640 1148.000 496.780 ;
        RECT 1147.310 496.500 1148.000 496.640 ;
        RECT 1147.310 496.440 1147.630 496.500 ;
        RECT 1147.770 400.760 1148.090 400.820 ;
        RECT 1147.575 400.620 1148.090 400.760 ;
        RECT 1147.770 400.560 1148.090 400.620 ;
        RECT 1147.310 386.820 1147.630 386.880 ;
        RECT 1147.785 386.820 1148.075 386.865 ;
        RECT 1147.310 386.680 1148.075 386.820 ;
        RECT 1147.310 386.620 1147.630 386.680 ;
        RECT 1147.785 386.635 1148.075 386.680 ;
        RECT 1147.770 386.140 1148.090 386.200 ;
        RECT 1147.575 386.000 1148.090 386.140 ;
        RECT 1147.770 385.940 1148.090 386.000 ;
        RECT 1147.785 338.200 1148.075 338.245 ;
        RECT 1148.230 338.200 1148.550 338.260 ;
        RECT 1147.785 338.060 1148.550 338.200 ;
        RECT 1147.785 338.015 1148.075 338.060 ;
        RECT 1148.230 338.000 1148.550 338.060 ;
        RECT 1147.785 289.580 1148.075 289.625 ;
        RECT 1148.230 289.580 1148.550 289.640 ;
        RECT 1147.785 289.440 1148.550 289.580 ;
        RECT 1147.785 289.395 1148.075 289.440 ;
        RECT 1148.230 289.380 1148.550 289.440 ;
        RECT 1147.770 241.640 1148.090 241.700 ;
        RECT 1147.575 241.500 1148.090 241.640 ;
        RECT 1147.770 241.440 1148.090 241.500 ;
        RECT 1147.310 206.960 1147.630 207.020 ;
        RECT 1148.230 206.960 1148.550 207.020 ;
        RECT 1147.310 206.820 1148.550 206.960 ;
        RECT 1147.310 206.760 1147.630 206.820 ;
        RECT 1148.230 206.760 1148.550 206.820 ;
        RECT 1147.785 193.020 1148.075 193.065 ;
        RECT 1148.230 193.020 1148.550 193.080 ;
        RECT 1147.785 192.880 1148.550 193.020 ;
        RECT 1147.785 192.835 1148.075 192.880 ;
        RECT 1148.230 192.820 1148.550 192.880 ;
        RECT 1147.770 145.080 1148.090 145.140 ;
        RECT 1147.575 144.940 1148.090 145.080 ;
        RECT 1147.770 144.880 1148.090 144.940 ;
        RECT 1147.770 110.540 1148.090 110.800 ;
        RECT 1147.860 110.120 1148.000 110.540 ;
        RECT 1147.770 109.860 1148.090 110.120 ;
        RECT 19.850 51.580 20.170 51.640 ;
        RECT 1147.770 51.580 1148.090 51.640 ;
        RECT 19.850 51.440 1148.090 51.580 ;
        RECT 19.850 51.380 20.170 51.440 ;
        RECT 1147.770 51.380 1148.090 51.440 ;
      LAYER via ;
        RECT 1151.480 1670.800 1151.740 1671.060 ;
        RECT 1147.800 1642.240 1148.060 1642.500 ;
        RECT 1147.800 1593.620 1148.060 1593.880 ;
        RECT 1147.340 1546.020 1147.600 1546.280 ;
        RECT 1147.340 1545.340 1147.600 1545.600 ;
        RECT 1147.800 1497.400 1148.060 1497.660 ;
        RECT 1147.800 1400.500 1148.060 1400.760 ;
        RECT 1148.260 1352.560 1148.520 1352.820 ;
        RECT 1147.800 1303.940 1148.060 1304.200 ;
        RECT 1148.260 1256.000 1148.520 1256.260 ;
        RECT 1148.260 1159.100 1148.520 1159.360 ;
        RECT 1149.180 1159.100 1149.440 1159.360 ;
        RECT 1148.260 1062.540 1148.520 1062.800 ;
        RECT 1149.180 1062.540 1149.440 1062.800 ;
        RECT 1148.260 965.980 1148.520 966.240 ;
        RECT 1149.180 965.980 1149.440 966.240 ;
        RECT 1148.260 869.420 1148.520 869.680 ;
        RECT 1149.180 869.420 1149.440 869.680 ;
        RECT 1147.800 820.800 1148.060 821.060 ;
        RECT 1149.180 820.800 1149.440 821.060 ;
        RECT 1147.800 689.900 1148.060 690.160 ;
        RECT 1147.340 689.560 1147.600 689.820 ;
        RECT 1147.800 593.340 1148.060 593.600 ;
        RECT 1147.340 593.000 1147.600 593.260 ;
        RECT 1147.800 496.780 1148.060 497.040 ;
        RECT 1147.340 496.440 1147.600 496.700 ;
        RECT 1147.800 400.560 1148.060 400.820 ;
        RECT 1147.340 386.620 1147.600 386.880 ;
        RECT 1147.800 385.940 1148.060 386.200 ;
        RECT 1148.260 338.000 1148.520 338.260 ;
        RECT 1148.260 289.380 1148.520 289.640 ;
        RECT 1147.800 241.440 1148.060 241.700 ;
        RECT 1147.340 206.760 1147.600 207.020 ;
        RECT 1148.260 206.760 1148.520 207.020 ;
        RECT 1148.260 192.820 1148.520 193.080 ;
        RECT 1147.800 144.880 1148.060 145.140 ;
        RECT 1147.800 110.540 1148.060 110.800 ;
        RECT 1147.800 109.860 1148.060 110.120 ;
        RECT 19.880 51.380 20.140 51.640 ;
        RECT 1147.800 51.380 1148.060 51.640 ;
      LAYER met2 ;
        RECT 1151.380 1700.340 1151.660 1704.000 ;
        RECT 1151.380 1700.000 1151.680 1700.340 ;
        RECT 1151.540 1671.090 1151.680 1700.000 ;
        RECT 1151.480 1670.770 1151.740 1671.090 ;
        RECT 1147.800 1642.210 1148.060 1642.530 ;
        RECT 1147.860 1593.910 1148.000 1642.210 ;
        RECT 1147.800 1593.590 1148.060 1593.910 ;
        RECT 1147.340 1545.990 1147.600 1546.310 ;
        RECT 1147.400 1545.630 1147.540 1545.990 ;
        RECT 1147.340 1545.310 1147.600 1545.630 ;
        RECT 1147.800 1497.370 1148.060 1497.690 ;
        RECT 1147.860 1472.610 1148.000 1497.370 ;
        RECT 1147.860 1472.470 1148.460 1472.610 ;
        RECT 1148.320 1414.130 1148.460 1472.470 ;
        RECT 1147.860 1413.990 1148.460 1414.130 ;
        RECT 1147.860 1400.790 1148.000 1413.990 ;
        RECT 1147.800 1400.470 1148.060 1400.790 ;
        RECT 1148.260 1352.530 1148.520 1352.850 ;
        RECT 1148.320 1317.570 1148.460 1352.530 ;
        RECT 1147.860 1317.430 1148.460 1317.570 ;
        RECT 1147.860 1304.230 1148.000 1317.430 ;
        RECT 1147.800 1303.910 1148.060 1304.230 ;
        RECT 1148.260 1255.970 1148.520 1256.290 ;
        RECT 1148.320 1221.010 1148.460 1255.970 ;
        RECT 1147.860 1220.870 1148.460 1221.010 ;
        RECT 1147.860 1207.525 1148.000 1220.870 ;
        RECT 1147.790 1207.155 1148.070 1207.525 ;
        RECT 1149.170 1207.155 1149.450 1207.525 ;
        RECT 1149.240 1159.390 1149.380 1207.155 ;
        RECT 1148.260 1159.070 1148.520 1159.390 ;
        RECT 1149.180 1159.070 1149.440 1159.390 ;
        RECT 1148.320 1124.450 1148.460 1159.070 ;
        RECT 1147.860 1124.310 1148.460 1124.450 ;
        RECT 1147.860 1110.965 1148.000 1124.310 ;
        RECT 1147.790 1110.595 1148.070 1110.965 ;
        RECT 1149.170 1110.595 1149.450 1110.965 ;
        RECT 1149.240 1062.830 1149.380 1110.595 ;
        RECT 1148.260 1062.510 1148.520 1062.830 ;
        RECT 1149.180 1062.510 1149.440 1062.830 ;
        RECT 1148.320 1027.890 1148.460 1062.510 ;
        RECT 1147.860 1027.750 1148.460 1027.890 ;
        RECT 1147.860 1014.405 1148.000 1027.750 ;
        RECT 1147.790 1014.035 1148.070 1014.405 ;
        RECT 1149.170 1014.035 1149.450 1014.405 ;
        RECT 1149.240 966.270 1149.380 1014.035 ;
        RECT 1148.260 965.950 1148.520 966.270 ;
        RECT 1149.180 965.950 1149.440 966.270 ;
        RECT 1148.320 931.330 1148.460 965.950 ;
        RECT 1147.860 931.190 1148.460 931.330 ;
        RECT 1147.860 917.845 1148.000 931.190 ;
        RECT 1147.790 917.475 1148.070 917.845 ;
        RECT 1149.170 917.475 1149.450 917.845 ;
        RECT 1149.240 869.710 1149.380 917.475 ;
        RECT 1148.260 869.390 1148.520 869.710 ;
        RECT 1149.180 869.390 1149.440 869.710 ;
        RECT 1148.320 834.770 1148.460 869.390 ;
        RECT 1147.860 834.630 1148.460 834.770 ;
        RECT 1147.860 821.090 1148.000 834.630 ;
        RECT 1147.800 820.770 1148.060 821.090 ;
        RECT 1149.180 820.770 1149.440 821.090 ;
        RECT 1149.240 773.005 1149.380 820.770 ;
        RECT 1148.250 772.635 1148.530 773.005 ;
        RECT 1149.170 772.635 1149.450 773.005 ;
        RECT 1148.320 738.210 1148.460 772.635 ;
        RECT 1147.860 738.070 1148.460 738.210 ;
        RECT 1147.860 690.190 1148.000 738.070 ;
        RECT 1147.800 689.870 1148.060 690.190 ;
        RECT 1147.340 689.530 1147.600 689.850 ;
        RECT 1147.400 676.445 1147.540 689.530 ;
        RECT 1147.330 676.075 1147.610 676.445 ;
        RECT 1148.250 676.075 1148.530 676.445 ;
        RECT 1148.320 641.650 1148.460 676.075 ;
        RECT 1147.860 641.510 1148.460 641.650 ;
        RECT 1147.860 593.630 1148.000 641.510 ;
        RECT 1147.800 593.310 1148.060 593.630 ;
        RECT 1147.340 592.970 1147.600 593.290 ;
        RECT 1147.400 579.885 1147.540 592.970 ;
        RECT 1147.330 579.515 1147.610 579.885 ;
        RECT 1148.250 579.515 1148.530 579.885 ;
        RECT 1148.320 545.090 1148.460 579.515 ;
        RECT 1147.860 544.950 1148.460 545.090 ;
        RECT 1147.860 497.070 1148.000 544.950 ;
        RECT 1147.800 496.750 1148.060 497.070 ;
        RECT 1147.340 496.410 1147.600 496.730 ;
        RECT 1147.400 483.325 1147.540 496.410 ;
        RECT 1147.330 482.955 1147.610 483.325 ;
        RECT 1148.250 482.955 1148.530 483.325 ;
        RECT 1148.320 448.530 1148.460 482.955 ;
        RECT 1147.860 448.390 1148.460 448.530 ;
        RECT 1147.860 400.850 1148.000 448.390 ;
        RECT 1147.800 400.530 1148.060 400.850 ;
        RECT 1147.340 386.650 1147.600 386.910 ;
        RECT 1147.340 386.590 1148.000 386.650 ;
        RECT 1147.400 386.510 1148.000 386.590 ;
        RECT 1147.860 386.230 1148.000 386.510 ;
        RECT 1147.800 385.910 1148.060 386.230 ;
        RECT 1148.260 337.970 1148.520 338.290 ;
        RECT 1148.320 337.805 1148.460 337.970 ;
        RECT 1148.250 337.435 1148.530 337.805 ;
        RECT 1148.250 289.835 1148.530 290.205 ;
        RECT 1148.320 289.670 1148.460 289.835 ;
        RECT 1148.260 289.350 1148.520 289.670 ;
        RECT 1147.800 241.410 1148.060 241.730 ;
        RECT 1147.860 207.130 1148.000 241.410 ;
        RECT 1147.400 207.050 1148.000 207.130 ;
        RECT 1147.340 206.990 1148.000 207.050 ;
        RECT 1147.340 206.730 1147.600 206.990 ;
        RECT 1148.260 206.730 1148.520 207.050 ;
        RECT 1148.320 193.110 1148.460 206.730 ;
        RECT 1148.260 192.790 1148.520 193.110 ;
        RECT 1147.800 144.850 1148.060 145.170 ;
        RECT 1147.860 110.830 1148.000 144.850 ;
        RECT 1147.800 110.510 1148.060 110.830 ;
        RECT 1147.800 109.830 1148.060 110.150 ;
        RECT 1147.860 51.670 1148.000 109.830 ;
        RECT 19.880 51.350 20.140 51.670 ;
        RECT 1147.800 51.350 1148.060 51.670 ;
        RECT 19.940 3.130 20.080 51.350 ;
        RECT 19.940 2.990 20.540 3.130 ;
        RECT 20.400 2.400 20.540 2.990 ;
        RECT 20.190 -4.800 20.750 2.400 ;
      LAYER via2 ;
        RECT 1147.790 1207.200 1148.070 1207.480 ;
        RECT 1149.170 1207.200 1149.450 1207.480 ;
        RECT 1147.790 1110.640 1148.070 1110.920 ;
        RECT 1149.170 1110.640 1149.450 1110.920 ;
        RECT 1147.790 1014.080 1148.070 1014.360 ;
        RECT 1149.170 1014.080 1149.450 1014.360 ;
        RECT 1147.790 917.520 1148.070 917.800 ;
        RECT 1149.170 917.520 1149.450 917.800 ;
        RECT 1148.250 772.680 1148.530 772.960 ;
        RECT 1149.170 772.680 1149.450 772.960 ;
        RECT 1147.330 676.120 1147.610 676.400 ;
        RECT 1148.250 676.120 1148.530 676.400 ;
        RECT 1147.330 579.560 1147.610 579.840 ;
        RECT 1148.250 579.560 1148.530 579.840 ;
        RECT 1147.330 483.000 1147.610 483.280 ;
        RECT 1148.250 483.000 1148.530 483.280 ;
        RECT 1148.250 337.480 1148.530 337.760 ;
        RECT 1148.250 289.880 1148.530 290.160 ;
      LAYER met3 ;
        RECT 1147.765 1207.490 1148.095 1207.505 ;
        RECT 1149.145 1207.490 1149.475 1207.505 ;
        RECT 1147.765 1207.190 1149.475 1207.490 ;
        RECT 1147.765 1207.175 1148.095 1207.190 ;
        RECT 1149.145 1207.175 1149.475 1207.190 ;
        RECT 1147.765 1110.930 1148.095 1110.945 ;
        RECT 1149.145 1110.930 1149.475 1110.945 ;
        RECT 1147.765 1110.630 1149.475 1110.930 ;
        RECT 1147.765 1110.615 1148.095 1110.630 ;
        RECT 1149.145 1110.615 1149.475 1110.630 ;
        RECT 1147.765 1014.370 1148.095 1014.385 ;
        RECT 1149.145 1014.370 1149.475 1014.385 ;
        RECT 1147.765 1014.070 1149.475 1014.370 ;
        RECT 1147.765 1014.055 1148.095 1014.070 ;
        RECT 1149.145 1014.055 1149.475 1014.070 ;
        RECT 1147.765 917.810 1148.095 917.825 ;
        RECT 1149.145 917.810 1149.475 917.825 ;
        RECT 1147.765 917.510 1149.475 917.810 ;
        RECT 1147.765 917.495 1148.095 917.510 ;
        RECT 1149.145 917.495 1149.475 917.510 ;
        RECT 1148.225 772.970 1148.555 772.985 ;
        RECT 1149.145 772.970 1149.475 772.985 ;
        RECT 1148.225 772.670 1149.475 772.970 ;
        RECT 1148.225 772.655 1148.555 772.670 ;
        RECT 1149.145 772.655 1149.475 772.670 ;
        RECT 1147.305 676.410 1147.635 676.425 ;
        RECT 1148.225 676.410 1148.555 676.425 ;
        RECT 1147.305 676.110 1148.555 676.410 ;
        RECT 1147.305 676.095 1147.635 676.110 ;
        RECT 1148.225 676.095 1148.555 676.110 ;
        RECT 1147.305 579.850 1147.635 579.865 ;
        RECT 1148.225 579.850 1148.555 579.865 ;
        RECT 1147.305 579.550 1148.555 579.850 ;
        RECT 1147.305 579.535 1147.635 579.550 ;
        RECT 1148.225 579.535 1148.555 579.550 ;
        RECT 1147.305 483.290 1147.635 483.305 ;
        RECT 1148.225 483.290 1148.555 483.305 ;
        RECT 1147.305 482.990 1148.555 483.290 ;
        RECT 1147.305 482.975 1147.635 482.990 ;
        RECT 1148.225 482.975 1148.555 482.990 ;
        RECT 1147.510 337.770 1147.890 337.780 ;
        RECT 1148.225 337.770 1148.555 337.785 ;
        RECT 1147.510 337.470 1148.555 337.770 ;
        RECT 1147.510 337.460 1147.890 337.470 ;
        RECT 1148.225 337.455 1148.555 337.470 ;
        RECT 1148.225 290.180 1148.555 290.185 ;
        RECT 1148.225 290.170 1148.810 290.180 ;
        RECT 1148.225 289.870 1149.010 290.170 ;
        RECT 1148.225 289.860 1148.810 289.870 ;
        RECT 1148.225 289.855 1148.555 289.860 ;
      LAYER via3 ;
        RECT 1147.540 337.460 1147.860 337.780 ;
        RECT 1148.460 289.860 1148.780 290.180 ;
      LAYER met4 ;
        RECT 1147.535 337.455 1147.865 337.785 ;
        RECT 1147.550 290.850 1147.850 337.455 ;
        RECT 1147.550 290.550 1148.770 290.850 ;
        RECT 1148.470 290.185 1148.770 290.550 ;
        RECT 1148.455 289.855 1148.785 290.185 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 47.910 51.920 48.230 51.980 ;
        RECT 1154.670 51.920 1154.990 51.980 ;
        RECT 47.910 51.780 1154.990 51.920 ;
        RECT 47.910 51.720 48.230 51.780 ;
        RECT 1154.670 51.720 1154.990 51.780 ;
        RECT 44.230 17.580 44.550 17.640 ;
        RECT 47.910 17.580 48.230 17.640 ;
        RECT 44.230 17.440 48.230 17.580 ;
        RECT 44.230 17.380 44.550 17.440 ;
        RECT 47.910 17.380 48.230 17.440 ;
      LAYER via ;
        RECT 47.940 51.720 48.200 51.980 ;
        RECT 1154.700 51.720 1154.960 51.980 ;
        RECT 44.260 17.380 44.520 17.640 ;
        RECT 47.940 17.380 48.200 17.640 ;
      LAYER met2 ;
        RECT 1154.140 1700.340 1154.420 1704.000 ;
        RECT 1154.140 1700.000 1154.440 1700.340 ;
        RECT 1154.300 1666.410 1154.440 1700.000 ;
        RECT 1154.300 1666.270 1154.900 1666.410 ;
        RECT 1154.760 52.010 1154.900 1666.270 ;
        RECT 47.940 51.690 48.200 52.010 ;
        RECT 1154.700 51.690 1154.960 52.010 ;
        RECT 48.000 17.670 48.140 51.690 ;
        RECT 44.260 17.350 44.520 17.670 ;
        RECT 47.940 17.350 48.200 17.670 ;
        RECT 44.320 2.400 44.460 17.350 ;
        RECT 44.110 -4.800 44.670 2.400 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 248.010 1666.240 248.330 1666.300 ;
        RECT 1174.910 1666.240 1175.230 1666.300 ;
        RECT 248.010 1666.100 1175.230 1666.240 ;
        RECT 248.010 1666.040 248.330 1666.100 ;
        RECT 1174.910 1666.040 1175.230 1666.100 ;
      LAYER via ;
        RECT 248.040 1666.040 248.300 1666.300 ;
        RECT 1174.940 1666.040 1175.200 1666.300 ;
      LAYER met2 ;
        RECT 1174.840 1700.340 1175.120 1704.000 ;
        RECT 1174.840 1700.000 1175.140 1700.340 ;
        RECT 1175.000 1666.330 1175.140 1700.000 ;
        RECT 248.040 1666.010 248.300 1666.330 ;
        RECT 1174.940 1666.010 1175.200 1666.330 ;
        RECT 248.100 17.410 248.240 1666.010 ;
        RECT 246.720 17.270 248.240 17.410 ;
        RECT 246.720 2.400 246.860 17.270 ;
        RECT 246.510 -4.800 247.070 2.400 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 268.710 1631.900 269.030 1631.960 ;
        RECT 1176.750 1631.900 1177.070 1631.960 ;
        RECT 268.710 1631.760 1177.070 1631.900 ;
        RECT 268.710 1631.700 269.030 1631.760 ;
        RECT 1176.750 1631.700 1177.070 1631.760 ;
        RECT 264.110 17.920 264.430 17.980 ;
        RECT 268.710 17.920 269.030 17.980 ;
        RECT 264.110 17.780 269.030 17.920 ;
        RECT 264.110 17.720 264.430 17.780 ;
        RECT 268.710 17.720 269.030 17.780 ;
      LAYER via ;
        RECT 268.740 1631.700 269.000 1631.960 ;
        RECT 1176.780 1631.700 1177.040 1631.960 ;
        RECT 264.140 17.720 264.400 17.980 ;
        RECT 268.740 17.720 269.000 17.980 ;
      LAYER met2 ;
        RECT 1176.680 1700.340 1176.960 1704.000 ;
        RECT 1176.680 1700.000 1176.980 1700.340 ;
        RECT 1176.840 1631.990 1176.980 1700.000 ;
        RECT 268.740 1631.670 269.000 1631.990 ;
        RECT 1176.780 1631.670 1177.040 1631.990 ;
        RECT 268.800 18.010 268.940 1631.670 ;
        RECT 264.140 17.690 264.400 18.010 ;
        RECT 268.740 17.690 269.000 18.010 ;
        RECT 264.200 2.400 264.340 17.690 ;
        RECT 263.990 -4.800 264.550 2.400 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 282.050 1611.160 282.370 1611.220 ;
        RECT 1178.130 1611.160 1178.450 1611.220 ;
        RECT 282.050 1611.020 1178.450 1611.160 ;
        RECT 282.050 1610.960 282.370 1611.020 ;
        RECT 1178.130 1610.960 1178.450 1611.020 ;
      LAYER via ;
        RECT 282.080 1610.960 282.340 1611.220 ;
        RECT 1178.160 1610.960 1178.420 1611.220 ;
      LAYER met2 ;
        RECT 1178.520 1700.340 1178.800 1704.000 ;
        RECT 1178.520 1700.000 1178.820 1700.340 ;
        RECT 1178.680 1666.410 1178.820 1700.000 ;
        RECT 1178.220 1666.270 1178.820 1666.410 ;
        RECT 1178.220 1611.250 1178.360 1666.270 ;
        RECT 282.080 1610.930 282.340 1611.250 ;
        RECT 1178.160 1610.930 1178.420 1611.250 ;
        RECT 282.140 2.400 282.280 1610.930 ;
        RECT 281.930 -4.800 282.490 2.400 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1180.430 1678.140 1180.750 1678.200 ;
        RECT 1184.110 1678.140 1184.430 1678.200 ;
        RECT 1180.430 1678.000 1184.430 1678.140 ;
        RECT 1180.430 1677.940 1180.750 1678.000 ;
        RECT 1184.110 1677.940 1184.430 1678.000 ;
        RECT 303.210 53.280 303.530 53.340 ;
        RECT 1184.110 53.280 1184.430 53.340 ;
        RECT 303.210 53.140 1184.430 53.280 ;
        RECT 303.210 53.080 303.530 53.140 ;
        RECT 1184.110 53.080 1184.430 53.140 ;
        RECT 299.990 16.900 300.310 16.960 ;
        RECT 303.210 16.900 303.530 16.960 ;
        RECT 299.990 16.760 303.530 16.900 ;
        RECT 299.990 16.700 300.310 16.760 ;
        RECT 303.210 16.700 303.530 16.760 ;
      LAYER via ;
        RECT 1180.460 1677.940 1180.720 1678.200 ;
        RECT 1184.140 1677.940 1184.400 1678.200 ;
        RECT 303.240 53.080 303.500 53.340 ;
        RECT 1184.140 53.080 1184.400 53.340 ;
        RECT 300.020 16.700 300.280 16.960 ;
        RECT 303.240 16.700 303.500 16.960 ;
      LAYER met2 ;
        RECT 1180.360 1700.340 1180.640 1704.000 ;
        RECT 1180.360 1700.000 1180.660 1700.340 ;
        RECT 1180.520 1678.230 1180.660 1700.000 ;
        RECT 1180.460 1677.910 1180.720 1678.230 ;
        RECT 1184.140 1677.910 1184.400 1678.230 ;
        RECT 1184.200 53.370 1184.340 1677.910 ;
        RECT 303.240 53.050 303.500 53.370 ;
        RECT 1184.140 53.050 1184.400 53.370 ;
        RECT 303.300 16.990 303.440 53.050 ;
        RECT 300.020 16.670 300.280 16.990 ;
        RECT 303.240 16.670 303.500 16.990 ;
        RECT 300.080 2.400 300.220 16.670 ;
        RECT 299.870 -4.800 300.430 2.400 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1182.270 1678.820 1182.590 1678.880 ;
        RECT 1183.650 1678.820 1183.970 1678.880 ;
        RECT 1182.270 1678.680 1183.970 1678.820 ;
        RECT 1182.270 1678.620 1182.590 1678.680 ;
        RECT 1183.650 1678.620 1183.970 1678.680 ;
        RECT 323.910 53.620 324.230 53.680 ;
        RECT 1183.650 53.620 1183.970 53.680 ;
        RECT 323.910 53.480 1183.970 53.620 ;
        RECT 323.910 53.420 324.230 53.480 ;
        RECT 1183.650 53.420 1183.970 53.480 ;
        RECT 317.930 16.900 318.250 16.960 ;
        RECT 323.910 16.900 324.230 16.960 ;
        RECT 317.930 16.760 324.230 16.900 ;
        RECT 317.930 16.700 318.250 16.760 ;
        RECT 323.910 16.700 324.230 16.760 ;
      LAYER via ;
        RECT 1182.300 1678.620 1182.560 1678.880 ;
        RECT 1183.680 1678.620 1183.940 1678.880 ;
        RECT 323.940 53.420 324.200 53.680 ;
        RECT 1183.680 53.420 1183.940 53.680 ;
        RECT 317.960 16.700 318.220 16.960 ;
        RECT 323.940 16.700 324.200 16.960 ;
      LAYER met2 ;
        RECT 1182.200 1700.340 1182.480 1704.000 ;
        RECT 1182.200 1700.000 1182.500 1700.340 ;
        RECT 1182.360 1678.910 1182.500 1700.000 ;
        RECT 1182.300 1678.590 1182.560 1678.910 ;
        RECT 1183.680 1678.590 1183.940 1678.910 ;
        RECT 1183.740 53.710 1183.880 1678.590 ;
        RECT 323.940 53.390 324.200 53.710 ;
        RECT 1183.680 53.390 1183.940 53.710 ;
        RECT 324.000 16.990 324.140 53.390 ;
        RECT 317.960 16.670 318.220 16.990 ;
        RECT 323.940 16.670 324.200 16.990 ;
        RECT 318.020 2.400 318.160 16.670 ;
        RECT 317.810 -4.800 318.370 2.400 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1151.910 1684.940 1152.230 1685.000 ;
        RECT 1184.110 1684.940 1184.430 1685.000 ;
        RECT 1151.910 1684.800 1184.430 1684.940 ;
        RECT 1151.910 1684.740 1152.230 1684.800 ;
        RECT 1184.110 1684.740 1184.430 1684.800 ;
        RECT 337.710 1597.560 338.030 1597.620 ;
        RECT 1148.690 1597.560 1149.010 1597.620 ;
        RECT 337.710 1597.420 1149.010 1597.560 ;
        RECT 337.710 1597.360 338.030 1597.420 ;
        RECT 1148.690 1597.360 1149.010 1597.420 ;
      LAYER via ;
        RECT 1151.940 1684.740 1152.200 1685.000 ;
        RECT 1184.140 1684.740 1184.400 1685.000 ;
        RECT 337.740 1597.360 338.000 1597.620 ;
        RECT 1148.720 1597.360 1148.980 1597.620 ;
      LAYER met2 ;
        RECT 1184.040 1700.340 1184.320 1704.000 ;
        RECT 1184.040 1700.000 1184.340 1700.340 ;
        RECT 1184.200 1685.030 1184.340 1700.000 ;
        RECT 1151.940 1684.710 1152.200 1685.030 ;
        RECT 1184.140 1684.710 1184.400 1685.030 ;
        RECT 1152.000 1670.490 1152.140 1684.710 ;
        RECT 1148.780 1670.350 1152.140 1670.490 ;
        RECT 1148.780 1597.650 1148.920 1670.350 ;
        RECT 337.740 1597.330 338.000 1597.650 ;
        RECT 1148.720 1597.330 1148.980 1597.650 ;
        RECT 337.800 3.130 337.940 1597.330 ;
        RECT 335.960 2.990 337.940 3.130 ;
        RECT 335.960 2.400 336.100 2.990 ;
        RECT 335.750 -4.800 336.310 2.400 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 358.410 1652.640 358.730 1652.700 ;
        RECT 1185.950 1652.640 1186.270 1652.700 ;
        RECT 358.410 1652.500 1186.270 1652.640 ;
        RECT 358.410 1652.440 358.730 1652.500 ;
        RECT 1185.950 1652.440 1186.270 1652.500 ;
        RECT 353.350 16.900 353.670 16.960 ;
        RECT 358.410 16.900 358.730 16.960 ;
        RECT 353.350 16.760 358.730 16.900 ;
        RECT 353.350 16.700 353.670 16.760 ;
        RECT 358.410 16.700 358.730 16.760 ;
      LAYER via ;
        RECT 358.440 1652.440 358.700 1652.700 ;
        RECT 1185.980 1652.440 1186.240 1652.700 ;
        RECT 353.380 16.700 353.640 16.960 ;
        RECT 358.440 16.700 358.700 16.960 ;
      LAYER met2 ;
        RECT 1185.880 1700.340 1186.160 1704.000 ;
        RECT 1185.880 1700.000 1186.180 1700.340 ;
        RECT 1186.040 1652.730 1186.180 1700.000 ;
        RECT 358.440 1652.410 358.700 1652.730 ;
        RECT 1185.980 1652.410 1186.240 1652.730 ;
        RECT 358.500 16.990 358.640 1652.410 ;
        RECT 353.380 16.670 353.640 16.990 ;
        RECT 358.440 16.670 358.700 16.990 ;
        RECT 353.440 2.400 353.580 16.670 ;
        RECT 353.230 -4.800 353.790 2.400 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1169.390 1665.900 1169.710 1665.960 ;
        RECT 1187.790 1665.900 1188.110 1665.960 ;
        RECT 1169.390 1665.760 1188.110 1665.900 ;
        RECT 1169.390 1665.700 1169.710 1665.760 ;
        RECT 1187.790 1665.700 1188.110 1665.760 ;
        RECT 372.210 1604.360 372.530 1604.420 ;
        RECT 1169.390 1604.360 1169.710 1604.420 ;
        RECT 372.210 1604.220 1169.710 1604.360 ;
        RECT 372.210 1604.160 372.530 1604.220 ;
        RECT 1169.390 1604.160 1169.710 1604.220 ;
        RECT 371.290 2.960 371.610 3.020 ;
        RECT 372.210 2.960 372.530 3.020 ;
        RECT 371.290 2.820 372.530 2.960 ;
        RECT 371.290 2.760 371.610 2.820 ;
        RECT 372.210 2.760 372.530 2.820 ;
      LAYER via ;
        RECT 1169.420 1665.700 1169.680 1665.960 ;
        RECT 1187.820 1665.700 1188.080 1665.960 ;
        RECT 372.240 1604.160 372.500 1604.420 ;
        RECT 1169.420 1604.160 1169.680 1604.420 ;
        RECT 371.320 2.760 371.580 3.020 ;
        RECT 372.240 2.760 372.500 3.020 ;
      LAYER met2 ;
        RECT 1187.720 1700.340 1188.000 1704.000 ;
        RECT 1187.720 1700.000 1188.020 1700.340 ;
        RECT 1187.880 1665.990 1188.020 1700.000 ;
        RECT 1169.420 1665.670 1169.680 1665.990 ;
        RECT 1187.820 1665.670 1188.080 1665.990 ;
        RECT 1169.480 1604.450 1169.620 1665.670 ;
        RECT 372.240 1604.130 372.500 1604.450 ;
        RECT 1169.420 1604.130 1169.680 1604.450 ;
        RECT 372.300 3.050 372.440 1604.130 ;
        RECT 371.320 2.730 371.580 3.050 ;
        RECT 372.240 2.730 372.500 3.050 ;
        RECT 371.380 2.400 371.520 2.730 ;
        RECT 371.170 -4.800 371.730 2.400 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 392.910 1645.840 393.230 1645.900 ;
        RECT 1189.630 1645.840 1189.950 1645.900 ;
        RECT 392.910 1645.700 1189.950 1645.840 ;
        RECT 392.910 1645.640 393.230 1645.700 ;
        RECT 1189.630 1645.640 1189.950 1645.700 ;
        RECT 389.230 16.900 389.550 16.960 ;
        RECT 392.910 16.900 393.230 16.960 ;
        RECT 389.230 16.760 393.230 16.900 ;
        RECT 389.230 16.700 389.550 16.760 ;
        RECT 392.910 16.700 393.230 16.760 ;
      LAYER via ;
        RECT 392.940 1645.640 393.200 1645.900 ;
        RECT 1189.660 1645.640 1189.920 1645.900 ;
        RECT 389.260 16.700 389.520 16.960 ;
        RECT 392.940 16.700 393.200 16.960 ;
      LAYER met2 ;
        RECT 1189.560 1700.340 1189.840 1704.000 ;
        RECT 1189.560 1700.000 1189.860 1700.340 ;
        RECT 1189.720 1645.930 1189.860 1700.000 ;
        RECT 392.940 1645.610 393.200 1645.930 ;
        RECT 1189.660 1645.610 1189.920 1645.930 ;
        RECT 393.000 16.990 393.140 1645.610 ;
        RECT 389.260 16.670 389.520 16.990 ;
        RECT 392.940 16.670 393.200 16.990 ;
        RECT 389.320 2.400 389.460 16.670 ;
        RECT 389.110 -4.800 389.670 2.400 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 413.610 1639.040 413.930 1639.100 ;
        RECT 1191.470 1639.040 1191.790 1639.100 ;
        RECT 413.610 1638.900 1191.790 1639.040 ;
        RECT 413.610 1638.840 413.930 1638.900 ;
        RECT 1191.470 1638.840 1191.790 1638.900 ;
        RECT 407.170 16.900 407.490 16.960 ;
        RECT 413.610 16.900 413.930 16.960 ;
        RECT 407.170 16.760 413.930 16.900 ;
        RECT 407.170 16.700 407.490 16.760 ;
        RECT 413.610 16.700 413.930 16.760 ;
      LAYER via ;
        RECT 413.640 1638.840 413.900 1639.100 ;
        RECT 1191.500 1638.840 1191.760 1639.100 ;
        RECT 407.200 16.700 407.460 16.960 ;
        RECT 413.640 16.700 413.900 16.960 ;
      LAYER met2 ;
        RECT 1191.400 1700.340 1191.680 1704.000 ;
        RECT 1191.400 1700.000 1191.700 1700.340 ;
        RECT 1191.560 1639.130 1191.700 1700.000 ;
        RECT 413.640 1638.810 413.900 1639.130 ;
        RECT 1191.500 1638.810 1191.760 1639.130 ;
        RECT 413.700 16.990 413.840 1638.810 ;
        RECT 407.200 16.670 407.460 16.990 ;
        RECT 413.640 16.670 413.900 16.990 ;
        RECT 407.260 2.400 407.400 16.670 ;
        RECT 407.050 -4.800 407.610 2.400 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 86.090 1659.440 86.410 1659.500 ;
        RECT 1156.510 1659.440 1156.830 1659.500 ;
        RECT 86.090 1659.300 1156.830 1659.440 ;
        RECT 86.090 1659.240 86.410 1659.300 ;
        RECT 1156.510 1659.240 1156.830 1659.300 ;
        RECT 68.150 20.300 68.470 20.360 ;
        RECT 86.090 20.300 86.410 20.360 ;
        RECT 68.150 20.160 86.410 20.300 ;
        RECT 68.150 20.100 68.470 20.160 ;
        RECT 86.090 20.100 86.410 20.160 ;
      LAYER via ;
        RECT 86.120 1659.240 86.380 1659.500 ;
        RECT 1156.540 1659.240 1156.800 1659.500 ;
        RECT 68.180 20.100 68.440 20.360 ;
        RECT 86.120 20.100 86.380 20.360 ;
      LAYER met2 ;
        RECT 1156.440 1700.340 1156.720 1704.000 ;
        RECT 1156.440 1700.000 1156.740 1700.340 ;
        RECT 1156.600 1659.530 1156.740 1700.000 ;
        RECT 86.120 1659.210 86.380 1659.530 ;
        RECT 1156.540 1659.210 1156.800 1659.530 ;
        RECT 86.180 20.390 86.320 1659.210 ;
        RECT 68.180 20.070 68.440 20.390 ;
        RECT 86.120 20.070 86.380 20.390 ;
        RECT 68.240 2.400 68.380 20.070 ;
        RECT 68.030 -4.800 68.590 2.400 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 427.410 1590.420 427.730 1590.480 ;
        RECT 1193.310 1590.420 1193.630 1590.480 ;
        RECT 427.410 1590.280 1193.630 1590.420 ;
        RECT 427.410 1590.220 427.730 1590.280 ;
        RECT 1193.310 1590.220 1193.630 1590.280 ;
        RECT 424.650 16.560 424.970 16.620 ;
        RECT 427.410 16.560 427.730 16.620 ;
        RECT 424.650 16.420 427.730 16.560 ;
        RECT 424.650 16.360 424.970 16.420 ;
        RECT 427.410 16.360 427.730 16.420 ;
      LAYER via ;
        RECT 427.440 1590.220 427.700 1590.480 ;
        RECT 1193.340 1590.220 1193.600 1590.480 ;
        RECT 424.680 16.360 424.940 16.620 ;
        RECT 427.440 16.360 427.700 16.620 ;
      LAYER met2 ;
        RECT 1193.240 1700.340 1193.520 1704.000 ;
        RECT 1193.240 1700.000 1193.540 1700.340 ;
        RECT 1193.400 1590.510 1193.540 1700.000 ;
        RECT 427.440 1590.190 427.700 1590.510 ;
        RECT 1193.340 1590.190 1193.600 1590.510 ;
        RECT 427.500 16.650 427.640 1590.190 ;
        RECT 424.680 16.330 424.940 16.650 ;
        RECT 427.440 16.330 427.700 16.650 ;
        RECT 424.740 2.400 424.880 16.330 ;
        RECT 424.530 -4.800 425.090 2.400 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 482.685 1680.195 482.855 1680.535 ;
        RECT 524.545 1680.365 524.715 1681.895 ;
        RECT 572.385 1681.045 572.555 1681.895 ;
        RECT 579.285 1681.045 579.915 1681.215 ;
        RECT 579.745 1680.705 579.915 1681.045 ;
        RECT 662.545 1680.365 662.715 1681.215 ;
        RECT 710.385 1680.365 710.555 1681.215 ;
        RECT 717.745 1680.365 717.915 1681.215 ;
        RECT 1159.345 1680.365 1159.515 1682.915 ;
        RECT 482.225 1680.025 482.855 1680.195 ;
      LAYER mcon ;
        RECT 1159.345 1682.745 1159.515 1682.915 ;
        RECT 524.545 1681.725 524.715 1681.895 ;
        RECT 572.385 1681.725 572.555 1681.895 ;
        RECT 662.545 1681.045 662.715 1681.215 ;
        RECT 482.685 1680.365 482.855 1680.535 ;
        RECT 710.385 1681.045 710.555 1681.215 ;
        RECT 717.745 1681.045 717.915 1681.215 ;
      LAYER met1 ;
        RECT 1159.285 1682.900 1159.575 1682.945 ;
        RECT 1195.150 1682.900 1195.470 1682.960 ;
        RECT 1159.285 1682.760 1195.470 1682.900 ;
        RECT 1159.285 1682.715 1159.575 1682.760 ;
        RECT 1195.150 1682.700 1195.470 1682.760 ;
        RECT 524.485 1681.880 524.775 1681.925 ;
        RECT 572.325 1681.880 572.615 1681.925 ;
        RECT 524.485 1681.740 572.615 1681.880 ;
        RECT 524.485 1681.695 524.775 1681.740 ;
        RECT 572.325 1681.695 572.615 1681.740 ;
        RECT 572.325 1681.200 572.615 1681.245 ;
        RECT 579.225 1681.200 579.515 1681.245 ;
        RECT 572.325 1681.060 579.515 1681.200 ;
        RECT 572.325 1681.015 572.615 1681.060 ;
        RECT 579.225 1681.015 579.515 1681.060 ;
        RECT 662.485 1681.200 662.775 1681.245 ;
        RECT 710.325 1681.200 710.615 1681.245 ;
        RECT 662.485 1681.060 710.615 1681.200 ;
        RECT 662.485 1681.015 662.775 1681.060 ;
        RECT 710.325 1681.015 710.615 1681.060 ;
        RECT 717.685 1681.200 717.975 1681.245 ;
        RECT 717.685 1681.060 765.740 1681.200 ;
        RECT 717.685 1681.015 717.975 1681.060 ;
        RECT 579.685 1680.860 579.975 1680.905 ;
        RECT 579.685 1680.720 644.300 1680.860 ;
        RECT 579.685 1680.675 579.975 1680.720 ;
        RECT 482.625 1680.520 482.915 1680.565 ;
        RECT 524.485 1680.520 524.775 1680.565 ;
        RECT 482.625 1680.380 524.775 1680.520 ;
        RECT 644.160 1680.520 644.300 1680.720 ;
        RECT 662.485 1680.520 662.775 1680.565 ;
        RECT 644.160 1680.380 662.775 1680.520 ;
        RECT 482.625 1680.335 482.915 1680.380 ;
        RECT 524.485 1680.335 524.775 1680.380 ;
        RECT 662.485 1680.335 662.775 1680.380 ;
        RECT 710.325 1680.520 710.615 1680.565 ;
        RECT 717.685 1680.520 717.975 1680.565 ;
        RECT 710.325 1680.380 717.975 1680.520 ;
        RECT 765.600 1680.520 765.740 1681.060 ;
        RECT 765.970 1680.520 766.290 1680.580 ;
        RECT 765.600 1680.380 766.290 1680.520 ;
        RECT 710.325 1680.335 710.615 1680.380 ;
        RECT 717.685 1680.335 717.975 1680.380 ;
        RECT 765.970 1680.320 766.290 1680.380 ;
        RECT 766.430 1680.520 766.750 1680.580 ;
        RECT 1056.230 1680.520 1056.550 1680.580 ;
        RECT 766.430 1680.380 1056.550 1680.520 ;
        RECT 766.430 1680.320 766.750 1680.380 ;
        RECT 1056.230 1680.320 1056.550 1680.380 ;
        RECT 1056.690 1680.520 1057.010 1680.580 ;
        RECT 1159.285 1680.520 1159.575 1680.565 ;
        RECT 1056.690 1680.380 1159.575 1680.520 ;
        RECT 1056.690 1680.320 1057.010 1680.380 ;
        RECT 1159.285 1680.335 1159.575 1680.380 ;
        RECT 448.110 1680.180 448.430 1680.240 ;
        RECT 482.165 1680.180 482.455 1680.225 ;
        RECT 448.110 1680.040 482.455 1680.180 ;
        RECT 448.110 1679.980 448.430 1680.040 ;
        RECT 482.165 1679.995 482.455 1680.040 ;
        RECT 442.590 15.880 442.910 15.940 ;
        RECT 448.110 15.880 448.430 15.940 ;
        RECT 442.590 15.740 448.430 15.880 ;
        RECT 442.590 15.680 442.910 15.740 ;
        RECT 448.110 15.680 448.430 15.740 ;
      LAYER via ;
        RECT 1195.180 1682.700 1195.440 1682.960 ;
        RECT 766.000 1680.320 766.260 1680.580 ;
        RECT 766.460 1680.320 766.720 1680.580 ;
        RECT 1056.260 1680.320 1056.520 1680.580 ;
        RECT 1056.720 1680.320 1056.980 1680.580 ;
        RECT 448.140 1679.980 448.400 1680.240 ;
        RECT 442.620 15.680 442.880 15.940 ;
        RECT 448.140 15.680 448.400 15.940 ;
      LAYER met2 ;
        RECT 1195.080 1700.340 1195.360 1704.000 ;
        RECT 1195.080 1700.000 1195.380 1700.340 ;
        RECT 1195.240 1682.990 1195.380 1700.000 ;
        RECT 1195.180 1682.670 1195.440 1682.990 ;
        RECT 766.060 1681.060 766.660 1681.200 ;
        RECT 766.060 1680.610 766.200 1681.060 ;
        RECT 766.520 1680.610 766.660 1681.060 ;
        RECT 1056.320 1680.610 1056.920 1680.690 ;
        RECT 766.000 1680.290 766.260 1680.610 ;
        RECT 766.460 1680.290 766.720 1680.610 ;
        RECT 1056.260 1680.550 1056.980 1680.610 ;
        RECT 1056.260 1680.290 1056.520 1680.550 ;
        RECT 1056.720 1680.290 1056.980 1680.550 ;
        RECT 448.140 1679.950 448.400 1680.270 ;
        RECT 448.200 15.970 448.340 1679.950 ;
        RECT 442.620 15.650 442.880 15.970 ;
        RECT 448.140 15.650 448.400 15.970 ;
        RECT 442.680 2.400 442.820 15.650 ;
        RECT 442.470 -4.800 443.030 2.400 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1196.990 1656.180 1197.310 1656.440 ;
        RECT 1197.080 1656.040 1197.220 1656.180 ;
        RECT 1197.910 1656.040 1198.230 1656.100 ;
        RECT 1197.080 1655.900 1198.230 1656.040 ;
        RECT 1197.910 1655.840 1198.230 1655.900 ;
        RECT 461.910 1625.100 462.230 1625.160 ;
        RECT 1197.910 1625.100 1198.230 1625.160 ;
        RECT 461.910 1624.960 1198.230 1625.100 ;
        RECT 461.910 1624.900 462.230 1624.960 ;
        RECT 1197.910 1624.900 1198.230 1624.960 ;
        RECT 460.530 2.960 460.850 3.020 ;
        RECT 461.910 2.960 462.230 3.020 ;
        RECT 460.530 2.820 462.230 2.960 ;
        RECT 460.530 2.760 460.850 2.820 ;
        RECT 461.910 2.760 462.230 2.820 ;
      LAYER via ;
        RECT 1197.020 1656.180 1197.280 1656.440 ;
        RECT 1197.940 1655.840 1198.200 1656.100 ;
        RECT 461.940 1624.900 462.200 1625.160 ;
        RECT 1197.940 1624.900 1198.200 1625.160 ;
        RECT 460.560 2.760 460.820 3.020 ;
        RECT 461.940 2.760 462.200 3.020 ;
      LAYER met2 ;
        RECT 1196.920 1700.340 1197.200 1704.000 ;
        RECT 1196.920 1700.000 1197.220 1700.340 ;
        RECT 1197.080 1656.470 1197.220 1700.000 ;
        RECT 1197.020 1656.150 1197.280 1656.470 ;
        RECT 1197.940 1655.810 1198.200 1656.130 ;
        RECT 1198.000 1625.190 1198.140 1655.810 ;
        RECT 461.940 1624.870 462.200 1625.190 ;
        RECT 1197.940 1624.870 1198.200 1625.190 ;
        RECT 462.000 3.050 462.140 1624.870 ;
        RECT 460.560 2.730 460.820 3.050 ;
        RECT 461.940 2.730 462.200 3.050 ;
        RECT 460.620 2.400 460.760 2.730 ;
        RECT 460.410 -4.800 460.970 2.400 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1194.230 1678.140 1194.550 1678.200 ;
        RECT 1198.830 1678.140 1199.150 1678.200 ;
        RECT 1194.230 1678.000 1199.150 1678.140 ;
        RECT 1194.230 1677.940 1194.550 1678.000 ;
        RECT 1198.830 1677.940 1199.150 1678.000 ;
        RECT 482.610 1632.240 482.930 1632.300 ;
        RECT 1194.230 1632.240 1194.550 1632.300 ;
        RECT 482.610 1632.100 1194.550 1632.240 ;
        RECT 482.610 1632.040 482.930 1632.100 ;
        RECT 1194.230 1632.040 1194.550 1632.100 ;
        RECT 478.470 15.540 478.790 15.600 ;
        RECT 482.610 15.540 482.930 15.600 ;
        RECT 478.470 15.400 482.930 15.540 ;
        RECT 478.470 15.340 478.790 15.400 ;
        RECT 482.610 15.340 482.930 15.400 ;
      LAYER via ;
        RECT 1194.260 1677.940 1194.520 1678.200 ;
        RECT 1198.860 1677.940 1199.120 1678.200 ;
        RECT 482.640 1632.040 482.900 1632.300 ;
        RECT 1194.260 1632.040 1194.520 1632.300 ;
        RECT 478.500 15.340 478.760 15.600 ;
        RECT 482.640 15.340 482.900 15.600 ;
      LAYER met2 ;
        RECT 1198.760 1700.340 1199.040 1704.000 ;
        RECT 1198.760 1700.000 1199.060 1700.340 ;
        RECT 1198.920 1678.230 1199.060 1700.000 ;
        RECT 1194.260 1677.910 1194.520 1678.230 ;
        RECT 1198.860 1677.910 1199.120 1678.230 ;
        RECT 1194.320 1632.330 1194.460 1677.910 ;
        RECT 482.640 1632.010 482.900 1632.330 ;
        RECT 1194.260 1632.010 1194.520 1632.330 ;
        RECT 482.700 15.630 482.840 1632.010 ;
        RECT 478.500 15.310 478.760 15.630 ;
        RECT 482.640 15.310 482.900 15.630 ;
        RECT 478.560 2.400 478.700 15.310 ;
        RECT 478.350 -4.800 478.910 2.400 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 496.410 1618.300 496.730 1618.360 ;
        RECT 1201.130 1618.300 1201.450 1618.360 ;
        RECT 496.410 1618.160 1201.450 1618.300 ;
        RECT 496.410 1618.100 496.730 1618.160 ;
        RECT 1201.130 1618.100 1201.450 1618.160 ;
      LAYER via ;
        RECT 496.440 1618.100 496.700 1618.360 ;
        RECT 1201.160 1618.100 1201.420 1618.360 ;
      LAYER met2 ;
        RECT 1200.600 1700.340 1200.880 1704.000 ;
        RECT 1200.600 1700.000 1200.900 1700.340 ;
        RECT 1200.760 1665.900 1200.900 1700.000 ;
        RECT 1200.760 1665.760 1201.360 1665.900 ;
        RECT 1201.220 1618.390 1201.360 1665.760 ;
        RECT 496.440 1618.070 496.700 1618.390 ;
        RECT 1201.160 1618.070 1201.420 1618.390 ;
        RECT 496.500 2.400 496.640 1618.070 ;
        RECT 496.290 -4.800 496.850 2.400 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1202.510 1679.160 1202.830 1679.220 ;
        RECT 1207.110 1679.160 1207.430 1679.220 ;
        RECT 1202.510 1679.020 1207.430 1679.160 ;
        RECT 1202.510 1678.960 1202.830 1679.020 ;
        RECT 1207.110 1678.960 1207.430 1679.020 ;
        RECT 517.110 1611.500 517.430 1611.560 ;
        RECT 1207.110 1611.500 1207.430 1611.560 ;
        RECT 517.110 1611.360 1207.430 1611.500 ;
        RECT 517.110 1611.300 517.430 1611.360 ;
        RECT 1207.110 1611.300 1207.430 1611.360 ;
        RECT 513.890 15.540 514.210 15.600 ;
        RECT 517.110 15.540 517.430 15.600 ;
        RECT 513.890 15.400 517.430 15.540 ;
        RECT 513.890 15.340 514.210 15.400 ;
        RECT 517.110 15.340 517.430 15.400 ;
      LAYER via ;
        RECT 1202.540 1678.960 1202.800 1679.220 ;
        RECT 1207.140 1678.960 1207.400 1679.220 ;
        RECT 517.140 1611.300 517.400 1611.560 ;
        RECT 1207.140 1611.300 1207.400 1611.560 ;
        RECT 513.920 15.340 514.180 15.600 ;
        RECT 517.140 15.340 517.400 15.600 ;
      LAYER met2 ;
        RECT 1202.440 1700.340 1202.720 1704.000 ;
        RECT 1202.440 1700.000 1202.740 1700.340 ;
        RECT 1202.600 1679.250 1202.740 1700.000 ;
        RECT 1202.540 1678.930 1202.800 1679.250 ;
        RECT 1207.140 1678.930 1207.400 1679.250 ;
        RECT 1207.200 1611.590 1207.340 1678.930 ;
        RECT 517.140 1611.270 517.400 1611.590 ;
        RECT 1207.140 1611.270 1207.400 1611.590 ;
        RECT 517.200 15.630 517.340 1611.270 ;
        RECT 513.920 15.310 514.180 15.630 ;
        RECT 517.140 15.310 517.400 15.630 ;
        RECT 513.980 2.400 514.120 15.310 ;
        RECT 513.770 -4.800 514.330 2.400 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1203.505 1642.285 1203.675 1690.395 ;
      LAYER mcon ;
        RECT 1203.505 1690.225 1203.675 1690.395 ;
      LAYER met1 ;
        RECT 1203.445 1690.380 1203.735 1690.425 ;
        RECT 1204.350 1690.380 1204.670 1690.440 ;
        RECT 1203.445 1690.240 1204.670 1690.380 ;
        RECT 1203.445 1690.195 1203.735 1690.240 ;
        RECT 1204.350 1690.180 1204.670 1690.240 ;
        RECT 1203.430 1642.440 1203.750 1642.500 ;
        RECT 1203.235 1642.300 1203.750 1642.440 ;
        RECT 1203.430 1642.240 1203.750 1642.300 ;
        RECT 537.350 1583.620 537.670 1583.680 ;
        RECT 1203.430 1583.620 1203.750 1583.680 ;
        RECT 537.350 1583.480 1203.750 1583.620 ;
        RECT 537.350 1583.420 537.670 1583.480 ;
        RECT 1203.430 1583.420 1203.750 1583.480 ;
        RECT 531.830 15.540 532.150 15.600 ;
        RECT 537.350 15.540 537.670 15.600 ;
        RECT 531.830 15.400 537.670 15.540 ;
        RECT 531.830 15.340 532.150 15.400 ;
        RECT 537.350 15.340 537.670 15.400 ;
      LAYER via ;
        RECT 1204.380 1690.180 1204.640 1690.440 ;
        RECT 1203.460 1642.240 1203.720 1642.500 ;
        RECT 537.380 1583.420 537.640 1583.680 ;
        RECT 1203.460 1583.420 1203.720 1583.680 ;
        RECT 531.860 15.340 532.120 15.600 ;
        RECT 537.380 15.340 537.640 15.600 ;
      LAYER met2 ;
        RECT 1204.280 1700.340 1204.560 1704.000 ;
        RECT 1204.280 1700.000 1204.580 1700.340 ;
        RECT 1204.440 1690.470 1204.580 1700.000 ;
        RECT 1204.380 1690.150 1204.640 1690.470 ;
        RECT 1203.460 1642.210 1203.720 1642.530 ;
        RECT 1203.520 1583.710 1203.660 1642.210 ;
        RECT 537.380 1583.390 537.640 1583.710 ;
        RECT 1203.460 1583.390 1203.720 1583.710 ;
        RECT 537.440 15.630 537.580 1583.390 ;
        RECT 531.860 15.310 532.120 15.630 ;
        RECT 537.380 15.310 537.640 15.630 ;
        RECT 531.920 2.400 532.060 15.310 ;
        RECT 531.710 -4.800 532.270 2.400 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 551.610 1555.740 551.930 1555.800 ;
        RECT 1205.730 1555.740 1206.050 1555.800 ;
        RECT 551.610 1555.600 1206.050 1555.740 ;
        RECT 551.610 1555.540 551.930 1555.600 ;
        RECT 1205.730 1555.540 1206.050 1555.600 ;
        RECT 549.770 2.960 550.090 3.020 ;
        RECT 551.610 2.960 551.930 3.020 ;
        RECT 549.770 2.820 551.930 2.960 ;
        RECT 549.770 2.760 550.090 2.820 ;
        RECT 551.610 2.760 551.930 2.820 ;
      LAYER via ;
        RECT 551.640 1555.540 551.900 1555.800 ;
        RECT 1205.760 1555.540 1206.020 1555.800 ;
        RECT 549.800 2.760 550.060 3.020 ;
        RECT 551.640 2.760 551.900 3.020 ;
      LAYER met2 ;
        RECT 1206.120 1700.340 1206.400 1704.000 ;
        RECT 1206.120 1700.000 1206.420 1700.340 ;
        RECT 1206.280 1560.330 1206.420 1700.000 ;
        RECT 1205.820 1560.190 1206.420 1560.330 ;
        RECT 1205.820 1555.830 1205.960 1560.190 ;
        RECT 551.640 1555.510 551.900 1555.830 ;
        RECT 1205.760 1555.510 1206.020 1555.830 ;
        RECT 551.700 3.050 551.840 1555.510 ;
        RECT 549.800 2.730 550.060 3.050 ;
        RECT 551.640 2.730 551.900 3.050 ;
        RECT 549.860 2.400 550.000 2.730 ;
        RECT 549.650 -4.800 550.210 2.400 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1201.130 1683.920 1201.450 1683.980 ;
        RECT 1208.030 1683.920 1208.350 1683.980 ;
        RECT 1201.130 1683.780 1208.350 1683.920 ;
        RECT 1201.130 1683.720 1201.450 1683.780 ;
        RECT 1208.030 1683.720 1208.350 1683.780 ;
        RECT 572.310 1666.580 572.630 1666.640 ;
        RECT 1201.130 1666.580 1201.450 1666.640 ;
        RECT 572.310 1666.440 1201.450 1666.580 ;
        RECT 572.310 1666.380 572.630 1666.440 ;
        RECT 1201.130 1666.380 1201.450 1666.440 ;
        RECT 567.710 14.860 568.030 14.920 ;
        RECT 572.310 14.860 572.630 14.920 ;
        RECT 567.710 14.720 572.630 14.860 ;
        RECT 567.710 14.660 568.030 14.720 ;
        RECT 572.310 14.660 572.630 14.720 ;
      LAYER via ;
        RECT 1201.160 1683.720 1201.420 1683.980 ;
        RECT 1208.060 1683.720 1208.320 1683.980 ;
        RECT 572.340 1666.380 572.600 1666.640 ;
        RECT 1201.160 1666.380 1201.420 1666.640 ;
        RECT 567.740 14.660 568.000 14.920 ;
        RECT 572.340 14.660 572.600 14.920 ;
      LAYER met2 ;
        RECT 1207.960 1700.340 1208.240 1704.000 ;
        RECT 1207.960 1700.000 1208.260 1700.340 ;
        RECT 1208.120 1684.010 1208.260 1700.000 ;
        RECT 1201.160 1683.690 1201.420 1684.010 ;
        RECT 1208.060 1683.690 1208.320 1684.010 ;
        RECT 1201.220 1666.670 1201.360 1683.690 ;
        RECT 572.340 1666.350 572.600 1666.670 ;
        RECT 1201.160 1666.350 1201.420 1666.670 ;
        RECT 572.400 14.950 572.540 1666.350 ;
        RECT 567.740 14.630 568.000 14.950 ;
        RECT 572.340 14.630 572.600 14.950 ;
        RECT 567.800 2.400 567.940 14.630 ;
        RECT 567.590 -4.800 568.150 2.400 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 586.110 1673.380 586.430 1673.440 ;
        RECT 1209.870 1673.380 1210.190 1673.440 ;
        RECT 586.110 1673.240 1210.190 1673.380 ;
        RECT 586.110 1673.180 586.430 1673.240 ;
        RECT 1209.870 1673.180 1210.190 1673.240 ;
      LAYER via ;
        RECT 586.140 1673.180 586.400 1673.440 ;
        RECT 1209.900 1673.180 1210.160 1673.440 ;
      LAYER met2 ;
        RECT 1209.800 1700.340 1210.080 1704.000 ;
        RECT 1209.800 1700.000 1210.100 1700.340 ;
        RECT 1209.960 1673.470 1210.100 1700.000 ;
        RECT 586.140 1673.150 586.400 1673.470 ;
        RECT 1209.900 1673.150 1210.160 1673.470 ;
        RECT 586.200 24.210 586.340 1673.150 ;
        RECT 585.740 24.070 586.340 24.210 ;
        RECT 585.740 2.400 585.880 24.070 ;
        RECT 585.530 -4.800 586.090 2.400 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1157.505 1594.005 1157.675 1642.115 ;
      LAYER mcon ;
        RECT 1157.505 1641.945 1157.675 1642.115 ;
      LAYER met1 ;
        RECT 1157.890 1665.900 1158.210 1665.960 ;
        RECT 1158.810 1665.900 1159.130 1665.960 ;
        RECT 1157.890 1665.760 1159.130 1665.900 ;
        RECT 1157.890 1665.700 1158.210 1665.760 ;
        RECT 1158.810 1665.700 1159.130 1665.760 ;
        RECT 1157.445 1642.100 1157.735 1642.145 ;
        RECT 1157.890 1642.100 1158.210 1642.160 ;
        RECT 1157.445 1641.960 1158.210 1642.100 ;
        RECT 1157.445 1641.915 1157.735 1641.960 ;
        RECT 1157.890 1641.900 1158.210 1641.960 ;
        RECT 1157.430 1594.160 1157.750 1594.220 ;
        RECT 1157.235 1594.020 1157.750 1594.160 ;
        RECT 1157.430 1593.960 1157.750 1594.020 ;
        RECT 99.890 1576.480 100.210 1576.540 ;
        RECT 1157.890 1576.480 1158.210 1576.540 ;
        RECT 99.890 1576.340 1158.210 1576.480 ;
        RECT 99.890 1576.280 100.210 1576.340 ;
        RECT 1157.890 1576.280 1158.210 1576.340 ;
        RECT 91.610 17.580 91.930 17.640 ;
        RECT 99.890 17.580 100.210 17.640 ;
        RECT 91.610 17.440 100.210 17.580 ;
        RECT 91.610 17.380 91.930 17.440 ;
        RECT 99.890 17.380 100.210 17.440 ;
      LAYER via ;
        RECT 1157.920 1665.700 1158.180 1665.960 ;
        RECT 1158.840 1665.700 1159.100 1665.960 ;
        RECT 1157.920 1641.900 1158.180 1642.160 ;
        RECT 1157.460 1593.960 1157.720 1594.220 ;
        RECT 99.920 1576.280 100.180 1576.540 ;
        RECT 1157.920 1576.280 1158.180 1576.540 ;
        RECT 91.640 17.380 91.900 17.640 ;
        RECT 99.920 17.380 100.180 17.640 ;
      LAYER met2 ;
        RECT 1158.740 1700.340 1159.020 1704.000 ;
        RECT 1158.740 1700.000 1159.040 1700.340 ;
        RECT 1158.900 1665.990 1159.040 1700.000 ;
        RECT 1157.920 1665.670 1158.180 1665.990 ;
        RECT 1158.840 1665.670 1159.100 1665.990 ;
        RECT 1157.980 1642.190 1158.120 1665.670 ;
        RECT 1157.920 1641.870 1158.180 1642.190 ;
        RECT 1157.460 1593.930 1157.720 1594.250 ;
        RECT 1157.520 1593.650 1157.660 1593.930 ;
        RECT 1157.520 1593.510 1158.120 1593.650 ;
        RECT 1157.980 1576.570 1158.120 1593.510 ;
        RECT 99.920 1576.250 100.180 1576.570 ;
        RECT 1157.920 1576.250 1158.180 1576.570 ;
        RECT 99.980 17.670 100.120 1576.250 ;
        RECT 91.640 17.350 91.900 17.670 ;
        RECT 99.920 17.350 100.180 17.670 ;
        RECT 91.700 2.400 91.840 17.350 ;
        RECT 91.490 -4.800 92.050 2.400 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 606.810 1652.980 607.130 1653.040 ;
        RECT 1211.710 1652.980 1212.030 1653.040 ;
        RECT 606.810 1652.840 1212.030 1652.980 ;
        RECT 606.810 1652.780 607.130 1652.840 ;
        RECT 1211.710 1652.780 1212.030 1652.840 ;
        RECT 603.130 14.520 603.450 14.580 ;
        RECT 606.810 14.520 607.130 14.580 ;
        RECT 603.130 14.380 607.130 14.520 ;
        RECT 603.130 14.320 603.450 14.380 ;
        RECT 606.810 14.320 607.130 14.380 ;
      LAYER via ;
        RECT 606.840 1652.780 607.100 1653.040 ;
        RECT 1211.740 1652.780 1212.000 1653.040 ;
        RECT 603.160 14.320 603.420 14.580 ;
        RECT 606.840 14.320 607.100 14.580 ;
      LAYER met2 ;
        RECT 1211.640 1700.340 1211.920 1704.000 ;
        RECT 1211.640 1700.000 1211.940 1700.340 ;
        RECT 1211.800 1653.070 1211.940 1700.000 ;
        RECT 606.840 1652.750 607.100 1653.070 ;
        RECT 1211.740 1652.750 1212.000 1653.070 ;
        RECT 606.900 14.610 607.040 1652.750 ;
        RECT 603.160 14.290 603.420 14.610 ;
        RECT 606.840 14.290 607.100 14.610 ;
        RECT 603.220 2.400 603.360 14.290 ;
        RECT 603.010 -4.800 603.570 2.400 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1212.630 1678.140 1212.950 1678.200 ;
        RECT 1213.550 1678.140 1213.870 1678.200 ;
        RECT 1212.630 1678.000 1213.870 1678.140 ;
        RECT 1212.630 1677.940 1212.950 1678.000 ;
        RECT 1213.550 1677.940 1213.870 1678.000 ;
        RECT 627.050 1604.700 627.370 1604.760 ;
        RECT 1212.630 1604.700 1212.950 1604.760 ;
        RECT 627.050 1604.560 1212.950 1604.700 ;
        RECT 627.050 1604.500 627.370 1604.560 ;
        RECT 1212.630 1604.500 1212.950 1604.560 ;
        RECT 621.070 20.980 621.390 21.040 ;
        RECT 627.050 20.980 627.370 21.040 ;
        RECT 621.070 20.840 627.370 20.980 ;
        RECT 621.070 20.780 621.390 20.840 ;
        RECT 627.050 20.780 627.370 20.840 ;
      LAYER via ;
        RECT 1212.660 1677.940 1212.920 1678.200 ;
        RECT 1213.580 1677.940 1213.840 1678.200 ;
        RECT 627.080 1604.500 627.340 1604.760 ;
        RECT 1212.660 1604.500 1212.920 1604.760 ;
        RECT 621.100 20.780 621.360 21.040 ;
        RECT 627.080 20.780 627.340 21.040 ;
      LAYER met2 ;
        RECT 1213.480 1700.340 1213.760 1704.000 ;
        RECT 1213.480 1700.000 1213.780 1700.340 ;
        RECT 1213.640 1678.230 1213.780 1700.000 ;
        RECT 1212.660 1677.910 1212.920 1678.230 ;
        RECT 1213.580 1677.910 1213.840 1678.230 ;
        RECT 1212.720 1604.790 1212.860 1677.910 ;
        RECT 627.080 1604.470 627.340 1604.790 ;
        RECT 1212.660 1604.470 1212.920 1604.790 ;
        RECT 627.140 21.070 627.280 1604.470 ;
        RECT 621.100 20.750 621.360 21.070 ;
        RECT 627.080 20.750 627.340 21.070 ;
        RECT 621.160 2.400 621.300 20.750 ;
        RECT 620.950 -4.800 621.510 2.400 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 120.590 1569.680 120.910 1569.740 ;
        RECT 1162.030 1569.680 1162.350 1569.740 ;
        RECT 120.590 1569.540 1162.350 1569.680 ;
        RECT 120.590 1569.480 120.910 1569.540 ;
        RECT 1162.030 1569.480 1162.350 1569.540 ;
        RECT 115.530 17.580 115.850 17.640 ;
        RECT 120.590 17.580 120.910 17.640 ;
        RECT 115.530 17.440 120.910 17.580 ;
        RECT 115.530 17.380 115.850 17.440 ;
        RECT 120.590 17.380 120.910 17.440 ;
      LAYER via ;
        RECT 120.620 1569.480 120.880 1569.740 ;
        RECT 1162.060 1569.480 1162.320 1569.740 ;
        RECT 115.560 17.380 115.820 17.640 ;
        RECT 120.620 17.380 120.880 17.640 ;
      LAYER met2 ;
        RECT 1161.500 1700.340 1161.780 1704.000 ;
        RECT 1161.500 1700.000 1161.800 1700.340 ;
        RECT 1161.660 1677.970 1161.800 1700.000 ;
        RECT 1161.660 1677.830 1162.260 1677.970 ;
        RECT 1162.120 1569.770 1162.260 1677.830 ;
        RECT 120.620 1569.450 120.880 1569.770 ;
        RECT 1162.060 1569.450 1162.320 1569.770 ;
        RECT 120.680 17.670 120.820 1569.450 ;
        RECT 115.560 17.350 115.820 17.670 ;
        RECT 120.620 17.350 120.880 17.670 ;
        RECT 115.620 2.400 115.760 17.350 ;
        RECT 115.410 -4.800 115.970 2.400 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1161.110 1679.840 1161.430 1679.900 ;
        RECT 1163.870 1679.840 1164.190 1679.900 ;
        RECT 1161.110 1679.700 1164.190 1679.840 ;
        RECT 1161.110 1679.640 1161.430 1679.700 ;
        RECT 1163.870 1679.640 1164.190 1679.700 ;
        RECT 155.090 1548.940 155.410 1549.000 ;
        RECT 1161.570 1548.940 1161.890 1549.000 ;
        RECT 155.090 1548.800 1161.890 1548.940 ;
        RECT 155.090 1548.740 155.410 1548.800 ;
        RECT 1161.570 1548.740 1161.890 1548.800 ;
        RECT 139.450 16.220 139.770 16.280 ;
        RECT 155.090 16.220 155.410 16.280 ;
        RECT 139.450 16.080 155.410 16.220 ;
        RECT 139.450 16.020 139.770 16.080 ;
        RECT 155.090 16.020 155.410 16.080 ;
      LAYER via ;
        RECT 1161.140 1679.640 1161.400 1679.900 ;
        RECT 1163.900 1679.640 1164.160 1679.900 ;
        RECT 155.120 1548.740 155.380 1549.000 ;
        RECT 1161.600 1548.740 1161.860 1549.000 ;
        RECT 139.480 16.020 139.740 16.280 ;
        RECT 155.120 16.020 155.380 16.280 ;
      LAYER met2 ;
        RECT 1163.800 1700.340 1164.080 1704.000 ;
        RECT 1163.800 1700.000 1164.100 1700.340 ;
        RECT 1163.960 1679.930 1164.100 1700.000 ;
        RECT 1161.140 1679.610 1161.400 1679.930 ;
        RECT 1163.900 1679.610 1164.160 1679.930 ;
        RECT 1161.200 1677.290 1161.340 1679.610 ;
        RECT 1161.200 1677.150 1161.800 1677.290 ;
        RECT 1161.660 1549.030 1161.800 1677.150 ;
        RECT 155.120 1548.710 155.380 1549.030 ;
        RECT 1161.600 1548.710 1161.860 1549.030 ;
        RECT 155.180 16.310 155.320 1548.710 ;
        RECT 139.480 15.990 139.740 16.310 ;
        RECT 155.120 15.990 155.380 16.310 ;
        RECT 139.540 2.400 139.680 15.990 ;
        RECT 139.330 -4.800 139.890 2.400 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 158.310 1562.880 158.630 1562.940 ;
        RECT 1165.710 1562.880 1166.030 1562.940 ;
        RECT 158.310 1562.740 1166.030 1562.880 ;
        RECT 158.310 1562.680 158.630 1562.740 ;
        RECT 1165.710 1562.680 1166.030 1562.740 ;
      LAYER via ;
        RECT 158.340 1562.680 158.600 1562.940 ;
        RECT 1165.740 1562.680 1166.000 1562.940 ;
      LAYER met2 ;
        RECT 1165.640 1700.340 1165.920 1704.000 ;
        RECT 1165.640 1700.000 1165.940 1700.340 ;
        RECT 1165.800 1562.970 1165.940 1700.000 ;
        RECT 158.340 1562.650 158.600 1562.970 ;
        RECT 1165.740 1562.650 1166.000 1562.970 ;
        RECT 158.400 17.410 158.540 1562.650 ;
        RECT 157.480 17.270 158.540 17.410 ;
        RECT 157.480 2.400 157.620 17.270 ;
        RECT 157.270 -4.800 157.830 2.400 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 217.190 1535.340 217.510 1535.400 ;
        RECT 1168.470 1535.340 1168.790 1535.400 ;
        RECT 217.190 1535.200 1168.790 1535.340 ;
        RECT 217.190 1535.140 217.510 1535.200 ;
        RECT 1168.470 1535.140 1168.790 1535.200 ;
        RECT 174.870 17.920 175.190 17.980 ;
        RECT 217.190 17.920 217.510 17.980 ;
        RECT 174.870 17.780 186.600 17.920 ;
        RECT 174.870 17.720 175.190 17.780 ;
        RECT 186.460 17.580 186.600 17.780 ;
        RECT 193.360 17.780 217.510 17.920 ;
        RECT 193.360 17.580 193.500 17.780 ;
        RECT 217.190 17.720 217.510 17.780 ;
        RECT 186.460 17.440 193.500 17.580 ;
      LAYER via ;
        RECT 217.220 1535.140 217.480 1535.400 ;
        RECT 1168.500 1535.140 1168.760 1535.400 ;
        RECT 174.900 17.720 175.160 17.980 ;
        RECT 217.220 17.720 217.480 17.980 ;
      LAYER met2 ;
        RECT 1167.480 1700.340 1167.760 1704.000 ;
        RECT 1167.480 1700.000 1167.780 1700.340 ;
        RECT 1167.640 1679.840 1167.780 1700.000 ;
        RECT 1167.640 1679.700 1168.240 1679.840 ;
        RECT 1168.100 1678.650 1168.240 1679.700 ;
        RECT 1168.100 1678.510 1168.700 1678.650 ;
        RECT 1168.560 1535.430 1168.700 1678.510 ;
        RECT 217.220 1535.110 217.480 1535.430 ;
        RECT 1168.500 1535.110 1168.760 1535.430 ;
        RECT 217.280 18.010 217.420 1535.110 ;
        RECT 174.900 17.690 175.160 18.010 ;
        RECT 217.220 17.690 217.480 18.010 ;
        RECT 174.960 2.400 175.100 17.690 ;
        RECT 174.750 -4.800 175.310 2.400 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER li1 ;
        RECT 1167.625 1587.205 1167.795 1635.315 ;
        RECT 1167.625 1528.045 1167.795 1545.555 ;
      LAYER mcon ;
        RECT 1167.625 1635.145 1167.795 1635.315 ;
        RECT 1167.625 1545.385 1167.795 1545.555 ;
      LAYER met1 ;
        RECT 1168.010 1668.620 1168.330 1668.680 ;
        RECT 1169.390 1668.620 1169.710 1668.680 ;
        RECT 1168.010 1668.480 1169.710 1668.620 ;
        RECT 1168.010 1668.420 1168.330 1668.480 ;
        RECT 1169.390 1668.420 1169.710 1668.480 ;
        RECT 1167.565 1635.300 1167.855 1635.345 ;
        RECT 1168.010 1635.300 1168.330 1635.360 ;
        RECT 1167.565 1635.160 1168.330 1635.300 ;
        RECT 1167.565 1635.115 1167.855 1635.160 ;
        RECT 1168.010 1635.100 1168.330 1635.160 ;
        RECT 1167.550 1587.360 1167.870 1587.420 ;
        RECT 1167.355 1587.220 1167.870 1587.360 ;
        RECT 1167.550 1587.160 1167.870 1587.220 ;
        RECT 1167.550 1545.540 1167.870 1545.600 ;
        RECT 1167.355 1545.400 1167.870 1545.540 ;
        RECT 1167.550 1545.340 1167.870 1545.400 ;
        RECT 192.350 1528.200 192.670 1528.260 ;
        RECT 1167.565 1528.200 1167.855 1528.245 ;
        RECT 192.350 1528.060 1167.855 1528.200 ;
        RECT 192.350 1528.000 192.670 1528.060 ;
        RECT 1167.565 1528.015 1167.855 1528.060 ;
      LAYER via ;
        RECT 1168.040 1668.420 1168.300 1668.680 ;
        RECT 1169.420 1668.420 1169.680 1668.680 ;
        RECT 1168.040 1635.100 1168.300 1635.360 ;
        RECT 1167.580 1587.160 1167.840 1587.420 ;
        RECT 1167.580 1545.340 1167.840 1545.600 ;
        RECT 192.380 1528.000 192.640 1528.260 ;
      LAYER met2 ;
        RECT 1169.320 1700.340 1169.600 1704.000 ;
        RECT 1169.320 1700.000 1169.620 1700.340 ;
        RECT 1169.480 1668.710 1169.620 1700.000 ;
        RECT 1168.040 1668.390 1168.300 1668.710 ;
        RECT 1169.420 1668.390 1169.680 1668.710 ;
        RECT 1168.100 1635.390 1168.240 1668.390 ;
        RECT 1168.040 1635.070 1168.300 1635.390 ;
        RECT 1167.580 1587.130 1167.840 1587.450 ;
        RECT 1167.640 1545.630 1167.780 1587.130 ;
        RECT 1167.580 1545.310 1167.840 1545.630 ;
        RECT 192.380 1527.970 192.640 1528.290 ;
        RECT 192.440 17.410 192.580 1527.970 ;
        RECT 192.440 17.270 193.040 17.410 ;
        RECT 192.900 2.400 193.040 17.270 ;
        RECT 192.690 -4.800 193.250 2.400 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 213.510 1521.400 213.830 1521.460 ;
        RECT 1171.230 1521.400 1171.550 1521.460 ;
        RECT 213.510 1521.260 1171.550 1521.400 ;
        RECT 213.510 1521.200 213.830 1521.260 ;
        RECT 1171.230 1521.200 1171.550 1521.260 ;
        RECT 210.750 17.580 211.070 17.640 ;
        RECT 213.510 17.580 213.830 17.640 ;
        RECT 210.750 17.440 213.830 17.580 ;
        RECT 210.750 17.380 211.070 17.440 ;
        RECT 213.510 17.380 213.830 17.440 ;
      LAYER via ;
        RECT 213.540 1521.200 213.800 1521.460 ;
        RECT 1171.260 1521.200 1171.520 1521.460 ;
        RECT 210.780 17.380 211.040 17.640 ;
        RECT 213.540 17.380 213.800 17.640 ;
      LAYER met2 ;
        RECT 1171.160 1700.340 1171.440 1704.000 ;
        RECT 1171.160 1700.000 1171.460 1700.340 ;
        RECT 1171.320 1521.490 1171.460 1700.000 ;
        RECT 213.540 1521.170 213.800 1521.490 ;
        RECT 1171.260 1521.170 1171.520 1521.490 ;
        RECT 213.600 17.670 213.740 1521.170 ;
        RECT 210.780 17.350 211.040 17.670 ;
        RECT 213.540 17.350 213.800 17.670 ;
        RECT 210.840 2.400 210.980 17.350 ;
        RECT 210.630 -4.800 211.190 2.400 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 1173.070 1665.560 1173.390 1665.620 ;
        RECT 1174.910 1665.560 1175.230 1665.620 ;
        RECT 1173.070 1665.420 1175.230 1665.560 ;
        RECT 1173.070 1665.360 1173.390 1665.420 ;
        RECT 1174.910 1665.360 1175.230 1665.420 ;
        RECT 251.690 1597.220 252.010 1597.280 ;
        RECT 1174.910 1597.220 1175.230 1597.280 ;
        RECT 251.690 1597.080 1175.230 1597.220 ;
        RECT 251.690 1597.020 252.010 1597.080 ;
        RECT 1174.910 1597.020 1175.230 1597.080 ;
        RECT 228.690 14.520 229.010 14.580 ;
        RECT 251.690 14.520 252.010 14.580 ;
        RECT 228.690 14.380 252.010 14.520 ;
        RECT 228.690 14.320 229.010 14.380 ;
        RECT 251.690 14.320 252.010 14.380 ;
      LAYER via ;
        RECT 1173.100 1665.360 1173.360 1665.620 ;
        RECT 1174.940 1665.360 1175.200 1665.620 ;
        RECT 251.720 1597.020 251.980 1597.280 ;
        RECT 1174.940 1597.020 1175.200 1597.280 ;
        RECT 228.720 14.320 228.980 14.580 ;
        RECT 251.720 14.320 251.980 14.580 ;
      LAYER met2 ;
        RECT 1173.000 1700.340 1173.280 1704.000 ;
        RECT 1173.000 1700.000 1173.300 1700.340 ;
        RECT 1173.160 1665.650 1173.300 1700.000 ;
        RECT 1173.100 1665.330 1173.360 1665.650 ;
        RECT 1174.940 1665.330 1175.200 1665.650 ;
        RECT 1175.000 1597.310 1175.140 1665.330 ;
        RECT 251.720 1596.990 251.980 1597.310 ;
        RECT 1174.940 1596.990 1175.200 1597.310 ;
        RECT 251.780 14.610 251.920 1596.990 ;
        RECT 228.720 14.290 228.980 14.610 ;
        RECT 251.720 14.290 251.980 14.610 ;
        RECT 228.780 2.400 228.920 14.290 ;
        RECT 228.570 -4.800 229.130 2.400 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 72.290 1687.320 72.610 1687.380 ;
        RECT 1154.670 1687.320 1154.990 1687.380 ;
        RECT 72.290 1687.180 1154.990 1687.320 ;
        RECT 72.290 1687.120 72.610 1687.180 ;
        RECT 1154.670 1687.120 1154.990 1687.180 ;
        RECT 50.210 17.580 50.530 17.640 ;
        RECT 72.290 17.580 72.610 17.640 ;
        RECT 50.210 17.440 72.610 17.580 ;
        RECT 50.210 17.380 50.530 17.440 ;
        RECT 72.290 17.380 72.610 17.440 ;
      LAYER via ;
        RECT 72.320 1687.120 72.580 1687.380 ;
        RECT 1154.700 1687.120 1154.960 1687.380 ;
        RECT 50.240 17.380 50.500 17.640 ;
        RECT 72.320 17.380 72.580 17.640 ;
      LAYER met2 ;
        RECT 1154.600 1700.340 1154.880 1704.000 ;
        RECT 1154.600 1700.000 1154.900 1700.340 ;
        RECT 1154.760 1687.410 1154.900 1700.000 ;
        RECT 72.320 1687.090 72.580 1687.410 ;
        RECT 1154.700 1687.090 1154.960 1687.410 ;
        RECT 72.380 17.670 72.520 1687.090 ;
        RECT 50.240 17.350 50.500 17.670 ;
        RECT 72.320 17.350 72.580 17.670 ;
        RECT 50.300 2.400 50.440 17.350 ;
        RECT 50.090 -4.800 50.650 2.400 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 254.910 1514.600 255.230 1514.660 ;
        RECT 1175.370 1514.600 1175.690 1514.660 ;
        RECT 254.910 1514.460 1175.690 1514.600 ;
        RECT 254.910 1514.400 255.230 1514.460 ;
        RECT 1175.370 1514.400 1175.690 1514.460 ;
        RECT 252.610 17.920 252.930 17.980 ;
        RECT 254.910 17.920 255.230 17.980 ;
        RECT 252.610 17.780 255.230 17.920 ;
        RECT 252.610 17.720 252.930 17.780 ;
        RECT 254.910 17.720 255.230 17.780 ;
      LAYER via ;
        RECT 254.940 1514.400 255.200 1514.660 ;
        RECT 1175.400 1514.400 1175.660 1514.660 ;
        RECT 252.640 17.720 252.900 17.980 ;
        RECT 254.940 17.720 255.200 17.980 ;
      LAYER met2 ;
        RECT 1175.300 1700.340 1175.580 1704.000 ;
        RECT 1175.300 1700.000 1175.600 1700.340 ;
        RECT 1175.460 1514.690 1175.600 1700.000 ;
        RECT 254.940 1514.370 255.200 1514.690 ;
        RECT 1175.400 1514.370 1175.660 1514.690 ;
        RECT 255.000 18.010 255.140 1514.370 ;
        RECT 252.640 17.690 252.900 18.010 ;
        RECT 254.940 17.690 255.200 18.010 ;
        RECT 252.700 2.400 252.840 17.690 ;
        RECT 252.490 -4.800 253.050 2.400 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1175.830 1664.880 1176.150 1664.940 ;
        RECT 1177.210 1664.880 1177.530 1664.940 ;
        RECT 1175.830 1664.740 1177.530 1664.880 ;
        RECT 1175.830 1664.680 1176.150 1664.740 ;
        RECT 1177.210 1664.680 1177.530 1664.740 ;
        RECT 270.090 18.260 270.410 18.320 ;
        RECT 1175.830 18.260 1176.150 18.320 ;
        RECT 270.090 18.120 1176.150 18.260 ;
        RECT 270.090 18.060 270.410 18.120 ;
        RECT 1175.830 18.060 1176.150 18.120 ;
      LAYER via ;
        RECT 1175.860 1664.680 1176.120 1664.940 ;
        RECT 1177.240 1664.680 1177.500 1664.940 ;
        RECT 270.120 18.060 270.380 18.320 ;
        RECT 1175.860 18.060 1176.120 18.320 ;
      LAYER met2 ;
        RECT 1177.140 1700.340 1177.420 1704.000 ;
        RECT 1177.140 1700.000 1177.440 1700.340 ;
        RECT 1177.300 1664.970 1177.440 1700.000 ;
        RECT 1175.860 1664.650 1176.120 1664.970 ;
        RECT 1177.240 1664.650 1177.500 1664.970 ;
        RECT 1175.920 18.350 1176.060 1664.650 ;
        RECT 270.120 18.030 270.380 18.350 ;
        RECT 1175.860 18.030 1176.120 18.350 ;
        RECT 270.180 2.400 270.320 18.030 ;
        RECT 269.970 -4.800 270.530 2.400 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1162.105 18.445 1162.275 20.315 ;
      LAYER mcon ;
        RECT 1162.105 20.145 1162.275 20.315 ;
      LAYER met1 ;
        RECT 1162.045 20.300 1162.335 20.345 ;
        RECT 1179.050 20.300 1179.370 20.360 ;
        RECT 1162.045 20.160 1179.370 20.300 ;
        RECT 1162.045 20.115 1162.335 20.160 ;
        RECT 1179.050 20.100 1179.370 20.160 ;
        RECT 288.030 18.600 288.350 18.660 ;
        RECT 1162.045 18.600 1162.335 18.645 ;
        RECT 288.030 18.460 1162.335 18.600 ;
        RECT 288.030 18.400 288.350 18.460 ;
        RECT 1162.045 18.415 1162.335 18.460 ;
      LAYER via ;
        RECT 1179.080 20.100 1179.340 20.360 ;
        RECT 288.060 18.400 288.320 18.660 ;
      LAYER met2 ;
        RECT 1178.980 1700.340 1179.260 1704.000 ;
        RECT 1178.980 1700.000 1179.280 1700.340 ;
        RECT 1179.140 20.390 1179.280 1700.000 ;
        RECT 1179.080 20.070 1179.340 20.390 ;
        RECT 288.060 18.370 288.320 18.690 ;
        RECT 288.120 2.400 288.260 18.370 ;
        RECT 287.910 -4.800 288.470 2.400 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 305.970 18.940 306.290 19.000 ;
        RECT 1180.430 18.940 1180.750 19.000 ;
        RECT 305.970 18.800 1180.750 18.940 ;
        RECT 305.970 18.740 306.290 18.800 ;
        RECT 1180.430 18.740 1180.750 18.800 ;
      LAYER via ;
        RECT 306.000 18.740 306.260 19.000 ;
        RECT 1180.460 18.740 1180.720 19.000 ;
      LAYER met2 ;
        RECT 1180.820 1700.340 1181.100 1704.000 ;
        RECT 1180.820 1700.000 1181.120 1700.340 ;
        RECT 1180.980 1669.810 1181.120 1700.000 ;
        RECT 1180.520 1669.670 1181.120 1669.810 ;
        RECT 1180.520 19.030 1180.660 1669.670 ;
        RECT 306.000 18.710 306.260 19.030 ;
        RECT 1180.460 18.710 1180.720 19.030 ;
        RECT 306.060 2.400 306.200 18.710 ;
        RECT 305.850 -4.800 306.410 2.400 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1181.350 1680.520 1181.670 1680.580 ;
        RECT 1182.730 1680.520 1183.050 1680.580 ;
        RECT 1181.350 1680.380 1183.050 1680.520 ;
        RECT 1181.350 1680.320 1181.670 1680.380 ;
        RECT 1182.730 1680.320 1183.050 1680.380 ;
        RECT 323.450 19.280 323.770 19.340 ;
        RECT 1180.890 19.280 1181.210 19.340 ;
        RECT 323.450 19.140 1181.210 19.280 ;
        RECT 323.450 19.080 323.770 19.140 ;
        RECT 1180.890 19.080 1181.210 19.140 ;
      LAYER via ;
        RECT 1181.380 1680.320 1181.640 1680.580 ;
        RECT 1182.760 1680.320 1183.020 1680.580 ;
        RECT 323.480 19.080 323.740 19.340 ;
        RECT 1180.920 19.080 1181.180 19.340 ;
      LAYER met2 ;
        RECT 1182.660 1700.340 1182.940 1704.000 ;
        RECT 1182.660 1700.000 1182.960 1700.340 ;
        RECT 1182.820 1680.610 1182.960 1700.000 ;
        RECT 1181.380 1680.290 1181.640 1680.610 ;
        RECT 1182.760 1680.290 1183.020 1680.610 ;
        RECT 1181.440 1669.130 1181.580 1680.290 ;
        RECT 1180.980 1668.990 1181.580 1669.130 ;
        RECT 1180.980 19.370 1181.120 1668.990 ;
        RECT 323.480 19.050 323.740 19.370 ;
        RECT 1180.920 19.050 1181.180 19.370 ;
        RECT 323.540 9.930 323.680 19.050 ;
        RECT 323.540 9.790 324.140 9.930 ;
        RECT 324.000 2.400 324.140 9.790 ;
        RECT 323.790 -4.800 324.350 2.400 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1181.350 1668.620 1181.670 1668.680 ;
        RECT 1184.570 1668.620 1184.890 1668.680 ;
        RECT 1181.350 1668.480 1184.890 1668.620 ;
        RECT 1181.350 1668.420 1181.670 1668.480 ;
        RECT 1184.570 1668.420 1184.890 1668.480 ;
        RECT 341.390 19.620 341.710 19.680 ;
        RECT 1181.350 19.620 1181.670 19.680 ;
        RECT 341.390 19.480 1181.670 19.620 ;
        RECT 341.390 19.420 341.710 19.480 ;
        RECT 1181.350 19.420 1181.670 19.480 ;
      LAYER via ;
        RECT 1181.380 1668.420 1181.640 1668.680 ;
        RECT 1184.600 1668.420 1184.860 1668.680 ;
        RECT 341.420 19.420 341.680 19.680 ;
        RECT 1181.380 19.420 1181.640 19.680 ;
      LAYER met2 ;
        RECT 1184.500 1700.340 1184.780 1704.000 ;
        RECT 1184.500 1700.000 1184.800 1700.340 ;
        RECT 1184.660 1668.710 1184.800 1700.000 ;
        RECT 1181.380 1668.390 1181.640 1668.710 ;
        RECT 1184.600 1668.390 1184.860 1668.710 ;
        RECT 1181.440 19.710 1181.580 1668.390 ;
        RECT 341.420 19.390 341.680 19.710 ;
        RECT 1181.380 19.390 1181.640 19.710 ;
        RECT 341.480 2.400 341.620 19.390 ;
        RECT 341.270 -4.800 341.830 2.400 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 372.745 15.385 372.915 19.975 ;
        RECT 420.125 15.385 420.295 19.975 ;
        RECT 469.345 14.705 469.515 19.975 ;
        RECT 517.185 14.705 517.355 19.975 ;
      LAYER mcon ;
        RECT 372.745 19.805 372.915 19.975 ;
        RECT 420.125 19.805 420.295 19.975 ;
        RECT 469.345 19.805 469.515 19.975 ;
        RECT 517.185 19.805 517.355 19.975 ;
      LAYER met1 ;
        RECT 1185.030 1656.380 1185.350 1656.440 ;
        RECT 1186.410 1656.380 1186.730 1656.440 ;
        RECT 1185.030 1656.240 1186.730 1656.380 ;
        RECT 1185.030 1656.180 1185.350 1656.240 ;
        RECT 1186.410 1656.180 1186.730 1656.240 ;
        RECT 359.330 19.960 359.650 20.020 ;
        RECT 372.685 19.960 372.975 20.005 ;
        RECT 359.330 19.820 372.975 19.960 ;
        RECT 359.330 19.760 359.650 19.820 ;
        RECT 372.685 19.775 372.975 19.820 ;
        RECT 420.065 19.960 420.355 20.005 ;
        RECT 469.285 19.960 469.575 20.005 ;
        RECT 420.065 19.820 469.575 19.960 ;
        RECT 420.065 19.775 420.355 19.820 ;
        RECT 469.285 19.775 469.575 19.820 ;
        RECT 517.125 19.960 517.415 20.005 ;
        RECT 1185.030 19.960 1185.350 20.020 ;
        RECT 517.125 19.820 1185.350 19.960 ;
        RECT 517.125 19.775 517.415 19.820 ;
        RECT 1185.030 19.760 1185.350 19.820 ;
        RECT 372.685 15.540 372.975 15.585 ;
        RECT 420.065 15.540 420.355 15.585 ;
        RECT 372.685 15.400 420.355 15.540 ;
        RECT 372.685 15.355 372.975 15.400 ;
        RECT 420.065 15.355 420.355 15.400 ;
        RECT 469.285 14.860 469.575 14.905 ;
        RECT 517.125 14.860 517.415 14.905 ;
        RECT 469.285 14.720 517.415 14.860 ;
        RECT 469.285 14.675 469.575 14.720 ;
        RECT 517.125 14.675 517.415 14.720 ;
      LAYER via ;
        RECT 1185.060 1656.180 1185.320 1656.440 ;
        RECT 1186.440 1656.180 1186.700 1656.440 ;
        RECT 359.360 19.760 359.620 20.020 ;
        RECT 1185.060 19.760 1185.320 20.020 ;
      LAYER met2 ;
        RECT 1186.340 1700.340 1186.620 1704.000 ;
        RECT 1186.340 1700.000 1186.640 1700.340 ;
        RECT 1186.500 1656.470 1186.640 1700.000 ;
        RECT 1185.060 1656.150 1185.320 1656.470 ;
        RECT 1186.440 1656.150 1186.700 1656.470 ;
        RECT 1185.120 20.050 1185.260 1656.150 ;
        RECT 359.360 19.730 359.620 20.050 ;
        RECT 1185.060 19.730 1185.320 20.050 ;
        RECT 359.420 2.400 359.560 19.730 ;
        RECT 359.210 -4.800 359.770 2.400 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 469.805 14.365 469.975 20.315 ;
        RECT 516.725 14.365 516.895 20.315 ;
        RECT 1161.645 17.085 1161.815 20.315 ;
      LAYER mcon ;
        RECT 469.805 20.145 469.975 20.315 ;
        RECT 516.725 20.145 516.895 20.315 ;
        RECT 1161.645 20.145 1161.815 20.315 ;
      LAYER met1 ;
        RECT 1188.710 1678.820 1189.030 1678.880 ;
        RECT 1192.390 1678.820 1192.710 1678.880 ;
        RECT 1188.710 1678.680 1192.710 1678.820 ;
        RECT 1188.710 1678.620 1189.030 1678.680 ;
        RECT 1192.390 1678.620 1192.710 1678.680 ;
        RECT 420.510 20.300 420.830 20.360 ;
        RECT 469.745 20.300 470.035 20.345 ;
        RECT 420.510 20.160 470.035 20.300 ;
        RECT 420.510 20.100 420.830 20.160 ;
        RECT 469.745 20.115 470.035 20.160 ;
        RECT 516.665 20.300 516.955 20.345 ;
        RECT 1161.585 20.300 1161.875 20.345 ;
        RECT 516.665 20.160 1161.875 20.300 ;
        RECT 516.665 20.115 516.955 20.160 ;
        RECT 1161.585 20.115 1161.875 20.160 ;
        RECT 1161.585 17.240 1161.875 17.285 ;
        RECT 1192.390 17.240 1192.710 17.300 ;
        RECT 1161.585 17.100 1192.710 17.240 ;
        RECT 1161.585 17.055 1161.875 17.100 ;
        RECT 1192.390 17.040 1192.710 17.100 ;
        RECT 377.270 15.880 377.590 15.940 ;
        RECT 420.510 15.880 420.830 15.940 ;
        RECT 377.270 15.740 420.830 15.880 ;
        RECT 377.270 15.680 377.590 15.740 ;
        RECT 420.510 15.680 420.830 15.740 ;
        RECT 469.745 14.520 470.035 14.565 ;
        RECT 516.665 14.520 516.955 14.565 ;
        RECT 469.745 14.380 516.955 14.520 ;
        RECT 469.745 14.335 470.035 14.380 ;
        RECT 516.665 14.335 516.955 14.380 ;
      LAYER via ;
        RECT 1188.740 1678.620 1189.000 1678.880 ;
        RECT 1192.420 1678.620 1192.680 1678.880 ;
        RECT 420.540 20.100 420.800 20.360 ;
        RECT 1192.420 17.040 1192.680 17.300 ;
        RECT 377.300 15.680 377.560 15.940 ;
        RECT 420.540 15.680 420.800 15.940 ;
      LAYER met2 ;
        RECT 1188.180 1700.410 1188.460 1704.000 ;
        RECT 1188.180 1700.270 1188.940 1700.410 ;
        RECT 1188.180 1700.000 1188.460 1700.270 ;
        RECT 1188.800 1678.910 1188.940 1700.270 ;
        RECT 1188.740 1678.590 1189.000 1678.910 ;
        RECT 1192.420 1678.590 1192.680 1678.910 ;
        RECT 420.540 20.070 420.800 20.390 ;
        RECT 420.600 15.970 420.740 20.070 ;
        RECT 1192.480 17.330 1192.620 1678.590 ;
        RECT 1192.420 17.010 1192.680 17.330 ;
        RECT 377.300 15.650 377.560 15.970 ;
        RECT 420.540 15.650 420.800 15.970 ;
        RECT 377.360 2.400 377.500 15.650 ;
        RECT 377.150 -4.800 377.710 2.400 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 395.210 20.640 395.530 20.700 ;
        RECT 1190.090 20.640 1190.410 20.700 ;
        RECT 395.210 20.500 1190.410 20.640 ;
        RECT 395.210 20.440 395.530 20.500 ;
        RECT 1190.090 20.440 1190.410 20.500 ;
      LAYER via ;
        RECT 395.240 20.440 395.500 20.700 ;
        RECT 1190.120 20.440 1190.380 20.700 ;
      LAYER met2 ;
        RECT 1190.020 1700.340 1190.300 1704.000 ;
        RECT 1190.020 1700.000 1190.320 1700.340 ;
        RECT 1190.180 20.730 1190.320 1700.000 ;
        RECT 395.240 20.410 395.500 20.730 ;
        RECT 1190.120 20.410 1190.380 20.730 ;
        RECT 395.300 2.400 395.440 20.410 ;
        RECT 395.090 -4.800 395.650 2.400 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1191.085 814.385 1191.255 862.495 ;
        RECT 1191.085 717.825 1191.255 765.935 ;
        RECT 1190.625 614.125 1190.795 669.375 ;
        RECT 1190.165 565.505 1190.335 607.155 ;
        RECT 1190.625 462.485 1190.795 510.595 ;
        RECT 1191.085 276.165 1191.255 324.275 ;
        RECT 1191.085 234.685 1191.255 255.595 ;
        RECT 1191.545 179.945 1191.715 227.715 ;
        RECT 1190.625 131.325 1190.795 179.435 ;
      LAYER mcon ;
        RECT 1191.085 862.325 1191.255 862.495 ;
        RECT 1191.085 765.765 1191.255 765.935 ;
        RECT 1190.625 669.205 1190.795 669.375 ;
        RECT 1190.165 606.985 1190.335 607.155 ;
        RECT 1190.625 510.425 1190.795 510.595 ;
        RECT 1191.085 324.105 1191.255 324.275 ;
        RECT 1191.085 255.425 1191.255 255.595 ;
        RECT 1191.545 227.545 1191.715 227.715 ;
        RECT 1190.625 179.265 1190.795 179.435 ;
      LAYER met1 ;
        RECT 1190.550 1648.900 1190.870 1648.960 ;
        RECT 1191.930 1648.900 1192.250 1648.960 ;
        RECT 1190.550 1648.760 1192.250 1648.900 ;
        RECT 1190.550 1648.700 1190.870 1648.760 ;
        RECT 1191.930 1648.700 1192.250 1648.760 ;
        RECT 1190.550 1511.340 1190.870 1511.600 ;
        RECT 1190.640 1510.520 1190.780 1511.340 ;
        RECT 1191.010 1510.520 1191.330 1510.580 ;
        RECT 1190.640 1510.380 1191.330 1510.520 ;
        RECT 1191.010 1510.320 1191.330 1510.380 ;
        RECT 1190.550 1448.980 1190.870 1449.040 ;
        RECT 1191.010 1448.980 1191.330 1449.040 ;
        RECT 1190.550 1448.840 1191.330 1448.980 ;
        RECT 1190.550 1448.780 1190.870 1448.840 ;
        RECT 1191.010 1448.780 1191.330 1448.840 ;
        RECT 1190.550 1186.840 1190.870 1186.900 ;
        RECT 1191.470 1186.840 1191.790 1186.900 ;
        RECT 1190.550 1186.700 1191.790 1186.840 ;
        RECT 1190.550 1186.640 1190.870 1186.700 ;
        RECT 1191.470 1186.640 1191.790 1186.700 ;
        RECT 1191.010 862.480 1191.330 862.540 ;
        RECT 1190.815 862.340 1191.330 862.480 ;
        RECT 1191.010 862.280 1191.330 862.340 ;
        RECT 1191.010 814.540 1191.330 814.600 ;
        RECT 1190.815 814.400 1191.330 814.540 ;
        RECT 1191.010 814.340 1191.330 814.400 ;
        RECT 1191.010 765.920 1191.330 765.980 ;
        RECT 1190.815 765.780 1191.330 765.920 ;
        RECT 1191.010 765.720 1191.330 765.780 ;
        RECT 1191.010 717.980 1191.330 718.040 ;
        RECT 1190.815 717.840 1191.330 717.980 ;
        RECT 1191.010 717.780 1191.330 717.840 ;
        RECT 1190.550 669.360 1190.870 669.420 ;
        RECT 1190.355 669.220 1190.870 669.360 ;
        RECT 1190.550 669.160 1190.870 669.220 ;
        RECT 1190.550 614.280 1190.870 614.340 ;
        RECT 1190.355 614.140 1190.870 614.280 ;
        RECT 1190.550 614.080 1190.870 614.140 ;
        RECT 1190.105 607.140 1190.395 607.185 ;
        RECT 1190.550 607.140 1190.870 607.200 ;
        RECT 1190.105 607.000 1190.870 607.140 ;
        RECT 1190.105 606.955 1190.395 607.000 ;
        RECT 1190.550 606.940 1190.870 607.000 ;
        RECT 1190.105 565.660 1190.395 565.705 ;
        RECT 1190.550 565.660 1190.870 565.720 ;
        RECT 1190.105 565.520 1190.870 565.660 ;
        RECT 1190.105 565.475 1190.395 565.520 ;
        RECT 1190.550 565.460 1190.870 565.520 ;
        RECT 1190.550 517.720 1190.870 517.780 ;
        RECT 1191.010 517.720 1191.330 517.780 ;
        RECT 1190.550 517.580 1191.330 517.720 ;
        RECT 1190.550 517.520 1190.870 517.580 ;
        RECT 1191.010 517.520 1191.330 517.580 ;
        RECT 1190.565 510.580 1190.855 510.625 ;
        RECT 1191.010 510.580 1191.330 510.640 ;
        RECT 1190.565 510.440 1191.330 510.580 ;
        RECT 1190.565 510.395 1190.855 510.440 ;
        RECT 1191.010 510.380 1191.330 510.440 ;
        RECT 1190.550 462.640 1190.870 462.700 ;
        RECT 1190.355 462.500 1190.870 462.640 ;
        RECT 1190.550 462.440 1190.870 462.500 ;
        RECT 1190.550 427.960 1190.870 428.020 ;
        RECT 1191.010 427.960 1191.330 428.020 ;
        RECT 1190.550 427.820 1191.330 427.960 ;
        RECT 1190.550 427.760 1190.870 427.820 ;
        RECT 1191.010 427.760 1191.330 427.820 ;
        RECT 1191.010 324.260 1191.330 324.320 ;
        RECT 1190.815 324.120 1191.330 324.260 ;
        RECT 1191.010 324.060 1191.330 324.120 ;
        RECT 1191.010 276.320 1191.330 276.380 ;
        RECT 1190.815 276.180 1191.330 276.320 ;
        RECT 1191.010 276.120 1191.330 276.180 ;
        RECT 1191.010 255.580 1191.330 255.640 ;
        RECT 1190.815 255.440 1191.330 255.580 ;
        RECT 1191.010 255.380 1191.330 255.440 ;
        RECT 1191.010 234.840 1191.330 234.900 ;
        RECT 1190.815 234.700 1191.330 234.840 ;
        RECT 1191.010 234.640 1191.330 234.700 ;
        RECT 1191.010 227.700 1191.330 227.760 ;
        RECT 1191.485 227.700 1191.775 227.745 ;
        RECT 1191.010 227.560 1191.775 227.700 ;
        RECT 1191.010 227.500 1191.330 227.560 ;
        RECT 1191.485 227.515 1191.775 227.560 ;
        RECT 1191.010 180.100 1191.330 180.160 ;
        RECT 1191.485 180.100 1191.775 180.145 ;
        RECT 1191.010 179.960 1191.775 180.100 ;
        RECT 1191.010 179.900 1191.330 179.960 ;
        RECT 1191.485 179.915 1191.775 179.960 ;
        RECT 1190.565 179.420 1190.855 179.465 ;
        RECT 1191.010 179.420 1191.330 179.480 ;
        RECT 1190.565 179.280 1191.330 179.420 ;
        RECT 1190.565 179.235 1190.855 179.280 ;
        RECT 1191.010 179.220 1191.330 179.280 ;
        RECT 1190.550 131.480 1190.870 131.540 ;
        RECT 1190.355 131.340 1190.870 131.480 ;
        RECT 1190.550 131.280 1190.870 131.340 ;
        RECT 1190.550 17.920 1190.870 17.980 ;
        RECT 1170.860 17.780 1190.870 17.920 ;
        RECT 1166.170 17.580 1166.490 17.640 ;
        RECT 1170.860 17.580 1171.000 17.780 ;
        RECT 1190.550 17.720 1190.870 17.780 ;
        RECT 1166.170 17.440 1171.000 17.580 ;
        RECT 1166.170 17.380 1166.490 17.440 ;
        RECT 1154.670 16.900 1154.990 16.960 ;
        RECT 414.160 16.760 1154.990 16.900 ;
        RECT 413.150 16.220 413.470 16.280 ;
        RECT 414.160 16.220 414.300 16.760 ;
        RECT 1154.670 16.700 1154.990 16.760 ;
        RECT 413.150 16.080 414.300 16.220 ;
        RECT 413.150 16.020 413.470 16.080 ;
      LAYER via ;
        RECT 1190.580 1648.700 1190.840 1648.960 ;
        RECT 1191.960 1648.700 1192.220 1648.960 ;
        RECT 1190.580 1511.340 1190.840 1511.600 ;
        RECT 1191.040 1510.320 1191.300 1510.580 ;
        RECT 1190.580 1448.780 1190.840 1449.040 ;
        RECT 1191.040 1448.780 1191.300 1449.040 ;
        RECT 1190.580 1186.640 1190.840 1186.900 ;
        RECT 1191.500 1186.640 1191.760 1186.900 ;
        RECT 1191.040 862.280 1191.300 862.540 ;
        RECT 1191.040 814.340 1191.300 814.600 ;
        RECT 1191.040 765.720 1191.300 765.980 ;
        RECT 1191.040 717.780 1191.300 718.040 ;
        RECT 1190.580 669.160 1190.840 669.420 ;
        RECT 1190.580 614.080 1190.840 614.340 ;
        RECT 1190.580 606.940 1190.840 607.200 ;
        RECT 1190.580 565.460 1190.840 565.720 ;
        RECT 1190.580 517.520 1190.840 517.780 ;
        RECT 1191.040 517.520 1191.300 517.780 ;
        RECT 1191.040 510.380 1191.300 510.640 ;
        RECT 1190.580 462.440 1190.840 462.700 ;
        RECT 1190.580 427.760 1190.840 428.020 ;
        RECT 1191.040 427.760 1191.300 428.020 ;
        RECT 1191.040 324.060 1191.300 324.320 ;
        RECT 1191.040 276.120 1191.300 276.380 ;
        RECT 1191.040 255.380 1191.300 255.640 ;
        RECT 1191.040 234.640 1191.300 234.900 ;
        RECT 1191.040 227.500 1191.300 227.760 ;
        RECT 1191.040 179.900 1191.300 180.160 ;
        RECT 1191.040 179.220 1191.300 179.480 ;
        RECT 1190.580 131.280 1190.840 131.540 ;
        RECT 1166.200 17.380 1166.460 17.640 ;
        RECT 1190.580 17.720 1190.840 17.980 ;
        RECT 413.180 16.020 413.440 16.280 ;
        RECT 1154.700 16.700 1154.960 16.960 ;
      LAYER met2 ;
        RECT 1191.860 1700.340 1192.140 1704.000 ;
        RECT 1191.860 1700.000 1192.160 1700.340 ;
        RECT 1192.020 1648.990 1192.160 1700.000 ;
        RECT 1190.580 1648.670 1190.840 1648.990 ;
        RECT 1191.960 1648.670 1192.220 1648.990 ;
        RECT 1190.640 1511.630 1190.780 1648.670 ;
        RECT 1190.580 1511.310 1190.840 1511.630 ;
        RECT 1191.040 1510.290 1191.300 1510.610 ;
        RECT 1191.100 1449.070 1191.240 1510.290 ;
        RECT 1190.580 1448.750 1190.840 1449.070 ;
        RECT 1191.040 1448.750 1191.300 1449.070 ;
        RECT 1190.640 1425.010 1190.780 1448.750 ;
        RECT 1190.640 1424.870 1191.240 1425.010 ;
        RECT 1191.100 1366.530 1191.240 1424.870 ;
        RECT 1190.640 1366.390 1191.240 1366.530 ;
        RECT 1190.640 1365.850 1190.780 1366.390 ;
        RECT 1190.640 1365.710 1191.240 1365.850 ;
        RECT 1191.100 1269.970 1191.240 1365.710 ;
        RECT 1190.640 1269.830 1191.240 1269.970 ;
        RECT 1190.640 1269.290 1190.780 1269.830 ;
        RECT 1190.640 1269.150 1191.240 1269.290 ;
        RECT 1191.100 1221.690 1191.240 1269.150 ;
        RECT 1191.100 1221.550 1191.700 1221.690 ;
        RECT 1191.560 1194.605 1191.700 1221.550 ;
        RECT 1191.490 1194.235 1191.770 1194.605 ;
        RECT 1190.570 1193.555 1190.850 1193.925 ;
        RECT 1190.640 1186.930 1190.780 1193.555 ;
        RECT 1190.580 1186.610 1190.840 1186.930 ;
        RECT 1191.500 1186.610 1191.760 1186.930 ;
        RECT 1191.560 1072.770 1191.700 1186.610 ;
        RECT 1191.100 1072.630 1191.700 1072.770 ;
        RECT 1191.100 883.050 1191.240 1072.630 ;
        RECT 1190.640 882.910 1191.240 883.050 ;
        RECT 1190.640 881.690 1190.780 882.910 ;
        RECT 1190.640 881.550 1191.240 881.690 ;
        RECT 1191.100 862.570 1191.240 881.550 ;
        RECT 1191.040 862.250 1191.300 862.570 ;
        RECT 1191.040 814.310 1191.300 814.630 ;
        RECT 1191.100 766.010 1191.240 814.310 ;
        RECT 1191.040 765.690 1191.300 766.010 ;
        RECT 1191.040 717.750 1191.300 718.070 ;
        RECT 1191.100 669.530 1191.240 717.750 ;
        RECT 1190.640 669.450 1191.240 669.530 ;
        RECT 1190.580 669.390 1191.240 669.450 ;
        RECT 1190.580 669.130 1190.840 669.390 ;
        RECT 1190.640 668.975 1190.780 669.130 ;
        RECT 1190.580 614.050 1190.840 614.370 ;
        RECT 1190.640 607.230 1190.780 614.050 ;
        RECT 1190.580 606.910 1190.840 607.230 ;
        RECT 1190.580 565.430 1190.840 565.750 ;
        RECT 1190.640 517.810 1190.780 565.430 ;
        RECT 1190.580 517.490 1190.840 517.810 ;
        RECT 1191.040 517.490 1191.300 517.810 ;
        RECT 1191.100 510.670 1191.240 517.490 ;
        RECT 1191.040 510.350 1191.300 510.670 ;
        RECT 1190.580 462.410 1190.840 462.730 ;
        RECT 1190.640 428.050 1190.780 462.410 ;
        RECT 1190.580 427.730 1190.840 428.050 ;
        RECT 1191.040 427.730 1191.300 428.050 ;
        RECT 1191.100 400.930 1191.240 427.730 ;
        RECT 1190.640 400.790 1191.240 400.930 ;
        RECT 1190.640 400.250 1190.780 400.790 ;
        RECT 1190.640 400.110 1191.240 400.250 ;
        RECT 1191.100 345.170 1191.240 400.110 ;
        RECT 1190.640 345.030 1191.240 345.170 ;
        RECT 1190.640 338.200 1190.780 345.030 ;
        RECT 1190.640 338.060 1191.240 338.200 ;
        RECT 1191.100 324.350 1191.240 338.060 ;
        RECT 1191.040 324.030 1191.300 324.350 ;
        RECT 1191.040 276.090 1191.300 276.410 ;
        RECT 1191.100 255.670 1191.240 276.090 ;
        RECT 1191.040 255.350 1191.300 255.670 ;
        RECT 1191.040 234.610 1191.300 234.930 ;
        RECT 1191.100 227.790 1191.240 234.610 ;
        RECT 1191.040 227.470 1191.300 227.790 ;
        RECT 1191.040 179.870 1191.300 180.190 ;
        RECT 1191.100 179.510 1191.240 179.870 ;
        RECT 1191.040 179.190 1191.300 179.510 ;
        RECT 1190.580 131.250 1190.840 131.570 ;
        RECT 1190.640 18.010 1190.780 131.250 ;
        RECT 1190.580 17.690 1190.840 18.010 ;
        RECT 1166.200 17.525 1166.460 17.670 ;
        RECT 1154.690 17.155 1154.970 17.525 ;
        RECT 1166.190 17.155 1166.470 17.525 ;
        RECT 1154.760 16.990 1154.900 17.155 ;
        RECT 1154.700 16.670 1154.960 16.990 ;
        RECT 413.180 15.990 413.440 16.310 ;
        RECT 413.240 2.400 413.380 15.990 ;
        RECT 413.030 -4.800 413.590 2.400 ;
      LAYER via2 ;
        RECT 1191.490 1194.280 1191.770 1194.560 ;
        RECT 1190.570 1193.600 1190.850 1193.880 ;
        RECT 1154.690 17.200 1154.970 17.480 ;
        RECT 1166.190 17.200 1166.470 17.480 ;
      LAYER met3 ;
        RECT 1191.465 1194.570 1191.795 1194.585 ;
        RECT 1189.870 1194.270 1191.795 1194.570 ;
        RECT 1189.870 1193.890 1190.170 1194.270 ;
        RECT 1191.465 1194.255 1191.795 1194.270 ;
        RECT 1190.545 1193.890 1190.875 1193.905 ;
        RECT 1189.870 1193.590 1190.875 1193.890 ;
        RECT 1190.545 1193.575 1190.875 1193.590 ;
        RECT 1154.665 17.490 1154.995 17.505 ;
        RECT 1166.165 17.490 1166.495 17.505 ;
        RECT 1154.665 17.190 1166.495 17.490 ;
        RECT 1154.665 17.175 1154.995 17.190 ;
        RECT 1166.165 17.175 1166.495 17.190 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1153.290 1678.140 1153.610 1678.200 ;
        RECT 1156.970 1678.140 1157.290 1678.200 ;
        RECT 1153.290 1678.000 1157.290 1678.140 ;
        RECT 1153.290 1677.940 1153.610 1678.000 ;
        RECT 1156.970 1677.940 1157.290 1678.000 ;
      LAYER via ;
        RECT 1153.320 1677.940 1153.580 1678.200 ;
        RECT 1157.000 1677.940 1157.260 1678.200 ;
      LAYER met2 ;
        RECT 1156.900 1700.340 1157.180 1704.000 ;
        RECT 1156.900 1700.000 1157.200 1700.340 ;
        RECT 1157.060 1678.230 1157.200 1700.000 ;
        RECT 1153.320 1677.910 1153.580 1678.230 ;
        RECT 1157.000 1677.910 1157.260 1678.230 ;
        RECT 1153.380 17.525 1153.520 1677.910 ;
        RECT 74.150 17.155 74.430 17.525 ;
        RECT 1153.310 17.155 1153.590 17.525 ;
        RECT 74.220 2.400 74.360 17.155 ;
        RECT 74.010 -4.800 74.570 2.400 ;
      LAYER via2 ;
        RECT 74.150 17.200 74.430 17.480 ;
        RECT 1153.310 17.200 1153.590 17.480 ;
      LAYER met3 ;
        RECT 74.125 17.490 74.455 17.505 ;
        RECT 1153.285 17.490 1153.615 17.505 ;
        RECT 74.125 17.190 1153.615 17.490 ;
        RECT 74.125 17.175 74.455 17.190 ;
        RECT 1153.285 17.175 1153.615 17.190 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1145.470 16.560 1145.790 16.620 ;
        RECT 448.200 16.420 1145.790 16.560 ;
        RECT 430.630 16.220 430.950 16.280 ;
        RECT 448.200 16.220 448.340 16.420 ;
        RECT 1145.470 16.360 1145.790 16.420 ;
        RECT 430.630 16.080 448.340 16.220 ;
        RECT 1168.930 16.220 1169.250 16.280 ;
        RECT 1193.770 16.220 1194.090 16.280 ;
        RECT 1168.930 16.080 1194.090 16.220 ;
        RECT 430.630 16.020 430.950 16.080 ;
        RECT 1168.930 16.020 1169.250 16.080 ;
        RECT 1193.770 16.020 1194.090 16.080 ;
      LAYER via ;
        RECT 430.660 16.020 430.920 16.280 ;
        RECT 1145.500 16.360 1145.760 16.620 ;
        RECT 1168.960 16.020 1169.220 16.280 ;
        RECT 1193.800 16.020 1194.060 16.280 ;
      LAYER met2 ;
        RECT 1193.700 1700.340 1193.980 1704.000 ;
        RECT 1193.700 1700.000 1194.000 1700.340 ;
        RECT 1145.500 16.330 1145.760 16.650 ;
        RECT 430.660 15.990 430.920 16.310 ;
        RECT 1145.560 16.165 1145.700 16.330 ;
        RECT 1193.860 16.310 1194.000 1700.000 ;
        RECT 1168.960 16.165 1169.220 16.310 ;
        RECT 430.720 2.400 430.860 15.990 ;
        RECT 1145.490 15.795 1145.770 16.165 ;
        RECT 1168.950 15.795 1169.230 16.165 ;
        RECT 1193.800 15.990 1194.060 16.310 ;
        RECT 430.510 -4.800 431.070 2.400 ;
      LAYER via2 ;
        RECT 1145.490 15.840 1145.770 16.120 ;
        RECT 1168.950 15.840 1169.230 16.120 ;
      LAYER met3 ;
        RECT 1145.465 16.130 1145.795 16.145 ;
        RECT 1168.925 16.130 1169.255 16.145 ;
        RECT 1145.465 15.830 1169.255 16.130 ;
        RECT 1145.465 15.815 1145.795 15.830 ;
        RECT 1168.925 15.815 1169.255 15.830 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1194.765 1587.205 1194.935 1597.575 ;
        RECT 1194.765 1497.445 1194.935 1545.555 ;
        RECT 1194.765 1026.545 1194.935 1094.375 ;
        RECT 1194.765 735.845 1194.935 765.935 ;
        RECT 1193.845 576.725 1194.015 607.155 ;
        RECT 1194.765 324.445 1194.935 372.555 ;
        RECT 1194.765 227.885 1194.935 275.995 ;
        RECT 1194.305 83.045 1194.475 107.355 ;
      LAYER mcon ;
        RECT 1194.765 1597.405 1194.935 1597.575 ;
        RECT 1194.765 1545.385 1194.935 1545.555 ;
        RECT 1194.765 1094.205 1194.935 1094.375 ;
        RECT 1194.765 765.765 1194.935 765.935 ;
        RECT 1193.845 606.985 1194.015 607.155 ;
        RECT 1194.765 372.385 1194.935 372.555 ;
        RECT 1194.765 275.825 1194.935 275.995 ;
        RECT 1194.305 107.185 1194.475 107.355 ;
      LAYER met1 ;
        RECT 1194.690 1666.240 1195.010 1666.300 ;
        RECT 1195.610 1666.240 1195.930 1666.300 ;
        RECT 1194.690 1666.100 1195.930 1666.240 ;
        RECT 1194.690 1666.040 1195.010 1666.100 ;
        RECT 1195.610 1666.040 1195.930 1666.100 ;
        RECT 1194.690 1597.560 1195.010 1597.620 ;
        RECT 1194.495 1597.420 1195.010 1597.560 ;
        RECT 1194.690 1597.360 1195.010 1597.420 ;
        RECT 1194.690 1587.360 1195.010 1587.420 ;
        RECT 1194.495 1587.220 1195.010 1587.360 ;
        RECT 1194.690 1587.160 1195.010 1587.220 ;
        RECT 1194.690 1545.540 1195.010 1545.600 ;
        RECT 1194.495 1545.400 1195.010 1545.540 ;
        RECT 1194.690 1545.340 1195.010 1545.400 ;
        RECT 1194.690 1497.600 1195.010 1497.660 ;
        RECT 1194.495 1497.460 1195.010 1497.600 ;
        RECT 1194.690 1497.400 1195.010 1497.460 ;
        RECT 1194.690 1145.360 1195.010 1145.420 ;
        RECT 1195.610 1145.360 1195.930 1145.420 ;
        RECT 1194.690 1145.220 1195.930 1145.360 ;
        RECT 1194.690 1145.160 1195.010 1145.220 ;
        RECT 1195.610 1145.160 1195.930 1145.220 ;
        RECT 1194.230 1094.360 1194.550 1094.420 ;
        RECT 1194.705 1094.360 1194.995 1094.405 ;
        RECT 1194.230 1094.220 1194.995 1094.360 ;
        RECT 1194.230 1094.160 1194.550 1094.220 ;
        RECT 1194.705 1094.175 1194.995 1094.220 ;
        RECT 1194.690 1026.700 1195.010 1026.760 ;
        RECT 1194.495 1026.560 1195.010 1026.700 ;
        RECT 1194.690 1026.500 1195.010 1026.560 ;
        RECT 1194.690 814.200 1195.010 814.260 ;
        RECT 1195.610 814.200 1195.930 814.260 ;
        RECT 1194.690 814.060 1195.930 814.200 ;
        RECT 1194.690 814.000 1195.010 814.060 ;
        RECT 1195.610 814.000 1195.930 814.060 ;
        RECT 1194.690 765.920 1195.010 765.980 ;
        RECT 1194.495 765.780 1195.010 765.920 ;
        RECT 1194.690 765.720 1195.010 765.780 ;
        RECT 1194.690 736.000 1195.010 736.060 ;
        RECT 1194.495 735.860 1195.010 736.000 ;
        RECT 1194.690 735.800 1195.010 735.860 ;
        RECT 1193.310 669.360 1193.630 669.420 ;
        RECT 1194.690 669.360 1195.010 669.420 ;
        RECT 1193.310 669.220 1195.010 669.360 ;
        RECT 1193.310 669.160 1193.630 669.220 ;
        RECT 1194.690 669.160 1195.010 669.220 ;
        RECT 1193.785 607.140 1194.075 607.185 ;
        RECT 1194.230 607.140 1194.550 607.200 ;
        RECT 1193.785 607.000 1194.550 607.140 ;
        RECT 1193.785 606.955 1194.075 607.000 ;
        RECT 1194.230 606.940 1194.550 607.000 ;
        RECT 1193.785 576.880 1194.075 576.925 ;
        RECT 1194.230 576.880 1194.550 576.940 ;
        RECT 1193.785 576.740 1194.550 576.880 ;
        RECT 1193.785 576.695 1194.075 576.740 ;
        RECT 1194.230 576.680 1194.550 576.740 ;
        RECT 1194.230 531.460 1194.550 531.720 ;
        RECT 1194.320 531.040 1194.460 531.460 ;
        RECT 1194.230 530.780 1194.550 531.040 ;
        RECT 1194.230 475.700 1194.550 475.960 ;
        RECT 1194.320 475.560 1194.460 475.700 ;
        RECT 1194.690 475.560 1195.010 475.620 ;
        RECT 1194.320 475.420 1195.010 475.560 ;
        RECT 1194.690 475.360 1195.010 475.420 ;
        RECT 1194.690 372.540 1195.010 372.600 ;
        RECT 1194.495 372.400 1195.010 372.540 ;
        RECT 1194.690 372.340 1195.010 372.400 ;
        RECT 1194.690 324.600 1195.010 324.660 ;
        RECT 1194.690 324.460 1195.205 324.600 ;
        RECT 1194.690 324.400 1195.010 324.460 ;
        RECT 1194.690 275.980 1195.010 276.040 ;
        RECT 1194.495 275.840 1195.010 275.980 ;
        RECT 1194.690 275.780 1195.010 275.840 ;
        RECT 1194.690 228.040 1195.010 228.100 ;
        RECT 1194.690 227.900 1195.205 228.040 ;
        RECT 1194.690 227.840 1195.010 227.900 ;
        RECT 1194.690 193.360 1195.010 193.420 ;
        RECT 1194.320 193.220 1195.010 193.360 ;
        RECT 1194.320 193.080 1194.460 193.220 ;
        RECT 1194.690 193.160 1195.010 193.220 ;
        RECT 1194.230 192.820 1194.550 193.080 ;
        RECT 1194.230 145.080 1194.550 145.140 ;
        RECT 1194.690 145.080 1195.010 145.140 ;
        RECT 1194.230 144.940 1195.010 145.080 ;
        RECT 1194.230 144.880 1194.550 144.940 ;
        RECT 1194.690 144.880 1195.010 144.940 ;
        RECT 1194.245 107.340 1194.535 107.385 ;
        RECT 1194.690 107.340 1195.010 107.400 ;
        RECT 1194.245 107.200 1195.010 107.340 ;
        RECT 1194.245 107.155 1194.535 107.200 ;
        RECT 1194.690 107.140 1195.010 107.200 ;
        RECT 1194.230 83.200 1194.550 83.260 ;
        RECT 1194.035 83.060 1194.550 83.200 ;
        RECT 1194.230 83.000 1194.550 83.060 ;
        RECT 448.570 16.220 448.890 16.280 ;
        RECT 448.570 16.080 1168.700 16.220 ;
        RECT 448.570 16.020 448.890 16.080 ;
        RECT 1168.560 15.880 1168.700 16.080 ;
        RECT 1194.230 15.880 1194.550 15.940 ;
        RECT 1168.560 15.740 1194.550 15.880 ;
        RECT 1194.230 15.680 1194.550 15.740 ;
      LAYER via ;
        RECT 1194.720 1666.040 1194.980 1666.300 ;
        RECT 1195.640 1666.040 1195.900 1666.300 ;
        RECT 1194.720 1597.360 1194.980 1597.620 ;
        RECT 1194.720 1587.160 1194.980 1587.420 ;
        RECT 1194.720 1545.340 1194.980 1545.600 ;
        RECT 1194.720 1497.400 1194.980 1497.660 ;
        RECT 1194.720 1145.160 1194.980 1145.420 ;
        RECT 1195.640 1145.160 1195.900 1145.420 ;
        RECT 1194.260 1094.160 1194.520 1094.420 ;
        RECT 1194.720 1026.500 1194.980 1026.760 ;
        RECT 1194.720 814.000 1194.980 814.260 ;
        RECT 1195.640 814.000 1195.900 814.260 ;
        RECT 1194.720 765.720 1194.980 765.980 ;
        RECT 1194.720 735.800 1194.980 736.060 ;
        RECT 1193.340 669.160 1193.600 669.420 ;
        RECT 1194.720 669.160 1194.980 669.420 ;
        RECT 1194.260 606.940 1194.520 607.200 ;
        RECT 1194.260 576.680 1194.520 576.940 ;
        RECT 1194.260 531.460 1194.520 531.720 ;
        RECT 1194.260 530.780 1194.520 531.040 ;
        RECT 1194.260 475.700 1194.520 475.960 ;
        RECT 1194.720 475.360 1194.980 475.620 ;
        RECT 1194.720 372.340 1194.980 372.600 ;
        RECT 1194.720 324.400 1194.980 324.660 ;
        RECT 1194.720 275.780 1194.980 276.040 ;
        RECT 1194.720 227.840 1194.980 228.100 ;
        RECT 1194.720 193.160 1194.980 193.420 ;
        RECT 1194.260 192.820 1194.520 193.080 ;
        RECT 1194.260 144.880 1194.520 145.140 ;
        RECT 1194.720 144.880 1194.980 145.140 ;
        RECT 1194.720 107.140 1194.980 107.400 ;
        RECT 1194.260 83.000 1194.520 83.260 ;
        RECT 448.600 16.020 448.860 16.280 ;
        RECT 1194.260 15.680 1194.520 15.940 ;
      LAYER met2 ;
        RECT 1195.540 1700.340 1195.820 1704.000 ;
        RECT 1195.540 1700.000 1195.840 1700.340 ;
        RECT 1195.700 1666.330 1195.840 1700.000 ;
        RECT 1194.720 1666.010 1194.980 1666.330 ;
        RECT 1195.640 1666.010 1195.900 1666.330 ;
        RECT 1194.780 1597.650 1194.920 1666.010 ;
        RECT 1194.720 1597.330 1194.980 1597.650 ;
        RECT 1194.720 1587.130 1194.980 1587.450 ;
        RECT 1194.780 1545.630 1194.920 1587.130 ;
        RECT 1194.720 1545.310 1194.980 1545.630 ;
        RECT 1194.720 1497.370 1194.980 1497.690 ;
        RECT 1194.780 1318.250 1194.920 1497.370 ;
        RECT 1194.320 1318.110 1194.920 1318.250 ;
        RECT 1194.320 1317.570 1194.460 1318.110 ;
        RECT 1194.320 1317.430 1194.920 1317.570 ;
        RECT 1194.780 1221.690 1194.920 1317.430 ;
        RECT 1194.320 1221.550 1194.920 1221.690 ;
        RECT 1194.320 1221.010 1194.460 1221.550 ;
        RECT 1194.320 1220.870 1194.920 1221.010 ;
        RECT 1194.780 1145.450 1194.920 1220.870 ;
        RECT 1194.720 1145.130 1194.980 1145.450 ;
        RECT 1195.640 1145.130 1195.900 1145.450 ;
        RECT 1195.700 1097.365 1195.840 1145.130 ;
        RECT 1194.250 1096.995 1194.530 1097.365 ;
        RECT 1195.630 1096.995 1195.910 1097.365 ;
        RECT 1194.320 1094.450 1194.460 1096.995 ;
        RECT 1194.260 1094.130 1194.520 1094.450 ;
        RECT 1194.720 1026.470 1194.980 1026.790 ;
        RECT 1194.780 932.010 1194.920 1026.470 ;
        RECT 1194.320 931.870 1194.920 932.010 ;
        RECT 1194.320 931.330 1194.460 931.870 ;
        RECT 1194.320 931.190 1194.920 931.330 ;
        RECT 1194.780 835.450 1194.920 931.190 ;
        RECT 1194.320 835.310 1194.920 835.450 ;
        RECT 1194.320 834.770 1194.460 835.310 ;
        RECT 1194.320 834.630 1194.920 834.770 ;
        RECT 1194.780 814.290 1194.920 834.630 ;
        RECT 1194.720 813.970 1194.980 814.290 ;
        RECT 1195.640 813.970 1195.900 814.290 ;
        RECT 1195.700 766.205 1195.840 813.970 ;
        RECT 1194.710 765.835 1194.990 766.205 ;
        RECT 1195.630 765.835 1195.910 766.205 ;
        RECT 1194.720 765.690 1194.980 765.835 ;
        RECT 1194.720 735.770 1194.980 736.090 ;
        RECT 1194.780 669.450 1194.920 735.770 ;
        RECT 1193.340 669.130 1193.600 669.450 ;
        RECT 1194.720 669.130 1194.980 669.450 ;
        RECT 1193.400 621.365 1193.540 669.130 ;
        RECT 1193.330 620.995 1193.610 621.365 ;
        RECT 1194.710 620.995 1194.990 621.365 ;
        RECT 1194.780 614.450 1194.920 620.995 ;
        RECT 1194.320 614.310 1194.920 614.450 ;
        RECT 1194.320 607.230 1194.460 614.310 ;
        RECT 1194.260 606.910 1194.520 607.230 ;
        RECT 1194.260 576.650 1194.520 576.970 ;
        RECT 1194.320 531.750 1194.460 576.650 ;
        RECT 1194.260 531.430 1194.520 531.750 ;
        RECT 1194.260 530.750 1194.520 531.070 ;
        RECT 1194.320 475.990 1194.460 530.750 ;
        RECT 1194.260 475.670 1194.520 475.990 ;
        RECT 1194.720 475.330 1194.980 475.650 ;
        RECT 1194.780 400.930 1194.920 475.330 ;
        RECT 1194.320 400.790 1194.920 400.930 ;
        RECT 1194.320 373.050 1194.460 400.790 ;
        RECT 1194.320 372.910 1194.920 373.050 ;
        RECT 1194.780 372.630 1194.920 372.910 ;
        RECT 1194.720 372.310 1194.980 372.630 ;
        RECT 1194.720 324.370 1194.980 324.690 ;
        RECT 1194.780 276.070 1194.920 324.370 ;
        RECT 1194.720 275.750 1194.980 276.070 ;
        RECT 1194.720 227.810 1194.980 228.130 ;
        RECT 1194.780 193.450 1194.920 227.810 ;
        RECT 1194.720 193.130 1194.980 193.450 ;
        RECT 1194.260 192.790 1194.520 193.110 ;
        RECT 1194.320 145.170 1194.460 192.790 ;
        RECT 1194.260 144.850 1194.520 145.170 ;
        RECT 1194.720 144.850 1194.980 145.170 ;
        RECT 1194.780 107.430 1194.920 144.850 ;
        RECT 1194.720 107.110 1194.980 107.430 ;
        RECT 1194.260 82.970 1194.520 83.290 ;
        RECT 448.600 15.990 448.860 16.310 ;
        RECT 448.660 2.400 448.800 15.990 ;
        RECT 1194.320 15.970 1194.460 82.970 ;
        RECT 1194.260 15.650 1194.520 15.970 ;
        RECT 448.450 -4.800 449.010 2.400 ;
      LAYER via2 ;
        RECT 1194.250 1097.040 1194.530 1097.320 ;
        RECT 1195.630 1097.040 1195.910 1097.320 ;
        RECT 1194.710 765.880 1194.990 766.160 ;
        RECT 1195.630 765.880 1195.910 766.160 ;
        RECT 1193.330 621.040 1193.610 621.320 ;
        RECT 1194.710 621.040 1194.990 621.320 ;
      LAYER met3 ;
        RECT 1194.225 1097.330 1194.555 1097.345 ;
        RECT 1195.605 1097.330 1195.935 1097.345 ;
        RECT 1194.225 1097.030 1195.935 1097.330 ;
        RECT 1194.225 1097.015 1194.555 1097.030 ;
        RECT 1195.605 1097.015 1195.935 1097.030 ;
        RECT 1194.685 766.170 1195.015 766.185 ;
        RECT 1195.605 766.170 1195.935 766.185 ;
        RECT 1194.685 765.870 1195.935 766.170 ;
        RECT 1194.685 765.855 1195.015 765.870 ;
        RECT 1195.605 765.855 1195.935 765.870 ;
        RECT 1193.305 621.330 1193.635 621.345 ;
        RECT 1194.685 621.330 1195.015 621.345 ;
        RECT 1193.305 621.030 1195.015 621.330 ;
        RECT 1193.305 621.015 1193.635 621.030 ;
        RECT 1194.685 621.015 1195.015 621.030 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 466.510 15.880 466.830 15.940 ;
        RECT 466.510 15.740 1166.860 15.880 ;
        RECT 466.510 15.680 466.830 15.740 ;
        RECT 1166.720 15.540 1166.860 15.740 ;
        RECT 1197.450 15.540 1197.770 15.600 ;
        RECT 1166.720 15.400 1197.770 15.540 ;
        RECT 1197.450 15.340 1197.770 15.400 ;
      LAYER via ;
        RECT 466.540 15.680 466.800 15.940 ;
        RECT 1197.480 15.340 1197.740 15.600 ;
      LAYER met2 ;
        RECT 1197.380 1700.340 1197.660 1704.000 ;
        RECT 1197.380 1700.000 1197.680 1700.340 ;
        RECT 466.540 15.650 466.800 15.970 ;
        RECT 466.600 2.400 466.740 15.650 ;
        RECT 1197.540 15.630 1197.680 1700.000 ;
        RECT 1197.480 15.310 1197.740 15.630 ;
        RECT 466.390 -4.800 466.950 2.400 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 541.580 15.400 1166.400 15.540 ;
        RECT 484.450 15.200 484.770 15.260 ;
        RECT 541.580 15.200 541.720 15.400 ;
        RECT 484.450 15.060 541.720 15.200 ;
        RECT 1166.260 15.200 1166.400 15.400 ;
        RECT 1199.290 15.200 1199.610 15.260 ;
        RECT 1166.260 15.060 1199.610 15.200 ;
        RECT 484.450 15.000 484.770 15.060 ;
        RECT 1199.290 15.000 1199.610 15.060 ;
      LAYER via ;
        RECT 484.480 15.000 484.740 15.260 ;
        RECT 1199.320 15.000 1199.580 15.260 ;
      LAYER met2 ;
        RECT 1199.220 1700.340 1199.500 1704.000 ;
        RECT 1199.220 1700.000 1199.520 1700.340 ;
        RECT 1199.380 15.290 1199.520 1700.000 ;
        RECT 484.480 14.970 484.740 15.290 ;
        RECT 1199.320 14.970 1199.580 15.290 ;
        RECT 484.540 2.400 484.680 14.970 ;
        RECT 484.330 -4.800 484.890 2.400 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1179.585 1689.205 1179.755 1690.395 ;
      LAYER mcon ;
        RECT 1179.585 1690.225 1179.755 1690.395 ;
      LAYER met1 ;
        RECT 1179.525 1690.380 1179.815 1690.425 ;
        RECT 1201.130 1690.380 1201.450 1690.440 ;
        RECT 1179.525 1690.240 1201.450 1690.380 ;
        RECT 1179.525 1690.195 1179.815 1690.240 ;
        RECT 1201.130 1690.180 1201.450 1690.240 ;
        RECT 503.310 1689.360 503.630 1689.420 ;
        RECT 1179.525 1689.360 1179.815 1689.405 ;
        RECT 503.310 1689.220 1179.815 1689.360 ;
        RECT 503.310 1689.160 503.630 1689.220 ;
        RECT 1179.525 1689.175 1179.815 1689.220 ;
      LAYER via ;
        RECT 1201.160 1690.180 1201.420 1690.440 ;
        RECT 503.340 1689.160 503.600 1689.420 ;
      LAYER met2 ;
        RECT 1201.060 1700.340 1201.340 1704.000 ;
        RECT 1201.060 1700.000 1201.360 1700.340 ;
        RECT 1201.220 1690.470 1201.360 1700.000 ;
        RECT 1201.160 1690.150 1201.420 1690.470 ;
        RECT 503.340 1689.130 503.600 1689.450 ;
        RECT 503.400 3.130 503.540 1689.130 ;
        RECT 502.480 2.990 503.540 3.130 ;
        RECT 502.480 2.400 502.620 2.990 ;
        RECT 502.270 -4.800 502.830 2.400 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1203.430 1678.140 1203.750 1678.200 ;
        RECT 1204.810 1678.140 1205.130 1678.200 ;
        RECT 1203.430 1678.000 1205.130 1678.140 ;
        RECT 1203.430 1677.940 1203.750 1678.000 ;
        RECT 1204.810 1677.940 1205.130 1678.000 ;
        RECT 542.040 15.060 1165.940 15.200 ;
        RECT 519.870 14.520 520.190 14.580 ;
        RECT 542.040 14.520 542.180 15.060 ;
        RECT 1165.800 14.860 1165.940 15.060 ;
        RECT 1204.810 14.860 1205.130 14.920 ;
        RECT 1165.800 14.720 1205.130 14.860 ;
        RECT 1204.810 14.660 1205.130 14.720 ;
        RECT 519.870 14.380 542.180 14.520 ;
        RECT 519.870 14.320 520.190 14.380 ;
      LAYER via ;
        RECT 1203.460 1677.940 1203.720 1678.200 ;
        RECT 1204.840 1677.940 1205.100 1678.200 ;
        RECT 519.900 14.320 520.160 14.580 ;
        RECT 1204.840 14.660 1205.100 14.920 ;
      LAYER met2 ;
        RECT 1202.900 1700.410 1203.180 1704.000 ;
        RECT 1202.900 1700.270 1203.660 1700.410 ;
        RECT 1202.900 1700.000 1203.180 1700.270 ;
        RECT 1203.520 1678.230 1203.660 1700.270 ;
        RECT 1203.460 1677.910 1203.720 1678.230 ;
        RECT 1204.840 1677.910 1205.100 1678.230 ;
        RECT 1204.900 14.950 1205.040 1677.910 ;
        RECT 1204.840 14.630 1205.100 14.950 ;
        RECT 519.900 14.290 520.160 14.610 ;
        RECT 519.960 2.400 520.100 14.290 ;
        RECT 519.750 -4.800 520.310 2.400 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1178.205 1688.525 1178.375 1690.055 ;
      LAYER mcon ;
        RECT 1178.205 1689.885 1178.375 1690.055 ;
      LAYER met1 ;
        RECT 537.810 1690.040 538.130 1690.100 ;
        RECT 1178.145 1690.040 1178.435 1690.085 ;
        RECT 537.810 1689.900 1178.435 1690.040 ;
        RECT 537.810 1689.840 538.130 1689.900 ;
        RECT 1178.145 1689.855 1178.435 1689.900 ;
        RECT 1178.145 1688.680 1178.435 1688.725 ;
        RECT 1204.810 1688.680 1205.130 1688.740 ;
        RECT 1178.145 1688.540 1205.130 1688.680 ;
        RECT 1178.145 1688.495 1178.435 1688.540 ;
        RECT 1204.810 1688.480 1205.130 1688.540 ;
      LAYER via ;
        RECT 537.840 1689.840 538.100 1690.100 ;
        RECT 1204.840 1688.480 1205.100 1688.740 ;
      LAYER met2 ;
        RECT 1204.740 1700.340 1205.020 1704.000 ;
        RECT 1204.740 1700.000 1205.040 1700.340 ;
        RECT 537.840 1689.810 538.100 1690.130 ;
        RECT 537.900 2.400 538.040 1689.810 ;
        RECT 1204.900 1688.770 1205.040 1700.000 ;
        RECT 1204.840 1688.450 1205.100 1688.770 ;
        RECT 537.690 -4.800 538.250 2.400 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1205.805 1304.325 1205.975 1352.435 ;
        RECT 1205.805 766.105 1205.975 814.215 ;
        RECT 1205.345 572.645 1205.515 620.755 ;
        RECT 1205.805 276.165 1205.975 324.275 ;
        RECT 1206.265 179.605 1206.435 227.715 ;
        RECT 1165.325 14.705 1165.495 18.615 ;
      LAYER mcon ;
        RECT 1205.805 1352.265 1205.975 1352.435 ;
        RECT 1205.805 814.045 1205.975 814.215 ;
        RECT 1205.345 620.585 1205.515 620.755 ;
        RECT 1205.805 324.105 1205.975 324.275 ;
        RECT 1206.265 227.545 1206.435 227.715 ;
        RECT 1165.325 18.445 1165.495 18.615 ;
      LAYER met1 ;
        RECT 1205.270 1666.580 1205.590 1666.640 ;
        RECT 1206.650 1666.580 1206.970 1666.640 ;
        RECT 1205.270 1666.440 1206.970 1666.580 ;
        RECT 1205.270 1666.380 1205.590 1666.440 ;
        RECT 1206.650 1666.380 1206.970 1666.440 ;
        RECT 1205.270 1448.980 1205.590 1449.040 ;
        RECT 1205.730 1448.980 1206.050 1449.040 ;
        RECT 1205.270 1448.840 1206.050 1448.980 ;
        RECT 1205.270 1448.780 1205.590 1448.840 ;
        RECT 1205.730 1448.780 1206.050 1448.840 ;
        RECT 1205.730 1352.420 1206.050 1352.480 ;
        RECT 1205.535 1352.280 1206.050 1352.420 ;
        RECT 1205.730 1352.220 1206.050 1352.280 ;
        RECT 1205.730 1304.480 1206.050 1304.540 ;
        RECT 1205.535 1304.340 1206.050 1304.480 ;
        RECT 1205.730 1304.280 1206.050 1304.340 ;
        RECT 1204.350 1235.120 1204.670 1235.180 ;
        RECT 1205.730 1235.120 1206.050 1235.180 ;
        RECT 1204.350 1234.980 1206.050 1235.120 ;
        RECT 1204.350 1234.920 1204.670 1234.980 ;
        RECT 1205.730 1234.920 1206.050 1234.980 ;
        RECT 1204.350 1145.360 1204.670 1145.420 ;
        RECT 1205.730 1145.360 1206.050 1145.420 ;
        RECT 1204.350 1145.220 1206.050 1145.360 ;
        RECT 1204.350 1145.160 1204.670 1145.220 ;
        RECT 1205.730 1145.160 1206.050 1145.220 ;
        RECT 1205.730 1007.320 1206.050 1007.380 ;
        RECT 1206.650 1007.320 1206.970 1007.380 ;
        RECT 1205.730 1007.180 1206.970 1007.320 ;
        RECT 1205.730 1007.120 1206.050 1007.180 ;
        RECT 1206.650 1007.120 1206.970 1007.180 ;
        RECT 1205.730 910.760 1206.050 910.820 ;
        RECT 1206.650 910.760 1206.970 910.820 ;
        RECT 1205.730 910.620 1206.970 910.760 ;
        RECT 1205.730 910.560 1206.050 910.620 ;
        RECT 1206.650 910.560 1206.970 910.620 ;
        RECT 1205.730 814.200 1206.050 814.260 ;
        RECT 1205.535 814.060 1206.050 814.200 ;
        RECT 1205.730 814.000 1206.050 814.060 ;
        RECT 1205.730 766.260 1206.050 766.320 ;
        RECT 1205.535 766.120 1206.050 766.260 ;
        RECT 1205.730 766.060 1206.050 766.120 ;
        RECT 1205.270 620.740 1205.590 620.800 ;
        RECT 1205.075 620.600 1205.590 620.740 ;
        RECT 1205.270 620.540 1205.590 620.600 ;
        RECT 1205.285 572.800 1205.575 572.845 ;
        RECT 1205.730 572.800 1206.050 572.860 ;
        RECT 1205.285 572.660 1206.050 572.800 ;
        RECT 1205.285 572.615 1205.575 572.660 ;
        RECT 1205.730 572.600 1206.050 572.660 ;
        RECT 1205.730 324.260 1206.050 324.320 ;
        RECT 1205.535 324.120 1206.050 324.260 ;
        RECT 1205.730 324.060 1206.050 324.120 ;
        RECT 1205.730 276.320 1206.050 276.380 ;
        RECT 1205.535 276.180 1206.050 276.320 ;
        RECT 1205.730 276.120 1206.050 276.180 ;
        RECT 1205.730 255.380 1206.050 255.640 ;
        RECT 1205.820 254.900 1205.960 255.380 ;
        RECT 1206.190 254.900 1206.510 254.960 ;
        RECT 1205.820 254.760 1206.510 254.900 ;
        RECT 1206.190 254.700 1206.510 254.760 ;
        RECT 1206.190 227.700 1206.510 227.760 ;
        RECT 1205.995 227.560 1206.510 227.700 ;
        RECT 1206.190 227.500 1206.510 227.560 ;
        RECT 1206.190 179.760 1206.510 179.820 ;
        RECT 1205.995 179.620 1206.510 179.760 ;
        RECT 1206.190 179.560 1206.510 179.620 ;
        RECT 1204.350 90.000 1204.670 90.060 ;
        RECT 1205.270 90.000 1205.590 90.060 ;
        RECT 1204.350 89.860 1205.590 90.000 ;
        RECT 1204.350 89.800 1204.670 89.860 ;
        RECT 1205.270 89.800 1205.590 89.860 ;
        RECT 1165.265 18.600 1165.555 18.645 ;
        RECT 1205.270 18.600 1205.590 18.660 ;
        RECT 1165.265 18.460 1205.590 18.600 ;
        RECT 1165.265 18.415 1165.555 18.460 ;
        RECT 1205.270 18.400 1205.590 18.460 ;
        RECT 1165.265 14.860 1165.555 14.905 ;
        RECT 572.860 14.720 1165.555 14.860 ;
        RECT 555.750 14.520 556.070 14.580 ;
        RECT 572.860 14.520 573.000 14.720 ;
        RECT 1165.265 14.675 1165.555 14.720 ;
        RECT 555.750 14.380 573.000 14.520 ;
        RECT 555.750 14.320 556.070 14.380 ;
      LAYER via ;
        RECT 1205.300 1666.380 1205.560 1666.640 ;
        RECT 1206.680 1666.380 1206.940 1666.640 ;
        RECT 1205.300 1448.780 1205.560 1449.040 ;
        RECT 1205.760 1448.780 1206.020 1449.040 ;
        RECT 1205.760 1352.220 1206.020 1352.480 ;
        RECT 1205.760 1304.280 1206.020 1304.540 ;
        RECT 1204.380 1234.920 1204.640 1235.180 ;
        RECT 1205.760 1234.920 1206.020 1235.180 ;
        RECT 1204.380 1145.160 1204.640 1145.420 ;
        RECT 1205.760 1145.160 1206.020 1145.420 ;
        RECT 1205.760 1007.120 1206.020 1007.380 ;
        RECT 1206.680 1007.120 1206.940 1007.380 ;
        RECT 1205.760 910.560 1206.020 910.820 ;
        RECT 1206.680 910.560 1206.940 910.820 ;
        RECT 1205.760 814.000 1206.020 814.260 ;
        RECT 1205.760 766.060 1206.020 766.320 ;
        RECT 1205.300 620.540 1205.560 620.800 ;
        RECT 1205.760 572.600 1206.020 572.860 ;
        RECT 1205.760 324.060 1206.020 324.320 ;
        RECT 1205.760 276.120 1206.020 276.380 ;
        RECT 1205.760 255.380 1206.020 255.640 ;
        RECT 1206.220 254.700 1206.480 254.960 ;
        RECT 1206.220 227.500 1206.480 227.760 ;
        RECT 1206.220 179.560 1206.480 179.820 ;
        RECT 1204.380 89.800 1204.640 90.060 ;
        RECT 1205.300 89.800 1205.560 90.060 ;
        RECT 1205.300 18.400 1205.560 18.660 ;
        RECT 555.780 14.320 556.040 14.580 ;
      LAYER met2 ;
        RECT 1206.580 1700.340 1206.860 1704.000 ;
        RECT 1206.580 1700.000 1206.880 1700.340 ;
        RECT 1206.740 1666.670 1206.880 1700.000 ;
        RECT 1205.300 1666.350 1205.560 1666.670 ;
        RECT 1206.680 1666.350 1206.940 1666.670 ;
        RECT 1205.360 1510.010 1205.500 1666.350 ;
        RECT 1205.360 1509.870 1205.960 1510.010 ;
        RECT 1205.820 1449.070 1205.960 1509.870 ;
        RECT 1205.300 1448.750 1205.560 1449.070 ;
        RECT 1205.760 1448.750 1206.020 1449.070 ;
        RECT 1205.360 1425.010 1205.500 1448.750 ;
        RECT 1205.360 1424.870 1205.960 1425.010 ;
        RECT 1205.820 1366.530 1205.960 1424.870 ;
        RECT 1205.360 1366.390 1205.960 1366.530 ;
        RECT 1205.360 1365.850 1205.500 1366.390 ;
        RECT 1205.360 1365.710 1205.960 1365.850 ;
        RECT 1205.820 1352.510 1205.960 1365.710 ;
        RECT 1205.760 1352.190 1206.020 1352.510 ;
        RECT 1205.760 1304.250 1206.020 1304.570 ;
        RECT 1205.820 1269.970 1205.960 1304.250 ;
        RECT 1205.360 1269.830 1205.960 1269.970 ;
        RECT 1205.360 1269.290 1205.500 1269.830 ;
        RECT 1205.360 1269.150 1205.960 1269.290 ;
        RECT 1205.820 1235.210 1205.960 1269.150 ;
        RECT 1204.380 1234.890 1204.640 1235.210 ;
        RECT 1205.760 1234.890 1206.020 1235.210 ;
        RECT 1204.440 1187.125 1204.580 1234.890 ;
        RECT 1204.370 1186.755 1204.650 1187.125 ;
        RECT 1205.290 1186.755 1205.570 1187.125 ;
        RECT 1205.360 1152.330 1205.500 1186.755 ;
        RECT 1205.360 1152.190 1205.960 1152.330 ;
        RECT 1205.820 1145.450 1205.960 1152.190 ;
        RECT 1204.380 1145.130 1204.640 1145.450 ;
        RECT 1205.760 1145.130 1206.020 1145.450 ;
        RECT 1204.440 1097.365 1204.580 1145.130 ;
        RECT 1204.370 1096.995 1204.650 1097.365 ;
        RECT 1205.290 1096.995 1205.570 1097.365 ;
        RECT 1205.360 1076.850 1205.500 1096.995 ;
        RECT 1205.360 1076.710 1205.960 1076.850 ;
        RECT 1205.820 1007.410 1205.960 1076.710 ;
        RECT 1205.760 1007.090 1206.020 1007.410 ;
        RECT 1206.680 1007.090 1206.940 1007.410 ;
        RECT 1206.740 959.325 1206.880 1007.090 ;
        RECT 1205.750 958.955 1206.030 959.325 ;
        RECT 1206.670 958.955 1206.950 959.325 ;
        RECT 1205.820 910.850 1205.960 958.955 ;
        RECT 1205.760 910.530 1206.020 910.850 ;
        RECT 1206.680 910.530 1206.940 910.850 ;
        RECT 1206.740 862.765 1206.880 910.530 ;
        RECT 1205.750 862.395 1206.030 862.765 ;
        RECT 1206.670 862.395 1206.950 862.765 ;
        RECT 1205.820 814.290 1205.960 862.395 ;
        RECT 1205.760 813.970 1206.020 814.290 ;
        RECT 1205.760 766.030 1206.020 766.350 ;
        RECT 1205.820 628.845 1205.960 766.030 ;
        RECT 1205.750 628.475 1206.030 628.845 ;
        RECT 1205.290 627.795 1205.570 628.165 ;
        RECT 1205.360 620.830 1205.500 627.795 ;
        RECT 1205.300 620.510 1205.560 620.830 ;
        RECT 1205.760 572.570 1206.020 572.890 ;
        RECT 1205.820 324.350 1205.960 572.570 ;
        RECT 1205.760 324.030 1206.020 324.350 ;
        RECT 1205.760 276.090 1206.020 276.410 ;
        RECT 1205.820 255.670 1205.960 276.090 ;
        RECT 1205.760 255.350 1206.020 255.670 ;
        RECT 1206.220 254.670 1206.480 254.990 ;
        RECT 1206.280 227.790 1206.420 254.670 ;
        RECT 1206.220 227.470 1206.480 227.790 ;
        RECT 1206.220 179.530 1206.480 179.850 ;
        RECT 1206.280 145.250 1206.420 179.530 ;
        RECT 1206.280 145.110 1206.880 145.250 ;
        RECT 1206.740 144.570 1206.880 145.110 ;
        RECT 1205.360 144.430 1206.880 144.570 ;
        RECT 1205.360 137.885 1205.500 144.430 ;
        RECT 1204.370 137.515 1204.650 137.885 ;
        RECT 1205.290 137.515 1205.570 137.885 ;
        RECT 1204.440 90.090 1204.580 137.515 ;
        RECT 1204.380 89.770 1204.640 90.090 ;
        RECT 1205.300 89.770 1205.560 90.090 ;
        RECT 1205.360 18.690 1205.500 89.770 ;
        RECT 1205.300 18.370 1205.560 18.690 ;
        RECT 555.780 14.290 556.040 14.610 ;
        RECT 555.840 2.400 555.980 14.290 ;
        RECT 555.630 -4.800 556.190 2.400 ;
      LAYER via2 ;
        RECT 1204.370 1186.800 1204.650 1187.080 ;
        RECT 1205.290 1186.800 1205.570 1187.080 ;
        RECT 1204.370 1097.040 1204.650 1097.320 ;
        RECT 1205.290 1097.040 1205.570 1097.320 ;
        RECT 1205.750 959.000 1206.030 959.280 ;
        RECT 1206.670 959.000 1206.950 959.280 ;
        RECT 1205.750 862.440 1206.030 862.720 ;
        RECT 1206.670 862.440 1206.950 862.720 ;
        RECT 1205.750 628.520 1206.030 628.800 ;
        RECT 1205.290 627.840 1205.570 628.120 ;
        RECT 1204.370 137.560 1204.650 137.840 ;
        RECT 1205.290 137.560 1205.570 137.840 ;
      LAYER met3 ;
        RECT 1204.345 1187.090 1204.675 1187.105 ;
        RECT 1205.265 1187.090 1205.595 1187.105 ;
        RECT 1204.345 1186.790 1205.595 1187.090 ;
        RECT 1204.345 1186.775 1204.675 1186.790 ;
        RECT 1205.265 1186.775 1205.595 1186.790 ;
        RECT 1204.345 1097.330 1204.675 1097.345 ;
        RECT 1205.265 1097.330 1205.595 1097.345 ;
        RECT 1204.345 1097.030 1205.595 1097.330 ;
        RECT 1204.345 1097.015 1204.675 1097.030 ;
        RECT 1205.265 1097.015 1205.595 1097.030 ;
        RECT 1205.725 959.290 1206.055 959.305 ;
        RECT 1206.645 959.290 1206.975 959.305 ;
        RECT 1205.725 958.990 1206.975 959.290 ;
        RECT 1205.725 958.975 1206.055 958.990 ;
        RECT 1206.645 958.975 1206.975 958.990 ;
        RECT 1205.725 862.730 1206.055 862.745 ;
        RECT 1206.645 862.730 1206.975 862.745 ;
        RECT 1205.725 862.430 1206.975 862.730 ;
        RECT 1205.725 862.415 1206.055 862.430 ;
        RECT 1206.645 862.415 1206.975 862.430 ;
        RECT 1205.725 628.810 1206.055 628.825 ;
        RECT 1205.510 628.495 1206.055 628.810 ;
        RECT 1205.510 628.145 1205.810 628.495 ;
        RECT 1205.265 627.830 1205.810 628.145 ;
        RECT 1205.265 627.815 1205.595 627.830 ;
        RECT 1204.345 137.850 1204.675 137.865 ;
        RECT 1205.265 137.850 1205.595 137.865 ;
        RECT 1204.345 137.550 1205.595 137.850 ;
        RECT 1204.345 137.535 1204.675 137.550 ;
        RECT 1205.265 137.535 1205.595 137.550 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1208.490 1690.040 1208.810 1690.100 ;
        RECT 1179.600 1689.900 1208.810 1690.040 ;
        RECT 579.210 1689.700 579.530 1689.760 ;
        RECT 1179.600 1689.700 1179.740 1689.900 ;
        RECT 1208.490 1689.840 1208.810 1689.900 ;
        RECT 579.210 1689.560 1179.740 1689.700 ;
        RECT 579.210 1689.500 579.530 1689.560 ;
        RECT 573.690 14.520 574.010 14.580 ;
        RECT 579.210 14.520 579.530 14.580 ;
        RECT 573.690 14.380 579.530 14.520 ;
        RECT 573.690 14.320 574.010 14.380 ;
        RECT 579.210 14.320 579.530 14.380 ;
      LAYER via ;
        RECT 579.240 1689.500 579.500 1689.760 ;
        RECT 1208.520 1689.840 1208.780 1690.100 ;
        RECT 573.720 14.320 573.980 14.580 ;
        RECT 579.240 14.320 579.500 14.580 ;
      LAYER met2 ;
        RECT 1208.420 1700.340 1208.700 1704.000 ;
        RECT 1208.420 1700.000 1208.720 1700.340 ;
        RECT 1208.580 1690.130 1208.720 1700.000 ;
        RECT 1208.520 1689.810 1208.780 1690.130 ;
        RECT 579.240 1689.470 579.500 1689.790 ;
        RECT 579.300 14.610 579.440 1689.470 ;
        RECT 573.720 14.290 573.980 14.610 ;
        RECT 579.240 14.290 579.500 14.610 ;
        RECT 573.780 2.400 573.920 14.290 ;
        RECT 573.570 -4.800 574.130 2.400 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1210.330 14.520 1210.650 14.580 ;
        RECT 607.360 14.380 1210.650 14.520 ;
        RECT 591.170 14.180 591.490 14.240 ;
        RECT 607.360 14.180 607.500 14.380 ;
        RECT 1210.330 14.320 1210.650 14.380 ;
        RECT 591.170 14.040 607.500 14.180 ;
        RECT 591.170 13.980 591.490 14.040 ;
      LAYER via ;
        RECT 591.200 13.980 591.460 14.240 ;
        RECT 1210.360 14.320 1210.620 14.580 ;
      LAYER met2 ;
        RECT 1210.260 1700.340 1210.540 1704.000 ;
        RECT 1210.260 1700.000 1210.560 1700.340 ;
        RECT 1210.420 14.610 1210.560 1700.000 ;
        RECT 1210.360 14.290 1210.620 14.610 ;
        RECT 591.200 13.950 591.460 14.270 ;
        RECT 591.260 2.400 591.400 13.950 ;
        RECT 591.050 -4.800 591.610 2.400 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 161.990 1688.680 162.310 1688.740 ;
        RECT 1159.730 1688.680 1160.050 1688.740 ;
        RECT 161.990 1688.540 1160.050 1688.680 ;
        RECT 161.990 1688.480 162.310 1688.540 ;
        RECT 1159.730 1688.480 1160.050 1688.540 ;
        RECT 161.990 17.580 162.310 17.640 ;
        RECT 143.680 17.440 162.310 17.580 ;
        RECT 97.590 17.240 97.910 17.300 ;
        RECT 143.680 17.240 143.820 17.440 ;
        RECT 161.990 17.380 162.310 17.440 ;
        RECT 97.590 17.100 143.820 17.240 ;
        RECT 97.590 17.040 97.910 17.100 ;
      LAYER via ;
        RECT 162.020 1688.480 162.280 1688.740 ;
        RECT 1159.760 1688.480 1160.020 1688.740 ;
        RECT 97.620 17.040 97.880 17.300 ;
        RECT 162.020 17.380 162.280 17.640 ;
      LAYER met2 ;
        RECT 1159.660 1700.340 1159.940 1704.000 ;
        RECT 1159.660 1700.000 1159.960 1700.340 ;
        RECT 1159.820 1688.770 1159.960 1700.000 ;
        RECT 162.020 1688.450 162.280 1688.770 ;
        RECT 1159.760 1688.450 1160.020 1688.770 ;
        RECT 162.080 17.670 162.220 1688.450 ;
        RECT 162.020 17.350 162.280 17.670 ;
        RECT 97.620 17.010 97.880 17.330 ;
        RECT 97.680 2.400 97.820 17.010 ;
        RECT 97.470 -4.800 98.030 2.400 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1210.790 1678.140 1211.110 1678.200 ;
        RECT 1212.170 1678.140 1212.490 1678.200 ;
        RECT 1210.790 1678.000 1212.490 1678.140 ;
        RECT 1210.790 1677.940 1211.110 1678.000 ;
        RECT 1212.170 1677.940 1212.490 1678.000 ;
        RECT 609.110 14.180 609.430 14.240 ;
        RECT 1210.790 14.180 1211.110 14.240 ;
        RECT 609.110 14.040 1211.110 14.180 ;
        RECT 609.110 13.980 609.430 14.040 ;
        RECT 1210.790 13.980 1211.110 14.040 ;
      LAYER via ;
        RECT 1210.820 1677.940 1211.080 1678.200 ;
        RECT 1212.200 1677.940 1212.460 1678.200 ;
        RECT 609.140 13.980 609.400 14.240 ;
        RECT 1210.820 13.980 1211.080 14.240 ;
      LAYER met2 ;
        RECT 1212.100 1700.340 1212.380 1704.000 ;
        RECT 1212.100 1700.000 1212.400 1700.340 ;
        RECT 1212.260 1678.230 1212.400 1700.000 ;
        RECT 1210.820 1677.910 1211.080 1678.230 ;
        RECT 1212.200 1677.910 1212.460 1678.230 ;
        RECT 1210.880 14.270 1211.020 1677.910 ;
        RECT 609.140 13.950 609.400 14.270 ;
        RECT 1210.820 13.950 1211.080 14.270 ;
        RECT 609.200 2.400 609.340 13.950 ;
        RECT 608.990 -4.800 609.550 2.400 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1178.665 1688.865 1178.835 1690.395 ;
      LAYER mcon ;
        RECT 1178.665 1690.225 1178.835 1690.395 ;
      LAYER met1 ;
        RECT 627.510 1690.380 627.830 1690.440 ;
        RECT 1178.605 1690.380 1178.895 1690.425 ;
        RECT 627.510 1690.240 1178.895 1690.380 ;
        RECT 627.510 1690.180 627.830 1690.240 ;
        RECT 1178.605 1690.195 1178.895 1690.240 ;
        RECT 1178.605 1689.020 1178.895 1689.065 ;
        RECT 1214.010 1689.020 1214.330 1689.080 ;
        RECT 1178.605 1688.880 1214.330 1689.020 ;
        RECT 1178.605 1688.835 1178.895 1688.880 ;
        RECT 1214.010 1688.820 1214.330 1688.880 ;
      LAYER via ;
        RECT 627.540 1690.180 627.800 1690.440 ;
        RECT 1214.040 1688.820 1214.300 1689.080 ;
      LAYER met2 ;
        RECT 1213.940 1700.340 1214.220 1704.000 ;
        RECT 1213.940 1700.000 1214.240 1700.340 ;
        RECT 627.540 1690.150 627.800 1690.470 ;
        RECT 627.600 17.410 627.740 1690.150 ;
        RECT 1214.100 1689.110 1214.240 1700.000 ;
        RECT 1214.040 1688.790 1214.300 1689.110 ;
        RECT 627.140 17.270 627.740 17.410 ;
        RECT 627.140 2.400 627.280 17.270 ;
        RECT 626.930 -4.800 627.490 2.400 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1161.960 1700.340 1162.240 1704.000 ;
        RECT 1161.960 1700.000 1162.260 1700.340 ;
        RECT 1162.120 1678.650 1162.260 1700.000 ;
        RECT 1162.120 1678.510 1164.100 1678.650 ;
        RECT 1163.960 18.885 1164.100 1678.510 ;
        RECT 121.530 18.515 121.810 18.885 ;
        RECT 1163.890 18.515 1164.170 18.885 ;
        RECT 121.600 2.400 121.740 18.515 ;
        RECT 121.390 -4.800 121.950 2.400 ;
      LAYER via2 ;
        RECT 121.530 18.560 121.810 18.840 ;
        RECT 1163.890 18.560 1164.170 18.840 ;
      LAYER met3 ;
        RECT 121.505 18.850 121.835 18.865 ;
        RECT 1163.865 18.850 1164.195 18.865 ;
        RECT 121.505 18.550 1164.195 18.850 ;
        RECT 121.505 18.535 121.835 18.550 ;
        RECT 1163.865 18.535 1164.195 18.550 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 175.790 1688.340 176.110 1688.400 ;
        RECT 1164.330 1688.340 1164.650 1688.400 ;
        RECT 175.790 1688.200 1164.650 1688.340 ;
        RECT 175.790 1688.140 176.110 1688.200 ;
        RECT 1164.330 1688.140 1164.650 1688.200 ;
        RECT 145.430 17.240 145.750 17.300 ;
        RECT 175.790 17.240 176.110 17.300 ;
        RECT 145.430 17.100 176.110 17.240 ;
        RECT 145.430 17.040 145.750 17.100 ;
        RECT 175.790 17.040 176.110 17.100 ;
      LAYER via ;
        RECT 175.820 1688.140 176.080 1688.400 ;
        RECT 1164.360 1688.140 1164.620 1688.400 ;
        RECT 145.460 17.040 145.720 17.300 ;
        RECT 175.820 17.040 176.080 17.300 ;
      LAYER met2 ;
        RECT 1164.260 1700.340 1164.540 1704.000 ;
        RECT 1164.260 1700.000 1164.560 1700.340 ;
        RECT 1164.420 1688.430 1164.560 1700.000 ;
        RECT 175.820 1688.110 176.080 1688.430 ;
        RECT 1164.360 1688.110 1164.620 1688.430 ;
        RECT 175.880 17.330 176.020 1688.110 ;
        RECT 145.460 17.010 145.720 17.330 ;
        RECT 175.820 17.010 176.080 17.330 ;
        RECT 145.520 2.400 145.660 17.010 ;
        RECT 145.310 -4.800 145.870 2.400 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1166.170 1684.600 1166.490 1684.660 ;
        RECT 1172.150 1684.600 1172.470 1684.660 ;
        RECT 1166.170 1684.460 1172.470 1684.600 ;
        RECT 1166.170 1684.400 1166.490 1684.460 ;
        RECT 1172.150 1684.400 1172.470 1684.460 ;
      LAYER via ;
        RECT 1166.200 1684.400 1166.460 1684.660 ;
        RECT 1172.180 1684.400 1172.440 1684.660 ;
      LAYER met2 ;
        RECT 1166.100 1700.340 1166.380 1704.000 ;
        RECT 1166.100 1700.000 1166.400 1700.340 ;
        RECT 1166.260 1684.690 1166.400 1700.000 ;
        RECT 1166.200 1684.370 1166.460 1684.690 ;
        RECT 1172.180 1684.370 1172.440 1684.690 ;
        RECT 1172.240 20.245 1172.380 1684.370 ;
        RECT 163.390 19.875 163.670 20.245 ;
        RECT 1172.170 19.875 1172.450 20.245 ;
        RECT 163.460 2.400 163.600 19.875 ;
        RECT 163.250 -4.800 163.810 2.400 ;
      LAYER via2 ;
        RECT 163.390 19.920 163.670 20.200 ;
        RECT 1172.170 19.920 1172.450 20.200 ;
      LAYER met3 ;
        RECT 163.365 20.210 163.695 20.225 ;
        RECT 1172.145 20.210 1172.475 20.225 ;
        RECT 163.365 19.910 1172.475 20.210 ;
        RECT 163.365 19.895 163.695 19.910 ;
        RECT 1172.145 19.895 1172.475 19.910 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 196.490 1689.020 196.810 1689.080 ;
        RECT 1168.010 1689.020 1168.330 1689.080 ;
        RECT 196.490 1688.880 1168.330 1689.020 ;
        RECT 196.490 1688.820 196.810 1688.880 ;
        RECT 1168.010 1688.820 1168.330 1688.880 ;
        RECT 180.850 16.220 181.170 16.280 ;
        RECT 196.490 16.220 196.810 16.280 ;
        RECT 180.850 16.080 196.810 16.220 ;
        RECT 180.850 16.020 181.170 16.080 ;
        RECT 196.490 16.020 196.810 16.080 ;
      LAYER via ;
        RECT 196.520 1688.820 196.780 1689.080 ;
        RECT 1168.040 1688.820 1168.300 1689.080 ;
        RECT 180.880 16.020 181.140 16.280 ;
        RECT 196.520 16.020 196.780 16.280 ;
      LAYER met2 ;
        RECT 1167.940 1700.340 1168.220 1704.000 ;
        RECT 1167.940 1700.000 1168.240 1700.340 ;
        RECT 1168.100 1689.110 1168.240 1700.000 ;
        RECT 196.520 1688.790 196.780 1689.110 ;
        RECT 1168.040 1688.790 1168.300 1689.110 ;
        RECT 196.580 16.310 196.720 1688.790 ;
        RECT 180.880 15.990 181.140 16.310 ;
        RECT 196.520 15.990 196.780 16.310 ;
        RECT 180.940 2.400 181.080 15.990 ;
        RECT 180.730 -4.800 181.290 2.400 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 198.790 17.240 199.110 17.300 ;
        RECT 198.790 17.100 1155.360 17.240 ;
        RECT 198.790 17.040 199.110 17.100 ;
        RECT 1155.220 16.560 1155.360 17.100 ;
        RECT 1170.770 16.560 1171.090 16.620 ;
        RECT 1155.220 16.420 1171.090 16.560 ;
        RECT 1170.770 16.360 1171.090 16.420 ;
      LAYER via ;
        RECT 198.820 17.040 199.080 17.300 ;
        RECT 1170.800 16.360 1171.060 16.620 ;
      LAYER met2 ;
        RECT 1169.780 1700.410 1170.060 1704.000 ;
        RECT 1169.780 1700.270 1170.540 1700.410 ;
        RECT 1169.780 1700.000 1170.060 1700.270 ;
        RECT 1170.400 1665.730 1170.540 1700.270 ;
        RECT 1170.400 1665.590 1171.000 1665.730 ;
        RECT 198.820 17.010 199.080 17.330 ;
        RECT 198.880 2.400 199.020 17.010 ;
        RECT 1170.860 16.650 1171.000 1665.590 ;
        RECT 1170.800 16.330 1171.060 16.650 ;
        RECT 198.670 -4.800 199.230 2.400 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met1 ;
        RECT 1170.310 1662.160 1170.630 1662.220 ;
        RECT 1171.690 1662.160 1172.010 1662.220 ;
        RECT 1170.310 1662.020 1172.010 1662.160 ;
        RECT 1170.310 1661.960 1170.630 1662.020 ;
        RECT 1171.690 1661.960 1172.010 1662.020 ;
        RECT 1170.310 17.920 1170.630 17.980 ;
        RECT 1156.140 17.780 1170.630 17.920 ;
        RECT 216.730 17.580 217.050 17.640 ;
        RECT 1156.140 17.580 1156.280 17.780 ;
        RECT 1170.310 17.720 1170.630 17.780 ;
        RECT 216.730 17.440 1156.280 17.580 ;
        RECT 216.730 17.380 217.050 17.440 ;
      LAYER via ;
        RECT 1170.340 1661.960 1170.600 1662.220 ;
        RECT 1171.720 1661.960 1171.980 1662.220 ;
        RECT 216.760 17.380 217.020 17.640 ;
        RECT 1170.340 17.720 1170.600 17.980 ;
      LAYER met2 ;
        RECT 1171.620 1700.340 1171.900 1704.000 ;
        RECT 1171.620 1700.000 1171.920 1700.340 ;
        RECT 1171.780 1662.250 1171.920 1700.000 ;
        RECT 1170.340 1661.930 1170.600 1662.250 ;
        RECT 1171.720 1661.930 1171.980 1662.250 ;
        RECT 1170.400 18.010 1170.540 1661.930 ;
        RECT 1170.340 17.690 1170.600 18.010 ;
        RECT 216.760 17.350 217.020 17.670 ;
        RECT 216.820 2.400 216.960 17.350 ;
        RECT 216.610 -4.800 217.170 2.400 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER li1 ;
        RECT 1155.665 16.745 1155.835 17.935 ;
      LAYER mcon ;
        RECT 1155.665 17.765 1155.835 17.935 ;
      LAYER met1 ;
        RECT 234.670 18.260 234.990 18.320 ;
        RECT 234.670 18.120 269.400 18.260 ;
        RECT 234.670 18.060 234.990 18.120 ;
        RECT 269.260 17.920 269.400 18.120 ;
        RECT 1155.605 17.920 1155.895 17.965 ;
        RECT 269.260 17.780 1155.895 17.920 ;
        RECT 1155.605 17.735 1155.895 17.780 ;
        RECT 1155.605 16.900 1155.895 16.945 ;
        RECT 1173.530 16.900 1173.850 16.960 ;
        RECT 1155.605 16.760 1173.850 16.900 ;
        RECT 1155.605 16.715 1155.895 16.760 ;
        RECT 1173.530 16.700 1173.850 16.760 ;
      LAYER via ;
        RECT 234.700 18.060 234.960 18.320 ;
        RECT 1173.560 16.700 1173.820 16.960 ;
      LAYER met2 ;
        RECT 1173.460 1700.410 1173.740 1704.000 ;
        RECT 1173.460 1700.270 1174.220 1700.410 ;
        RECT 1173.460 1700.000 1173.740 1700.270 ;
        RECT 1174.080 1666.410 1174.220 1700.270 ;
        RECT 1173.620 1666.270 1174.220 1666.410 ;
        RECT 234.700 18.030 234.960 18.350 ;
        RECT 234.760 2.400 234.900 18.030 ;
        RECT 1173.620 16.990 1173.760 1666.270 ;
        RECT 1173.560 16.670 1173.820 16.990 ;
        RECT 234.550 -4.800 235.110 2.400 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 79.190 1687.660 79.510 1687.720 ;
        RECT 1155.130 1687.660 1155.450 1687.720 ;
        RECT 79.190 1687.520 1155.450 1687.660 ;
        RECT 79.190 1687.460 79.510 1687.520 ;
        RECT 1155.130 1687.460 1155.450 1687.520 ;
        RECT 56.190 15.200 56.510 15.260 ;
        RECT 79.190 15.200 79.510 15.260 ;
        RECT 56.190 15.060 79.510 15.200 ;
        RECT 56.190 15.000 56.510 15.060 ;
        RECT 79.190 15.000 79.510 15.060 ;
      LAYER via ;
        RECT 79.220 1687.460 79.480 1687.720 ;
        RECT 1155.160 1687.460 1155.420 1687.720 ;
        RECT 56.220 15.000 56.480 15.260 ;
        RECT 79.220 15.000 79.480 15.260 ;
      LAYER met2 ;
        RECT 1155.060 1700.340 1155.340 1704.000 ;
        RECT 1155.060 1700.000 1155.360 1700.340 ;
        RECT 1155.220 1687.750 1155.360 1700.000 ;
        RECT 79.220 1687.430 79.480 1687.750 ;
        RECT 1155.160 1687.430 1155.420 1687.750 ;
        RECT 79.280 15.290 79.420 1687.430 ;
        RECT 56.220 14.970 56.480 15.290 ;
        RECT 79.220 14.970 79.480 15.290 ;
        RECT 56.280 2.400 56.420 14.970 ;
        RECT 56.070 -4.800 56.630 2.400 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1157.820 1700.410 1158.100 1704.000 ;
        RECT 1157.520 1700.270 1158.100 1700.410 ;
        RECT 1157.520 1658.930 1157.660 1700.270 ;
        RECT 1157.820 1700.000 1158.100 1700.270 ;
        RECT 1155.680 1658.790 1157.660 1658.930 ;
        RECT 1155.680 18.205 1155.820 1658.790 ;
        RECT 80.130 17.835 80.410 18.205 ;
        RECT 1155.610 17.835 1155.890 18.205 ;
        RECT 80.200 2.400 80.340 17.835 ;
        RECT 79.990 -4.800 80.550 2.400 ;
      LAYER via2 ;
        RECT 80.130 17.880 80.410 18.160 ;
        RECT 1155.610 17.880 1155.890 18.160 ;
      LAYER met3 ;
        RECT 80.105 18.170 80.435 18.185 ;
        RECT 1155.585 18.170 1155.915 18.185 ;
        RECT 80.105 17.870 1155.915 18.170 ;
        RECT 80.105 17.855 80.435 17.870 ;
        RECT 1155.585 17.855 1155.915 17.870 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 141.290 1688.000 141.610 1688.060 ;
        RECT 1160.190 1688.000 1160.510 1688.060 ;
        RECT 141.290 1687.860 1160.510 1688.000 ;
        RECT 141.290 1687.800 141.610 1687.860 ;
        RECT 1160.190 1687.800 1160.510 1687.860 ;
        RECT 103.570 20.640 103.890 20.700 ;
        RECT 141.290 20.640 141.610 20.700 ;
        RECT 103.570 20.500 141.610 20.640 ;
        RECT 103.570 20.440 103.890 20.500 ;
        RECT 141.290 20.440 141.610 20.500 ;
      LAYER via ;
        RECT 141.320 1687.800 141.580 1688.060 ;
        RECT 1160.220 1687.800 1160.480 1688.060 ;
        RECT 103.600 20.440 103.860 20.700 ;
        RECT 141.320 20.440 141.580 20.700 ;
      LAYER met2 ;
        RECT 1160.120 1700.340 1160.400 1704.000 ;
        RECT 1160.120 1700.000 1160.420 1700.340 ;
        RECT 1160.280 1688.090 1160.420 1700.000 ;
        RECT 141.320 1687.770 141.580 1688.090 ;
        RECT 1160.220 1687.770 1160.480 1688.090 ;
        RECT 141.380 20.730 141.520 1687.770 ;
        RECT 103.600 20.410 103.860 20.730 ;
        RECT 141.320 20.410 141.580 20.730 ;
        RECT 103.660 2.400 103.800 20.410 ;
        RECT 103.450 -4.800 104.010 2.400 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1162.420 1700.410 1162.700 1704.000 ;
        RECT 1162.420 1700.270 1163.180 1700.410 ;
        RECT 1162.420 1700.000 1162.700 1700.270 ;
        RECT 1163.040 1679.330 1163.180 1700.270 ;
        RECT 1163.040 1679.190 1165.020 1679.330 ;
        RECT 1164.880 19.565 1165.020 1679.190 ;
        RECT 127.510 19.195 127.790 19.565 ;
        RECT 1164.810 19.195 1165.090 19.565 ;
        RECT 127.580 2.400 127.720 19.195 ;
        RECT 127.370 -4.800 127.930 2.400 ;
      LAYER via2 ;
        RECT 127.510 19.240 127.790 19.520 ;
        RECT 1164.810 19.240 1165.090 19.520 ;
      LAYER met3 ;
        RECT 127.485 19.530 127.815 19.545 ;
        RECT 1164.785 19.530 1165.115 19.545 ;
        RECT 127.485 19.230 1165.115 19.530 ;
        RECT 127.485 19.215 127.815 19.230 ;
        RECT 1164.785 19.215 1165.115 19.230 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met1 ;
        RECT 51.590 1686.980 51.910 1687.040 ;
        RECT 1152.370 1686.980 1152.690 1687.040 ;
        RECT 51.590 1686.840 1152.690 1686.980 ;
        RECT 51.590 1686.780 51.910 1686.840 ;
        RECT 1152.370 1686.780 1152.690 1686.840 ;
        RECT 26.290 17.240 26.610 17.300 ;
        RECT 51.590 17.240 51.910 17.300 ;
        RECT 26.290 17.100 51.910 17.240 ;
        RECT 26.290 17.040 26.610 17.100 ;
        RECT 51.590 17.040 51.910 17.100 ;
      LAYER via ;
        RECT 51.620 1686.780 51.880 1687.040 ;
        RECT 1152.400 1686.780 1152.660 1687.040 ;
        RECT 26.320 17.040 26.580 17.300 ;
        RECT 51.620 17.040 51.880 17.300 ;
      LAYER met2 ;
        RECT 1152.300 1700.340 1152.580 1704.000 ;
        RECT 1152.300 1700.000 1152.600 1700.340 ;
        RECT 1152.460 1687.070 1152.600 1700.000 ;
        RECT 51.620 1686.750 51.880 1687.070 ;
        RECT 1152.400 1686.750 1152.660 1687.070 ;
        RECT 51.680 17.330 51.820 1686.750 ;
        RECT 26.320 17.010 26.580 17.330 ;
        RECT 51.620 17.010 51.880 17.330 ;
        RECT 26.380 2.400 26.520 17.010 ;
        RECT 26.170 -4.800 26.730 2.400 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1152.760 1700.340 1153.040 1704.000 ;
        RECT 1152.760 1700.000 1153.060 1700.340 ;
        RECT 1152.920 16.845 1153.060 1700.000 ;
        RECT 32.290 16.475 32.570 16.845 ;
        RECT 1152.850 16.475 1153.130 16.845 ;
        RECT 32.360 2.400 32.500 16.475 ;
        RECT 32.150 -4.800 32.710 2.400 ;
      LAYER via2 ;
        RECT 32.290 16.520 32.570 16.800 ;
        RECT 1152.850 16.520 1153.130 16.800 ;
      LAYER met3 ;
        RECT 32.265 16.810 32.595 16.825 ;
        RECT 1152.825 16.810 1153.155 16.825 ;
        RECT 32.265 16.510 1153.155 16.810 ;
        RECT 32.265 16.495 32.595 16.510 ;
        RECT 1152.825 16.495 1153.155 16.510 ;
    END
  END wbs_we_i
  PIN vccd1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -9.980 -4.620 -6.980 3524.300 ;
        RECT 4.020 -9.220 7.020 3528.900 ;
        RECT 184.020 -9.220 187.020 3528.900 ;
        RECT 364.020 -9.220 367.020 3528.900 ;
        RECT 544.020 -9.220 547.020 3528.900 ;
        RECT 724.020 -9.220 727.020 3528.900 ;
        RECT 904.020 -9.220 907.020 3528.900 ;
        RECT 1084.020 -9.220 1087.020 3528.900 ;
        RECT 1264.020 -9.220 1267.020 3528.900 ;
        RECT 1444.020 -9.220 1447.020 3528.900 ;
        RECT 1624.020 -9.220 1627.020 3528.900 ;
        RECT 1804.020 -9.220 1807.020 3528.900 ;
        RECT 1984.020 -9.220 1987.020 3528.900 ;
        RECT 2164.020 -9.220 2167.020 3528.900 ;
        RECT 2344.020 -9.220 2347.020 3528.900 ;
        RECT 2524.020 -9.220 2527.020 3528.900 ;
        RECT 2704.020 -9.220 2707.020 3528.900 ;
        RECT 2884.020 -9.220 2887.020 3528.900 ;
        RECT 2926.600 -4.620 2929.600 3524.300 ;
      LAYER via4 ;
        RECT -9.070 3523.010 -7.890 3524.190 ;
        RECT -9.070 3521.410 -7.890 3522.590 ;
        RECT -9.070 3431.090 -7.890 3432.270 ;
        RECT -9.070 3429.490 -7.890 3430.670 ;
        RECT -9.070 3251.090 -7.890 3252.270 ;
        RECT -9.070 3249.490 -7.890 3250.670 ;
        RECT -9.070 3071.090 -7.890 3072.270 ;
        RECT -9.070 3069.490 -7.890 3070.670 ;
        RECT -9.070 2891.090 -7.890 2892.270 ;
        RECT -9.070 2889.490 -7.890 2890.670 ;
        RECT -9.070 2711.090 -7.890 2712.270 ;
        RECT -9.070 2709.490 -7.890 2710.670 ;
        RECT -9.070 2531.090 -7.890 2532.270 ;
        RECT -9.070 2529.490 -7.890 2530.670 ;
        RECT -9.070 2351.090 -7.890 2352.270 ;
        RECT -9.070 2349.490 -7.890 2350.670 ;
        RECT -9.070 2171.090 -7.890 2172.270 ;
        RECT -9.070 2169.490 -7.890 2170.670 ;
        RECT -9.070 1991.090 -7.890 1992.270 ;
        RECT -9.070 1989.490 -7.890 1990.670 ;
        RECT -9.070 1811.090 -7.890 1812.270 ;
        RECT -9.070 1809.490 -7.890 1810.670 ;
        RECT -9.070 1631.090 -7.890 1632.270 ;
        RECT -9.070 1629.490 -7.890 1630.670 ;
        RECT -9.070 1451.090 -7.890 1452.270 ;
        RECT -9.070 1449.490 -7.890 1450.670 ;
        RECT -9.070 1271.090 -7.890 1272.270 ;
        RECT -9.070 1269.490 -7.890 1270.670 ;
        RECT -9.070 1091.090 -7.890 1092.270 ;
        RECT -9.070 1089.490 -7.890 1090.670 ;
        RECT -9.070 911.090 -7.890 912.270 ;
        RECT -9.070 909.490 -7.890 910.670 ;
        RECT -9.070 731.090 -7.890 732.270 ;
        RECT -9.070 729.490 -7.890 730.670 ;
        RECT -9.070 551.090 -7.890 552.270 ;
        RECT -9.070 549.490 -7.890 550.670 ;
        RECT -9.070 371.090 -7.890 372.270 ;
        RECT -9.070 369.490 -7.890 370.670 ;
        RECT -9.070 191.090 -7.890 192.270 ;
        RECT -9.070 189.490 -7.890 190.670 ;
        RECT -9.070 11.090 -7.890 12.270 ;
        RECT -9.070 9.490 -7.890 10.670 ;
        RECT -9.070 -2.910 -7.890 -1.730 ;
        RECT -9.070 -4.510 -7.890 -3.330 ;
        RECT 4.930 3523.010 6.110 3524.190 ;
        RECT 4.930 3521.410 6.110 3522.590 ;
        RECT 4.930 3431.090 6.110 3432.270 ;
        RECT 4.930 3429.490 6.110 3430.670 ;
        RECT 4.930 3251.090 6.110 3252.270 ;
        RECT 4.930 3249.490 6.110 3250.670 ;
        RECT 4.930 3071.090 6.110 3072.270 ;
        RECT 4.930 3069.490 6.110 3070.670 ;
        RECT 4.930 2891.090 6.110 2892.270 ;
        RECT 4.930 2889.490 6.110 2890.670 ;
        RECT 4.930 2711.090 6.110 2712.270 ;
        RECT 4.930 2709.490 6.110 2710.670 ;
        RECT 4.930 2531.090 6.110 2532.270 ;
        RECT 4.930 2529.490 6.110 2530.670 ;
        RECT 4.930 2351.090 6.110 2352.270 ;
        RECT 4.930 2349.490 6.110 2350.670 ;
        RECT 4.930 2171.090 6.110 2172.270 ;
        RECT 4.930 2169.490 6.110 2170.670 ;
        RECT 4.930 1991.090 6.110 1992.270 ;
        RECT 4.930 1989.490 6.110 1990.670 ;
        RECT 4.930 1811.090 6.110 1812.270 ;
        RECT 4.930 1809.490 6.110 1810.670 ;
        RECT 4.930 1631.090 6.110 1632.270 ;
        RECT 4.930 1629.490 6.110 1630.670 ;
        RECT 4.930 1451.090 6.110 1452.270 ;
        RECT 4.930 1449.490 6.110 1450.670 ;
        RECT 4.930 1271.090 6.110 1272.270 ;
        RECT 4.930 1269.490 6.110 1270.670 ;
        RECT 4.930 1091.090 6.110 1092.270 ;
        RECT 4.930 1089.490 6.110 1090.670 ;
        RECT 4.930 911.090 6.110 912.270 ;
        RECT 4.930 909.490 6.110 910.670 ;
        RECT 4.930 731.090 6.110 732.270 ;
        RECT 4.930 729.490 6.110 730.670 ;
        RECT 4.930 551.090 6.110 552.270 ;
        RECT 4.930 549.490 6.110 550.670 ;
        RECT 4.930 371.090 6.110 372.270 ;
        RECT 4.930 369.490 6.110 370.670 ;
        RECT 4.930 191.090 6.110 192.270 ;
        RECT 4.930 189.490 6.110 190.670 ;
        RECT 4.930 11.090 6.110 12.270 ;
        RECT 4.930 9.490 6.110 10.670 ;
        RECT 4.930 -2.910 6.110 -1.730 ;
        RECT 4.930 -4.510 6.110 -3.330 ;
        RECT 184.930 3523.010 186.110 3524.190 ;
        RECT 184.930 3521.410 186.110 3522.590 ;
        RECT 184.930 3431.090 186.110 3432.270 ;
        RECT 184.930 3429.490 186.110 3430.670 ;
        RECT 184.930 3251.090 186.110 3252.270 ;
        RECT 184.930 3249.490 186.110 3250.670 ;
        RECT 184.930 3071.090 186.110 3072.270 ;
        RECT 184.930 3069.490 186.110 3070.670 ;
        RECT 184.930 2891.090 186.110 2892.270 ;
        RECT 184.930 2889.490 186.110 2890.670 ;
        RECT 184.930 2711.090 186.110 2712.270 ;
        RECT 184.930 2709.490 186.110 2710.670 ;
        RECT 184.930 2531.090 186.110 2532.270 ;
        RECT 184.930 2529.490 186.110 2530.670 ;
        RECT 184.930 2351.090 186.110 2352.270 ;
        RECT 184.930 2349.490 186.110 2350.670 ;
        RECT 184.930 2171.090 186.110 2172.270 ;
        RECT 184.930 2169.490 186.110 2170.670 ;
        RECT 184.930 1991.090 186.110 1992.270 ;
        RECT 184.930 1989.490 186.110 1990.670 ;
        RECT 184.930 1811.090 186.110 1812.270 ;
        RECT 184.930 1809.490 186.110 1810.670 ;
        RECT 184.930 1631.090 186.110 1632.270 ;
        RECT 184.930 1629.490 186.110 1630.670 ;
        RECT 184.930 1451.090 186.110 1452.270 ;
        RECT 184.930 1449.490 186.110 1450.670 ;
        RECT 184.930 1271.090 186.110 1272.270 ;
        RECT 184.930 1269.490 186.110 1270.670 ;
        RECT 184.930 1091.090 186.110 1092.270 ;
        RECT 184.930 1089.490 186.110 1090.670 ;
        RECT 184.930 911.090 186.110 912.270 ;
        RECT 184.930 909.490 186.110 910.670 ;
        RECT 184.930 731.090 186.110 732.270 ;
        RECT 184.930 729.490 186.110 730.670 ;
        RECT 184.930 551.090 186.110 552.270 ;
        RECT 184.930 549.490 186.110 550.670 ;
        RECT 184.930 371.090 186.110 372.270 ;
        RECT 184.930 369.490 186.110 370.670 ;
        RECT 184.930 191.090 186.110 192.270 ;
        RECT 184.930 189.490 186.110 190.670 ;
        RECT 184.930 11.090 186.110 12.270 ;
        RECT 184.930 9.490 186.110 10.670 ;
        RECT 184.930 -2.910 186.110 -1.730 ;
        RECT 184.930 -4.510 186.110 -3.330 ;
        RECT 364.930 3523.010 366.110 3524.190 ;
        RECT 364.930 3521.410 366.110 3522.590 ;
        RECT 364.930 3431.090 366.110 3432.270 ;
        RECT 364.930 3429.490 366.110 3430.670 ;
        RECT 364.930 3251.090 366.110 3252.270 ;
        RECT 364.930 3249.490 366.110 3250.670 ;
        RECT 364.930 3071.090 366.110 3072.270 ;
        RECT 364.930 3069.490 366.110 3070.670 ;
        RECT 364.930 2891.090 366.110 2892.270 ;
        RECT 364.930 2889.490 366.110 2890.670 ;
        RECT 364.930 2711.090 366.110 2712.270 ;
        RECT 364.930 2709.490 366.110 2710.670 ;
        RECT 364.930 2531.090 366.110 2532.270 ;
        RECT 364.930 2529.490 366.110 2530.670 ;
        RECT 364.930 2351.090 366.110 2352.270 ;
        RECT 364.930 2349.490 366.110 2350.670 ;
        RECT 364.930 2171.090 366.110 2172.270 ;
        RECT 364.930 2169.490 366.110 2170.670 ;
        RECT 364.930 1991.090 366.110 1992.270 ;
        RECT 364.930 1989.490 366.110 1990.670 ;
        RECT 364.930 1811.090 366.110 1812.270 ;
        RECT 364.930 1809.490 366.110 1810.670 ;
        RECT 364.930 1631.090 366.110 1632.270 ;
        RECT 364.930 1629.490 366.110 1630.670 ;
        RECT 364.930 1451.090 366.110 1452.270 ;
        RECT 364.930 1449.490 366.110 1450.670 ;
        RECT 364.930 1271.090 366.110 1272.270 ;
        RECT 364.930 1269.490 366.110 1270.670 ;
        RECT 364.930 1091.090 366.110 1092.270 ;
        RECT 364.930 1089.490 366.110 1090.670 ;
        RECT 364.930 911.090 366.110 912.270 ;
        RECT 364.930 909.490 366.110 910.670 ;
        RECT 364.930 731.090 366.110 732.270 ;
        RECT 364.930 729.490 366.110 730.670 ;
        RECT 364.930 551.090 366.110 552.270 ;
        RECT 364.930 549.490 366.110 550.670 ;
        RECT 364.930 371.090 366.110 372.270 ;
        RECT 364.930 369.490 366.110 370.670 ;
        RECT 364.930 191.090 366.110 192.270 ;
        RECT 364.930 189.490 366.110 190.670 ;
        RECT 364.930 11.090 366.110 12.270 ;
        RECT 364.930 9.490 366.110 10.670 ;
        RECT 364.930 -2.910 366.110 -1.730 ;
        RECT 364.930 -4.510 366.110 -3.330 ;
        RECT 544.930 3523.010 546.110 3524.190 ;
        RECT 544.930 3521.410 546.110 3522.590 ;
        RECT 544.930 3431.090 546.110 3432.270 ;
        RECT 544.930 3429.490 546.110 3430.670 ;
        RECT 544.930 3251.090 546.110 3252.270 ;
        RECT 544.930 3249.490 546.110 3250.670 ;
        RECT 544.930 3071.090 546.110 3072.270 ;
        RECT 544.930 3069.490 546.110 3070.670 ;
        RECT 544.930 2891.090 546.110 2892.270 ;
        RECT 544.930 2889.490 546.110 2890.670 ;
        RECT 544.930 2711.090 546.110 2712.270 ;
        RECT 544.930 2709.490 546.110 2710.670 ;
        RECT 544.930 2531.090 546.110 2532.270 ;
        RECT 544.930 2529.490 546.110 2530.670 ;
        RECT 544.930 2351.090 546.110 2352.270 ;
        RECT 544.930 2349.490 546.110 2350.670 ;
        RECT 544.930 2171.090 546.110 2172.270 ;
        RECT 544.930 2169.490 546.110 2170.670 ;
        RECT 544.930 1991.090 546.110 1992.270 ;
        RECT 544.930 1989.490 546.110 1990.670 ;
        RECT 544.930 1811.090 546.110 1812.270 ;
        RECT 544.930 1809.490 546.110 1810.670 ;
        RECT 544.930 1631.090 546.110 1632.270 ;
        RECT 544.930 1629.490 546.110 1630.670 ;
        RECT 544.930 1451.090 546.110 1452.270 ;
        RECT 544.930 1449.490 546.110 1450.670 ;
        RECT 544.930 1271.090 546.110 1272.270 ;
        RECT 544.930 1269.490 546.110 1270.670 ;
        RECT 544.930 1091.090 546.110 1092.270 ;
        RECT 544.930 1089.490 546.110 1090.670 ;
        RECT 544.930 911.090 546.110 912.270 ;
        RECT 544.930 909.490 546.110 910.670 ;
        RECT 544.930 731.090 546.110 732.270 ;
        RECT 544.930 729.490 546.110 730.670 ;
        RECT 544.930 551.090 546.110 552.270 ;
        RECT 544.930 549.490 546.110 550.670 ;
        RECT 544.930 371.090 546.110 372.270 ;
        RECT 544.930 369.490 546.110 370.670 ;
        RECT 544.930 191.090 546.110 192.270 ;
        RECT 544.930 189.490 546.110 190.670 ;
        RECT 544.930 11.090 546.110 12.270 ;
        RECT 544.930 9.490 546.110 10.670 ;
        RECT 544.930 -2.910 546.110 -1.730 ;
        RECT 544.930 -4.510 546.110 -3.330 ;
        RECT 724.930 3523.010 726.110 3524.190 ;
        RECT 724.930 3521.410 726.110 3522.590 ;
        RECT 724.930 3431.090 726.110 3432.270 ;
        RECT 724.930 3429.490 726.110 3430.670 ;
        RECT 724.930 3251.090 726.110 3252.270 ;
        RECT 724.930 3249.490 726.110 3250.670 ;
        RECT 724.930 3071.090 726.110 3072.270 ;
        RECT 724.930 3069.490 726.110 3070.670 ;
        RECT 724.930 2891.090 726.110 2892.270 ;
        RECT 724.930 2889.490 726.110 2890.670 ;
        RECT 724.930 2711.090 726.110 2712.270 ;
        RECT 724.930 2709.490 726.110 2710.670 ;
        RECT 724.930 2531.090 726.110 2532.270 ;
        RECT 724.930 2529.490 726.110 2530.670 ;
        RECT 724.930 2351.090 726.110 2352.270 ;
        RECT 724.930 2349.490 726.110 2350.670 ;
        RECT 724.930 2171.090 726.110 2172.270 ;
        RECT 724.930 2169.490 726.110 2170.670 ;
        RECT 724.930 1991.090 726.110 1992.270 ;
        RECT 724.930 1989.490 726.110 1990.670 ;
        RECT 724.930 1811.090 726.110 1812.270 ;
        RECT 724.930 1809.490 726.110 1810.670 ;
        RECT 724.930 1631.090 726.110 1632.270 ;
        RECT 724.930 1629.490 726.110 1630.670 ;
        RECT 724.930 1451.090 726.110 1452.270 ;
        RECT 724.930 1449.490 726.110 1450.670 ;
        RECT 724.930 1271.090 726.110 1272.270 ;
        RECT 724.930 1269.490 726.110 1270.670 ;
        RECT 724.930 1091.090 726.110 1092.270 ;
        RECT 724.930 1089.490 726.110 1090.670 ;
        RECT 724.930 911.090 726.110 912.270 ;
        RECT 724.930 909.490 726.110 910.670 ;
        RECT 724.930 731.090 726.110 732.270 ;
        RECT 724.930 729.490 726.110 730.670 ;
        RECT 724.930 551.090 726.110 552.270 ;
        RECT 724.930 549.490 726.110 550.670 ;
        RECT 724.930 371.090 726.110 372.270 ;
        RECT 724.930 369.490 726.110 370.670 ;
        RECT 724.930 191.090 726.110 192.270 ;
        RECT 724.930 189.490 726.110 190.670 ;
        RECT 724.930 11.090 726.110 12.270 ;
        RECT 724.930 9.490 726.110 10.670 ;
        RECT 724.930 -2.910 726.110 -1.730 ;
        RECT 724.930 -4.510 726.110 -3.330 ;
        RECT 904.930 3523.010 906.110 3524.190 ;
        RECT 904.930 3521.410 906.110 3522.590 ;
        RECT 904.930 3431.090 906.110 3432.270 ;
        RECT 904.930 3429.490 906.110 3430.670 ;
        RECT 904.930 3251.090 906.110 3252.270 ;
        RECT 904.930 3249.490 906.110 3250.670 ;
        RECT 904.930 3071.090 906.110 3072.270 ;
        RECT 904.930 3069.490 906.110 3070.670 ;
        RECT 904.930 2891.090 906.110 2892.270 ;
        RECT 904.930 2889.490 906.110 2890.670 ;
        RECT 904.930 2711.090 906.110 2712.270 ;
        RECT 904.930 2709.490 906.110 2710.670 ;
        RECT 904.930 2531.090 906.110 2532.270 ;
        RECT 904.930 2529.490 906.110 2530.670 ;
        RECT 904.930 2351.090 906.110 2352.270 ;
        RECT 904.930 2349.490 906.110 2350.670 ;
        RECT 904.930 2171.090 906.110 2172.270 ;
        RECT 904.930 2169.490 906.110 2170.670 ;
        RECT 904.930 1991.090 906.110 1992.270 ;
        RECT 904.930 1989.490 906.110 1990.670 ;
        RECT 904.930 1811.090 906.110 1812.270 ;
        RECT 904.930 1809.490 906.110 1810.670 ;
        RECT 904.930 1631.090 906.110 1632.270 ;
        RECT 904.930 1629.490 906.110 1630.670 ;
        RECT 904.930 1451.090 906.110 1452.270 ;
        RECT 904.930 1449.490 906.110 1450.670 ;
        RECT 904.930 1271.090 906.110 1272.270 ;
        RECT 904.930 1269.490 906.110 1270.670 ;
        RECT 904.930 1091.090 906.110 1092.270 ;
        RECT 904.930 1089.490 906.110 1090.670 ;
        RECT 904.930 911.090 906.110 912.270 ;
        RECT 904.930 909.490 906.110 910.670 ;
        RECT 904.930 731.090 906.110 732.270 ;
        RECT 904.930 729.490 906.110 730.670 ;
        RECT 904.930 551.090 906.110 552.270 ;
        RECT 904.930 549.490 906.110 550.670 ;
        RECT 904.930 371.090 906.110 372.270 ;
        RECT 904.930 369.490 906.110 370.670 ;
        RECT 904.930 191.090 906.110 192.270 ;
        RECT 904.930 189.490 906.110 190.670 ;
        RECT 904.930 11.090 906.110 12.270 ;
        RECT 904.930 9.490 906.110 10.670 ;
        RECT 904.930 -2.910 906.110 -1.730 ;
        RECT 904.930 -4.510 906.110 -3.330 ;
        RECT 1084.930 3523.010 1086.110 3524.190 ;
        RECT 1084.930 3521.410 1086.110 3522.590 ;
        RECT 1084.930 3431.090 1086.110 3432.270 ;
        RECT 1084.930 3429.490 1086.110 3430.670 ;
        RECT 1084.930 3251.090 1086.110 3252.270 ;
        RECT 1084.930 3249.490 1086.110 3250.670 ;
        RECT 1084.930 3071.090 1086.110 3072.270 ;
        RECT 1084.930 3069.490 1086.110 3070.670 ;
        RECT 1084.930 2891.090 1086.110 2892.270 ;
        RECT 1084.930 2889.490 1086.110 2890.670 ;
        RECT 1084.930 2711.090 1086.110 2712.270 ;
        RECT 1084.930 2709.490 1086.110 2710.670 ;
        RECT 1084.930 2531.090 1086.110 2532.270 ;
        RECT 1084.930 2529.490 1086.110 2530.670 ;
        RECT 1084.930 2351.090 1086.110 2352.270 ;
        RECT 1084.930 2349.490 1086.110 2350.670 ;
        RECT 1084.930 2171.090 1086.110 2172.270 ;
        RECT 1084.930 2169.490 1086.110 2170.670 ;
        RECT 1084.930 1991.090 1086.110 1992.270 ;
        RECT 1084.930 1989.490 1086.110 1990.670 ;
        RECT 1084.930 1811.090 1086.110 1812.270 ;
        RECT 1084.930 1809.490 1086.110 1810.670 ;
        RECT 1084.930 1631.090 1086.110 1632.270 ;
        RECT 1084.930 1629.490 1086.110 1630.670 ;
        RECT 1084.930 1451.090 1086.110 1452.270 ;
        RECT 1084.930 1449.490 1086.110 1450.670 ;
        RECT 1084.930 1271.090 1086.110 1272.270 ;
        RECT 1084.930 1269.490 1086.110 1270.670 ;
        RECT 1084.930 1091.090 1086.110 1092.270 ;
        RECT 1084.930 1089.490 1086.110 1090.670 ;
        RECT 1084.930 911.090 1086.110 912.270 ;
        RECT 1084.930 909.490 1086.110 910.670 ;
        RECT 1084.930 731.090 1086.110 732.270 ;
        RECT 1084.930 729.490 1086.110 730.670 ;
        RECT 1084.930 551.090 1086.110 552.270 ;
        RECT 1084.930 549.490 1086.110 550.670 ;
        RECT 1084.930 371.090 1086.110 372.270 ;
        RECT 1084.930 369.490 1086.110 370.670 ;
        RECT 1084.930 191.090 1086.110 192.270 ;
        RECT 1084.930 189.490 1086.110 190.670 ;
        RECT 1084.930 11.090 1086.110 12.270 ;
        RECT 1084.930 9.490 1086.110 10.670 ;
        RECT 1084.930 -2.910 1086.110 -1.730 ;
        RECT 1084.930 -4.510 1086.110 -3.330 ;
        RECT 1264.930 3523.010 1266.110 3524.190 ;
        RECT 1264.930 3521.410 1266.110 3522.590 ;
        RECT 1264.930 3431.090 1266.110 3432.270 ;
        RECT 1264.930 3429.490 1266.110 3430.670 ;
        RECT 1264.930 3251.090 1266.110 3252.270 ;
        RECT 1264.930 3249.490 1266.110 3250.670 ;
        RECT 1264.930 3071.090 1266.110 3072.270 ;
        RECT 1264.930 3069.490 1266.110 3070.670 ;
        RECT 1264.930 2891.090 1266.110 2892.270 ;
        RECT 1264.930 2889.490 1266.110 2890.670 ;
        RECT 1264.930 2711.090 1266.110 2712.270 ;
        RECT 1264.930 2709.490 1266.110 2710.670 ;
        RECT 1264.930 2531.090 1266.110 2532.270 ;
        RECT 1264.930 2529.490 1266.110 2530.670 ;
        RECT 1264.930 2351.090 1266.110 2352.270 ;
        RECT 1264.930 2349.490 1266.110 2350.670 ;
        RECT 1264.930 2171.090 1266.110 2172.270 ;
        RECT 1264.930 2169.490 1266.110 2170.670 ;
        RECT 1264.930 1991.090 1266.110 1992.270 ;
        RECT 1264.930 1989.490 1266.110 1990.670 ;
        RECT 1264.930 1811.090 1266.110 1812.270 ;
        RECT 1264.930 1809.490 1266.110 1810.670 ;
        RECT 1264.930 1631.090 1266.110 1632.270 ;
        RECT 1264.930 1629.490 1266.110 1630.670 ;
        RECT 1264.930 1451.090 1266.110 1452.270 ;
        RECT 1264.930 1449.490 1266.110 1450.670 ;
        RECT 1264.930 1271.090 1266.110 1272.270 ;
        RECT 1264.930 1269.490 1266.110 1270.670 ;
        RECT 1264.930 1091.090 1266.110 1092.270 ;
        RECT 1264.930 1089.490 1266.110 1090.670 ;
        RECT 1264.930 911.090 1266.110 912.270 ;
        RECT 1264.930 909.490 1266.110 910.670 ;
        RECT 1264.930 731.090 1266.110 732.270 ;
        RECT 1264.930 729.490 1266.110 730.670 ;
        RECT 1264.930 551.090 1266.110 552.270 ;
        RECT 1264.930 549.490 1266.110 550.670 ;
        RECT 1264.930 371.090 1266.110 372.270 ;
        RECT 1264.930 369.490 1266.110 370.670 ;
        RECT 1264.930 191.090 1266.110 192.270 ;
        RECT 1264.930 189.490 1266.110 190.670 ;
        RECT 1264.930 11.090 1266.110 12.270 ;
        RECT 1264.930 9.490 1266.110 10.670 ;
        RECT 1264.930 -2.910 1266.110 -1.730 ;
        RECT 1264.930 -4.510 1266.110 -3.330 ;
        RECT 1444.930 3523.010 1446.110 3524.190 ;
        RECT 1444.930 3521.410 1446.110 3522.590 ;
        RECT 1444.930 3431.090 1446.110 3432.270 ;
        RECT 1444.930 3429.490 1446.110 3430.670 ;
        RECT 1444.930 3251.090 1446.110 3252.270 ;
        RECT 1444.930 3249.490 1446.110 3250.670 ;
        RECT 1444.930 3071.090 1446.110 3072.270 ;
        RECT 1444.930 3069.490 1446.110 3070.670 ;
        RECT 1444.930 2891.090 1446.110 2892.270 ;
        RECT 1444.930 2889.490 1446.110 2890.670 ;
        RECT 1444.930 2711.090 1446.110 2712.270 ;
        RECT 1444.930 2709.490 1446.110 2710.670 ;
        RECT 1444.930 2531.090 1446.110 2532.270 ;
        RECT 1444.930 2529.490 1446.110 2530.670 ;
        RECT 1444.930 2351.090 1446.110 2352.270 ;
        RECT 1444.930 2349.490 1446.110 2350.670 ;
        RECT 1444.930 2171.090 1446.110 2172.270 ;
        RECT 1444.930 2169.490 1446.110 2170.670 ;
        RECT 1444.930 1991.090 1446.110 1992.270 ;
        RECT 1444.930 1989.490 1446.110 1990.670 ;
        RECT 1444.930 1811.090 1446.110 1812.270 ;
        RECT 1444.930 1809.490 1446.110 1810.670 ;
        RECT 1444.930 1631.090 1446.110 1632.270 ;
        RECT 1444.930 1629.490 1446.110 1630.670 ;
        RECT 1444.930 1451.090 1446.110 1452.270 ;
        RECT 1444.930 1449.490 1446.110 1450.670 ;
        RECT 1444.930 1271.090 1446.110 1272.270 ;
        RECT 1444.930 1269.490 1446.110 1270.670 ;
        RECT 1444.930 1091.090 1446.110 1092.270 ;
        RECT 1444.930 1089.490 1446.110 1090.670 ;
        RECT 1444.930 911.090 1446.110 912.270 ;
        RECT 1444.930 909.490 1446.110 910.670 ;
        RECT 1444.930 731.090 1446.110 732.270 ;
        RECT 1444.930 729.490 1446.110 730.670 ;
        RECT 1444.930 551.090 1446.110 552.270 ;
        RECT 1444.930 549.490 1446.110 550.670 ;
        RECT 1444.930 371.090 1446.110 372.270 ;
        RECT 1444.930 369.490 1446.110 370.670 ;
        RECT 1444.930 191.090 1446.110 192.270 ;
        RECT 1444.930 189.490 1446.110 190.670 ;
        RECT 1444.930 11.090 1446.110 12.270 ;
        RECT 1444.930 9.490 1446.110 10.670 ;
        RECT 1444.930 -2.910 1446.110 -1.730 ;
        RECT 1444.930 -4.510 1446.110 -3.330 ;
        RECT 1624.930 3523.010 1626.110 3524.190 ;
        RECT 1624.930 3521.410 1626.110 3522.590 ;
        RECT 1624.930 3431.090 1626.110 3432.270 ;
        RECT 1624.930 3429.490 1626.110 3430.670 ;
        RECT 1624.930 3251.090 1626.110 3252.270 ;
        RECT 1624.930 3249.490 1626.110 3250.670 ;
        RECT 1624.930 3071.090 1626.110 3072.270 ;
        RECT 1624.930 3069.490 1626.110 3070.670 ;
        RECT 1624.930 2891.090 1626.110 2892.270 ;
        RECT 1624.930 2889.490 1626.110 2890.670 ;
        RECT 1624.930 2711.090 1626.110 2712.270 ;
        RECT 1624.930 2709.490 1626.110 2710.670 ;
        RECT 1624.930 2531.090 1626.110 2532.270 ;
        RECT 1624.930 2529.490 1626.110 2530.670 ;
        RECT 1624.930 2351.090 1626.110 2352.270 ;
        RECT 1624.930 2349.490 1626.110 2350.670 ;
        RECT 1624.930 2171.090 1626.110 2172.270 ;
        RECT 1624.930 2169.490 1626.110 2170.670 ;
        RECT 1624.930 1991.090 1626.110 1992.270 ;
        RECT 1624.930 1989.490 1626.110 1990.670 ;
        RECT 1624.930 1811.090 1626.110 1812.270 ;
        RECT 1624.930 1809.490 1626.110 1810.670 ;
        RECT 1624.930 1631.090 1626.110 1632.270 ;
        RECT 1624.930 1629.490 1626.110 1630.670 ;
        RECT 1624.930 1451.090 1626.110 1452.270 ;
        RECT 1624.930 1449.490 1626.110 1450.670 ;
        RECT 1624.930 1271.090 1626.110 1272.270 ;
        RECT 1624.930 1269.490 1626.110 1270.670 ;
        RECT 1624.930 1091.090 1626.110 1092.270 ;
        RECT 1624.930 1089.490 1626.110 1090.670 ;
        RECT 1624.930 911.090 1626.110 912.270 ;
        RECT 1624.930 909.490 1626.110 910.670 ;
        RECT 1624.930 731.090 1626.110 732.270 ;
        RECT 1624.930 729.490 1626.110 730.670 ;
        RECT 1624.930 551.090 1626.110 552.270 ;
        RECT 1624.930 549.490 1626.110 550.670 ;
        RECT 1624.930 371.090 1626.110 372.270 ;
        RECT 1624.930 369.490 1626.110 370.670 ;
        RECT 1624.930 191.090 1626.110 192.270 ;
        RECT 1624.930 189.490 1626.110 190.670 ;
        RECT 1624.930 11.090 1626.110 12.270 ;
        RECT 1624.930 9.490 1626.110 10.670 ;
        RECT 1624.930 -2.910 1626.110 -1.730 ;
        RECT 1624.930 -4.510 1626.110 -3.330 ;
        RECT 1804.930 3523.010 1806.110 3524.190 ;
        RECT 1804.930 3521.410 1806.110 3522.590 ;
        RECT 1804.930 3431.090 1806.110 3432.270 ;
        RECT 1804.930 3429.490 1806.110 3430.670 ;
        RECT 1804.930 3251.090 1806.110 3252.270 ;
        RECT 1804.930 3249.490 1806.110 3250.670 ;
        RECT 1804.930 3071.090 1806.110 3072.270 ;
        RECT 1804.930 3069.490 1806.110 3070.670 ;
        RECT 1804.930 2891.090 1806.110 2892.270 ;
        RECT 1804.930 2889.490 1806.110 2890.670 ;
        RECT 1804.930 2711.090 1806.110 2712.270 ;
        RECT 1804.930 2709.490 1806.110 2710.670 ;
        RECT 1804.930 2531.090 1806.110 2532.270 ;
        RECT 1804.930 2529.490 1806.110 2530.670 ;
        RECT 1804.930 2351.090 1806.110 2352.270 ;
        RECT 1804.930 2349.490 1806.110 2350.670 ;
        RECT 1804.930 2171.090 1806.110 2172.270 ;
        RECT 1804.930 2169.490 1806.110 2170.670 ;
        RECT 1804.930 1991.090 1806.110 1992.270 ;
        RECT 1804.930 1989.490 1806.110 1990.670 ;
        RECT 1804.930 1811.090 1806.110 1812.270 ;
        RECT 1804.930 1809.490 1806.110 1810.670 ;
        RECT 1804.930 1631.090 1806.110 1632.270 ;
        RECT 1804.930 1629.490 1806.110 1630.670 ;
        RECT 1804.930 1451.090 1806.110 1452.270 ;
        RECT 1804.930 1449.490 1806.110 1450.670 ;
        RECT 1804.930 1271.090 1806.110 1272.270 ;
        RECT 1804.930 1269.490 1806.110 1270.670 ;
        RECT 1804.930 1091.090 1806.110 1092.270 ;
        RECT 1804.930 1089.490 1806.110 1090.670 ;
        RECT 1804.930 911.090 1806.110 912.270 ;
        RECT 1804.930 909.490 1806.110 910.670 ;
        RECT 1804.930 731.090 1806.110 732.270 ;
        RECT 1804.930 729.490 1806.110 730.670 ;
        RECT 1804.930 551.090 1806.110 552.270 ;
        RECT 1804.930 549.490 1806.110 550.670 ;
        RECT 1804.930 371.090 1806.110 372.270 ;
        RECT 1804.930 369.490 1806.110 370.670 ;
        RECT 1804.930 191.090 1806.110 192.270 ;
        RECT 1804.930 189.490 1806.110 190.670 ;
        RECT 1804.930 11.090 1806.110 12.270 ;
        RECT 1804.930 9.490 1806.110 10.670 ;
        RECT 1804.930 -2.910 1806.110 -1.730 ;
        RECT 1804.930 -4.510 1806.110 -3.330 ;
        RECT 1984.930 3523.010 1986.110 3524.190 ;
        RECT 1984.930 3521.410 1986.110 3522.590 ;
        RECT 1984.930 3431.090 1986.110 3432.270 ;
        RECT 1984.930 3429.490 1986.110 3430.670 ;
        RECT 1984.930 3251.090 1986.110 3252.270 ;
        RECT 1984.930 3249.490 1986.110 3250.670 ;
        RECT 1984.930 3071.090 1986.110 3072.270 ;
        RECT 1984.930 3069.490 1986.110 3070.670 ;
        RECT 1984.930 2891.090 1986.110 2892.270 ;
        RECT 1984.930 2889.490 1986.110 2890.670 ;
        RECT 1984.930 2711.090 1986.110 2712.270 ;
        RECT 1984.930 2709.490 1986.110 2710.670 ;
        RECT 1984.930 2531.090 1986.110 2532.270 ;
        RECT 1984.930 2529.490 1986.110 2530.670 ;
        RECT 1984.930 2351.090 1986.110 2352.270 ;
        RECT 1984.930 2349.490 1986.110 2350.670 ;
        RECT 1984.930 2171.090 1986.110 2172.270 ;
        RECT 1984.930 2169.490 1986.110 2170.670 ;
        RECT 1984.930 1991.090 1986.110 1992.270 ;
        RECT 1984.930 1989.490 1986.110 1990.670 ;
        RECT 1984.930 1811.090 1986.110 1812.270 ;
        RECT 1984.930 1809.490 1986.110 1810.670 ;
        RECT 1984.930 1631.090 1986.110 1632.270 ;
        RECT 1984.930 1629.490 1986.110 1630.670 ;
        RECT 1984.930 1451.090 1986.110 1452.270 ;
        RECT 1984.930 1449.490 1986.110 1450.670 ;
        RECT 1984.930 1271.090 1986.110 1272.270 ;
        RECT 1984.930 1269.490 1986.110 1270.670 ;
        RECT 1984.930 1091.090 1986.110 1092.270 ;
        RECT 1984.930 1089.490 1986.110 1090.670 ;
        RECT 1984.930 911.090 1986.110 912.270 ;
        RECT 1984.930 909.490 1986.110 910.670 ;
        RECT 1984.930 731.090 1986.110 732.270 ;
        RECT 1984.930 729.490 1986.110 730.670 ;
        RECT 1984.930 551.090 1986.110 552.270 ;
        RECT 1984.930 549.490 1986.110 550.670 ;
        RECT 1984.930 371.090 1986.110 372.270 ;
        RECT 1984.930 369.490 1986.110 370.670 ;
        RECT 1984.930 191.090 1986.110 192.270 ;
        RECT 1984.930 189.490 1986.110 190.670 ;
        RECT 1984.930 11.090 1986.110 12.270 ;
        RECT 1984.930 9.490 1986.110 10.670 ;
        RECT 1984.930 -2.910 1986.110 -1.730 ;
        RECT 1984.930 -4.510 1986.110 -3.330 ;
        RECT 2164.930 3523.010 2166.110 3524.190 ;
        RECT 2164.930 3521.410 2166.110 3522.590 ;
        RECT 2164.930 3431.090 2166.110 3432.270 ;
        RECT 2164.930 3429.490 2166.110 3430.670 ;
        RECT 2164.930 3251.090 2166.110 3252.270 ;
        RECT 2164.930 3249.490 2166.110 3250.670 ;
        RECT 2164.930 3071.090 2166.110 3072.270 ;
        RECT 2164.930 3069.490 2166.110 3070.670 ;
        RECT 2164.930 2891.090 2166.110 2892.270 ;
        RECT 2164.930 2889.490 2166.110 2890.670 ;
        RECT 2164.930 2711.090 2166.110 2712.270 ;
        RECT 2164.930 2709.490 2166.110 2710.670 ;
        RECT 2164.930 2531.090 2166.110 2532.270 ;
        RECT 2164.930 2529.490 2166.110 2530.670 ;
        RECT 2164.930 2351.090 2166.110 2352.270 ;
        RECT 2164.930 2349.490 2166.110 2350.670 ;
        RECT 2164.930 2171.090 2166.110 2172.270 ;
        RECT 2164.930 2169.490 2166.110 2170.670 ;
        RECT 2164.930 1991.090 2166.110 1992.270 ;
        RECT 2164.930 1989.490 2166.110 1990.670 ;
        RECT 2164.930 1811.090 2166.110 1812.270 ;
        RECT 2164.930 1809.490 2166.110 1810.670 ;
        RECT 2164.930 1631.090 2166.110 1632.270 ;
        RECT 2164.930 1629.490 2166.110 1630.670 ;
        RECT 2164.930 1451.090 2166.110 1452.270 ;
        RECT 2164.930 1449.490 2166.110 1450.670 ;
        RECT 2164.930 1271.090 2166.110 1272.270 ;
        RECT 2164.930 1269.490 2166.110 1270.670 ;
        RECT 2164.930 1091.090 2166.110 1092.270 ;
        RECT 2164.930 1089.490 2166.110 1090.670 ;
        RECT 2164.930 911.090 2166.110 912.270 ;
        RECT 2164.930 909.490 2166.110 910.670 ;
        RECT 2164.930 731.090 2166.110 732.270 ;
        RECT 2164.930 729.490 2166.110 730.670 ;
        RECT 2164.930 551.090 2166.110 552.270 ;
        RECT 2164.930 549.490 2166.110 550.670 ;
        RECT 2164.930 371.090 2166.110 372.270 ;
        RECT 2164.930 369.490 2166.110 370.670 ;
        RECT 2164.930 191.090 2166.110 192.270 ;
        RECT 2164.930 189.490 2166.110 190.670 ;
        RECT 2164.930 11.090 2166.110 12.270 ;
        RECT 2164.930 9.490 2166.110 10.670 ;
        RECT 2164.930 -2.910 2166.110 -1.730 ;
        RECT 2164.930 -4.510 2166.110 -3.330 ;
        RECT 2344.930 3523.010 2346.110 3524.190 ;
        RECT 2344.930 3521.410 2346.110 3522.590 ;
        RECT 2344.930 3431.090 2346.110 3432.270 ;
        RECT 2344.930 3429.490 2346.110 3430.670 ;
        RECT 2344.930 3251.090 2346.110 3252.270 ;
        RECT 2344.930 3249.490 2346.110 3250.670 ;
        RECT 2344.930 3071.090 2346.110 3072.270 ;
        RECT 2344.930 3069.490 2346.110 3070.670 ;
        RECT 2344.930 2891.090 2346.110 2892.270 ;
        RECT 2344.930 2889.490 2346.110 2890.670 ;
        RECT 2344.930 2711.090 2346.110 2712.270 ;
        RECT 2344.930 2709.490 2346.110 2710.670 ;
        RECT 2344.930 2531.090 2346.110 2532.270 ;
        RECT 2344.930 2529.490 2346.110 2530.670 ;
        RECT 2344.930 2351.090 2346.110 2352.270 ;
        RECT 2344.930 2349.490 2346.110 2350.670 ;
        RECT 2344.930 2171.090 2346.110 2172.270 ;
        RECT 2344.930 2169.490 2346.110 2170.670 ;
        RECT 2344.930 1991.090 2346.110 1992.270 ;
        RECT 2344.930 1989.490 2346.110 1990.670 ;
        RECT 2344.930 1811.090 2346.110 1812.270 ;
        RECT 2344.930 1809.490 2346.110 1810.670 ;
        RECT 2344.930 1631.090 2346.110 1632.270 ;
        RECT 2344.930 1629.490 2346.110 1630.670 ;
        RECT 2344.930 1451.090 2346.110 1452.270 ;
        RECT 2344.930 1449.490 2346.110 1450.670 ;
        RECT 2344.930 1271.090 2346.110 1272.270 ;
        RECT 2344.930 1269.490 2346.110 1270.670 ;
        RECT 2344.930 1091.090 2346.110 1092.270 ;
        RECT 2344.930 1089.490 2346.110 1090.670 ;
        RECT 2344.930 911.090 2346.110 912.270 ;
        RECT 2344.930 909.490 2346.110 910.670 ;
        RECT 2344.930 731.090 2346.110 732.270 ;
        RECT 2344.930 729.490 2346.110 730.670 ;
        RECT 2344.930 551.090 2346.110 552.270 ;
        RECT 2344.930 549.490 2346.110 550.670 ;
        RECT 2344.930 371.090 2346.110 372.270 ;
        RECT 2344.930 369.490 2346.110 370.670 ;
        RECT 2344.930 191.090 2346.110 192.270 ;
        RECT 2344.930 189.490 2346.110 190.670 ;
        RECT 2344.930 11.090 2346.110 12.270 ;
        RECT 2344.930 9.490 2346.110 10.670 ;
        RECT 2344.930 -2.910 2346.110 -1.730 ;
        RECT 2344.930 -4.510 2346.110 -3.330 ;
        RECT 2524.930 3523.010 2526.110 3524.190 ;
        RECT 2524.930 3521.410 2526.110 3522.590 ;
        RECT 2524.930 3431.090 2526.110 3432.270 ;
        RECT 2524.930 3429.490 2526.110 3430.670 ;
        RECT 2524.930 3251.090 2526.110 3252.270 ;
        RECT 2524.930 3249.490 2526.110 3250.670 ;
        RECT 2524.930 3071.090 2526.110 3072.270 ;
        RECT 2524.930 3069.490 2526.110 3070.670 ;
        RECT 2524.930 2891.090 2526.110 2892.270 ;
        RECT 2524.930 2889.490 2526.110 2890.670 ;
        RECT 2524.930 2711.090 2526.110 2712.270 ;
        RECT 2524.930 2709.490 2526.110 2710.670 ;
        RECT 2524.930 2531.090 2526.110 2532.270 ;
        RECT 2524.930 2529.490 2526.110 2530.670 ;
        RECT 2524.930 2351.090 2526.110 2352.270 ;
        RECT 2524.930 2349.490 2526.110 2350.670 ;
        RECT 2524.930 2171.090 2526.110 2172.270 ;
        RECT 2524.930 2169.490 2526.110 2170.670 ;
        RECT 2524.930 1991.090 2526.110 1992.270 ;
        RECT 2524.930 1989.490 2526.110 1990.670 ;
        RECT 2524.930 1811.090 2526.110 1812.270 ;
        RECT 2524.930 1809.490 2526.110 1810.670 ;
        RECT 2524.930 1631.090 2526.110 1632.270 ;
        RECT 2524.930 1629.490 2526.110 1630.670 ;
        RECT 2524.930 1451.090 2526.110 1452.270 ;
        RECT 2524.930 1449.490 2526.110 1450.670 ;
        RECT 2524.930 1271.090 2526.110 1272.270 ;
        RECT 2524.930 1269.490 2526.110 1270.670 ;
        RECT 2524.930 1091.090 2526.110 1092.270 ;
        RECT 2524.930 1089.490 2526.110 1090.670 ;
        RECT 2524.930 911.090 2526.110 912.270 ;
        RECT 2524.930 909.490 2526.110 910.670 ;
        RECT 2524.930 731.090 2526.110 732.270 ;
        RECT 2524.930 729.490 2526.110 730.670 ;
        RECT 2524.930 551.090 2526.110 552.270 ;
        RECT 2524.930 549.490 2526.110 550.670 ;
        RECT 2524.930 371.090 2526.110 372.270 ;
        RECT 2524.930 369.490 2526.110 370.670 ;
        RECT 2524.930 191.090 2526.110 192.270 ;
        RECT 2524.930 189.490 2526.110 190.670 ;
        RECT 2524.930 11.090 2526.110 12.270 ;
        RECT 2524.930 9.490 2526.110 10.670 ;
        RECT 2524.930 -2.910 2526.110 -1.730 ;
        RECT 2524.930 -4.510 2526.110 -3.330 ;
        RECT 2704.930 3523.010 2706.110 3524.190 ;
        RECT 2704.930 3521.410 2706.110 3522.590 ;
        RECT 2704.930 3431.090 2706.110 3432.270 ;
        RECT 2704.930 3429.490 2706.110 3430.670 ;
        RECT 2704.930 3251.090 2706.110 3252.270 ;
        RECT 2704.930 3249.490 2706.110 3250.670 ;
        RECT 2704.930 3071.090 2706.110 3072.270 ;
        RECT 2704.930 3069.490 2706.110 3070.670 ;
        RECT 2704.930 2891.090 2706.110 2892.270 ;
        RECT 2704.930 2889.490 2706.110 2890.670 ;
        RECT 2704.930 2711.090 2706.110 2712.270 ;
        RECT 2704.930 2709.490 2706.110 2710.670 ;
        RECT 2704.930 2531.090 2706.110 2532.270 ;
        RECT 2704.930 2529.490 2706.110 2530.670 ;
        RECT 2704.930 2351.090 2706.110 2352.270 ;
        RECT 2704.930 2349.490 2706.110 2350.670 ;
        RECT 2704.930 2171.090 2706.110 2172.270 ;
        RECT 2704.930 2169.490 2706.110 2170.670 ;
        RECT 2704.930 1991.090 2706.110 1992.270 ;
        RECT 2704.930 1989.490 2706.110 1990.670 ;
        RECT 2704.930 1811.090 2706.110 1812.270 ;
        RECT 2704.930 1809.490 2706.110 1810.670 ;
        RECT 2704.930 1631.090 2706.110 1632.270 ;
        RECT 2704.930 1629.490 2706.110 1630.670 ;
        RECT 2704.930 1451.090 2706.110 1452.270 ;
        RECT 2704.930 1449.490 2706.110 1450.670 ;
        RECT 2704.930 1271.090 2706.110 1272.270 ;
        RECT 2704.930 1269.490 2706.110 1270.670 ;
        RECT 2704.930 1091.090 2706.110 1092.270 ;
        RECT 2704.930 1089.490 2706.110 1090.670 ;
        RECT 2704.930 911.090 2706.110 912.270 ;
        RECT 2704.930 909.490 2706.110 910.670 ;
        RECT 2704.930 731.090 2706.110 732.270 ;
        RECT 2704.930 729.490 2706.110 730.670 ;
        RECT 2704.930 551.090 2706.110 552.270 ;
        RECT 2704.930 549.490 2706.110 550.670 ;
        RECT 2704.930 371.090 2706.110 372.270 ;
        RECT 2704.930 369.490 2706.110 370.670 ;
        RECT 2704.930 191.090 2706.110 192.270 ;
        RECT 2704.930 189.490 2706.110 190.670 ;
        RECT 2704.930 11.090 2706.110 12.270 ;
        RECT 2704.930 9.490 2706.110 10.670 ;
        RECT 2704.930 -2.910 2706.110 -1.730 ;
        RECT 2704.930 -4.510 2706.110 -3.330 ;
        RECT 2884.930 3523.010 2886.110 3524.190 ;
        RECT 2884.930 3521.410 2886.110 3522.590 ;
        RECT 2884.930 3431.090 2886.110 3432.270 ;
        RECT 2884.930 3429.490 2886.110 3430.670 ;
        RECT 2884.930 3251.090 2886.110 3252.270 ;
        RECT 2884.930 3249.490 2886.110 3250.670 ;
        RECT 2884.930 3071.090 2886.110 3072.270 ;
        RECT 2884.930 3069.490 2886.110 3070.670 ;
        RECT 2884.930 2891.090 2886.110 2892.270 ;
        RECT 2884.930 2889.490 2886.110 2890.670 ;
        RECT 2884.930 2711.090 2886.110 2712.270 ;
        RECT 2884.930 2709.490 2886.110 2710.670 ;
        RECT 2884.930 2531.090 2886.110 2532.270 ;
        RECT 2884.930 2529.490 2886.110 2530.670 ;
        RECT 2884.930 2351.090 2886.110 2352.270 ;
        RECT 2884.930 2349.490 2886.110 2350.670 ;
        RECT 2884.930 2171.090 2886.110 2172.270 ;
        RECT 2884.930 2169.490 2886.110 2170.670 ;
        RECT 2884.930 1991.090 2886.110 1992.270 ;
        RECT 2884.930 1989.490 2886.110 1990.670 ;
        RECT 2884.930 1811.090 2886.110 1812.270 ;
        RECT 2884.930 1809.490 2886.110 1810.670 ;
        RECT 2884.930 1631.090 2886.110 1632.270 ;
        RECT 2884.930 1629.490 2886.110 1630.670 ;
        RECT 2884.930 1451.090 2886.110 1452.270 ;
        RECT 2884.930 1449.490 2886.110 1450.670 ;
        RECT 2884.930 1271.090 2886.110 1272.270 ;
        RECT 2884.930 1269.490 2886.110 1270.670 ;
        RECT 2884.930 1091.090 2886.110 1092.270 ;
        RECT 2884.930 1089.490 2886.110 1090.670 ;
        RECT 2884.930 911.090 2886.110 912.270 ;
        RECT 2884.930 909.490 2886.110 910.670 ;
        RECT 2884.930 731.090 2886.110 732.270 ;
        RECT 2884.930 729.490 2886.110 730.670 ;
        RECT 2884.930 551.090 2886.110 552.270 ;
        RECT 2884.930 549.490 2886.110 550.670 ;
        RECT 2884.930 371.090 2886.110 372.270 ;
        RECT 2884.930 369.490 2886.110 370.670 ;
        RECT 2884.930 191.090 2886.110 192.270 ;
        RECT 2884.930 189.490 2886.110 190.670 ;
        RECT 2884.930 11.090 2886.110 12.270 ;
        RECT 2884.930 9.490 2886.110 10.670 ;
        RECT 2884.930 -2.910 2886.110 -1.730 ;
        RECT 2884.930 -4.510 2886.110 -3.330 ;
        RECT 2927.510 3523.010 2928.690 3524.190 ;
        RECT 2927.510 3521.410 2928.690 3522.590 ;
        RECT 2927.510 3431.090 2928.690 3432.270 ;
        RECT 2927.510 3429.490 2928.690 3430.670 ;
        RECT 2927.510 3251.090 2928.690 3252.270 ;
        RECT 2927.510 3249.490 2928.690 3250.670 ;
        RECT 2927.510 3071.090 2928.690 3072.270 ;
        RECT 2927.510 3069.490 2928.690 3070.670 ;
        RECT 2927.510 2891.090 2928.690 2892.270 ;
        RECT 2927.510 2889.490 2928.690 2890.670 ;
        RECT 2927.510 2711.090 2928.690 2712.270 ;
        RECT 2927.510 2709.490 2928.690 2710.670 ;
        RECT 2927.510 2531.090 2928.690 2532.270 ;
        RECT 2927.510 2529.490 2928.690 2530.670 ;
        RECT 2927.510 2351.090 2928.690 2352.270 ;
        RECT 2927.510 2349.490 2928.690 2350.670 ;
        RECT 2927.510 2171.090 2928.690 2172.270 ;
        RECT 2927.510 2169.490 2928.690 2170.670 ;
        RECT 2927.510 1991.090 2928.690 1992.270 ;
        RECT 2927.510 1989.490 2928.690 1990.670 ;
        RECT 2927.510 1811.090 2928.690 1812.270 ;
        RECT 2927.510 1809.490 2928.690 1810.670 ;
        RECT 2927.510 1631.090 2928.690 1632.270 ;
        RECT 2927.510 1629.490 2928.690 1630.670 ;
        RECT 2927.510 1451.090 2928.690 1452.270 ;
        RECT 2927.510 1449.490 2928.690 1450.670 ;
        RECT 2927.510 1271.090 2928.690 1272.270 ;
        RECT 2927.510 1269.490 2928.690 1270.670 ;
        RECT 2927.510 1091.090 2928.690 1092.270 ;
        RECT 2927.510 1089.490 2928.690 1090.670 ;
        RECT 2927.510 911.090 2928.690 912.270 ;
        RECT 2927.510 909.490 2928.690 910.670 ;
        RECT 2927.510 731.090 2928.690 732.270 ;
        RECT 2927.510 729.490 2928.690 730.670 ;
        RECT 2927.510 551.090 2928.690 552.270 ;
        RECT 2927.510 549.490 2928.690 550.670 ;
        RECT 2927.510 371.090 2928.690 372.270 ;
        RECT 2927.510 369.490 2928.690 370.670 ;
        RECT 2927.510 191.090 2928.690 192.270 ;
        RECT 2927.510 189.490 2928.690 190.670 ;
        RECT 2927.510 11.090 2928.690 12.270 ;
        RECT 2927.510 9.490 2928.690 10.670 ;
        RECT 2927.510 -2.910 2928.690 -1.730 ;
        RECT 2927.510 -4.510 2928.690 -3.330 ;
      LAYER met5 ;
        RECT -9.980 3524.300 -6.980 3524.310 ;
        RECT 4.020 3524.300 7.020 3524.310 ;
        RECT 184.020 3524.300 187.020 3524.310 ;
        RECT 364.020 3524.300 367.020 3524.310 ;
        RECT 544.020 3524.300 547.020 3524.310 ;
        RECT 724.020 3524.300 727.020 3524.310 ;
        RECT 904.020 3524.300 907.020 3524.310 ;
        RECT 1084.020 3524.300 1087.020 3524.310 ;
        RECT 1264.020 3524.300 1267.020 3524.310 ;
        RECT 1444.020 3524.300 1447.020 3524.310 ;
        RECT 1624.020 3524.300 1627.020 3524.310 ;
        RECT 1804.020 3524.300 1807.020 3524.310 ;
        RECT 1984.020 3524.300 1987.020 3524.310 ;
        RECT 2164.020 3524.300 2167.020 3524.310 ;
        RECT 2344.020 3524.300 2347.020 3524.310 ;
        RECT 2524.020 3524.300 2527.020 3524.310 ;
        RECT 2704.020 3524.300 2707.020 3524.310 ;
        RECT 2884.020 3524.300 2887.020 3524.310 ;
        RECT 2926.600 3524.300 2929.600 3524.310 ;
        RECT -9.980 3521.300 2929.600 3524.300 ;
        RECT -9.980 3521.290 -6.980 3521.300 ;
        RECT 4.020 3521.290 7.020 3521.300 ;
        RECT 184.020 3521.290 187.020 3521.300 ;
        RECT 364.020 3521.290 367.020 3521.300 ;
        RECT 544.020 3521.290 547.020 3521.300 ;
        RECT 724.020 3521.290 727.020 3521.300 ;
        RECT 904.020 3521.290 907.020 3521.300 ;
        RECT 1084.020 3521.290 1087.020 3521.300 ;
        RECT 1264.020 3521.290 1267.020 3521.300 ;
        RECT 1444.020 3521.290 1447.020 3521.300 ;
        RECT 1624.020 3521.290 1627.020 3521.300 ;
        RECT 1804.020 3521.290 1807.020 3521.300 ;
        RECT 1984.020 3521.290 1987.020 3521.300 ;
        RECT 2164.020 3521.290 2167.020 3521.300 ;
        RECT 2344.020 3521.290 2347.020 3521.300 ;
        RECT 2524.020 3521.290 2527.020 3521.300 ;
        RECT 2704.020 3521.290 2707.020 3521.300 ;
        RECT 2884.020 3521.290 2887.020 3521.300 ;
        RECT 2926.600 3521.290 2929.600 3521.300 ;
        RECT -9.980 3432.380 -6.980 3432.390 ;
        RECT 4.020 3432.380 7.020 3432.390 ;
        RECT 184.020 3432.380 187.020 3432.390 ;
        RECT 364.020 3432.380 367.020 3432.390 ;
        RECT 544.020 3432.380 547.020 3432.390 ;
        RECT 724.020 3432.380 727.020 3432.390 ;
        RECT 904.020 3432.380 907.020 3432.390 ;
        RECT 1084.020 3432.380 1087.020 3432.390 ;
        RECT 1264.020 3432.380 1267.020 3432.390 ;
        RECT 1444.020 3432.380 1447.020 3432.390 ;
        RECT 1624.020 3432.380 1627.020 3432.390 ;
        RECT 1804.020 3432.380 1807.020 3432.390 ;
        RECT 1984.020 3432.380 1987.020 3432.390 ;
        RECT 2164.020 3432.380 2167.020 3432.390 ;
        RECT 2344.020 3432.380 2347.020 3432.390 ;
        RECT 2524.020 3432.380 2527.020 3432.390 ;
        RECT 2704.020 3432.380 2707.020 3432.390 ;
        RECT 2884.020 3432.380 2887.020 3432.390 ;
        RECT 2926.600 3432.380 2929.600 3432.390 ;
        RECT -14.580 3429.380 2934.200 3432.380 ;
        RECT -9.980 3429.370 -6.980 3429.380 ;
        RECT 4.020 3429.370 7.020 3429.380 ;
        RECT 184.020 3429.370 187.020 3429.380 ;
        RECT 364.020 3429.370 367.020 3429.380 ;
        RECT 544.020 3429.370 547.020 3429.380 ;
        RECT 724.020 3429.370 727.020 3429.380 ;
        RECT 904.020 3429.370 907.020 3429.380 ;
        RECT 1084.020 3429.370 1087.020 3429.380 ;
        RECT 1264.020 3429.370 1267.020 3429.380 ;
        RECT 1444.020 3429.370 1447.020 3429.380 ;
        RECT 1624.020 3429.370 1627.020 3429.380 ;
        RECT 1804.020 3429.370 1807.020 3429.380 ;
        RECT 1984.020 3429.370 1987.020 3429.380 ;
        RECT 2164.020 3429.370 2167.020 3429.380 ;
        RECT 2344.020 3429.370 2347.020 3429.380 ;
        RECT 2524.020 3429.370 2527.020 3429.380 ;
        RECT 2704.020 3429.370 2707.020 3429.380 ;
        RECT 2884.020 3429.370 2887.020 3429.380 ;
        RECT 2926.600 3429.370 2929.600 3429.380 ;
        RECT -9.980 3252.380 -6.980 3252.390 ;
        RECT 4.020 3252.380 7.020 3252.390 ;
        RECT 184.020 3252.380 187.020 3252.390 ;
        RECT 364.020 3252.380 367.020 3252.390 ;
        RECT 544.020 3252.380 547.020 3252.390 ;
        RECT 724.020 3252.380 727.020 3252.390 ;
        RECT 904.020 3252.380 907.020 3252.390 ;
        RECT 1084.020 3252.380 1087.020 3252.390 ;
        RECT 1264.020 3252.380 1267.020 3252.390 ;
        RECT 1444.020 3252.380 1447.020 3252.390 ;
        RECT 1624.020 3252.380 1627.020 3252.390 ;
        RECT 1804.020 3252.380 1807.020 3252.390 ;
        RECT 1984.020 3252.380 1987.020 3252.390 ;
        RECT 2164.020 3252.380 2167.020 3252.390 ;
        RECT 2344.020 3252.380 2347.020 3252.390 ;
        RECT 2524.020 3252.380 2527.020 3252.390 ;
        RECT 2704.020 3252.380 2707.020 3252.390 ;
        RECT 2884.020 3252.380 2887.020 3252.390 ;
        RECT 2926.600 3252.380 2929.600 3252.390 ;
        RECT -14.580 3249.380 2934.200 3252.380 ;
        RECT -9.980 3249.370 -6.980 3249.380 ;
        RECT 4.020 3249.370 7.020 3249.380 ;
        RECT 184.020 3249.370 187.020 3249.380 ;
        RECT 364.020 3249.370 367.020 3249.380 ;
        RECT 544.020 3249.370 547.020 3249.380 ;
        RECT 724.020 3249.370 727.020 3249.380 ;
        RECT 904.020 3249.370 907.020 3249.380 ;
        RECT 1084.020 3249.370 1087.020 3249.380 ;
        RECT 1264.020 3249.370 1267.020 3249.380 ;
        RECT 1444.020 3249.370 1447.020 3249.380 ;
        RECT 1624.020 3249.370 1627.020 3249.380 ;
        RECT 1804.020 3249.370 1807.020 3249.380 ;
        RECT 1984.020 3249.370 1987.020 3249.380 ;
        RECT 2164.020 3249.370 2167.020 3249.380 ;
        RECT 2344.020 3249.370 2347.020 3249.380 ;
        RECT 2524.020 3249.370 2527.020 3249.380 ;
        RECT 2704.020 3249.370 2707.020 3249.380 ;
        RECT 2884.020 3249.370 2887.020 3249.380 ;
        RECT 2926.600 3249.370 2929.600 3249.380 ;
        RECT -9.980 3072.380 -6.980 3072.390 ;
        RECT 4.020 3072.380 7.020 3072.390 ;
        RECT 184.020 3072.380 187.020 3072.390 ;
        RECT 364.020 3072.380 367.020 3072.390 ;
        RECT 544.020 3072.380 547.020 3072.390 ;
        RECT 724.020 3072.380 727.020 3072.390 ;
        RECT 904.020 3072.380 907.020 3072.390 ;
        RECT 1084.020 3072.380 1087.020 3072.390 ;
        RECT 1264.020 3072.380 1267.020 3072.390 ;
        RECT 1444.020 3072.380 1447.020 3072.390 ;
        RECT 1624.020 3072.380 1627.020 3072.390 ;
        RECT 1804.020 3072.380 1807.020 3072.390 ;
        RECT 1984.020 3072.380 1987.020 3072.390 ;
        RECT 2164.020 3072.380 2167.020 3072.390 ;
        RECT 2344.020 3072.380 2347.020 3072.390 ;
        RECT 2524.020 3072.380 2527.020 3072.390 ;
        RECT 2704.020 3072.380 2707.020 3072.390 ;
        RECT 2884.020 3072.380 2887.020 3072.390 ;
        RECT 2926.600 3072.380 2929.600 3072.390 ;
        RECT -14.580 3069.380 2934.200 3072.380 ;
        RECT -9.980 3069.370 -6.980 3069.380 ;
        RECT 4.020 3069.370 7.020 3069.380 ;
        RECT 184.020 3069.370 187.020 3069.380 ;
        RECT 364.020 3069.370 367.020 3069.380 ;
        RECT 544.020 3069.370 547.020 3069.380 ;
        RECT 724.020 3069.370 727.020 3069.380 ;
        RECT 904.020 3069.370 907.020 3069.380 ;
        RECT 1084.020 3069.370 1087.020 3069.380 ;
        RECT 1264.020 3069.370 1267.020 3069.380 ;
        RECT 1444.020 3069.370 1447.020 3069.380 ;
        RECT 1624.020 3069.370 1627.020 3069.380 ;
        RECT 1804.020 3069.370 1807.020 3069.380 ;
        RECT 1984.020 3069.370 1987.020 3069.380 ;
        RECT 2164.020 3069.370 2167.020 3069.380 ;
        RECT 2344.020 3069.370 2347.020 3069.380 ;
        RECT 2524.020 3069.370 2527.020 3069.380 ;
        RECT 2704.020 3069.370 2707.020 3069.380 ;
        RECT 2884.020 3069.370 2887.020 3069.380 ;
        RECT 2926.600 3069.370 2929.600 3069.380 ;
        RECT -9.980 2892.380 -6.980 2892.390 ;
        RECT 4.020 2892.380 7.020 2892.390 ;
        RECT 184.020 2892.380 187.020 2892.390 ;
        RECT 364.020 2892.380 367.020 2892.390 ;
        RECT 544.020 2892.380 547.020 2892.390 ;
        RECT 724.020 2892.380 727.020 2892.390 ;
        RECT 904.020 2892.380 907.020 2892.390 ;
        RECT 1084.020 2892.380 1087.020 2892.390 ;
        RECT 1264.020 2892.380 1267.020 2892.390 ;
        RECT 1444.020 2892.380 1447.020 2892.390 ;
        RECT 1624.020 2892.380 1627.020 2892.390 ;
        RECT 1804.020 2892.380 1807.020 2892.390 ;
        RECT 1984.020 2892.380 1987.020 2892.390 ;
        RECT 2164.020 2892.380 2167.020 2892.390 ;
        RECT 2344.020 2892.380 2347.020 2892.390 ;
        RECT 2524.020 2892.380 2527.020 2892.390 ;
        RECT 2704.020 2892.380 2707.020 2892.390 ;
        RECT 2884.020 2892.380 2887.020 2892.390 ;
        RECT 2926.600 2892.380 2929.600 2892.390 ;
        RECT -14.580 2889.380 2934.200 2892.380 ;
        RECT -9.980 2889.370 -6.980 2889.380 ;
        RECT 4.020 2889.370 7.020 2889.380 ;
        RECT 184.020 2889.370 187.020 2889.380 ;
        RECT 364.020 2889.370 367.020 2889.380 ;
        RECT 544.020 2889.370 547.020 2889.380 ;
        RECT 724.020 2889.370 727.020 2889.380 ;
        RECT 904.020 2889.370 907.020 2889.380 ;
        RECT 1084.020 2889.370 1087.020 2889.380 ;
        RECT 1264.020 2889.370 1267.020 2889.380 ;
        RECT 1444.020 2889.370 1447.020 2889.380 ;
        RECT 1624.020 2889.370 1627.020 2889.380 ;
        RECT 1804.020 2889.370 1807.020 2889.380 ;
        RECT 1984.020 2889.370 1987.020 2889.380 ;
        RECT 2164.020 2889.370 2167.020 2889.380 ;
        RECT 2344.020 2889.370 2347.020 2889.380 ;
        RECT 2524.020 2889.370 2527.020 2889.380 ;
        RECT 2704.020 2889.370 2707.020 2889.380 ;
        RECT 2884.020 2889.370 2887.020 2889.380 ;
        RECT 2926.600 2889.370 2929.600 2889.380 ;
        RECT -9.980 2712.380 -6.980 2712.390 ;
        RECT 4.020 2712.380 7.020 2712.390 ;
        RECT 184.020 2712.380 187.020 2712.390 ;
        RECT 364.020 2712.380 367.020 2712.390 ;
        RECT 544.020 2712.380 547.020 2712.390 ;
        RECT 724.020 2712.380 727.020 2712.390 ;
        RECT 904.020 2712.380 907.020 2712.390 ;
        RECT 1084.020 2712.380 1087.020 2712.390 ;
        RECT 1264.020 2712.380 1267.020 2712.390 ;
        RECT 1444.020 2712.380 1447.020 2712.390 ;
        RECT 1624.020 2712.380 1627.020 2712.390 ;
        RECT 1804.020 2712.380 1807.020 2712.390 ;
        RECT 1984.020 2712.380 1987.020 2712.390 ;
        RECT 2164.020 2712.380 2167.020 2712.390 ;
        RECT 2344.020 2712.380 2347.020 2712.390 ;
        RECT 2524.020 2712.380 2527.020 2712.390 ;
        RECT 2704.020 2712.380 2707.020 2712.390 ;
        RECT 2884.020 2712.380 2887.020 2712.390 ;
        RECT 2926.600 2712.380 2929.600 2712.390 ;
        RECT -14.580 2709.380 2934.200 2712.380 ;
        RECT -9.980 2709.370 -6.980 2709.380 ;
        RECT 4.020 2709.370 7.020 2709.380 ;
        RECT 184.020 2709.370 187.020 2709.380 ;
        RECT 364.020 2709.370 367.020 2709.380 ;
        RECT 544.020 2709.370 547.020 2709.380 ;
        RECT 724.020 2709.370 727.020 2709.380 ;
        RECT 904.020 2709.370 907.020 2709.380 ;
        RECT 1084.020 2709.370 1087.020 2709.380 ;
        RECT 1264.020 2709.370 1267.020 2709.380 ;
        RECT 1444.020 2709.370 1447.020 2709.380 ;
        RECT 1624.020 2709.370 1627.020 2709.380 ;
        RECT 1804.020 2709.370 1807.020 2709.380 ;
        RECT 1984.020 2709.370 1987.020 2709.380 ;
        RECT 2164.020 2709.370 2167.020 2709.380 ;
        RECT 2344.020 2709.370 2347.020 2709.380 ;
        RECT 2524.020 2709.370 2527.020 2709.380 ;
        RECT 2704.020 2709.370 2707.020 2709.380 ;
        RECT 2884.020 2709.370 2887.020 2709.380 ;
        RECT 2926.600 2709.370 2929.600 2709.380 ;
        RECT -9.980 2532.380 -6.980 2532.390 ;
        RECT 4.020 2532.380 7.020 2532.390 ;
        RECT 184.020 2532.380 187.020 2532.390 ;
        RECT 364.020 2532.380 367.020 2532.390 ;
        RECT 544.020 2532.380 547.020 2532.390 ;
        RECT 724.020 2532.380 727.020 2532.390 ;
        RECT 904.020 2532.380 907.020 2532.390 ;
        RECT 1084.020 2532.380 1087.020 2532.390 ;
        RECT 1264.020 2532.380 1267.020 2532.390 ;
        RECT 1444.020 2532.380 1447.020 2532.390 ;
        RECT 1624.020 2532.380 1627.020 2532.390 ;
        RECT 1804.020 2532.380 1807.020 2532.390 ;
        RECT 1984.020 2532.380 1987.020 2532.390 ;
        RECT 2164.020 2532.380 2167.020 2532.390 ;
        RECT 2344.020 2532.380 2347.020 2532.390 ;
        RECT 2524.020 2532.380 2527.020 2532.390 ;
        RECT 2704.020 2532.380 2707.020 2532.390 ;
        RECT 2884.020 2532.380 2887.020 2532.390 ;
        RECT 2926.600 2532.380 2929.600 2532.390 ;
        RECT -14.580 2529.380 2934.200 2532.380 ;
        RECT -9.980 2529.370 -6.980 2529.380 ;
        RECT 4.020 2529.370 7.020 2529.380 ;
        RECT 184.020 2529.370 187.020 2529.380 ;
        RECT 364.020 2529.370 367.020 2529.380 ;
        RECT 544.020 2529.370 547.020 2529.380 ;
        RECT 724.020 2529.370 727.020 2529.380 ;
        RECT 904.020 2529.370 907.020 2529.380 ;
        RECT 1084.020 2529.370 1087.020 2529.380 ;
        RECT 1264.020 2529.370 1267.020 2529.380 ;
        RECT 1444.020 2529.370 1447.020 2529.380 ;
        RECT 1624.020 2529.370 1627.020 2529.380 ;
        RECT 1804.020 2529.370 1807.020 2529.380 ;
        RECT 1984.020 2529.370 1987.020 2529.380 ;
        RECT 2164.020 2529.370 2167.020 2529.380 ;
        RECT 2344.020 2529.370 2347.020 2529.380 ;
        RECT 2524.020 2529.370 2527.020 2529.380 ;
        RECT 2704.020 2529.370 2707.020 2529.380 ;
        RECT 2884.020 2529.370 2887.020 2529.380 ;
        RECT 2926.600 2529.370 2929.600 2529.380 ;
        RECT -9.980 2352.380 -6.980 2352.390 ;
        RECT 4.020 2352.380 7.020 2352.390 ;
        RECT 184.020 2352.380 187.020 2352.390 ;
        RECT 364.020 2352.380 367.020 2352.390 ;
        RECT 544.020 2352.380 547.020 2352.390 ;
        RECT 724.020 2352.380 727.020 2352.390 ;
        RECT 904.020 2352.380 907.020 2352.390 ;
        RECT 1084.020 2352.380 1087.020 2352.390 ;
        RECT 1264.020 2352.380 1267.020 2352.390 ;
        RECT 1444.020 2352.380 1447.020 2352.390 ;
        RECT 1624.020 2352.380 1627.020 2352.390 ;
        RECT 1804.020 2352.380 1807.020 2352.390 ;
        RECT 1984.020 2352.380 1987.020 2352.390 ;
        RECT 2164.020 2352.380 2167.020 2352.390 ;
        RECT 2344.020 2352.380 2347.020 2352.390 ;
        RECT 2524.020 2352.380 2527.020 2352.390 ;
        RECT 2704.020 2352.380 2707.020 2352.390 ;
        RECT 2884.020 2352.380 2887.020 2352.390 ;
        RECT 2926.600 2352.380 2929.600 2352.390 ;
        RECT -14.580 2349.380 2934.200 2352.380 ;
        RECT -9.980 2349.370 -6.980 2349.380 ;
        RECT 4.020 2349.370 7.020 2349.380 ;
        RECT 184.020 2349.370 187.020 2349.380 ;
        RECT 364.020 2349.370 367.020 2349.380 ;
        RECT 544.020 2349.370 547.020 2349.380 ;
        RECT 724.020 2349.370 727.020 2349.380 ;
        RECT 904.020 2349.370 907.020 2349.380 ;
        RECT 1084.020 2349.370 1087.020 2349.380 ;
        RECT 1264.020 2349.370 1267.020 2349.380 ;
        RECT 1444.020 2349.370 1447.020 2349.380 ;
        RECT 1624.020 2349.370 1627.020 2349.380 ;
        RECT 1804.020 2349.370 1807.020 2349.380 ;
        RECT 1984.020 2349.370 1987.020 2349.380 ;
        RECT 2164.020 2349.370 2167.020 2349.380 ;
        RECT 2344.020 2349.370 2347.020 2349.380 ;
        RECT 2524.020 2349.370 2527.020 2349.380 ;
        RECT 2704.020 2349.370 2707.020 2349.380 ;
        RECT 2884.020 2349.370 2887.020 2349.380 ;
        RECT 2926.600 2349.370 2929.600 2349.380 ;
        RECT -9.980 2172.380 -6.980 2172.390 ;
        RECT 4.020 2172.380 7.020 2172.390 ;
        RECT 184.020 2172.380 187.020 2172.390 ;
        RECT 364.020 2172.380 367.020 2172.390 ;
        RECT 544.020 2172.380 547.020 2172.390 ;
        RECT 724.020 2172.380 727.020 2172.390 ;
        RECT 904.020 2172.380 907.020 2172.390 ;
        RECT 1084.020 2172.380 1087.020 2172.390 ;
        RECT 1264.020 2172.380 1267.020 2172.390 ;
        RECT 1444.020 2172.380 1447.020 2172.390 ;
        RECT 1624.020 2172.380 1627.020 2172.390 ;
        RECT 1804.020 2172.380 1807.020 2172.390 ;
        RECT 1984.020 2172.380 1987.020 2172.390 ;
        RECT 2164.020 2172.380 2167.020 2172.390 ;
        RECT 2344.020 2172.380 2347.020 2172.390 ;
        RECT 2524.020 2172.380 2527.020 2172.390 ;
        RECT 2704.020 2172.380 2707.020 2172.390 ;
        RECT 2884.020 2172.380 2887.020 2172.390 ;
        RECT 2926.600 2172.380 2929.600 2172.390 ;
        RECT -14.580 2169.380 2934.200 2172.380 ;
        RECT -9.980 2169.370 -6.980 2169.380 ;
        RECT 4.020 2169.370 7.020 2169.380 ;
        RECT 184.020 2169.370 187.020 2169.380 ;
        RECT 364.020 2169.370 367.020 2169.380 ;
        RECT 544.020 2169.370 547.020 2169.380 ;
        RECT 724.020 2169.370 727.020 2169.380 ;
        RECT 904.020 2169.370 907.020 2169.380 ;
        RECT 1084.020 2169.370 1087.020 2169.380 ;
        RECT 1264.020 2169.370 1267.020 2169.380 ;
        RECT 1444.020 2169.370 1447.020 2169.380 ;
        RECT 1624.020 2169.370 1627.020 2169.380 ;
        RECT 1804.020 2169.370 1807.020 2169.380 ;
        RECT 1984.020 2169.370 1987.020 2169.380 ;
        RECT 2164.020 2169.370 2167.020 2169.380 ;
        RECT 2344.020 2169.370 2347.020 2169.380 ;
        RECT 2524.020 2169.370 2527.020 2169.380 ;
        RECT 2704.020 2169.370 2707.020 2169.380 ;
        RECT 2884.020 2169.370 2887.020 2169.380 ;
        RECT 2926.600 2169.370 2929.600 2169.380 ;
        RECT -9.980 1992.380 -6.980 1992.390 ;
        RECT 4.020 1992.380 7.020 1992.390 ;
        RECT 184.020 1992.380 187.020 1992.390 ;
        RECT 364.020 1992.380 367.020 1992.390 ;
        RECT 544.020 1992.380 547.020 1992.390 ;
        RECT 724.020 1992.380 727.020 1992.390 ;
        RECT 904.020 1992.380 907.020 1992.390 ;
        RECT 1084.020 1992.380 1087.020 1992.390 ;
        RECT 1264.020 1992.380 1267.020 1992.390 ;
        RECT 1444.020 1992.380 1447.020 1992.390 ;
        RECT 1624.020 1992.380 1627.020 1992.390 ;
        RECT 1804.020 1992.380 1807.020 1992.390 ;
        RECT 1984.020 1992.380 1987.020 1992.390 ;
        RECT 2164.020 1992.380 2167.020 1992.390 ;
        RECT 2344.020 1992.380 2347.020 1992.390 ;
        RECT 2524.020 1992.380 2527.020 1992.390 ;
        RECT 2704.020 1992.380 2707.020 1992.390 ;
        RECT 2884.020 1992.380 2887.020 1992.390 ;
        RECT 2926.600 1992.380 2929.600 1992.390 ;
        RECT -14.580 1989.380 2934.200 1992.380 ;
        RECT -9.980 1989.370 -6.980 1989.380 ;
        RECT 4.020 1989.370 7.020 1989.380 ;
        RECT 184.020 1989.370 187.020 1989.380 ;
        RECT 364.020 1989.370 367.020 1989.380 ;
        RECT 544.020 1989.370 547.020 1989.380 ;
        RECT 724.020 1989.370 727.020 1989.380 ;
        RECT 904.020 1989.370 907.020 1989.380 ;
        RECT 1084.020 1989.370 1087.020 1989.380 ;
        RECT 1264.020 1989.370 1267.020 1989.380 ;
        RECT 1444.020 1989.370 1447.020 1989.380 ;
        RECT 1624.020 1989.370 1627.020 1989.380 ;
        RECT 1804.020 1989.370 1807.020 1989.380 ;
        RECT 1984.020 1989.370 1987.020 1989.380 ;
        RECT 2164.020 1989.370 2167.020 1989.380 ;
        RECT 2344.020 1989.370 2347.020 1989.380 ;
        RECT 2524.020 1989.370 2527.020 1989.380 ;
        RECT 2704.020 1989.370 2707.020 1989.380 ;
        RECT 2884.020 1989.370 2887.020 1989.380 ;
        RECT 2926.600 1989.370 2929.600 1989.380 ;
        RECT -9.980 1812.380 -6.980 1812.390 ;
        RECT 4.020 1812.380 7.020 1812.390 ;
        RECT 184.020 1812.380 187.020 1812.390 ;
        RECT 364.020 1812.380 367.020 1812.390 ;
        RECT 544.020 1812.380 547.020 1812.390 ;
        RECT 724.020 1812.380 727.020 1812.390 ;
        RECT 904.020 1812.380 907.020 1812.390 ;
        RECT 1084.020 1812.380 1087.020 1812.390 ;
        RECT 1264.020 1812.380 1267.020 1812.390 ;
        RECT 1444.020 1812.380 1447.020 1812.390 ;
        RECT 1624.020 1812.380 1627.020 1812.390 ;
        RECT 1804.020 1812.380 1807.020 1812.390 ;
        RECT 1984.020 1812.380 1987.020 1812.390 ;
        RECT 2164.020 1812.380 2167.020 1812.390 ;
        RECT 2344.020 1812.380 2347.020 1812.390 ;
        RECT 2524.020 1812.380 2527.020 1812.390 ;
        RECT 2704.020 1812.380 2707.020 1812.390 ;
        RECT 2884.020 1812.380 2887.020 1812.390 ;
        RECT 2926.600 1812.380 2929.600 1812.390 ;
        RECT -14.580 1809.380 2934.200 1812.380 ;
        RECT -9.980 1809.370 -6.980 1809.380 ;
        RECT 4.020 1809.370 7.020 1809.380 ;
        RECT 184.020 1809.370 187.020 1809.380 ;
        RECT 364.020 1809.370 367.020 1809.380 ;
        RECT 544.020 1809.370 547.020 1809.380 ;
        RECT 724.020 1809.370 727.020 1809.380 ;
        RECT 904.020 1809.370 907.020 1809.380 ;
        RECT 1084.020 1809.370 1087.020 1809.380 ;
        RECT 1264.020 1809.370 1267.020 1809.380 ;
        RECT 1444.020 1809.370 1447.020 1809.380 ;
        RECT 1624.020 1809.370 1627.020 1809.380 ;
        RECT 1804.020 1809.370 1807.020 1809.380 ;
        RECT 1984.020 1809.370 1987.020 1809.380 ;
        RECT 2164.020 1809.370 2167.020 1809.380 ;
        RECT 2344.020 1809.370 2347.020 1809.380 ;
        RECT 2524.020 1809.370 2527.020 1809.380 ;
        RECT 2704.020 1809.370 2707.020 1809.380 ;
        RECT 2884.020 1809.370 2887.020 1809.380 ;
        RECT 2926.600 1809.370 2929.600 1809.380 ;
        RECT -9.980 1632.380 -6.980 1632.390 ;
        RECT 4.020 1632.380 7.020 1632.390 ;
        RECT 184.020 1632.380 187.020 1632.390 ;
        RECT 364.020 1632.380 367.020 1632.390 ;
        RECT 544.020 1632.380 547.020 1632.390 ;
        RECT 724.020 1632.380 727.020 1632.390 ;
        RECT 904.020 1632.380 907.020 1632.390 ;
        RECT 1084.020 1632.380 1087.020 1632.390 ;
        RECT 1264.020 1632.380 1267.020 1632.390 ;
        RECT 1444.020 1632.380 1447.020 1632.390 ;
        RECT 1624.020 1632.380 1627.020 1632.390 ;
        RECT 1804.020 1632.380 1807.020 1632.390 ;
        RECT 1984.020 1632.380 1987.020 1632.390 ;
        RECT 2164.020 1632.380 2167.020 1632.390 ;
        RECT 2344.020 1632.380 2347.020 1632.390 ;
        RECT 2524.020 1632.380 2527.020 1632.390 ;
        RECT 2704.020 1632.380 2707.020 1632.390 ;
        RECT 2884.020 1632.380 2887.020 1632.390 ;
        RECT 2926.600 1632.380 2929.600 1632.390 ;
        RECT -14.580 1629.380 2934.200 1632.380 ;
        RECT -9.980 1629.370 -6.980 1629.380 ;
        RECT 4.020 1629.370 7.020 1629.380 ;
        RECT 184.020 1629.370 187.020 1629.380 ;
        RECT 364.020 1629.370 367.020 1629.380 ;
        RECT 544.020 1629.370 547.020 1629.380 ;
        RECT 724.020 1629.370 727.020 1629.380 ;
        RECT 904.020 1629.370 907.020 1629.380 ;
        RECT 1084.020 1629.370 1087.020 1629.380 ;
        RECT 1264.020 1629.370 1267.020 1629.380 ;
        RECT 1444.020 1629.370 1447.020 1629.380 ;
        RECT 1624.020 1629.370 1627.020 1629.380 ;
        RECT 1804.020 1629.370 1807.020 1629.380 ;
        RECT 1984.020 1629.370 1987.020 1629.380 ;
        RECT 2164.020 1629.370 2167.020 1629.380 ;
        RECT 2344.020 1629.370 2347.020 1629.380 ;
        RECT 2524.020 1629.370 2527.020 1629.380 ;
        RECT 2704.020 1629.370 2707.020 1629.380 ;
        RECT 2884.020 1629.370 2887.020 1629.380 ;
        RECT 2926.600 1629.370 2929.600 1629.380 ;
        RECT -9.980 1452.380 -6.980 1452.390 ;
        RECT 4.020 1452.380 7.020 1452.390 ;
        RECT 184.020 1452.380 187.020 1452.390 ;
        RECT 364.020 1452.380 367.020 1452.390 ;
        RECT 544.020 1452.380 547.020 1452.390 ;
        RECT 724.020 1452.380 727.020 1452.390 ;
        RECT 904.020 1452.380 907.020 1452.390 ;
        RECT 1084.020 1452.380 1087.020 1452.390 ;
        RECT 1264.020 1452.380 1267.020 1452.390 ;
        RECT 1444.020 1452.380 1447.020 1452.390 ;
        RECT 1624.020 1452.380 1627.020 1452.390 ;
        RECT 1804.020 1452.380 1807.020 1452.390 ;
        RECT 1984.020 1452.380 1987.020 1452.390 ;
        RECT 2164.020 1452.380 2167.020 1452.390 ;
        RECT 2344.020 1452.380 2347.020 1452.390 ;
        RECT 2524.020 1452.380 2527.020 1452.390 ;
        RECT 2704.020 1452.380 2707.020 1452.390 ;
        RECT 2884.020 1452.380 2887.020 1452.390 ;
        RECT 2926.600 1452.380 2929.600 1452.390 ;
        RECT -14.580 1449.380 2934.200 1452.380 ;
        RECT -9.980 1449.370 -6.980 1449.380 ;
        RECT 4.020 1449.370 7.020 1449.380 ;
        RECT 184.020 1449.370 187.020 1449.380 ;
        RECT 364.020 1449.370 367.020 1449.380 ;
        RECT 544.020 1449.370 547.020 1449.380 ;
        RECT 724.020 1449.370 727.020 1449.380 ;
        RECT 904.020 1449.370 907.020 1449.380 ;
        RECT 1084.020 1449.370 1087.020 1449.380 ;
        RECT 1264.020 1449.370 1267.020 1449.380 ;
        RECT 1444.020 1449.370 1447.020 1449.380 ;
        RECT 1624.020 1449.370 1627.020 1449.380 ;
        RECT 1804.020 1449.370 1807.020 1449.380 ;
        RECT 1984.020 1449.370 1987.020 1449.380 ;
        RECT 2164.020 1449.370 2167.020 1449.380 ;
        RECT 2344.020 1449.370 2347.020 1449.380 ;
        RECT 2524.020 1449.370 2527.020 1449.380 ;
        RECT 2704.020 1449.370 2707.020 1449.380 ;
        RECT 2884.020 1449.370 2887.020 1449.380 ;
        RECT 2926.600 1449.370 2929.600 1449.380 ;
        RECT -9.980 1272.380 -6.980 1272.390 ;
        RECT 4.020 1272.380 7.020 1272.390 ;
        RECT 184.020 1272.380 187.020 1272.390 ;
        RECT 364.020 1272.380 367.020 1272.390 ;
        RECT 544.020 1272.380 547.020 1272.390 ;
        RECT 724.020 1272.380 727.020 1272.390 ;
        RECT 904.020 1272.380 907.020 1272.390 ;
        RECT 1084.020 1272.380 1087.020 1272.390 ;
        RECT 1264.020 1272.380 1267.020 1272.390 ;
        RECT 1444.020 1272.380 1447.020 1272.390 ;
        RECT 1624.020 1272.380 1627.020 1272.390 ;
        RECT 1804.020 1272.380 1807.020 1272.390 ;
        RECT 1984.020 1272.380 1987.020 1272.390 ;
        RECT 2164.020 1272.380 2167.020 1272.390 ;
        RECT 2344.020 1272.380 2347.020 1272.390 ;
        RECT 2524.020 1272.380 2527.020 1272.390 ;
        RECT 2704.020 1272.380 2707.020 1272.390 ;
        RECT 2884.020 1272.380 2887.020 1272.390 ;
        RECT 2926.600 1272.380 2929.600 1272.390 ;
        RECT -14.580 1269.380 2934.200 1272.380 ;
        RECT -9.980 1269.370 -6.980 1269.380 ;
        RECT 4.020 1269.370 7.020 1269.380 ;
        RECT 184.020 1269.370 187.020 1269.380 ;
        RECT 364.020 1269.370 367.020 1269.380 ;
        RECT 544.020 1269.370 547.020 1269.380 ;
        RECT 724.020 1269.370 727.020 1269.380 ;
        RECT 904.020 1269.370 907.020 1269.380 ;
        RECT 1084.020 1269.370 1087.020 1269.380 ;
        RECT 1264.020 1269.370 1267.020 1269.380 ;
        RECT 1444.020 1269.370 1447.020 1269.380 ;
        RECT 1624.020 1269.370 1627.020 1269.380 ;
        RECT 1804.020 1269.370 1807.020 1269.380 ;
        RECT 1984.020 1269.370 1987.020 1269.380 ;
        RECT 2164.020 1269.370 2167.020 1269.380 ;
        RECT 2344.020 1269.370 2347.020 1269.380 ;
        RECT 2524.020 1269.370 2527.020 1269.380 ;
        RECT 2704.020 1269.370 2707.020 1269.380 ;
        RECT 2884.020 1269.370 2887.020 1269.380 ;
        RECT 2926.600 1269.370 2929.600 1269.380 ;
        RECT -9.980 1092.380 -6.980 1092.390 ;
        RECT 4.020 1092.380 7.020 1092.390 ;
        RECT 184.020 1092.380 187.020 1092.390 ;
        RECT 364.020 1092.380 367.020 1092.390 ;
        RECT 544.020 1092.380 547.020 1092.390 ;
        RECT 724.020 1092.380 727.020 1092.390 ;
        RECT 904.020 1092.380 907.020 1092.390 ;
        RECT 1084.020 1092.380 1087.020 1092.390 ;
        RECT 1264.020 1092.380 1267.020 1092.390 ;
        RECT 1444.020 1092.380 1447.020 1092.390 ;
        RECT 1624.020 1092.380 1627.020 1092.390 ;
        RECT 1804.020 1092.380 1807.020 1092.390 ;
        RECT 1984.020 1092.380 1987.020 1092.390 ;
        RECT 2164.020 1092.380 2167.020 1092.390 ;
        RECT 2344.020 1092.380 2347.020 1092.390 ;
        RECT 2524.020 1092.380 2527.020 1092.390 ;
        RECT 2704.020 1092.380 2707.020 1092.390 ;
        RECT 2884.020 1092.380 2887.020 1092.390 ;
        RECT 2926.600 1092.380 2929.600 1092.390 ;
        RECT -14.580 1089.380 2934.200 1092.380 ;
        RECT -9.980 1089.370 -6.980 1089.380 ;
        RECT 4.020 1089.370 7.020 1089.380 ;
        RECT 184.020 1089.370 187.020 1089.380 ;
        RECT 364.020 1089.370 367.020 1089.380 ;
        RECT 544.020 1089.370 547.020 1089.380 ;
        RECT 724.020 1089.370 727.020 1089.380 ;
        RECT 904.020 1089.370 907.020 1089.380 ;
        RECT 1084.020 1089.370 1087.020 1089.380 ;
        RECT 1264.020 1089.370 1267.020 1089.380 ;
        RECT 1444.020 1089.370 1447.020 1089.380 ;
        RECT 1624.020 1089.370 1627.020 1089.380 ;
        RECT 1804.020 1089.370 1807.020 1089.380 ;
        RECT 1984.020 1089.370 1987.020 1089.380 ;
        RECT 2164.020 1089.370 2167.020 1089.380 ;
        RECT 2344.020 1089.370 2347.020 1089.380 ;
        RECT 2524.020 1089.370 2527.020 1089.380 ;
        RECT 2704.020 1089.370 2707.020 1089.380 ;
        RECT 2884.020 1089.370 2887.020 1089.380 ;
        RECT 2926.600 1089.370 2929.600 1089.380 ;
        RECT -9.980 912.380 -6.980 912.390 ;
        RECT 4.020 912.380 7.020 912.390 ;
        RECT 184.020 912.380 187.020 912.390 ;
        RECT 364.020 912.380 367.020 912.390 ;
        RECT 544.020 912.380 547.020 912.390 ;
        RECT 724.020 912.380 727.020 912.390 ;
        RECT 904.020 912.380 907.020 912.390 ;
        RECT 1084.020 912.380 1087.020 912.390 ;
        RECT 1264.020 912.380 1267.020 912.390 ;
        RECT 1444.020 912.380 1447.020 912.390 ;
        RECT 1624.020 912.380 1627.020 912.390 ;
        RECT 1804.020 912.380 1807.020 912.390 ;
        RECT 1984.020 912.380 1987.020 912.390 ;
        RECT 2164.020 912.380 2167.020 912.390 ;
        RECT 2344.020 912.380 2347.020 912.390 ;
        RECT 2524.020 912.380 2527.020 912.390 ;
        RECT 2704.020 912.380 2707.020 912.390 ;
        RECT 2884.020 912.380 2887.020 912.390 ;
        RECT 2926.600 912.380 2929.600 912.390 ;
        RECT -14.580 909.380 2934.200 912.380 ;
        RECT -9.980 909.370 -6.980 909.380 ;
        RECT 4.020 909.370 7.020 909.380 ;
        RECT 184.020 909.370 187.020 909.380 ;
        RECT 364.020 909.370 367.020 909.380 ;
        RECT 544.020 909.370 547.020 909.380 ;
        RECT 724.020 909.370 727.020 909.380 ;
        RECT 904.020 909.370 907.020 909.380 ;
        RECT 1084.020 909.370 1087.020 909.380 ;
        RECT 1264.020 909.370 1267.020 909.380 ;
        RECT 1444.020 909.370 1447.020 909.380 ;
        RECT 1624.020 909.370 1627.020 909.380 ;
        RECT 1804.020 909.370 1807.020 909.380 ;
        RECT 1984.020 909.370 1987.020 909.380 ;
        RECT 2164.020 909.370 2167.020 909.380 ;
        RECT 2344.020 909.370 2347.020 909.380 ;
        RECT 2524.020 909.370 2527.020 909.380 ;
        RECT 2704.020 909.370 2707.020 909.380 ;
        RECT 2884.020 909.370 2887.020 909.380 ;
        RECT 2926.600 909.370 2929.600 909.380 ;
        RECT -9.980 732.380 -6.980 732.390 ;
        RECT 4.020 732.380 7.020 732.390 ;
        RECT 184.020 732.380 187.020 732.390 ;
        RECT 364.020 732.380 367.020 732.390 ;
        RECT 544.020 732.380 547.020 732.390 ;
        RECT 724.020 732.380 727.020 732.390 ;
        RECT 904.020 732.380 907.020 732.390 ;
        RECT 1084.020 732.380 1087.020 732.390 ;
        RECT 1264.020 732.380 1267.020 732.390 ;
        RECT 1444.020 732.380 1447.020 732.390 ;
        RECT 1624.020 732.380 1627.020 732.390 ;
        RECT 1804.020 732.380 1807.020 732.390 ;
        RECT 1984.020 732.380 1987.020 732.390 ;
        RECT 2164.020 732.380 2167.020 732.390 ;
        RECT 2344.020 732.380 2347.020 732.390 ;
        RECT 2524.020 732.380 2527.020 732.390 ;
        RECT 2704.020 732.380 2707.020 732.390 ;
        RECT 2884.020 732.380 2887.020 732.390 ;
        RECT 2926.600 732.380 2929.600 732.390 ;
        RECT -14.580 729.380 2934.200 732.380 ;
        RECT -9.980 729.370 -6.980 729.380 ;
        RECT 4.020 729.370 7.020 729.380 ;
        RECT 184.020 729.370 187.020 729.380 ;
        RECT 364.020 729.370 367.020 729.380 ;
        RECT 544.020 729.370 547.020 729.380 ;
        RECT 724.020 729.370 727.020 729.380 ;
        RECT 904.020 729.370 907.020 729.380 ;
        RECT 1084.020 729.370 1087.020 729.380 ;
        RECT 1264.020 729.370 1267.020 729.380 ;
        RECT 1444.020 729.370 1447.020 729.380 ;
        RECT 1624.020 729.370 1627.020 729.380 ;
        RECT 1804.020 729.370 1807.020 729.380 ;
        RECT 1984.020 729.370 1987.020 729.380 ;
        RECT 2164.020 729.370 2167.020 729.380 ;
        RECT 2344.020 729.370 2347.020 729.380 ;
        RECT 2524.020 729.370 2527.020 729.380 ;
        RECT 2704.020 729.370 2707.020 729.380 ;
        RECT 2884.020 729.370 2887.020 729.380 ;
        RECT 2926.600 729.370 2929.600 729.380 ;
        RECT -9.980 552.380 -6.980 552.390 ;
        RECT 4.020 552.380 7.020 552.390 ;
        RECT 184.020 552.380 187.020 552.390 ;
        RECT 364.020 552.380 367.020 552.390 ;
        RECT 544.020 552.380 547.020 552.390 ;
        RECT 724.020 552.380 727.020 552.390 ;
        RECT 904.020 552.380 907.020 552.390 ;
        RECT 1084.020 552.380 1087.020 552.390 ;
        RECT 1264.020 552.380 1267.020 552.390 ;
        RECT 1444.020 552.380 1447.020 552.390 ;
        RECT 1624.020 552.380 1627.020 552.390 ;
        RECT 1804.020 552.380 1807.020 552.390 ;
        RECT 1984.020 552.380 1987.020 552.390 ;
        RECT 2164.020 552.380 2167.020 552.390 ;
        RECT 2344.020 552.380 2347.020 552.390 ;
        RECT 2524.020 552.380 2527.020 552.390 ;
        RECT 2704.020 552.380 2707.020 552.390 ;
        RECT 2884.020 552.380 2887.020 552.390 ;
        RECT 2926.600 552.380 2929.600 552.390 ;
        RECT -14.580 549.380 2934.200 552.380 ;
        RECT -9.980 549.370 -6.980 549.380 ;
        RECT 4.020 549.370 7.020 549.380 ;
        RECT 184.020 549.370 187.020 549.380 ;
        RECT 364.020 549.370 367.020 549.380 ;
        RECT 544.020 549.370 547.020 549.380 ;
        RECT 724.020 549.370 727.020 549.380 ;
        RECT 904.020 549.370 907.020 549.380 ;
        RECT 1084.020 549.370 1087.020 549.380 ;
        RECT 1264.020 549.370 1267.020 549.380 ;
        RECT 1444.020 549.370 1447.020 549.380 ;
        RECT 1624.020 549.370 1627.020 549.380 ;
        RECT 1804.020 549.370 1807.020 549.380 ;
        RECT 1984.020 549.370 1987.020 549.380 ;
        RECT 2164.020 549.370 2167.020 549.380 ;
        RECT 2344.020 549.370 2347.020 549.380 ;
        RECT 2524.020 549.370 2527.020 549.380 ;
        RECT 2704.020 549.370 2707.020 549.380 ;
        RECT 2884.020 549.370 2887.020 549.380 ;
        RECT 2926.600 549.370 2929.600 549.380 ;
        RECT -9.980 372.380 -6.980 372.390 ;
        RECT 4.020 372.380 7.020 372.390 ;
        RECT 184.020 372.380 187.020 372.390 ;
        RECT 364.020 372.380 367.020 372.390 ;
        RECT 544.020 372.380 547.020 372.390 ;
        RECT 724.020 372.380 727.020 372.390 ;
        RECT 904.020 372.380 907.020 372.390 ;
        RECT 1084.020 372.380 1087.020 372.390 ;
        RECT 1264.020 372.380 1267.020 372.390 ;
        RECT 1444.020 372.380 1447.020 372.390 ;
        RECT 1624.020 372.380 1627.020 372.390 ;
        RECT 1804.020 372.380 1807.020 372.390 ;
        RECT 1984.020 372.380 1987.020 372.390 ;
        RECT 2164.020 372.380 2167.020 372.390 ;
        RECT 2344.020 372.380 2347.020 372.390 ;
        RECT 2524.020 372.380 2527.020 372.390 ;
        RECT 2704.020 372.380 2707.020 372.390 ;
        RECT 2884.020 372.380 2887.020 372.390 ;
        RECT 2926.600 372.380 2929.600 372.390 ;
        RECT -14.580 369.380 2934.200 372.380 ;
        RECT -9.980 369.370 -6.980 369.380 ;
        RECT 4.020 369.370 7.020 369.380 ;
        RECT 184.020 369.370 187.020 369.380 ;
        RECT 364.020 369.370 367.020 369.380 ;
        RECT 544.020 369.370 547.020 369.380 ;
        RECT 724.020 369.370 727.020 369.380 ;
        RECT 904.020 369.370 907.020 369.380 ;
        RECT 1084.020 369.370 1087.020 369.380 ;
        RECT 1264.020 369.370 1267.020 369.380 ;
        RECT 1444.020 369.370 1447.020 369.380 ;
        RECT 1624.020 369.370 1627.020 369.380 ;
        RECT 1804.020 369.370 1807.020 369.380 ;
        RECT 1984.020 369.370 1987.020 369.380 ;
        RECT 2164.020 369.370 2167.020 369.380 ;
        RECT 2344.020 369.370 2347.020 369.380 ;
        RECT 2524.020 369.370 2527.020 369.380 ;
        RECT 2704.020 369.370 2707.020 369.380 ;
        RECT 2884.020 369.370 2887.020 369.380 ;
        RECT 2926.600 369.370 2929.600 369.380 ;
        RECT -9.980 192.380 -6.980 192.390 ;
        RECT 4.020 192.380 7.020 192.390 ;
        RECT 184.020 192.380 187.020 192.390 ;
        RECT 364.020 192.380 367.020 192.390 ;
        RECT 544.020 192.380 547.020 192.390 ;
        RECT 724.020 192.380 727.020 192.390 ;
        RECT 904.020 192.380 907.020 192.390 ;
        RECT 1084.020 192.380 1087.020 192.390 ;
        RECT 1264.020 192.380 1267.020 192.390 ;
        RECT 1444.020 192.380 1447.020 192.390 ;
        RECT 1624.020 192.380 1627.020 192.390 ;
        RECT 1804.020 192.380 1807.020 192.390 ;
        RECT 1984.020 192.380 1987.020 192.390 ;
        RECT 2164.020 192.380 2167.020 192.390 ;
        RECT 2344.020 192.380 2347.020 192.390 ;
        RECT 2524.020 192.380 2527.020 192.390 ;
        RECT 2704.020 192.380 2707.020 192.390 ;
        RECT 2884.020 192.380 2887.020 192.390 ;
        RECT 2926.600 192.380 2929.600 192.390 ;
        RECT -14.580 189.380 2934.200 192.380 ;
        RECT -9.980 189.370 -6.980 189.380 ;
        RECT 4.020 189.370 7.020 189.380 ;
        RECT 184.020 189.370 187.020 189.380 ;
        RECT 364.020 189.370 367.020 189.380 ;
        RECT 544.020 189.370 547.020 189.380 ;
        RECT 724.020 189.370 727.020 189.380 ;
        RECT 904.020 189.370 907.020 189.380 ;
        RECT 1084.020 189.370 1087.020 189.380 ;
        RECT 1264.020 189.370 1267.020 189.380 ;
        RECT 1444.020 189.370 1447.020 189.380 ;
        RECT 1624.020 189.370 1627.020 189.380 ;
        RECT 1804.020 189.370 1807.020 189.380 ;
        RECT 1984.020 189.370 1987.020 189.380 ;
        RECT 2164.020 189.370 2167.020 189.380 ;
        RECT 2344.020 189.370 2347.020 189.380 ;
        RECT 2524.020 189.370 2527.020 189.380 ;
        RECT 2704.020 189.370 2707.020 189.380 ;
        RECT 2884.020 189.370 2887.020 189.380 ;
        RECT 2926.600 189.370 2929.600 189.380 ;
        RECT -9.980 12.380 -6.980 12.390 ;
        RECT 4.020 12.380 7.020 12.390 ;
        RECT 184.020 12.380 187.020 12.390 ;
        RECT 364.020 12.380 367.020 12.390 ;
        RECT 544.020 12.380 547.020 12.390 ;
        RECT 724.020 12.380 727.020 12.390 ;
        RECT 904.020 12.380 907.020 12.390 ;
        RECT 1084.020 12.380 1087.020 12.390 ;
        RECT 1264.020 12.380 1267.020 12.390 ;
        RECT 1444.020 12.380 1447.020 12.390 ;
        RECT 1624.020 12.380 1627.020 12.390 ;
        RECT 1804.020 12.380 1807.020 12.390 ;
        RECT 1984.020 12.380 1987.020 12.390 ;
        RECT 2164.020 12.380 2167.020 12.390 ;
        RECT 2344.020 12.380 2347.020 12.390 ;
        RECT 2524.020 12.380 2527.020 12.390 ;
        RECT 2704.020 12.380 2707.020 12.390 ;
        RECT 2884.020 12.380 2887.020 12.390 ;
        RECT 2926.600 12.380 2929.600 12.390 ;
        RECT -14.580 9.380 2934.200 12.380 ;
        RECT -9.980 9.370 -6.980 9.380 ;
        RECT 4.020 9.370 7.020 9.380 ;
        RECT 184.020 9.370 187.020 9.380 ;
        RECT 364.020 9.370 367.020 9.380 ;
        RECT 544.020 9.370 547.020 9.380 ;
        RECT 724.020 9.370 727.020 9.380 ;
        RECT 904.020 9.370 907.020 9.380 ;
        RECT 1084.020 9.370 1087.020 9.380 ;
        RECT 1264.020 9.370 1267.020 9.380 ;
        RECT 1444.020 9.370 1447.020 9.380 ;
        RECT 1624.020 9.370 1627.020 9.380 ;
        RECT 1804.020 9.370 1807.020 9.380 ;
        RECT 1984.020 9.370 1987.020 9.380 ;
        RECT 2164.020 9.370 2167.020 9.380 ;
        RECT 2344.020 9.370 2347.020 9.380 ;
        RECT 2524.020 9.370 2527.020 9.380 ;
        RECT 2704.020 9.370 2707.020 9.380 ;
        RECT 2884.020 9.370 2887.020 9.380 ;
        RECT 2926.600 9.370 2929.600 9.380 ;
        RECT -9.980 -1.620 -6.980 -1.610 ;
        RECT 4.020 -1.620 7.020 -1.610 ;
        RECT 184.020 -1.620 187.020 -1.610 ;
        RECT 364.020 -1.620 367.020 -1.610 ;
        RECT 544.020 -1.620 547.020 -1.610 ;
        RECT 724.020 -1.620 727.020 -1.610 ;
        RECT 904.020 -1.620 907.020 -1.610 ;
        RECT 1084.020 -1.620 1087.020 -1.610 ;
        RECT 1264.020 -1.620 1267.020 -1.610 ;
        RECT 1444.020 -1.620 1447.020 -1.610 ;
        RECT 1624.020 -1.620 1627.020 -1.610 ;
        RECT 1804.020 -1.620 1807.020 -1.610 ;
        RECT 1984.020 -1.620 1987.020 -1.610 ;
        RECT 2164.020 -1.620 2167.020 -1.610 ;
        RECT 2344.020 -1.620 2347.020 -1.610 ;
        RECT 2524.020 -1.620 2527.020 -1.610 ;
        RECT 2704.020 -1.620 2707.020 -1.610 ;
        RECT 2884.020 -1.620 2887.020 -1.610 ;
        RECT 2926.600 -1.620 2929.600 -1.610 ;
        RECT -9.980 -4.620 2929.600 -1.620 ;
        RECT -9.980 -4.630 -6.980 -4.620 ;
        RECT 4.020 -4.630 7.020 -4.620 ;
        RECT 184.020 -4.630 187.020 -4.620 ;
        RECT 364.020 -4.630 367.020 -4.620 ;
        RECT 544.020 -4.630 547.020 -4.620 ;
        RECT 724.020 -4.630 727.020 -4.620 ;
        RECT 904.020 -4.630 907.020 -4.620 ;
        RECT 1084.020 -4.630 1087.020 -4.620 ;
        RECT 1264.020 -4.630 1267.020 -4.620 ;
        RECT 1444.020 -4.630 1447.020 -4.620 ;
        RECT 1624.020 -4.630 1627.020 -4.620 ;
        RECT 1804.020 -4.630 1807.020 -4.620 ;
        RECT 1984.020 -4.630 1987.020 -4.620 ;
        RECT 2164.020 -4.630 2167.020 -4.620 ;
        RECT 2344.020 -4.630 2347.020 -4.620 ;
        RECT 2524.020 -4.630 2527.020 -4.620 ;
        RECT 2704.020 -4.630 2707.020 -4.620 ;
        RECT 2884.020 -4.630 2887.020 -4.620 ;
        RECT 2926.600 -4.630 2929.600 -4.620 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -14.580 -9.220 -11.580 3528.900 ;
        RECT 94.020 -9.220 97.020 3528.900 ;
        RECT 274.020 -9.220 277.020 3528.900 ;
        RECT 454.020 -9.220 457.020 3528.900 ;
        RECT 634.020 -9.220 637.020 3528.900 ;
        RECT 814.020 -9.220 817.020 3528.900 ;
        RECT 994.020 -9.220 997.020 3528.900 ;
        RECT 1174.020 -9.220 1177.020 3528.900 ;
        RECT 1354.020 -9.220 1357.020 3528.900 ;
        RECT 1534.020 -9.220 1537.020 3528.900 ;
        RECT 1714.020 -9.220 1717.020 3528.900 ;
        RECT 1894.020 -9.220 1897.020 3528.900 ;
        RECT 2074.020 -9.220 2077.020 3528.900 ;
        RECT 2254.020 -9.220 2257.020 3528.900 ;
        RECT 2434.020 -9.220 2437.020 3528.900 ;
        RECT 2614.020 -9.220 2617.020 3528.900 ;
        RECT 2794.020 -9.220 2797.020 3528.900 ;
        RECT 2931.200 -9.220 2934.200 3528.900 ;
      LAYER via4 ;
        RECT -13.670 3527.610 -12.490 3528.790 ;
        RECT -13.670 3526.010 -12.490 3527.190 ;
        RECT -13.670 3341.090 -12.490 3342.270 ;
        RECT -13.670 3339.490 -12.490 3340.670 ;
        RECT -13.670 3161.090 -12.490 3162.270 ;
        RECT -13.670 3159.490 -12.490 3160.670 ;
        RECT -13.670 2981.090 -12.490 2982.270 ;
        RECT -13.670 2979.490 -12.490 2980.670 ;
        RECT -13.670 2801.090 -12.490 2802.270 ;
        RECT -13.670 2799.490 -12.490 2800.670 ;
        RECT -13.670 2621.090 -12.490 2622.270 ;
        RECT -13.670 2619.490 -12.490 2620.670 ;
        RECT -13.670 2441.090 -12.490 2442.270 ;
        RECT -13.670 2439.490 -12.490 2440.670 ;
        RECT -13.670 2261.090 -12.490 2262.270 ;
        RECT -13.670 2259.490 -12.490 2260.670 ;
        RECT -13.670 2081.090 -12.490 2082.270 ;
        RECT -13.670 2079.490 -12.490 2080.670 ;
        RECT -13.670 1901.090 -12.490 1902.270 ;
        RECT -13.670 1899.490 -12.490 1900.670 ;
        RECT -13.670 1721.090 -12.490 1722.270 ;
        RECT -13.670 1719.490 -12.490 1720.670 ;
        RECT -13.670 1541.090 -12.490 1542.270 ;
        RECT -13.670 1539.490 -12.490 1540.670 ;
        RECT -13.670 1361.090 -12.490 1362.270 ;
        RECT -13.670 1359.490 -12.490 1360.670 ;
        RECT -13.670 1181.090 -12.490 1182.270 ;
        RECT -13.670 1179.490 -12.490 1180.670 ;
        RECT -13.670 1001.090 -12.490 1002.270 ;
        RECT -13.670 999.490 -12.490 1000.670 ;
        RECT -13.670 821.090 -12.490 822.270 ;
        RECT -13.670 819.490 -12.490 820.670 ;
        RECT -13.670 641.090 -12.490 642.270 ;
        RECT -13.670 639.490 -12.490 640.670 ;
        RECT -13.670 461.090 -12.490 462.270 ;
        RECT -13.670 459.490 -12.490 460.670 ;
        RECT -13.670 281.090 -12.490 282.270 ;
        RECT -13.670 279.490 -12.490 280.670 ;
        RECT -13.670 101.090 -12.490 102.270 ;
        RECT -13.670 99.490 -12.490 100.670 ;
        RECT -13.670 -7.510 -12.490 -6.330 ;
        RECT -13.670 -9.110 -12.490 -7.930 ;
        RECT 94.930 3527.610 96.110 3528.790 ;
        RECT 94.930 3526.010 96.110 3527.190 ;
        RECT 94.930 3341.090 96.110 3342.270 ;
        RECT 94.930 3339.490 96.110 3340.670 ;
        RECT 94.930 3161.090 96.110 3162.270 ;
        RECT 94.930 3159.490 96.110 3160.670 ;
        RECT 94.930 2981.090 96.110 2982.270 ;
        RECT 94.930 2979.490 96.110 2980.670 ;
        RECT 94.930 2801.090 96.110 2802.270 ;
        RECT 94.930 2799.490 96.110 2800.670 ;
        RECT 94.930 2621.090 96.110 2622.270 ;
        RECT 94.930 2619.490 96.110 2620.670 ;
        RECT 94.930 2441.090 96.110 2442.270 ;
        RECT 94.930 2439.490 96.110 2440.670 ;
        RECT 94.930 2261.090 96.110 2262.270 ;
        RECT 94.930 2259.490 96.110 2260.670 ;
        RECT 94.930 2081.090 96.110 2082.270 ;
        RECT 94.930 2079.490 96.110 2080.670 ;
        RECT 94.930 1901.090 96.110 1902.270 ;
        RECT 94.930 1899.490 96.110 1900.670 ;
        RECT 94.930 1721.090 96.110 1722.270 ;
        RECT 94.930 1719.490 96.110 1720.670 ;
        RECT 94.930 1541.090 96.110 1542.270 ;
        RECT 94.930 1539.490 96.110 1540.670 ;
        RECT 94.930 1361.090 96.110 1362.270 ;
        RECT 94.930 1359.490 96.110 1360.670 ;
        RECT 94.930 1181.090 96.110 1182.270 ;
        RECT 94.930 1179.490 96.110 1180.670 ;
        RECT 94.930 1001.090 96.110 1002.270 ;
        RECT 94.930 999.490 96.110 1000.670 ;
        RECT 94.930 821.090 96.110 822.270 ;
        RECT 94.930 819.490 96.110 820.670 ;
        RECT 94.930 641.090 96.110 642.270 ;
        RECT 94.930 639.490 96.110 640.670 ;
        RECT 94.930 461.090 96.110 462.270 ;
        RECT 94.930 459.490 96.110 460.670 ;
        RECT 94.930 281.090 96.110 282.270 ;
        RECT 94.930 279.490 96.110 280.670 ;
        RECT 94.930 101.090 96.110 102.270 ;
        RECT 94.930 99.490 96.110 100.670 ;
        RECT 94.930 -7.510 96.110 -6.330 ;
        RECT 94.930 -9.110 96.110 -7.930 ;
        RECT 274.930 3527.610 276.110 3528.790 ;
        RECT 274.930 3526.010 276.110 3527.190 ;
        RECT 274.930 3341.090 276.110 3342.270 ;
        RECT 274.930 3339.490 276.110 3340.670 ;
        RECT 274.930 3161.090 276.110 3162.270 ;
        RECT 274.930 3159.490 276.110 3160.670 ;
        RECT 274.930 2981.090 276.110 2982.270 ;
        RECT 274.930 2979.490 276.110 2980.670 ;
        RECT 274.930 2801.090 276.110 2802.270 ;
        RECT 274.930 2799.490 276.110 2800.670 ;
        RECT 274.930 2621.090 276.110 2622.270 ;
        RECT 274.930 2619.490 276.110 2620.670 ;
        RECT 274.930 2441.090 276.110 2442.270 ;
        RECT 274.930 2439.490 276.110 2440.670 ;
        RECT 274.930 2261.090 276.110 2262.270 ;
        RECT 274.930 2259.490 276.110 2260.670 ;
        RECT 274.930 2081.090 276.110 2082.270 ;
        RECT 274.930 2079.490 276.110 2080.670 ;
        RECT 274.930 1901.090 276.110 1902.270 ;
        RECT 274.930 1899.490 276.110 1900.670 ;
        RECT 274.930 1721.090 276.110 1722.270 ;
        RECT 274.930 1719.490 276.110 1720.670 ;
        RECT 274.930 1541.090 276.110 1542.270 ;
        RECT 274.930 1539.490 276.110 1540.670 ;
        RECT 274.930 1361.090 276.110 1362.270 ;
        RECT 274.930 1359.490 276.110 1360.670 ;
        RECT 274.930 1181.090 276.110 1182.270 ;
        RECT 274.930 1179.490 276.110 1180.670 ;
        RECT 274.930 1001.090 276.110 1002.270 ;
        RECT 274.930 999.490 276.110 1000.670 ;
        RECT 274.930 821.090 276.110 822.270 ;
        RECT 274.930 819.490 276.110 820.670 ;
        RECT 274.930 641.090 276.110 642.270 ;
        RECT 274.930 639.490 276.110 640.670 ;
        RECT 274.930 461.090 276.110 462.270 ;
        RECT 274.930 459.490 276.110 460.670 ;
        RECT 274.930 281.090 276.110 282.270 ;
        RECT 274.930 279.490 276.110 280.670 ;
        RECT 274.930 101.090 276.110 102.270 ;
        RECT 274.930 99.490 276.110 100.670 ;
        RECT 274.930 -7.510 276.110 -6.330 ;
        RECT 274.930 -9.110 276.110 -7.930 ;
        RECT 454.930 3527.610 456.110 3528.790 ;
        RECT 454.930 3526.010 456.110 3527.190 ;
        RECT 454.930 3341.090 456.110 3342.270 ;
        RECT 454.930 3339.490 456.110 3340.670 ;
        RECT 454.930 3161.090 456.110 3162.270 ;
        RECT 454.930 3159.490 456.110 3160.670 ;
        RECT 454.930 2981.090 456.110 2982.270 ;
        RECT 454.930 2979.490 456.110 2980.670 ;
        RECT 454.930 2801.090 456.110 2802.270 ;
        RECT 454.930 2799.490 456.110 2800.670 ;
        RECT 454.930 2621.090 456.110 2622.270 ;
        RECT 454.930 2619.490 456.110 2620.670 ;
        RECT 454.930 2441.090 456.110 2442.270 ;
        RECT 454.930 2439.490 456.110 2440.670 ;
        RECT 454.930 2261.090 456.110 2262.270 ;
        RECT 454.930 2259.490 456.110 2260.670 ;
        RECT 454.930 2081.090 456.110 2082.270 ;
        RECT 454.930 2079.490 456.110 2080.670 ;
        RECT 454.930 1901.090 456.110 1902.270 ;
        RECT 454.930 1899.490 456.110 1900.670 ;
        RECT 454.930 1721.090 456.110 1722.270 ;
        RECT 454.930 1719.490 456.110 1720.670 ;
        RECT 454.930 1541.090 456.110 1542.270 ;
        RECT 454.930 1539.490 456.110 1540.670 ;
        RECT 454.930 1361.090 456.110 1362.270 ;
        RECT 454.930 1359.490 456.110 1360.670 ;
        RECT 454.930 1181.090 456.110 1182.270 ;
        RECT 454.930 1179.490 456.110 1180.670 ;
        RECT 454.930 1001.090 456.110 1002.270 ;
        RECT 454.930 999.490 456.110 1000.670 ;
        RECT 454.930 821.090 456.110 822.270 ;
        RECT 454.930 819.490 456.110 820.670 ;
        RECT 454.930 641.090 456.110 642.270 ;
        RECT 454.930 639.490 456.110 640.670 ;
        RECT 454.930 461.090 456.110 462.270 ;
        RECT 454.930 459.490 456.110 460.670 ;
        RECT 454.930 281.090 456.110 282.270 ;
        RECT 454.930 279.490 456.110 280.670 ;
        RECT 454.930 101.090 456.110 102.270 ;
        RECT 454.930 99.490 456.110 100.670 ;
        RECT 454.930 -7.510 456.110 -6.330 ;
        RECT 454.930 -9.110 456.110 -7.930 ;
        RECT 634.930 3527.610 636.110 3528.790 ;
        RECT 634.930 3526.010 636.110 3527.190 ;
        RECT 634.930 3341.090 636.110 3342.270 ;
        RECT 634.930 3339.490 636.110 3340.670 ;
        RECT 634.930 3161.090 636.110 3162.270 ;
        RECT 634.930 3159.490 636.110 3160.670 ;
        RECT 634.930 2981.090 636.110 2982.270 ;
        RECT 634.930 2979.490 636.110 2980.670 ;
        RECT 634.930 2801.090 636.110 2802.270 ;
        RECT 634.930 2799.490 636.110 2800.670 ;
        RECT 634.930 2621.090 636.110 2622.270 ;
        RECT 634.930 2619.490 636.110 2620.670 ;
        RECT 634.930 2441.090 636.110 2442.270 ;
        RECT 634.930 2439.490 636.110 2440.670 ;
        RECT 634.930 2261.090 636.110 2262.270 ;
        RECT 634.930 2259.490 636.110 2260.670 ;
        RECT 634.930 2081.090 636.110 2082.270 ;
        RECT 634.930 2079.490 636.110 2080.670 ;
        RECT 634.930 1901.090 636.110 1902.270 ;
        RECT 634.930 1899.490 636.110 1900.670 ;
        RECT 634.930 1721.090 636.110 1722.270 ;
        RECT 634.930 1719.490 636.110 1720.670 ;
        RECT 634.930 1541.090 636.110 1542.270 ;
        RECT 634.930 1539.490 636.110 1540.670 ;
        RECT 634.930 1361.090 636.110 1362.270 ;
        RECT 634.930 1359.490 636.110 1360.670 ;
        RECT 634.930 1181.090 636.110 1182.270 ;
        RECT 634.930 1179.490 636.110 1180.670 ;
        RECT 634.930 1001.090 636.110 1002.270 ;
        RECT 634.930 999.490 636.110 1000.670 ;
        RECT 634.930 821.090 636.110 822.270 ;
        RECT 634.930 819.490 636.110 820.670 ;
        RECT 634.930 641.090 636.110 642.270 ;
        RECT 634.930 639.490 636.110 640.670 ;
        RECT 634.930 461.090 636.110 462.270 ;
        RECT 634.930 459.490 636.110 460.670 ;
        RECT 634.930 281.090 636.110 282.270 ;
        RECT 634.930 279.490 636.110 280.670 ;
        RECT 634.930 101.090 636.110 102.270 ;
        RECT 634.930 99.490 636.110 100.670 ;
        RECT 634.930 -7.510 636.110 -6.330 ;
        RECT 634.930 -9.110 636.110 -7.930 ;
        RECT 814.930 3527.610 816.110 3528.790 ;
        RECT 814.930 3526.010 816.110 3527.190 ;
        RECT 814.930 3341.090 816.110 3342.270 ;
        RECT 814.930 3339.490 816.110 3340.670 ;
        RECT 814.930 3161.090 816.110 3162.270 ;
        RECT 814.930 3159.490 816.110 3160.670 ;
        RECT 814.930 2981.090 816.110 2982.270 ;
        RECT 814.930 2979.490 816.110 2980.670 ;
        RECT 814.930 2801.090 816.110 2802.270 ;
        RECT 814.930 2799.490 816.110 2800.670 ;
        RECT 814.930 2621.090 816.110 2622.270 ;
        RECT 814.930 2619.490 816.110 2620.670 ;
        RECT 814.930 2441.090 816.110 2442.270 ;
        RECT 814.930 2439.490 816.110 2440.670 ;
        RECT 814.930 2261.090 816.110 2262.270 ;
        RECT 814.930 2259.490 816.110 2260.670 ;
        RECT 814.930 2081.090 816.110 2082.270 ;
        RECT 814.930 2079.490 816.110 2080.670 ;
        RECT 814.930 1901.090 816.110 1902.270 ;
        RECT 814.930 1899.490 816.110 1900.670 ;
        RECT 814.930 1721.090 816.110 1722.270 ;
        RECT 814.930 1719.490 816.110 1720.670 ;
        RECT 814.930 1541.090 816.110 1542.270 ;
        RECT 814.930 1539.490 816.110 1540.670 ;
        RECT 814.930 1361.090 816.110 1362.270 ;
        RECT 814.930 1359.490 816.110 1360.670 ;
        RECT 814.930 1181.090 816.110 1182.270 ;
        RECT 814.930 1179.490 816.110 1180.670 ;
        RECT 814.930 1001.090 816.110 1002.270 ;
        RECT 814.930 999.490 816.110 1000.670 ;
        RECT 814.930 821.090 816.110 822.270 ;
        RECT 814.930 819.490 816.110 820.670 ;
        RECT 814.930 641.090 816.110 642.270 ;
        RECT 814.930 639.490 816.110 640.670 ;
        RECT 814.930 461.090 816.110 462.270 ;
        RECT 814.930 459.490 816.110 460.670 ;
        RECT 814.930 281.090 816.110 282.270 ;
        RECT 814.930 279.490 816.110 280.670 ;
        RECT 814.930 101.090 816.110 102.270 ;
        RECT 814.930 99.490 816.110 100.670 ;
        RECT 814.930 -7.510 816.110 -6.330 ;
        RECT 814.930 -9.110 816.110 -7.930 ;
        RECT 994.930 3527.610 996.110 3528.790 ;
        RECT 994.930 3526.010 996.110 3527.190 ;
        RECT 994.930 3341.090 996.110 3342.270 ;
        RECT 994.930 3339.490 996.110 3340.670 ;
        RECT 994.930 3161.090 996.110 3162.270 ;
        RECT 994.930 3159.490 996.110 3160.670 ;
        RECT 994.930 2981.090 996.110 2982.270 ;
        RECT 994.930 2979.490 996.110 2980.670 ;
        RECT 994.930 2801.090 996.110 2802.270 ;
        RECT 994.930 2799.490 996.110 2800.670 ;
        RECT 994.930 2621.090 996.110 2622.270 ;
        RECT 994.930 2619.490 996.110 2620.670 ;
        RECT 994.930 2441.090 996.110 2442.270 ;
        RECT 994.930 2439.490 996.110 2440.670 ;
        RECT 994.930 2261.090 996.110 2262.270 ;
        RECT 994.930 2259.490 996.110 2260.670 ;
        RECT 994.930 2081.090 996.110 2082.270 ;
        RECT 994.930 2079.490 996.110 2080.670 ;
        RECT 994.930 1901.090 996.110 1902.270 ;
        RECT 994.930 1899.490 996.110 1900.670 ;
        RECT 994.930 1721.090 996.110 1722.270 ;
        RECT 994.930 1719.490 996.110 1720.670 ;
        RECT 994.930 1541.090 996.110 1542.270 ;
        RECT 994.930 1539.490 996.110 1540.670 ;
        RECT 994.930 1361.090 996.110 1362.270 ;
        RECT 994.930 1359.490 996.110 1360.670 ;
        RECT 994.930 1181.090 996.110 1182.270 ;
        RECT 994.930 1179.490 996.110 1180.670 ;
        RECT 994.930 1001.090 996.110 1002.270 ;
        RECT 994.930 999.490 996.110 1000.670 ;
        RECT 994.930 821.090 996.110 822.270 ;
        RECT 994.930 819.490 996.110 820.670 ;
        RECT 994.930 641.090 996.110 642.270 ;
        RECT 994.930 639.490 996.110 640.670 ;
        RECT 994.930 461.090 996.110 462.270 ;
        RECT 994.930 459.490 996.110 460.670 ;
        RECT 994.930 281.090 996.110 282.270 ;
        RECT 994.930 279.490 996.110 280.670 ;
        RECT 994.930 101.090 996.110 102.270 ;
        RECT 994.930 99.490 996.110 100.670 ;
        RECT 994.930 -7.510 996.110 -6.330 ;
        RECT 994.930 -9.110 996.110 -7.930 ;
        RECT 1174.930 3527.610 1176.110 3528.790 ;
        RECT 1174.930 3526.010 1176.110 3527.190 ;
        RECT 1174.930 3341.090 1176.110 3342.270 ;
        RECT 1174.930 3339.490 1176.110 3340.670 ;
        RECT 1174.930 3161.090 1176.110 3162.270 ;
        RECT 1174.930 3159.490 1176.110 3160.670 ;
        RECT 1174.930 2981.090 1176.110 2982.270 ;
        RECT 1174.930 2979.490 1176.110 2980.670 ;
        RECT 1174.930 2801.090 1176.110 2802.270 ;
        RECT 1174.930 2799.490 1176.110 2800.670 ;
        RECT 1174.930 2621.090 1176.110 2622.270 ;
        RECT 1174.930 2619.490 1176.110 2620.670 ;
        RECT 1174.930 2441.090 1176.110 2442.270 ;
        RECT 1174.930 2439.490 1176.110 2440.670 ;
        RECT 1174.930 2261.090 1176.110 2262.270 ;
        RECT 1174.930 2259.490 1176.110 2260.670 ;
        RECT 1174.930 2081.090 1176.110 2082.270 ;
        RECT 1174.930 2079.490 1176.110 2080.670 ;
        RECT 1174.930 1901.090 1176.110 1902.270 ;
        RECT 1174.930 1899.490 1176.110 1900.670 ;
        RECT 1174.930 1721.090 1176.110 1722.270 ;
        RECT 1174.930 1719.490 1176.110 1720.670 ;
        RECT 1174.930 1541.090 1176.110 1542.270 ;
        RECT 1174.930 1539.490 1176.110 1540.670 ;
        RECT 1174.930 1361.090 1176.110 1362.270 ;
        RECT 1174.930 1359.490 1176.110 1360.670 ;
        RECT 1174.930 1181.090 1176.110 1182.270 ;
        RECT 1174.930 1179.490 1176.110 1180.670 ;
        RECT 1174.930 1001.090 1176.110 1002.270 ;
        RECT 1174.930 999.490 1176.110 1000.670 ;
        RECT 1174.930 821.090 1176.110 822.270 ;
        RECT 1174.930 819.490 1176.110 820.670 ;
        RECT 1174.930 641.090 1176.110 642.270 ;
        RECT 1174.930 639.490 1176.110 640.670 ;
        RECT 1174.930 461.090 1176.110 462.270 ;
        RECT 1174.930 459.490 1176.110 460.670 ;
        RECT 1174.930 281.090 1176.110 282.270 ;
        RECT 1174.930 279.490 1176.110 280.670 ;
        RECT 1174.930 101.090 1176.110 102.270 ;
        RECT 1174.930 99.490 1176.110 100.670 ;
        RECT 1174.930 -7.510 1176.110 -6.330 ;
        RECT 1174.930 -9.110 1176.110 -7.930 ;
        RECT 1354.930 3527.610 1356.110 3528.790 ;
        RECT 1354.930 3526.010 1356.110 3527.190 ;
        RECT 1354.930 3341.090 1356.110 3342.270 ;
        RECT 1354.930 3339.490 1356.110 3340.670 ;
        RECT 1354.930 3161.090 1356.110 3162.270 ;
        RECT 1354.930 3159.490 1356.110 3160.670 ;
        RECT 1354.930 2981.090 1356.110 2982.270 ;
        RECT 1354.930 2979.490 1356.110 2980.670 ;
        RECT 1354.930 2801.090 1356.110 2802.270 ;
        RECT 1354.930 2799.490 1356.110 2800.670 ;
        RECT 1354.930 2621.090 1356.110 2622.270 ;
        RECT 1354.930 2619.490 1356.110 2620.670 ;
        RECT 1354.930 2441.090 1356.110 2442.270 ;
        RECT 1354.930 2439.490 1356.110 2440.670 ;
        RECT 1354.930 2261.090 1356.110 2262.270 ;
        RECT 1354.930 2259.490 1356.110 2260.670 ;
        RECT 1354.930 2081.090 1356.110 2082.270 ;
        RECT 1354.930 2079.490 1356.110 2080.670 ;
        RECT 1354.930 1901.090 1356.110 1902.270 ;
        RECT 1354.930 1899.490 1356.110 1900.670 ;
        RECT 1354.930 1721.090 1356.110 1722.270 ;
        RECT 1354.930 1719.490 1356.110 1720.670 ;
        RECT 1354.930 1541.090 1356.110 1542.270 ;
        RECT 1354.930 1539.490 1356.110 1540.670 ;
        RECT 1354.930 1361.090 1356.110 1362.270 ;
        RECT 1354.930 1359.490 1356.110 1360.670 ;
        RECT 1354.930 1181.090 1356.110 1182.270 ;
        RECT 1354.930 1179.490 1356.110 1180.670 ;
        RECT 1354.930 1001.090 1356.110 1002.270 ;
        RECT 1354.930 999.490 1356.110 1000.670 ;
        RECT 1354.930 821.090 1356.110 822.270 ;
        RECT 1354.930 819.490 1356.110 820.670 ;
        RECT 1354.930 641.090 1356.110 642.270 ;
        RECT 1354.930 639.490 1356.110 640.670 ;
        RECT 1354.930 461.090 1356.110 462.270 ;
        RECT 1354.930 459.490 1356.110 460.670 ;
        RECT 1354.930 281.090 1356.110 282.270 ;
        RECT 1354.930 279.490 1356.110 280.670 ;
        RECT 1354.930 101.090 1356.110 102.270 ;
        RECT 1354.930 99.490 1356.110 100.670 ;
        RECT 1354.930 -7.510 1356.110 -6.330 ;
        RECT 1354.930 -9.110 1356.110 -7.930 ;
        RECT 1534.930 3527.610 1536.110 3528.790 ;
        RECT 1534.930 3526.010 1536.110 3527.190 ;
        RECT 1534.930 3341.090 1536.110 3342.270 ;
        RECT 1534.930 3339.490 1536.110 3340.670 ;
        RECT 1534.930 3161.090 1536.110 3162.270 ;
        RECT 1534.930 3159.490 1536.110 3160.670 ;
        RECT 1534.930 2981.090 1536.110 2982.270 ;
        RECT 1534.930 2979.490 1536.110 2980.670 ;
        RECT 1534.930 2801.090 1536.110 2802.270 ;
        RECT 1534.930 2799.490 1536.110 2800.670 ;
        RECT 1534.930 2621.090 1536.110 2622.270 ;
        RECT 1534.930 2619.490 1536.110 2620.670 ;
        RECT 1534.930 2441.090 1536.110 2442.270 ;
        RECT 1534.930 2439.490 1536.110 2440.670 ;
        RECT 1534.930 2261.090 1536.110 2262.270 ;
        RECT 1534.930 2259.490 1536.110 2260.670 ;
        RECT 1534.930 2081.090 1536.110 2082.270 ;
        RECT 1534.930 2079.490 1536.110 2080.670 ;
        RECT 1534.930 1901.090 1536.110 1902.270 ;
        RECT 1534.930 1899.490 1536.110 1900.670 ;
        RECT 1534.930 1721.090 1536.110 1722.270 ;
        RECT 1534.930 1719.490 1536.110 1720.670 ;
        RECT 1534.930 1541.090 1536.110 1542.270 ;
        RECT 1534.930 1539.490 1536.110 1540.670 ;
        RECT 1534.930 1361.090 1536.110 1362.270 ;
        RECT 1534.930 1359.490 1536.110 1360.670 ;
        RECT 1534.930 1181.090 1536.110 1182.270 ;
        RECT 1534.930 1179.490 1536.110 1180.670 ;
        RECT 1534.930 1001.090 1536.110 1002.270 ;
        RECT 1534.930 999.490 1536.110 1000.670 ;
        RECT 1534.930 821.090 1536.110 822.270 ;
        RECT 1534.930 819.490 1536.110 820.670 ;
        RECT 1534.930 641.090 1536.110 642.270 ;
        RECT 1534.930 639.490 1536.110 640.670 ;
        RECT 1534.930 461.090 1536.110 462.270 ;
        RECT 1534.930 459.490 1536.110 460.670 ;
        RECT 1534.930 281.090 1536.110 282.270 ;
        RECT 1534.930 279.490 1536.110 280.670 ;
        RECT 1534.930 101.090 1536.110 102.270 ;
        RECT 1534.930 99.490 1536.110 100.670 ;
        RECT 1534.930 -7.510 1536.110 -6.330 ;
        RECT 1534.930 -9.110 1536.110 -7.930 ;
        RECT 1714.930 3527.610 1716.110 3528.790 ;
        RECT 1714.930 3526.010 1716.110 3527.190 ;
        RECT 1714.930 3341.090 1716.110 3342.270 ;
        RECT 1714.930 3339.490 1716.110 3340.670 ;
        RECT 1714.930 3161.090 1716.110 3162.270 ;
        RECT 1714.930 3159.490 1716.110 3160.670 ;
        RECT 1714.930 2981.090 1716.110 2982.270 ;
        RECT 1714.930 2979.490 1716.110 2980.670 ;
        RECT 1714.930 2801.090 1716.110 2802.270 ;
        RECT 1714.930 2799.490 1716.110 2800.670 ;
        RECT 1714.930 2621.090 1716.110 2622.270 ;
        RECT 1714.930 2619.490 1716.110 2620.670 ;
        RECT 1714.930 2441.090 1716.110 2442.270 ;
        RECT 1714.930 2439.490 1716.110 2440.670 ;
        RECT 1714.930 2261.090 1716.110 2262.270 ;
        RECT 1714.930 2259.490 1716.110 2260.670 ;
        RECT 1714.930 2081.090 1716.110 2082.270 ;
        RECT 1714.930 2079.490 1716.110 2080.670 ;
        RECT 1714.930 1901.090 1716.110 1902.270 ;
        RECT 1714.930 1899.490 1716.110 1900.670 ;
        RECT 1714.930 1721.090 1716.110 1722.270 ;
        RECT 1714.930 1719.490 1716.110 1720.670 ;
        RECT 1714.930 1541.090 1716.110 1542.270 ;
        RECT 1714.930 1539.490 1716.110 1540.670 ;
        RECT 1714.930 1361.090 1716.110 1362.270 ;
        RECT 1714.930 1359.490 1716.110 1360.670 ;
        RECT 1714.930 1181.090 1716.110 1182.270 ;
        RECT 1714.930 1179.490 1716.110 1180.670 ;
        RECT 1714.930 1001.090 1716.110 1002.270 ;
        RECT 1714.930 999.490 1716.110 1000.670 ;
        RECT 1714.930 821.090 1716.110 822.270 ;
        RECT 1714.930 819.490 1716.110 820.670 ;
        RECT 1714.930 641.090 1716.110 642.270 ;
        RECT 1714.930 639.490 1716.110 640.670 ;
        RECT 1714.930 461.090 1716.110 462.270 ;
        RECT 1714.930 459.490 1716.110 460.670 ;
        RECT 1714.930 281.090 1716.110 282.270 ;
        RECT 1714.930 279.490 1716.110 280.670 ;
        RECT 1714.930 101.090 1716.110 102.270 ;
        RECT 1714.930 99.490 1716.110 100.670 ;
        RECT 1714.930 -7.510 1716.110 -6.330 ;
        RECT 1714.930 -9.110 1716.110 -7.930 ;
        RECT 1894.930 3527.610 1896.110 3528.790 ;
        RECT 1894.930 3526.010 1896.110 3527.190 ;
        RECT 1894.930 3341.090 1896.110 3342.270 ;
        RECT 1894.930 3339.490 1896.110 3340.670 ;
        RECT 1894.930 3161.090 1896.110 3162.270 ;
        RECT 1894.930 3159.490 1896.110 3160.670 ;
        RECT 1894.930 2981.090 1896.110 2982.270 ;
        RECT 1894.930 2979.490 1896.110 2980.670 ;
        RECT 1894.930 2801.090 1896.110 2802.270 ;
        RECT 1894.930 2799.490 1896.110 2800.670 ;
        RECT 1894.930 2621.090 1896.110 2622.270 ;
        RECT 1894.930 2619.490 1896.110 2620.670 ;
        RECT 1894.930 2441.090 1896.110 2442.270 ;
        RECT 1894.930 2439.490 1896.110 2440.670 ;
        RECT 1894.930 2261.090 1896.110 2262.270 ;
        RECT 1894.930 2259.490 1896.110 2260.670 ;
        RECT 1894.930 2081.090 1896.110 2082.270 ;
        RECT 1894.930 2079.490 1896.110 2080.670 ;
        RECT 1894.930 1901.090 1896.110 1902.270 ;
        RECT 1894.930 1899.490 1896.110 1900.670 ;
        RECT 1894.930 1721.090 1896.110 1722.270 ;
        RECT 1894.930 1719.490 1896.110 1720.670 ;
        RECT 1894.930 1541.090 1896.110 1542.270 ;
        RECT 1894.930 1539.490 1896.110 1540.670 ;
        RECT 1894.930 1361.090 1896.110 1362.270 ;
        RECT 1894.930 1359.490 1896.110 1360.670 ;
        RECT 1894.930 1181.090 1896.110 1182.270 ;
        RECT 1894.930 1179.490 1896.110 1180.670 ;
        RECT 1894.930 1001.090 1896.110 1002.270 ;
        RECT 1894.930 999.490 1896.110 1000.670 ;
        RECT 1894.930 821.090 1896.110 822.270 ;
        RECT 1894.930 819.490 1896.110 820.670 ;
        RECT 1894.930 641.090 1896.110 642.270 ;
        RECT 1894.930 639.490 1896.110 640.670 ;
        RECT 1894.930 461.090 1896.110 462.270 ;
        RECT 1894.930 459.490 1896.110 460.670 ;
        RECT 1894.930 281.090 1896.110 282.270 ;
        RECT 1894.930 279.490 1896.110 280.670 ;
        RECT 1894.930 101.090 1896.110 102.270 ;
        RECT 1894.930 99.490 1896.110 100.670 ;
        RECT 1894.930 -7.510 1896.110 -6.330 ;
        RECT 1894.930 -9.110 1896.110 -7.930 ;
        RECT 2074.930 3527.610 2076.110 3528.790 ;
        RECT 2074.930 3526.010 2076.110 3527.190 ;
        RECT 2074.930 3341.090 2076.110 3342.270 ;
        RECT 2074.930 3339.490 2076.110 3340.670 ;
        RECT 2074.930 3161.090 2076.110 3162.270 ;
        RECT 2074.930 3159.490 2076.110 3160.670 ;
        RECT 2074.930 2981.090 2076.110 2982.270 ;
        RECT 2074.930 2979.490 2076.110 2980.670 ;
        RECT 2074.930 2801.090 2076.110 2802.270 ;
        RECT 2074.930 2799.490 2076.110 2800.670 ;
        RECT 2074.930 2621.090 2076.110 2622.270 ;
        RECT 2074.930 2619.490 2076.110 2620.670 ;
        RECT 2074.930 2441.090 2076.110 2442.270 ;
        RECT 2074.930 2439.490 2076.110 2440.670 ;
        RECT 2074.930 2261.090 2076.110 2262.270 ;
        RECT 2074.930 2259.490 2076.110 2260.670 ;
        RECT 2074.930 2081.090 2076.110 2082.270 ;
        RECT 2074.930 2079.490 2076.110 2080.670 ;
        RECT 2074.930 1901.090 2076.110 1902.270 ;
        RECT 2074.930 1899.490 2076.110 1900.670 ;
        RECT 2074.930 1721.090 2076.110 1722.270 ;
        RECT 2074.930 1719.490 2076.110 1720.670 ;
        RECT 2074.930 1541.090 2076.110 1542.270 ;
        RECT 2074.930 1539.490 2076.110 1540.670 ;
        RECT 2074.930 1361.090 2076.110 1362.270 ;
        RECT 2074.930 1359.490 2076.110 1360.670 ;
        RECT 2074.930 1181.090 2076.110 1182.270 ;
        RECT 2074.930 1179.490 2076.110 1180.670 ;
        RECT 2074.930 1001.090 2076.110 1002.270 ;
        RECT 2074.930 999.490 2076.110 1000.670 ;
        RECT 2074.930 821.090 2076.110 822.270 ;
        RECT 2074.930 819.490 2076.110 820.670 ;
        RECT 2074.930 641.090 2076.110 642.270 ;
        RECT 2074.930 639.490 2076.110 640.670 ;
        RECT 2074.930 461.090 2076.110 462.270 ;
        RECT 2074.930 459.490 2076.110 460.670 ;
        RECT 2074.930 281.090 2076.110 282.270 ;
        RECT 2074.930 279.490 2076.110 280.670 ;
        RECT 2074.930 101.090 2076.110 102.270 ;
        RECT 2074.930 99.490 2076.110 100.670 ;
        RECT 2074.930 -7.510 2076.110 -6.330 ;
        RECT 2074.930 -9.110 2076.110 -7.930 ;
        RECT 2254.930 3527.610 2256.110 3528.790 ;
        RECT 2254.930 3526.010 2256.110 3527.190 ;
        RECT 2254.930 3341.090 2256.110 3342.270 ;
        RECT 2254.930 3339.490 2256.110 3340.670 ;
        RECT 2254.930 3161.090 2256.110 3162.270 ;
        RECT 2254.930 3159.490 2256.110 3160.670 ;
        RECT 2254.930 2981.090 2256.110 2982.270 ;
        RECT 2254.930 2979.490 2256.110 2980.670 ;
        RECT 2254.930 2801.090 2256.110 2802.270 ;
        RECT 2254.930 2799.490 2256.110 2800.670 ;
        RECT 2254.930 2621.090 2256.110 2622.270 ;
        RECT 2254.930 2619.490 2256.110 2620.670 ;
        RECT 2254.930 2441.090 2256.110 2442.270 ;
        RECT 2254.930 2439.490 2256.110 2440.670 ;
        RECT 2254.930 2261.090 2256.110 2262.270 ;
        RECT 2254.930 2259.490 2256.110 2260.670 ;
        RECT 2254.930 2081.090 2256.110 2082.270 ;
        RECT 2254.930 2079.490 2256.110 2080.670 ;
        RECT 2254.930 1901.090 2256.110 1902.270 ;
        RECT 2254.930 1899.490 2256.110 1900.670 ;
        RECT 2254.930 1721.090 2256.110 1722.270 ;
        RECT 2254.930 1719.490 2256.110 1720.670 ;
        RECT 2254.930 1541.090 2256.110 1542.270 ;
        RECT 2254.930 1539.490 2256.110 1540.670 ;
        RECT 2254.930 1361.090 2256.110 1362.270 ;
        RECT 2254.930 1359.490 2256.110 1360.670 ;
        RECT 2254.930 1181.090 2256.110 1182.270 ;
        RECT 2254.930 1179.490 2256.110 1180.670 ;
        RECT 2254.930 1001.090 2256.110 1002.270 ;
        RECT 2254.930 999.490 2256.110 1000.670 ;
        RECT 2254.930 821.090 2256.110 822.270 ;
        RECT 2254.930 819.490 2256.110 820.670 ;
        RECT 2254.930 641.090 2256.110 642.270 ;
        RECT 2254.930 639.490 2256.110 640.670 ;
        RECT 2254.930 461.090 2256.110 462.270 ;
        RECT 2254.930 459.490 2256.110 460.670 ;
        RECT 2254.930 281.090 2256.110 282.270 ;
        RECT 2254.930 279.490 2256.110 280.670 ;
        RECT 2254.930 101.090 2256.110 102.270 ;
        RECT 2254.930 99.490 2256.110 100.670 ;
        RECT 2254.930 -7.510 2256.110 -6.330 ;
        RECT 2254.930 -9.110 2256.110 -7.930 ;
        RECT 2434.930 3527.610 2436.110 3528.790 ;
        RECT 2434.930 3526.010 2436.110 3527.190 ;
        RECT 2434.930 3341.090 2436.110 3342.270 ;
        RECT 2434.930 3339.490 2436.110 3340.670 ;
        RECT 2434.930 3161.090 2436.110 3162.270 ;
        RECT 2434.930 3159.490 2436.110 3160.670 ;
        RECT 2434.930 2981.090 2436.110 2982.270 ;
        RECT 2434.930 2979.490 2436.110 2980.670 ;
        RECT 2434.930 2801.090 2436.110 2802.270 ;
        RECT 2434.930 2799.490 2436.110 2800.670 ;
        RECT 2434.930 2621.090 2436.110 2622.270 ;
        RECT 2434.930 2619.490 2436.110 2620.670 ;
        RECT 2434.930 2441.090 2436.110 2442.270 ;
        RECT 2434.930 2439.490 2436.110 2440.670 ;
        RECT 2434.930 2261.090 2436.110 2262.270 ;
        RECT 2434.930 2259.490 2436.110 2260.670 ;
        RECT 2434.930 2081.090 2436.110 2082.270 ;
        RECT 2434.930 2079.490 2436.110 2080.670 ;
        RECT 2434.930 1901.090 2436.110 1902.270 ;
        RECT 2434.930 1899.490 2436.110 1900.670 ;
        RECT 2434.930 1721.090 2436.110 1722.270 ;
        RECT 2434.930 1719.490 2436.110 1720.670 ;
        RECT 2434.930 1541.090 2436.110 1542.270 ;
        RECT 2434.930 1539.490 2436.110 1540.670 ;
        RECT 2434.930 1361.090 2436.110 1362.270 ;
        RECT 2434.930 1359.490 2436.110 1360.670 ;
        RECT 2434.930 1181.090 2436.110 1182.270 ;
        RECT 2434.930 1179.490 2436.110 1180.670 ;
        RECT 2434.930 1001.090 2436.110 1002.270 ;
        RECT 2434.930 999.490 2436.110 1000.670 ;
        RECT 2434.930 821.090 2436.110 822.270 ;
        RECT 2434.930 819.490 2436.110 820.670 ;
        RECT 2434.930 641.090 2436.110 642.270 ;
        RECT 2434.930 639.490 2436.110 640.670 ;
        RECT 2434.930 461.090 2436.110 462.270 ;
        RECT 2434.930 459.490 2436.110 460.670 ;
        RECT 2434.930 281.090 2436.110 282.270 ;
        RECT 2434.930 279.490 2436.110 280.670 ;
        RECT 2434.930 101.090 2436.110 102.270 ;
        RECT 2434.930 99.490 2436.110 100.670 ;
        RECT 2434.930 -7.510 2436.110 -6.330 ;
        RECT 2434.930 -9.110 2436.110 -7.930 ;
        RECT 2614.930 3527.610 2616.110 3528.790 ;
        RECT 2614.930 3526.010 2616.110 3527.190 ;
        RECT 2614.930 3341.090 2616.110 3342.270 ;
        RECT 2614.930 3339.490 2616.110 3340.670 ;
        RECT 2614.930 3161.090 2616.110 3162.270 ;
        RECT 2614.930 3159.490 2616.110 3160.670 ;
        RECT 2614.930 2981.090 2616.110 2982.270 ;
        RECT 2614.930 2979.490 2616.110 2980.670 ;
        RECT 2614.930 2801.090 2616.110 2802.270 ;
        RECT 2614.930 2799.490 2616.110 2800.670 ;
        RECT 2614.930 2621.090 2616.110 2622.270 ;
        RECT 2614.930 2619.490 2616.110 2620.670 ;
        RECT 2614.930 2441.090 2616.110 2442.270 ;
        RECT 2614.930 2439.490 2616.110 2440.670 ;
        RECT 2614.930 2261.090 2616.110 2262.270 ;
        RECT 2614.930 2259.490 2616.110 2260.670 ;
        RECT 2614.930 2081.090 2616.110 2082.270 ;
        RECT 2614.930 2079.490 2616.110 2080.670 ;
        RECT 2614.930 1901.090 2616.110 1902.270 ;
        RECT 2614.930 1899.490 2616.110 1900.670 ;
        RECT 2614.930 1721.090 2616.110 1722.270 ;
        RECT 2614.930 1719.490 2616.110 1720.670 ;
        RECT 2614.930 1541.090 2616.110 1542.270 ;
        RECT 2614.930 1539.490 2616.110 1540.670 ;
        RECT 2614.930 1361.090 2616.110 1362.270 ;
        RECT 2614.930 1359.490 2616.110 1360.670 ;
        RECT 2614.930 1181.090 2616.110 1182.270 ;
        RECT 2614.930 1179.490 2616.110 1180.670 ;
        RECT 2614.930 1001.090 2616.110 1002.270 ;
        RECT 2614.930 999.490 2616.110 1000.670 ;
        RECT 2614.930 821.090 2616.110 822.270 ;
        RECT 2614.930 819.490 2616.110 820.670 ;
        RECT 2614.930 641.090 2616.110 642.270 ;
        RECT 2614.930 639.490 2616.110 640.670 ;
        RECT 2614.930 461.090 2616.110 462.270 ;
        RECT 2614.930 459.490 2616.110 460.670 ;
        RECT 2614.930 281.090 2616.110 282.270 ;
        RECT 2614.930 279.490 2616.110 280.670 ;
        RECT 2614.930 101.090 2616.110 102.270 ;
        RECT 2614.930 99.490 2616.110 100.670 ;
        RECT 2614.930 -7.510 2616.110 -6.330 ;
        RECT 2614.930 -9.110 2616.110 -7.930 ;
        RECT 2794.930 3527.610 2796.110 3528.790 ;
        RECT 2794.930 3526.010 2796.110 3527.190 ;
        RECT 2794.930 3341.090 2796.110 3342.270 ;
        RECT 2794.930 3339.490 2796.110 3340.670 ;
        RECT 2794.930 3161.090 2796.110 3162.270 ;
        RECT 2794.930 3159.490 2796.110 3160.670 ;
        RECT 2794.930 2981.090 2796.110 2982.270 ;
        RECT 2794.930 2979.490 2796.110 2980.670 ;
        RECT 2794.930 2801.090 2796.110 2802.270 ;
        RECT 2794.930 2799.490 2796.110 2800.670 ;
        RECT 2794.930 2621.090 2796.110 2622.270 ;
        RECT 2794.930 2619.490 2796.110 2620.670 ;
        RECT 2794.930 2441.090 2796.110 2442.270 ;
        RECT 2794.930 2439.490 2796.110 2440.670 ;
        RECT 2794.930 2261.090 2796.110 2262.270 ;
        RECT 2794.930 2259.490 2796.110 2260.670 ;
        RECT 2794.930 2081.090 2796.110 2082.270 ;
        RECT 2794.930 2079.490 2796.110 2080.670 ;
        RECT 2794.930 1901.090 2796.110 1902.270 ;
        RECT 2794.930 1899.490 2796.110 1900.670 ;
        RECT 2794.930 1721.090 2796.110 1722.270 ;
        RECT 2794.930 1719.490 2796.110 1720.670 ;
        RECT 2794.930 1541.090 2796.110 1542.270 ;
        RECT 2794.930 1539.490 2796.110 1540.670 ;
        RECT 2794.930 1361.090 2796.110 1362.270 ;
        RECT 2794.930 1359.490 2796.110 1360.670 ;
        RECT 2794.930 1181.090 2796.110 1182.270 ;
        RECT 2794.930 1179.490 2796.110 1180.670 ;
        RECT 2794.930 1001.090 2796.110 1002.270 ;
        RECT 2794.930 999.490 2796.110 1000.670 ;
        RECT 2794.930 821.090 2796.110 822.270 ;
        RECT 2794.930 819.490 2796.110 820.670 ;
        RECT 2794.930 641.090 2796.110 642.270 ;
        RECT 2794.930 639.490 2796.110 640.670 ;
        RECT 2794.930 461.090 2796.110 462.270 ;
        RECT 2794.930 459.490 2796.110 460.670 ;
        RECT 2794.930 281.090 2796.110 282.270 ;
        RECT 2794.930 279.490 2796.110 280.670 ;
        RECT 2794.930 101.090 2796.110 102.270 ;
        RECT 2794.930 99.490 2796.110 100.670 ;
        RECT 2794.930 -7.510 2796.110 -6.330 ;
        RECT 2794.930 -9.110 2796.110 -7.930 ;
        RECT 2932.110 3527.610 2933.290 3528.790 ;
        RECT 2932.110 3526.010 2933.290 3527.190 ;
        RECT 2932.110 3341.090 2933.290 3342.270 ;
        RECT 2932.110 3339.490 2933.290 3340.670 ;
        RECT 2932.110 3161.090 2933.290 3162.270 ;
        RECT 2932.110 3159.490 2933.290 3160.670 ;
        RECT 2932.110 2981.090 2933.290 2982.270 ;
        RECT 2932.110 2979.490 2933.290 2980.670 ;
        RECT 2932.110 2801.090 2933.290 2802.270 ;
        RECT 2932.110 2799.490 2933.290 2800.670 ;
        RECT 2932.110 2621.090 2933.290 2622.270 ;
        RECT 2932.110 2619.490 2933.290 2620.670 ;
        RECT 2932.110 2441.090 2933.290 2442.270 ;
        RECT 2932.110 2439.490 2933.290 2440.670 ;
        RECT 2932.110 2261.090 2933.290 2262.270 ;
        RECT 2932.110 2259.490 2933.290 2260.670 ;
        RECT 2932.110 2081.090 2933.290 2082.270 ;
        RECT 2932.110 2079.490 2933.290 2080.670 ;
        RECT 2932.110 1901.090 2933.290 1902.270 ;
        RECT 2932.110 1899.490 2933.290 1900.670 ;
        RECT 2932.110 1721.090 2933.290 1722.270 ;
        RECT 2932.110 1719.490 2933.290 1720.670 ;
        RECT 2932.110 1541.090 2933.290 1542.270 ;
        RECT 2932.110 1539.490 2933.290 1540.670 ;
        RECT 2932.110 1361.090 2933.290 1362.270 ;
        RECT 2932.110 1359.490 2933.290 1360.670 ;
        RECT 2932.110 1181.090 2933.290 1182.270 ;
        RECT 2932.110 1179.490 2933.290 1180.670 ;
        RECT 2932.110 1001.090 2933.290 1002.270 ;
        RECT 2932.110 999.490 2933.290 1000.670 ;
        RECT 2932.110 821.090 2933.290 822.270 ;
        RECT 2932.110 819.490 2933.290 820.670 ;
        RECT 2932.110 641.090 2933.290 642.270 ;
        RECT 2932.110 639.490 2933.290 640.670 ;
        RECT 2932.110 461.090 2933.290 462.270 ;
        RECT 2932.110 459.490 2933.290 460.670 ;
        RECT 2932.110 281.090 2933.290 282.270 ;
        RECT 2932.110 279.490 2933.290 280.670 ;
        RECT 2932.110 101.090 2933.290 102.270 ;
        RECT 2932.110 99.490 2933.290 100.670 ;
        RECT 2932.110 -7.510 2933.290 -6.330 ;
        RECT 2932.110 -9.110 2933.290 -7.930 ;
      LAYER met5 ;
        RECT -14.580 3528.900 -11.580 3528.910 ;
        RECT 94.020 3528.900 97.020 3528.910 ;
        RECT 274.020 3528.900 277.020 3528.910 ;
        RECT 454.020 3528.900 457.020 3528.910 ;
        RECT 634.020 3528.900 637.020 3528.910 ;
        RECT 814.020 3528.900 817.020 3528.910 ;
        RECT 994.020 3528.900 997.020 3528.910 ;
        RECT 1174.020 3528.900 1177.020 3528.910 ;
        RECT 1354.020 3528.900 1357.020 3528.910 ;
        RECT 1534.020 3528.900 1537.020 3528.910 ;
        RECT 1714.020 3528.900 1717.020 3528.910 ;
        RECT 1894.020 3528.900 1897.020 3528.910 ;
        RECT 2074.020 3528.900 2077.020 3528.910 ;
        RECT 2254.020 3528.900 2257.020 3528.910 ;
        RECT 2434.020 3528.900 2437.020 3528.910 ;
        RECT 2614.020 3528.900 2617.020 3528.910 ;
        RECT 2794.020 3528.900 2797.020 3528.910 ;
        RECT 2931.200 3528.900 2934.200 3528.910 ;
        RECT -14.580 3525.900 2934.200 3528.900 ;
        RECT -14.580 3525.890 -11.580 3525.900 ;
        RECT 94.020 3525.890 97.020 3525.900 ;
        RECT 274.020 3525.890 277.020 3525.900 ;
        RECT 454.020 3525.890 457.020 3525.900 ;
        RECT 634.020 3525.890 637.020 3525.900 ;
        RECT 814.020 3525.890 817.020 3525.900 ;
        RECT 994.020 3525.890 997.020 3525.900 ;
        RECT 1174.020 3525.890 1177.020 3525.900 ;
        RECT 1354.020 3525.890 1357.020 3525.900 ;
        RECT 1534.020 3525.890 1537.020 3525.900 ;
        RECT 1714.020 3525.890 1717.020 3525.900 ;
        RECT 1894.020 3525.890 1897.020 3525.900 ;
        RECT 2074.020 3525.890 2077.020 3525.900 ;
        RECT 2254.020 3525.890 2257.020 3525.900 ;
        RECT 2434.020 3525.890 2437.020 3525.900 ;
        RECT 2614.020 3525.890 2617.020 3525.900 ;
        RECT 2794.020 3525.890 2797.020 3525.900 ;
        RECT 2931.200 3525.890 2934.200 3525.900 ;
        RECT -14.580 3342.380 -11.580 3342.390 ;
        RECT 94.020 3342.380 97.020 3342.390 ;
        RECT 274.020 3342.380 277.020 3342.390 ;
        RECT 454.020 3342.380 457.020 3342.390 ;
        RECT 634.020 3342.380 637.020 3342.390 ;
        RECT 814.020 3342.380 817.020 3342.390 ;
        RECT 994.020 3342.380 997.020 3342.390 ;
        RECT 1174.020 3342.380 1177.020 3342.390 ;
        RECT 1354.020 3342.380 1357.020 3342.390 ;
        RECT 1534.020 3342.380 1537.020 3342.390 ;
        RECT 1714.020 3342.380 1717.020 3342.390 ;
        RECT 1894.020 3342.380 1897.020 3342.390 ;
        RECT 2074.020 3342.380 2077.020 3342.390 ;
        RECT 2254.020 3342.380 2257.020 3342.390 ;
        RECT 2434.020 3342.380 2437.020 3342.390 ;
        RECT 2614.020 3342.380 2617.020 3342.390 ;
        RECT 2794.020 3342.380 2797.020 3342.390 ;
        RECT 2931.200 3342.380 2934.200 3342.390 ;
        RECT -14.580 3339.380 2934.200 3342.380 ;
        RECT -14.580 3339.370 -11.580 3339.380 ;
        RECT 94.020 3339.370 97.020 3339.380 ;
        RECT 274.020 3339.370 277.020 3339.380 ;
        RECT 454.020 3339.370 457.020 3339.380 ;
        RECT 634.020 3339.370 637.020 3339.380 ;
        RECT 814.020 3339.370 817.020 3339.380 ;
        RECT 994.020 3339.370 997.020 3339.380 ;
        RECT 1174.020 3339.370 1177.020 3339.380 ;
        RECT 1354.020 3339.370 1357.020 3339.380 ;
        RECT 1534.020 3339.370 1537.020 3339.380 ;
        RECT 1714.020 3339.370 1717.020 3339.380 ;
        RECT 1894.020 3339.370 1897.020 3339.380 ;
        RECT 2074.020 3339.370 2077.020 3339.380 ;
        RECT 2254.020 3339.370 2257.020 3339.380 ;
        RECT 2434.020 3339.370 2437.020 3339.380 ;
        RECT 2614.020 3339.370 2617.020 3339.380 ;
        RECT 2794.020 3339.370 2797.020 3339.380 ;
        RECT 2931.200 3339.370 2934.200 3339.380 ;
        RECT -14.580 3162.380 -11.580 3162.390 ;
        RECT 94.020 3162.380 97.020 3162.390 ;
        RECT 274.020 3162.380 277.020 3162.390 ;
        RECT 454.020 3162.380 457.020 3162.390 ;
        RECT 634.020 3162.380 637.020 3162.390 ;
        RECT 814.020 3162.380 817.020 3162.390 ;
        RECT 994.020 3162.380 997.020 3162.390 ;
        RECT 1174.020 3162.380 1177.020 3162.390 ;
        RECT 1354.020 3162.380 1357.020 3162.390 ;
        RECT 1534.020 3162.380 1537.020 3162.390 ;
        RECT 1714.020 3162.380 1717.020 3162.390 ;
        RECT 1894.020 3162.380 1897.020 3162.390 ;
        RECT 2074.020 3162.380 2077.020 3162.390 ;
        RECT 2254.020 3162.380 2257.020 3162.390 ;
        RECT 2434.020 3162.380 2437.020 3162.390 ;
        RECT 2614.020 3162.380 2617.020 3162.390 ;
        RECT 2794.020 3162.380 2797.020 3162.390 ;
        RECT 2931.200 3162.380 2934.200 3162.390 ;
        RECT -14.580 3159.380 2934.200 3162.380 ;
        RECT -14.580 3159.370 -11.580 3159.380 ;
        RECT 94.020 3159.370 97.020 3159.380 ;
        RECT 274.020 3159.370 277.020 3159.380 ;
        RECT 454.020 3159.370 457.020 3159.380 ;
        RECT 634.020 3159.370 637.020 3159.380 ;
        RECT 814.020 3159.370 817.020 3159.380 ;
        RECT 994.020 3159.370 997.020 3159.380 ;
        RECT 1174.020 3159.370 1177.020 3159.380 ;
        RECT 1354.020 3159.370 1357.020 3159.380 ;
        RECT 1534.020 3159.370 1537.020 3159.380 ;
        RECT 1714.020 3159.370 1717.020 3159.380 ;
        RECT 1894.020 3159.370 1897.020 3159.380 ;
        RECT 2074.020 3159.370 2077.020 3159.380 ;
        RECT 2254.020 3159.370 2257.020 3159.380 ;
        RECT 2434.020 3159.370 2437.020 3159.380 ;
        RECT 2614.020 3159.370 2617.020 3159.380 ;
        RECT 2794.020 3159.370 2797.020 3159.380 ;
        RECT 2931.200 3159.370 2934.200 3159.380 ;
        RECT -14.580 2982.380 -11.580 2982.390 ;
        RECT 94.020 2982.380 97.020 2982.390 ;
        RECT 274.020 2982.380 277.020 2982.390 ;
        RECT 454.020 2982.380 457.020 2982.390 ;
        RECT 634.020 2982.380 637.020 2982.390 ;
        RECT 814.020 2982.380 817.020 2982.390 ;
        RECT 994.020 2982.380 997.020 2982.390 ;
        RECT 1174.020 2982.380 1177.020 2982.390 ;
        RECT 1354.020 2982.380 1357.020 2982.390 ;
        RECT 1534.020 2982.380 1537.020 2982.390 ;
        RECT 1714.020 2982.380 1717.020 2982.390 ;
        RECT 1894.020 2982.380 1897.020 2982.390 ;
        RECT 2074.020 2982.380 2077.020 2982.390 ;
        RECT 2254.020 2982.380 2257.020 2982.390 ;
        RECT 2434.020 2982.380 2437.020 2982.390 ;
        RECT 2614.020 2982.380 2617.020 2982.390 ;
        RECT 2794.020 2982.380 2797.020 2982.390 ;
        RECT 2931.200 2982.380 2934.200 2982.390 ;
        RECT -14.580 2979.380 2934.200 2982.380 ;
        RECT -14.580 2979.370 -11.580 2979.380 ;
        RECT 94.020 2979.370 97.020 2979.380 ;
        RECT 274.020 2979.370 277.020 2979.380 ;
        RECT 454.020 2979.370 457.020 2979.380 ;
        RECT 634.020 2979.370 637.020 2979.380 ;
        RECT 814.020 2979.370 817.020 2979.380 ;
        RECT 994.020 2979.370 997.020 2979.380 ;
        RECT 1174.020 2979.370 1177.020 2979.380 ;
        RECT 1354.020 2979.370 1357.020 2979.380 ;
        RECT 1534.020 2979.370 1537.020 2979.380 ;
        RECT 1714.020 2979.370 1717.020 2979.380 ;
        RECT 1894.020 2979.370 1897.020 2979.380 ;
        RECT 2074.020 2979.370 2077.020 2979.380 ;
        RECT 2254.020 2979.370 2257.020 2979.380 ;
        RECT 2434.020 2979.370 2437.020 2979.380 ;
        RECT 2614.020 2979.370 2617.020 2979.380 ;
        RECT 2794.020 2979.370 2797.020 2979.380 ;
        RECT 2931.200 2979.370 2934.200 2979.380 ;
        RECT -14.580 2802.380 -11.580 2802.390 ;
        RECT 94.020 2802.380 97.020 2802.390 ;
        RECT 274.020 2802.380 277.020 2802.390 ;
        RECT 454.020 2802.380 457.020 2802.390 ;
        RECT 634.020 2802.380 637.020 2802.390 ;
        RECT 814.020 2802.380 817.020 2802.390 ;
        RECT 994.020 2802.380 997.020 2802.390 ;
        RECT 1174.020 2802.380 1177.020 2802.390 ;
        RECT 1354.020 2802.380 1357.020 2802.390 ;
        RECT 1534.020 2802.380 1537.020 2802.390 ;
        RECT 1714.020 2802.380 1717.020 2802.390 ;
        RECT 1894.020 2802.380 1897.020 2802.390 ;
        RECT 2074.020 2802.380 2077.020 2802.390 ;
        RECT 2254.020 2802.380 2257.020 2802.390 ;
        RECT 2434.020 2802.380 2437.020 2802.390 ;
        RECT 2614.020 2802.380 2617.020 2802.390 ;
        RECT 2794.020 2802.380 2797.020 2802.390 ;
        RECT 2931.200 2802.380 2934.200 2802.390 ;
        RECT -14.580 2799.380 2934.200 2802.380 ;
        RECT -14.580 2799.370 -11.580 2799.380 ;
        RECT 94.020 2799.370 97.020 2799.380 ;
        RECT 274.020 2799.370 277.020 2799.380 ;
        RECT 454.020 2799.370 457.020 2799.380 ;
        RECT 634.020 2799.370 637.020 2799.380 ;
        RECT 814.020 2799.370 817.020 2799.380 ;
        RECT 994.020 2799.370 997.020 2799.380 ;
        RECT 1174.020 2799.370 1177.020 2799.380 ;
        RECT 1354.020 2799.370 1357.020 2799.380 ;
        RECT 1534.020 2799.370 1537.020 2799.380 ;
        RECT 1714.020 2799.370 1717.020 2799.380 ;
        RECT 1894.020 2799.370 1897.020 2799.380 ;
        RECT 2074.020 2799.370 2077.020 2799.380 ;
        RECT 2254.020 2799.370 2257.020 2799.380 ;
        RECT 2434.020 2799.370 2437.020 2799.380 ;
        RECT 2614.020 2799.370 2617.020 2799.380 ;
        RECT 2794.020 2799.370 2797.020 2799.380 ;
        RECT 2931.200 2799.370 2934.200 2799.380 ;
        RECT -14.580 2622.380 -11.580 2622.390 ;
        RECT 94.020 2622.380 97.020 2622.390 ;
        RECT 274.020 2622.380 277.020 2622.390 ;
        RECT 454.020 2622.380 457.020 2622.390 ;
        RECT 634.020 2622.380 637.020 2622.390 ;
        RECT 814.020 2622.380 817.020 2622.390 ;
        RECT 994.020 2622.380 997.020 2622.390 ;
        RECT 1174.020 2622.380 1177.020 2622.390 ;
        RECT 1354.020 2622.380 1357.020 2622.390 ;
        RECT 1534.020 2622.380 1537.020 2622.390 ;
        RECT 1714.020 2622.380 1717.020 2622.390 ;
        RECT 1894.020 2622.380 1897.020 2622.390 ;
        RECT 2074.020 2622.380 2077.020 2622.390 ;
        RECT 2254.020 2622.380 2257.020 2622.390 ;
        RECT 2434.020 2622.380 2437.020 2622.390 ;
        RECT 2614.020 2622.380 2617.020 2622.390 ;
        RECT 2794.020 2622.380 2797.020 2622.390 ;
        RECT 2931.200 2622.380 2934.200 2622.390 ;
        RECT -14.580 2619.380 2934.200 2622.380 ;
        RECT -14.580 2619.370 -11.580 2619.380 ;
        RECT 94.020 2619.370 97.020 2619.380 ;
        RECT 274.020 2619.370 277.020 2619.380 ;
        RECT 454.020 2619.370 457.020 2619.380 ;
        RECT 634.020 2619.370 637.020 2619.380 ;
        RECT 814.020 2619.370 817.020 2619.380 ;
        RECT 994.020 2619.370 997.020 2619.380 ;
        RECT 1174.020 2619.370 1177.020 2619.380 ;
        RECT 1354.020 2619.370 1357.020 2619.380 ;
        RECT 1534.020 2619.370 1537.020 2619.380 ;
        RECT 1714.020 2619.370 1717.020 2619.380 ;
        RECT 1894.020 2619.370 1897.020 2619.380 ;
        RECT 2074.020 2619.370 2077.020 2619.380 ;
        RECT 2254.020 2619.370 2257.020 2619.380 ;
        RECT 2434.020 2619.370 2437.020 2619.380 ;
        RECT 2614.020 2619.370 2617.020 2619.380 ;
        RECT 2794.020 2619.370 2797.020 2619.380 ;
        RECT 2931.200 2619.370 2934.200 2619.380 ;
        RECT -14.580 2442.380 -11.580 2442.390 ;
        RECT 94.020 2442.380 97.020 2442.390 ;
        RECT 274.020 2442.380 277.020 2442.390 ;
        RECT 454.020 2442.380 457.020 2442.390 ;
        RECT 634.020 2442.380 637.020 2442.390 ;
        RECT 814.020 2442.380 817.020 2442.390 ;
        RECT 994.020 2442.380 997.020 2442.390 ;
        RECT 1174.020 2442.380 1177.020 2442.390 ;
        RECT 1354.020 2442.380 1357.020 2442.390 ;
        RECT 1534.020 2442.380 1537.020 2442.390 ;
        RECT 1714.020 2442.380 1717.020 2442.390 ;
        RECT 1894.020 2442.380 1897.020 2442.390 ;
        RECT 2074.020 2442.380 2077.020 2442.390 ;
        RECT 2254.020 2442.380 2257.020 2442.390 ;
        RECT 2434.020 2442.380 2437.020 2442.390 ;
        RECT 2614.020 2442.380 2617.020 2442.390 ;
        RECT 2794.020 2442.380 2797.020 2442.390 ;
        RECT 2931.200 2442.380 2934.200 2442.390 ;
        RECT -14.580 2439.380 2934.200 2442.380 ;
        RECT -14.580 2439.370 -11.580 2439.380 ;
        RECT 94.020 2439.370 97.020 2439.380 ;
        RECT 274.020 2439.370 277.020 2439.380 ;
        RECT 454.020 2439.370 457.020 2439.380 ;
        RECT 634.020 2439.370 637.020 2439.380 ;
        RECT 814.020 2439.370 817.020 2439.380 ;
        RECT 994.020 2439.370 997.020 2439.380 ;
        RECT 1174.020 2439.370 1177.020 2439.380 ;
        RECT 1354.020 2439.370 1357.020 2439.380 ;
        RECT 1534.020 2439.370 1537.020 2439.380 ;
        RECT 1714.020 2439.370 1717.020 2439.380 ;
        RECT 1894.020 2439.370 1897.020 2439.380 ;
        RECT 2074.020 2439.370 2077.020 2439.380 ;
        RECT 2254.020 2439.370 2257.020 2439.380 ;
        RECT 2434.020 2439.370 2437.020 2439.380 ;
        RECT 2614.020 2439.370 2617.020 2439.380 ;
        RECT 2794.020 2439.370 2797.020 2439.380 ;
        RECT 2931.200 2439.370 2934.200 2439.380 ;
        RECT -14.580 2262.380 -11.580 2262.390 ;
        RECT 94.020 2262.380 97.020 2262.390 ;
        RECT 274.020 2262.380 277.020 2262.390 ;
        RECT 454.020 2262.380 457.020 2262.390 ;
        RECT 634.020 2262.380 637.020 2262.390 ;
        RECT 814.020 2262.380 817.020 2262.390 ;
        RECT 994.020 2262.380 997.020 2262.390 ;
        RECT 1174.020 2262.380 1177.020 2262.390 ;
        RECT 1354.020 2262.380 1357.020 2262.390 ;
        RECT 1534.020 2262.380 1537.020 2262.390 ;
        RECT 1714.020 2262.380 1717.020 2262.390 ;
        RECT 1894.020 2262.380 1897.020 2262.390 ;
        RECT 2074.020 2262.380 2077.020 2262.390 ;
        RECT 2254.020 2262.380 2257.020 2262.390 ;
        RECT 2434.020 2262.380 2437.020 2262.390 ;
        RECT 2614.020 2262.380 2617.020 2262.390 ;
        RECT 2794.020 2262.380 2797.020 2262.390 ;
        RECT 2931.200 2262.380 2934.200 2262.390 ;
        RECT -14.580 2259.380 2934.200 2262.380 ;
        RECT -14.580 2259.370 -11.580 2259.380 ;
        RECT 94.020 2259.370 97.020 2259.380 ;
        RECT 274.020 2259.370 277.020 2259.380 ;
        RECT 454.020 2259.370 457.020 2259.380 ;
        RECT 634.020 2259.370 637.020 2259.380 ;
        RECT 814.020 2259.370 817.020 2259.380 ;
        RECT 994.020 2259.370 997.020 2259.380 ;
        RECT 1174.020 2259.370 1177.020 2259.380 ;
        RECT 1354.020 2259.370 1357.020 2259.380 ;
        RECT 1534.020 2259.370 1537.020 2259.380 ;
        RECT 1714.020 2259.370 1717.020 2259.380 ;
        RECT 1894.020 2259.370 1897.020 2259.380 ;
        RECT 2074.020 2259.370 2077.020 2259.380 ;
        RECT 2254.020 2259.370 2257.020 2259.380 ;
        RECT 2434.020 2259.370 2437.020 2259.380 ;
        RECT 2614.020 2259.370 2617.020 2259.380 ;
        RECT 2794.020 2259.370 2797.020 2259.380 ;
        RECT 2931.200 2259.370 2934.200 2259.380 ;
        RECT -14.580 2082.380 -11.580 2082.390 ;
        RECT 94.020 2082.380 97.020 2082.390 ;
        RECT 274.020 2082.380 277.020 2082.390 ;
        RECT 454.020 2082.380 457.020 2082.390 ;
        RECT 634.020 2082.380 637.020 2082.390 ;
        RECT 814.020 2082.380 817.020 2082.390 ;
        RECT 994.020 2082.380 997.020 2082.390 ;
        RECT 1174.020 2082.380 1177.020 2082.390 ;
        RECT 1354.020 2082.380 1357.020 2082.390 ;
        RECT 1534.020 2082.380 1537.020 2082.390 ;
        RECT 1714.020 2082.380 1717.020 2082.390 ;
        RECT 1894.020 2082.380 1897.020 2082.390 ;
        RECT 2074.020 2082.380 2077.020 2082.390 ;
        RECT 2254.020 2082.380 2257.020 2082.390 ;
        RECT 2434.020 2082.380 2437.020 2082.390 ;
        RECT 2614.020 2082.380 2617.020 2082.390 ;
        RECT 2794.020 2082.380 2797.020 2082.390 ;
        RECT 2931.200 2082.380 2934.200 2082.390 ;
        RECT -14.580 2079.380 2934.200 2082.380 ;
        RECT -14.580 2079.370 -11.580 2079.380 ;
        RECT 94.020 2079.370 97.020 2079.380 ;
        RECT 274.020 2079.370 277.020 2079.380 ;
        RECT 454.020 2079.370 457.020 2079.380 ;
        RECT 634.020 2079.370 637.020 2079.380 ;
        RECT 814.020 2079.370 817.020 2079.380 ;
        RECT 994.020 2079.370 997.020 2079.380 ;
        RECT 1174.020 2079.370 1177.020 2079.380 ;
        RECT 1354.020 2079.370 1357.020 2079.380 ;
        RECT 1534.020 2079.370 1537.020 2079.380 ;
        RECT 1714.020 2079.370 1717.020 2079.380 ;
        RECT 1894.020 2079.370 1897.020 2079.380 ;
        RECT 2074.020 2079.370 2077.020 2079.380 ;
        RECT 2254.020 2079.370 2257.020 2079.380 ;
        RECT 2434.020 2079.370 2437.020 2079.380 ;
        RECT 2614.020 2079.370 2617.020 2079.380 ;
        RECT 2794.020 2079.370 2797.020 2079.380 ;
        RECT 2931.200 2079.370 2934.200 2079.380 ;
        RECT -14.580 1902.380 -11.580 1902.390 ;
        RECT 94.020 1902.380 97.020 1902.390 ;
        RECT 274.020 1902.380 277.020 1902.390 ;
        RECT 454.020 1902.380 457.020 1902.390 ;
        RECT 634.020 1902.380 637.020 1902.390 ;
        RECT 814.020 1902.380 817.020 1902.390 ;
        RECT 994.020 1902.380 997.020 1902.390 ;
        RECT 1174.020 1902.380 1177.020 1902.390 ;
        RECT 1354.020 1902.380 1357.020 1902.390 ;
        RECT 1534.020 1902.380 1537.020 1902.390 ;
        RECT 1714.020 1902.380 1717.020 1902.390 ;
        RECT 1894.020 1902.380 1897.020 1902.390 ;
        RECT 2074.020 1902.380 2077.020 1902.390 ;
        RECT 2254.020 1902.380 2257.020 1902.390 ;
        RECT 2434.020 1902.380 2437.020 1902.390 ;
        RECT 2614.020 1902.380 2617.020 1902.390 ;
        RECT 2794.020 1902.380 2797.020 1902.390 ;
        RECT 2931.200 1902.380 2934.200 1902.390 ;
        RECT -14.580 1899.380 2934.200 1902.380 ;
        RECT -14.580 1899.370 -11.580 1899.380 ;
        RECT 94.020 1899.370 97.020 1899.380 ;
        RECT 274.020 1899.370 277.020 1899.380 ;
        RECT 454.020 1899.370 457.020 1899.380 ;
        RECT 634.020 1899.370 637.020 1899.380 ;
        RECT 814.020 1899.370 817.020 1899.380 ;
        RECT 994.020 1899.370 997.020 1899.380 ;
        RECT 1174.020 1899.370 1177.020 1899.380 ;
        RECT 1354.020 1899.370 1357.020 1899.380 ;
        RECT 1534.020 1899.370 1537.020 1899.380 ;
        RECT 1714.020 1899.370 1717.020 1899.380 ;
        RECT 1894.020 1899.370 1897.020 1899.380 ;
        RECT 2074.020 1899.370 2077.020 1899.380 ;
        RECT 2254.020 1899.370 2257.020 1899.380 ;
        RECT 2434.020 1899.370 2437.020 1899.380 ;
        RECT 2614.020 1899.370 2617.020 1899.380 ;
        RECT 2794.020 1899.370 2797.020 1899.380 ;
        RECT 2931.200 1899.370 2934.200 1899.380 ;
        RECT -14.580 1722.380 -11.580 1722.390 ;
        RECT 94.020 1722.380 97.020 1722.390 ;
        RECT 274.020 1722.380 277.020 1722.390 ;
        RECT 454.020 1722.380 457.020 1722.390 ;
        RECT 634.020 1722.380 637.020 1722.390 ;
        RECT 814.020 1722.380 817.020 1722.390 ;
        RECT 994.020 1722.380 997.020 1722.390 ;
        RECT 1174.020 1722.380 1177.020 1722.390 ;
        RECT 1354.020 1722.380 1357.020 1722.390 ;
        RECT 1534.020 1722.380 1537.020 1722.390 ;
        RECT 1714.020 1722.380 1717.020 1722.390 ;
        RECT 1894.020 1722.380 1897.020 1722.390 ;
        RECT 2074.020 1722.380 2077.020 1722.390 ;
        RECT 2254.020 1722.380 2257.020 1722.390 ;
        RECT 2434.020 1722.380 2437.020 1722.390 ;
        RECT 2614.020 1722.380 2617.020 1722.390 ;
        RECT 2794.020 1722.380 2797.020 1722.390 ;
        RECT 2931.200 1722.380 2934.200 1722.390 ;
        RECT -14.580 1719.380 2934.200 1722.380 ;
        RECT -14.580 1719.370 -11.580 1719.380 ;
        RECT 94.020 1719.370 97.020 1719.380 ;
        RECT 274.020 1719.370 277.020 1719.380 ;
        RECT 454.020 1719.370 457.020 1719.380 ;
        RECT 634.020 1719.370 637.020 1719.380 ;
        RECT 814.020 1719.370 817.020 1719.380 ;
        RECT 994.020 1719.370 997.020 1719.380 ;
        RECT 1174.020 1719.370 1177.020 1719.380 ;
        RECT 1354.020 1719.370 1357.020 1719.380 ;
        RECT 1534.020 1719.370 1537.020 1719.380 ;
        RECT 1714.020 1719.370 1717.020 1719.380 ;
        RECT 1894.020 1719.370 1897.020 1719.380 ;
        RECT 2074.020 1719.370 2077.020 1719.380 ;
        RECT 2254.020 1719.370 2257.020 1719.380 ;
        RECT 2434.020 1719.370 2437.020 1719.380 ;
        RECT 2614.020 1719.370 2617.020 1719.380 ;
        RECT 2794.020 1719.370 2797.020 1719.380 ;
        RECT 2931.200 1719.370 2934.200 1719.380 ;
        RECT -14.580 1542.380 -11.580 1542.390 ;
        RECT 94.020 1542.380 97.020 1542.390 ;
        RECT 274.020 1542.380 277.020 1542.390 ;
        RECT 454.020 1542.380 457.020 1542.390 ;
        RECT 634.020 1542.380 637.020 1542.390 ;
        RECT 814.020 1542.380 817.020 1542.390 ;
        RECT 994.020 1542.380 997.020 1542.390 ;
        RECT 1174.020 1542.380 1177.020 1542.390 ;
        RECT 1354.020 1542.380 1357.020 1542.390 ;
        RECT 1534.020 1542.380 1537.020 1542.390 ;
        RECT 1714.020 1542.380 1717.020 1542.390 ;
        RECT 1894.020 1542.380 1897.020 1542.390 ;
        RECT 2074.020 1542.380 2077.020 1542.390 ;
        RECT 2254.020 1542.380 2257.020 1542.390 ;
        RECT 2434.020 1542.380 2437.020 1542.390 ;
        RECT 2614.020 1542.380 2617.020 1542.390 ;
        RECT 2794.020 1542.380 2797.020 1542.390 ;
        RECT 2931.200 1542.380 2934.200 1542.390 ;
        RECT -14.580 1539.380 2934.200 1542.380 ;
        RECT -14.580 1539.370 -11.580 1539.380 ;
        RECT 94.020 1539.370 97.020 1539.380 ;
        RECT 274.020 1539.370 277.020 1539.380 ;
        RECT 454.020 1539.370 457.020 1539.380 ;
        RECT 634.020 1539.370 637.020 1539.380 ;
        RECT 814.020 1539.370 817.020 1539.380 ;
        RECT 994.020 1539.370 997.020 1539.380 ;
        RECT 1174.020 1539.370 1177.020 1539.380 ;
        RECT 1354.020 1539.370 1357.020 1539.380 ;
        RECT 1534.020 1539.370 1537.020 1539.380 ;
        RECT 1714.020 1539.370 1717.020 1539.380 ;
        RECT 1894.020 1539.370 1897.020 1539.380 ;
        RECT 2074.020 1539.370 2077.020 1539.380 ;
        RECT 2254.020 1539.370 2257.020 1539.380 ;
        RECT 2434.020 1539.370 2437.020 1539.380 ;
        RECT 2614.020 1539.370 2617.020 1539.380 ;
        RECT 2794.020 1539.370 2797.020 1539.380 ;
        RECT 2931.200 1539.370 2934.200 1539.380 ;
        RECT -14.580 1362.380 -11.580 1362.390 ;
        RECT 94.020 1362.380 97.020 1362.390 ;
        RECT 274.020 1362.380 277.020 1362.390 ;
        RECT 454.020 1362.380 457.020 1362.390 ;
        RECT 634.020 1362.380 637.020 1362.390 ;
        RECT 814.020 1362.380 817.020 1362.390 ;
        RECT 994.020 1362.380 997.020 1362.390 ;
        RECT 1174.020 1362.380 1177.020 1362.390 ;
        RECT 1354.020 1362.380 1357.020 1362.390 ;
        RECT 1534.020 1362.380 1537.020 1362.390 ;
        RECT 1714.020 1362.380 1717.020 1362.390 ;
        RECT 1894.020 1362.380 1897.020 1362.390 ;
        RECT 2074.020 1362.380 2077.020 1362.390 ;
        RECT 2254.020 1362.380 2257.020 1362.390 ;
        RECT 2434.020 1362.380 2437.020 1362.390 ;
        RECT 2614.020 1362.380 2617.020 1362.390 ;
        RECT 2794.020 1362.380 2797.020 1362.390 ;
        RECT 2931.200 1362.380 2934.200 1362.390 ;
        RECT -14.580 1359.380 2934.200 1362.380 ;
        RECT -14.580 1359.370 -11.580 1359.380 ;
        RECT 94.020 1359.370 97.020 1359.380 ;
        RECT 274.020 1359.370 277.020 1359.380 ;
        RECT 454.020 1359.370 457.020 1359.380 ;
        RECT 634.020 1359.370 637.020 1359.380 ;
        RECT 814.020 1359.370 817.020 1359.380 ;
        RECT 994.020 1359.370 997.020 1359.380 ;
        RECT 1174.020 1359.370 1177.020 1359.380 ;
        RECT 1354.020 1359.370 1357.020 1359.380 ;
        RECT 1534.020 1359.370 1537.020 1359.380 ;
        RECT 1714.020 1359.370 1717.020 1359.380 ;
        RECT 1894.020 1359.370 1897.020 1359.380 ;
        RECT 2074.020 1359.370 2077.020 1359.380 ;
        RECT 2254.020 1359.370 2257.020 1359.380 ;
        RECT 2434.020 1359.370 2437.020 1359.380 ;
        RECT 2614.020 1359.370 2617.020 1359.380 ;
        RECT 2794.020 1359.370 2797.020 1359.380 ;
        RECT 2931.200 1359.370 2934.200 1359.380 ;
        RECT -14.580 1182.380 -11.580 1182.390 ;
        RECT 94.020 1182.380 97.020 1182.390 ;
        RECT 274.020 1182.380 277.020 1182.390 ;
        RECT 454.020 1182.380 457.020 1182.390 ;
        RECT 634.020 1182.380 637.020 1182.390 ;
        RECT 814.020 1182.380 817.020 1182.390 ;
        RECT 994.020 1182.380 997.020 1182.390 ;
        RECT 1174.020 1182.380 1177.020 1182.390 ;
        RECT 1354.020 1182.380 1357.020 1182.390 ;
        RECT 1534.020 1182.380 1537.020 1182.390 ;
        RECT 1714.020 1182.380 1717.020 1182.390 ;
        RECT 1894.020 1182.380 1897.020 1182.390 ;
        RECT 2074.020 1182.380 2077.020 1182.390 ;
        RECT 2254.020 1182.380 2257.020 1182.390 ;
        RECT 2434.020 1182.380 2437.020 1182.390 ;
        RECT 2614.020 1182.380 2617.020 1182.390 ;
        RECT 2794.020 1182.380 2797.020 1182.390 ;
        RECT 2931.200 1182.380 2934.200 1182.390 ;
        RECT -14.580 1179.380 2934.200 1182.380 ;
        RECT -14.580 1179.370 -11.580 1179.380 ;
        RECT 94.020 1179.370 97.020 1179.380 ;
        RECT 274.020 1179.370 277.020 1179.380 ;
        RECT 454.020 1179.370 457.020 1179.380 ;
        RECT 634.020 1179.370 637.020 1179.380 ;
        RECT 814.020 1179.370 817.020 1179.380 ;
        RECT 994.020 1179.370 997.020 1179.380 ;
        RECT 1174.020 1179.370 1177.020 1179.380 ;
        RECT 1354.020 1179.370 1357.020 1179.380 ;
        RECT 1534.020 1179.370 1537.020 1179.380 ;
        RECT 1714.020 1179.370 1717.020 1179.380 ;
        RECT 1894.020 1179.370 1897.020 1179.380 ;
        RECT 2074.020 1179.370 2077.020 1179.380 ;
        RECT 2254.020 1179.370 2257.020 1179.380 ;
        RECT 2434.020 1179.370 2437.020 1179.380 ;
        RECT 2614.020 1179.370 2617.020 1179.380 ;
        RECT 2794.020 1179.370 2797.020 1179.380 ;
        RECT 2931.200 1179.370 2934.200 1179.380 ;
        RECT -14.580 1002.380 -11.580 1002.390 ;
        RECT 94.020 1002.380 97.020 1002.390 ;
        RECT 274.020 1002.380 277.020 1002.390 ;
        RECT 454.020 1002.380 457.020 1002.390 ;
        RECT 634.020 1002.380 637.020 1002.390 ;
        RECT 814.020 1002.380 817.020 1002.390 ;
        RECT 994.020 1002.380 997.020 1002.390 ;
        RECT 1174.020 1002.380 1177.020 1002.390 ;
        RECT 1354.020 1002.380 1357.020 1002.390 ;
        RECT 1534.020 1002.380 1537.020 1002.390 ;
        RECT 1714.020 1002.380 1717.020 1002.390 ;
        RECT 1894.020 1002.380 1897.020 1002.390 ;
        RECT 2074.020 1002.380 2077.020 1002.390 ;
        RECT 2254.020 1002.380 2257.020 1002.390 ;
        RECT 2434.020 1002.380 2437.020 1002.390 ;
        RECT 2614.020 1002.380 2617.020 1002.390 ;
        RECT 2794.020 1002.380 2797.020 1002.390 ;
        RECT 2931.200 1002.380 2934.200 1002.390 ;
        RECT -14.580 999.380 2934.200 1002.380 ;
        RECT -14.580 999.370 -11.580 999.380 ;
        RECT 94.020 999.370 97.020 999.380 ;
        RECT 274.020 999.370 277.020 999.380 ;
        RECT 454.020 999.370 457.020 999.380 ;
        RECT 634.020 999.370 637.020 999.380 ;
        RECT 814.020 999.370 817.020 999.380 ;
        RECT 994.020 999.370 997.020 999.380 ;
        RECT 1174.020 999.370 1177.020 999.380 ;
        RECT 1354.020 999.370 1357.020 999.380 ;
        RECT 1534.020 999.370 1537.020 999.380 ;
        RECT 1714.020 999.370 1717.020 999.380 ;
        RECT 1894.020 999.370 1897.020 999.380 ;
        RECT 2074.020 999.370 2077.020 999.380 ;
        RECT 2254.020 999.370 2257.020 999.380 ;
        RECT 2434.020 999.370 2437.020 999.380 ;
        RECT 2614.020 999.370 2617.020 999.380 ;
        RECT 2794.020 999.370 2797.020 999.380 ;
        RECT 2931.200 999.370 2934.200 999.380 ;
        RECT -14.580 822.380 -11.580 822.390 ;
        RECT 94.020 822.380 97.020 822.390 ;
        RECT 274.020 822.380 277.020 822.390 ;
        RECT 454.020 822.380 457.020 822.390 ;
        RECT 634.020 822.380 637.020 822.390 ;
        RECT 814.020 822.380 817.020 822.390 ;
        RECT 994.020 822.380 997.020 822.390 ;
        RECT 1174.020 822.380 1177.020 822.390 ;
        RECT 1354.020 822.380 1357.020 822.390 ;
        RECT 1534.020 822.380 1537.020 822.390 ;
        RECT 1714.020 822.380 1717.020 822.390 ;
        RECT 1894.020 822.380 1897.020 822.390 ;
        RECT 2074.020 822.380 2077.020 822.390 ;
        RECT 2254.020 822.380 2257.020 822.390 ;
        RECT 2434.020 822.380 2437.020 822.390 ;
        RECT 2614.020 822.380 2617.020 822.390 ;
        RECT 2794.020 822.380 2797.020 822.390 ;
        RECT 2931.200 822.380 2934.200 822.390 ;
        RECT -14.580 819.380 2934.200 822.380 ;
        RECT -14.580 819.370 -11.580 819.380 ;
        RECT 94.020 819.370 97.020 819.380 ;
        RECT 274.020 819.370 277.020 819.380 ;
        RECT 454.020 819.370 457.020 819.380 ;
        RECT 634.020 819.370 637.020 819.380 ;
        RECT 814.020 819.370 817.020 819.380 ;
        RECT 994.020 819.370 997.020 819.380 ;
        RECT 1174.020 819.370 1177.020 819.380 ;
        RECT 1354.020 819.370 1357.020 819.380 ;
        RECT 1534.020 819.370 1537.020 819.380 ;
        RECT 1714.020 819.370 1717.020 819.380 ;
        RECT 1894.020 819.370 1897.020 819.380 ;
        RECT 2074.020 819.370 2077.020 819.380 ;
        RECT 2254.020 819.370 2257.020 819.380 ;
        RECT 2434.020 819.370 2437.020 819.380 ;
        RECT 2614.020 819.370 2617.020 819.380 ;
        RECT 2794.020 819.370 2797.020 819.380 ;
        RECT 2931.200 819.370 2934.200 819.380 ;
        RECT -14.580 642.380 -11.580 642.390 ;
        RECT 94.020 642.380 97.020 642.390 ;
        RECT 274.020 642.380 277.020 642.390 ;
        RECT 454.020 642.380 457.020 642.390 ;
        RECT 634.020 642.380 637.020 642.390 ;
        RECT 814.020 642.380 817.020 642.390 ;
        RECT 994.020 642.380 997.020 642.390 ;
        RECT 1174.020 642.380 1177.020 642.390 ;
        RECT 1354.020 642.380 1357.020 642.390 ;
        RECT 1534.020 642.380 1537.020 642.390 ;
        RECT 1714.020 642.380 1717.020 642.390 ;
        RECT 1894.020 642.380 1897.020 642.390 ;
        RECT 2074.020 642.380 2077.020 642.390 ;
        RECT 2254.020 642.380 2257.020 642.390 ;
        RECT 2434.020 642.380 2437.020 642.390 ;
        RECT 2614.020 642.380 2617.020 642.390 ;
        RECT 2794.020 642.380 2797.020 642.390 ;
        RECT 2931.200 642.380 2934.200 642.390 ;
        RECT -14.580 639.380 2934.200 642.380 ;
        RECT -14.580 639.370 -11.580 639.380 ;
        RECT 94.020 639.370 97.020 639.380 ;
        RECT 274.020 639.370 277.020 639.380 ;
        RECT 454.020 639.370 457.020 639.380 ;
        RECT 634.020 639.370 637.020 639.380 ;
        RECT 814.020 639.370 817.020 639.380 ;
        RECT 994.020 639.370 997.020 639.380 ;
        RECT 1174.020 639.370 1177.020 639.380 ;
        RECT 1354.020 639.370 1357.020 639.380 ;
        RECT 1534.020 639.370 1537.020 639.380 ;
        RECT 1714.020 639.370 1717.020 639.380 ;
        RECT 1894.020 639.370 1897.020 639.380 ;
        RECT 2074.020 639.370 2077.020 639.380 ;
        RECT 2254.020 639.370 2257.020 639.380 ;
        RECT 2434.020 639.370 2437.020 639.380 ;
        RECT 2614.020 639.370 2617.020 639.380 ;
        RECT 2794.020 639.370 2797.020 639.380 ;
        RECT 2931.200 639.370 2934.200 639.380 ;
        RECT -14.580 462.380 -11.580 462.390 ;
        RECT 94.020 462.380 97.020 462.390 ;
        RECT 274.020 462.380 277.020 462.390 ;
        RECT 454.020 462.380 457.020 462.390 ;
        RECT 634.020 462.380 637.020 462.390 ;
        RECT 814.020 462.380 817.020 462.390 ;
        RECT 994.020 462.380 997.020 462.390 ;
        RECT 1174.020 462.380 1177.020 462.390 ;
        RECT 1354.020 462.380 1357.020 462.390 ;
        RECT 1534.020 462.380 1537.020 462.390 ;
        RECT 1714.020 462.380 1717.020 462.390 ;
        RECT 1894.020 462.380 1897.020 462.390 ;
        RECT 2074.020 462.380 2077.020 462.390 ;
        RECT 2254.020 462.380 2257.020 462.390 ;
        RECT 2434.020 462.380 2437.020 462.390 ;
        RECT 2614.020 462.380 2617.020 462.390 ;
        RECT 2794.020 462.380 2797.020 462.390 ;
        RECT 2931.200 462.380 2934.200 462.390 ;
        RECT -14.580 459.380 2934.200 462.380 ;
        RECT -14.580 459.370 -11.580 459.380 ;
        RECT 94.020 459.370 97.020 459.380 ;
        RECT 274.020 459.370 277.020 459.380 ;
        RECT 454.020 459.370 457.020 459.380 ;
        RECT 634.020 459.370 637.020 459.380 ;
        RECT 814.020 459.370 817.020 459.380 ;
        RECT 994.020 459.370 997.020 459.380 ;
        RECT 1174.020 459.370 1177.020 459.380 ;
        RECT 1354.020 459.370 1357.020 459.380 ;
        RECT 1534.020 459.370 1537.020 459.380 ;
        RECT 1714.020 459.370 1717.020 459.380 ;
        RECT 1894.020 459.370 1897.020 459.380 ;
        RECT 2074.020 459.370 2077.020 459.380 ;
        RECT 2254.020 459.370 2257.020 459.380 ;
        RECT 2434.020 459.370 2437.020 459.380 ;
        RECT 2614.020 459.370 2617.020 459.380 ;
        RECT 2794.020 459.370 2797.020 459.380 ;
        RECT 2931.200 459.370 2934.200 459.380 ;
        RECT -14.580 282.380 -11.580 282.390 ;
        RECT 94.020 282.380 97.020 282.390 ;
        RECT 274.020 282.380 277.020 282.390 ;
        RECT 454.020 282.380 457.020 282.390 ;
        RECT 634.020 282.380 637.020 282.390 ;
        RECT 814.020 282.380 817.020 282.390 ;
        RECT 994.020 282.380 997.020 282.390 ;
        RECT 1174.020 282.380 1177.020 282.390 ;
        RECT 1354.020 282.380 1357.020 282.390 ;
        RECT 1534.020 282.380 1537.020 282.390 ;
        RECT 1714.020 282.380 1717.020 282.390 ;
        RECT 1894.020 282.380 1897.020 282.390 ;
        RECT 2074.020 282.380 2077.020 282.390 ;
        RECT 2254.020 282.380 2257.020 282.390 ;
        RECT 2434.020 282.380 2437.020 282.390 ;
        RECT 2614.020 282.380 2617.020 282.390 ;
        RECT 2794.020 282.380 2797.020 282.390 ;
        RECT 2931.200 282.380 2934.200 282.390 ;
        RECT -14.580 279.380 2934.200 282.380 ;
        RECT -14.580 279.370 -11.580 279.380 ;
        RECT 94.020 279.370 97.020 279.380 ;
        RECT 274.020 279.370 277.020 279.380 ;
        RECT 454.020 279.370 457.020 279.380 ;
        RECT 634.020 279.370 637.020 279.380 ;
        RECT 814.020 279.370 817.020 279.380 ;
        RECT 994.020 279.370 997.020 279.380 ;
        RECT 1174.020 279.370 1177.020 279.380 ;
        RECT 1354.020 279.370 1357.020 279.380 ;
        RECT 1534.020 279.370 1537.020 279.380 ;
        RECT 1714.020 279.370 1717.020 279.380 ;
        RECT 1894.020 279.370 1897.020 279.380 ;
        RECT 2074.020 279.370 2077.020 279.380 ;
        RECT 2254.020 279.370 2257.020 279.380 ;
        RECT 2434.020 279.370 2437.020 279.380 ;
        RECT 2614.020 279.370 2617.020 279.380 ;
        RECT 2794.020 279.370 2797.020 279.380 ;
        RECT 2931.200 279.370 2934.200 279.380 ;
        RECT -14.580 102.380 -11.580 102.390 ;
        RECT 94.020 102.380 97.020 102.390 ;
        RECT 274.020 102.380 277.020 102.390 ;
        RECT 454.020 102.380 457.020 102.390 ;
        RECT 634.020 102.380 637.020 102.390 ;
        RECT 814.020 102.380 817.020 102.390 ;
        RECT 994.020 102.380 997.020 102.390 ;
        RECT 1174.020 102.380 1177.020 102.390 ;
        RECT 1354.020 102.380 1357.020 102.390 ;
        RECT 1534.020 102.380 1537.020 102.390 ;
        RECT 1714.020 102.380 1717.020 102.390 ;
        RECT 1894.020 102.380 1897.020 102.390 ;
        RECT 2074.020 102.380 2077.020 102.390 ;
        RECT 2254.020 102.380 2257.020 102.390 ;
        RECT 2434.020 102.380 2437.020 102.390 ;
        RECT 2614.020 102.380 2617.020 102.390 ;
        RECT 2794.020 102.380 2797.020 102.390 ;
        RECT 2931.200 102.380 2934.200 102.390 ;
        RECT -14.580 99.380 2934.200 102.380 ;
        RECT -14.580 99.370 -11.580 99.380 ;
        RECT 94.020 99.370 97.020 99.380 ;
        RECT 274.020 99.370 277.020 99.380 ;
        RECT 454.020 99.370 457.020 99.380 ;
        RECT 634.020 99.370 637.020 99.380 ;
        RECT 814.020 99.370 817.020 99.380 ;
        RECT 994.020 99.370 997.020 99.380 ;
        RECT 1174.020 99.370 1177.020 99.380 ;
        RECT 1354.020 99.370 1357.020 99.380 ;
        RECT 1534.020 99.370 1537.020 99.380 ;
        RECT 1714.020 99.370 1717.020 99.380 ;
        RECT 1894.020 99.370 1897.020 99.380 ;
        RECT 2074.020 99.370 2077.020 99.380 ;
        RECT 2254.020 99.370 2257.020 99.380 ;
        RECT 2434.020 99.370 2437.020 99.380 ;
        RECT 2614.020 99.370 2617.020 99.380 ;
        RECT 2794.020 99.370 2797.020 99.380 ;
        RECT 2931.200 99.370 2934.200 99.380 ;
        RECT -14.580 -6.220 -11.580 -6.210 ;
        RECT 94.020 -6.220 97.020 -6.210 ;
        RECT 274.020 -6.220 277.020 -6.210 ;
        RECT 454.020 -6.220 457.020 -6.210 ;
        RECT 634.020 -6.220 637.020 -6.210 ;
        RECT 814.020 -6.220 817.020 -6.210 ;
        RECT 994.020 -6.220 997.020 -6.210 ;
        RECT 1174.020 -6.220 1177.020 -6.210 ;
        RECT 1354.020 -6.220 1357.020 -6.210 ;
        RECT 1534.020 -6.220 1537.020 -6.210 ;
        RECT 1714.020 -6.220 1717.020 -6.210 ;
        RECT 1894.020 -6.220 1897.020 -6.210 ;
        RECT 2074.020 -6.220 2077.020 -6.210 ;
        RECT 2254.020 -6.220 2257.020 -6.210 ;
        RECT 2434.020 -6.220 2437.020 -6.210 ;
        RECT 2614.020 -6.220 2617.020 -6.210 ;
        RECT 2794.020 -6.220 2797.020 -6.210 ;
        RECT 2931.200 -6.220 2934.200 -6.210 ;
        RECT -14.580 -9.220 2934.200 -6.220 ;
        RECT -14.580 -9.230 -11.580 -9.220 ;
        RECT 94.020 -9.230 97.020 -9.220 ;
        RECT 274.020 -9.230 277.020 -9.220 ;
        RECT 454.020 -9.230 457.020 -9.220 ;
        RECT 634.020 -9.230 637.020 -9.220 ;
        RECT 814.020 -9.230 817.020 -9.220 ;
        RECT 994.020 -9.230 997.020 -9.220 ;
        RECT 1174.020 -9.230 1177.020 -9.220 ;
        RECT 1354.020 -9.230 1357.020 -9.220 ;
        RECT 1534.020 -9.230 1537.020 -9.220 ;
        RECT 1714.020 -9.230 1717.020 -9.220 ;
        RECT 1894.020 -9.230 1897.020 -9.220 ;
        RECT 2074.020 -9.230 2077.020 -9.220 ;
        RECT 2254.020 -9.230 2257.020 -9.220 ;
        RECT 2434.020 -9.230 2437.020 -9.220 ;
        RECT 2614.020 -9.230 2617.020 -9.220 ;
        RECT 2794.020 -9.230 2797.020 -9.220 ;
        RECT 2931.200 -9.230 2934.200 -9.220 ;
    END
  END vssd1
  PIN vccd2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -19.180 -13.820 -16.180 3533.500 ;
        RECT 22.020 -18.420 25.020 3538.100 ;
        RECT 202.020 -18.420 205.020 3538.100 ;
        RECT 382.020 -18.420 385.020 3538.100 ;
        RECT 562.020 -18.420 565.020 3538.100 ;
        RECT 742.020 -18.420 745.020 3538.100 ;
        RECT 922.020 -18.420 925.020 3538.100 ;
        RECT 1102.020 -18.420 1105.020 3538.100 ;
        RECT 1282.020 -18.420 1285.020 3538.100 ;
        RECT 1462.020 -18.420 1465.020 3538.100 ;
        RECT 1642.020 -18.420 1645.020 3538.100 ;
        RECT 1822.020 -18.420 1825.020 3538.100 ;
        RECT 2002.020 -18.420 2005.020 3538.100 ;
        RECT 2182.020 -18.420 2185.020 3538.100 ;
        RECT 2362.020 -18.420 2365.020 3538.100 ;
        RECT 2542.020 -18.420 2545.020 3538.100 ;
        RECT 2722.020 -18.420 2725.020 3538.100 ;
        RECT 2902.020 -18.420 2905.020 3538.100 ;
        RECT 2935.800 -13.820 2938.800 3533.500 ;
      LAYER via4 ;
        RECT -18.270 3532.210 -17.090 3533.390 ;
        RECT -18.270 3530.610 -17.090 3531.790 ;
        RECT -18.270 3449.090 -17.090 3450.270 ;
        RECT -18.270 3447.490 -17.090 3448.670 ;
        RECT -18.270 3269.090 -17.090 3270.270 ;
        RECT -18.270 3267.490 -17.090 3268.670 ;
        RECT -18.270 3089.090 -17.090 3090.270 ;
        RECT -18.270 3087.490 -17.090 3088.670 ;
        RECT -18.270 2909.090 -17.090 2910.270 ;
        RECT -18.270 2907.490 -17.090 2908.670 ;
        RECT -18.270 2729.090 -17.090 2730.270 ;
        RECT -18.270 2727.490 -17.090 2728.670 ;
        RECT -18.270 2549.090 -17.090 2550.270 ;
        RECT -18.270 2547.490 -17.090 2548.670 ;
        RECT -18.270 2369.090 -17.090 2370.270 ;
        RECT -18.270 2367.490 -17.090 2368.670 ;
        RECT -18.270 2189.090 -17.090 2190.270 ;
        RECT -18.270 2187.490 -17.090 2188.670 ;
        RECT -18.270 2009.090 -17.090 2010.270 ;
        RECT -18.270 2007.490 -17.090 2008.670 ;
        RECT -18.270 1829.090 -17.090 1830.270 ;
        RECT -18.270 1827.490 -17.090 1828.670 ;
        RECT -18.270 1649.090 -17.090 1650.270 ;
        RECT -18.270 1647.490 -17.090 1648.670 ;
        RECT -18.270 1469.090 -17.090 1470.270 ;
        RECT -18.270 1467.490 -17.090 1468.670 ;
        RECT -18.270 1289.090 -17.090 1290.270 ;
        RECT -18.270 1287.490 -17.090 1288.670 ;
        RECT -18.270 1109.090 -17.090 1110.270 ;
        RECT -18.270 1107.490 -17.090 1108.670 ;
        RECT -18.270 929.090 -17.090 930.270 ;
        RECT -18.270 927.490 -17.090 928.670 ;
        RECT -18.270 749.090 -17.090 750.270 ;
        RECT -18.270 747.490 -17.090 748.670 ;
        RECT -18.270 569.090 -17.090 570.270 ;
        RECT -18.270 567.490 -17.090 568.670 ;
        RECT -18.270 389.090 -17.090 390.270 ;
        RECT -18.270 387.490 -17.090 388.670 ;
        RECT -18.270 209.090 -17.090 210.270 ;
        RECT -18.270 207.490 -17.090 208.670 ;
        RECT -18.270 29.090 -17.090 30.270 ;
        RECT -18.270 27.490 -17.090 28.670 ;
        RECT -18.270 -12.110 -17.090 -10.930 ;
        RECT -18.270 -13.710 -17.090 -12.530 ;
        RECT 22.930 3532.210 24.110 3533.390 ;
        RECT 22.930 3530.610 24.110 3531.790 ;
        RECT 22.930 3449.090 24.110 3450.270 ;
        RECT 22.930 3447.490 24.110 3448.670 ;
        RECT 22.930 3269.090 24.110 3270.270 ;
        RECT 22.930 3267.490 24.110 3268.670 ;
        RECT 22.930 3089.090 24.110 3090.270 ;
        RECT 22.930 3087.490 24.110 3088.670 ;
        RECT 22.930 2909.090 24.110 2910.270 ;
        RECT 22.930 2907.490 24.110 2908.670 ;
        RECT 22.930 2729.090 24.110 2730.270 ;
        RECT 22.930 2727.490 24.110 2728.670 ;
        RECT 22.930 2549.090 24.110 2550.270 ;
        RECT 22.930 2547.490 24.110 2548.670 ;
        RECT 22.930 2369.090 24.110 2370.270 ;
        RECT 22.930 2367.490 24.110 2368.670 ;
        RECT 22.930 2189.090 24.110 2190.270 ;
        RECT 22.930 2187.490 24.110 2188.670 ;
        RECT 22.930 2009.090 24.110 2010.270 ;
        RECT 22.930 2007.490 24.110 2008.670 ;
        RECT 22.930 1829.090 24.110 1830.270 ;
        RECT 22.930 1827.490 24.110 1828.670 ;
        RECT 22.930 1649.090 24.110 1650.270 ;
        RECT 22.930 1647.490 24.110 1648.670 ;
        RECT 22.930 1469.090 24.110 1470.270 ;
        RECT 22.930 1467.490 24.110 1468.670 ;
        RECT 22.930 1289.090 24.110 1290.270 ;
        RECT 22.930 1287.490 24.110 1288.670 ;
        RECT 22.930 1109.090 24.110 1110.270 ;
        RECT 22.930 1107.490 24.110 1108.670 ;
        RECT 22.930 929.090 24.110 930.270 ;
        RECT 22.930 927.490 24.110 928.670 ;
        RECT 22.930 749.090 24.110 750.270 ;
        RECT 22.930 747.490 24.110 748.670 ;
        RECT 22.930 569.090 24.110 570.270 ;
        RECT 22.930 567.490 24.110 568.670 ;
        RECT 22.930 389.090 24.110 390.270 ;
        RECT 22.930 387.490 24.110 388.670 ;
        RECT 22.930 209.090 24.110 210.270 ;
        RECT 22.930 207.490 24.110 208.670 ;
        RECT 22.930 29.090 24.110 30.270 ;
        RECT 22.930 27.490 24.110 28.670 ;
        RECT 22.930 -12.110 24.110 -10.930 ;
        RECT 22.930 -13.710 24.110 -12.530 ;
        RECT 202.930 3532.210 204.110 3533.390 ;
        RECT 202.930 3530.610 204.110 3531.790 ;
        RECT 202.930 3449.090 204.110 3450.270 ;
        RECT 202.930 3447.490 204.110 3448.670 ;
        RECT 202.930 3269.090 204.110 3270.270 ;
        RECT 202.930 3267.490 204.110 3268.670 ;
        RECT 202.930 3089.090 204.110 3090.270 ;
        RECT 202.930 3087.490 204.110 3088.670 ;
        RECT 202.930 2909.090 204.110 2910.270 ;
        RECT 202.930 2907.490 204.110 2908.670 ;
        RECT 202.930 2729.090 204.110 2730.270 ;
        RECT 202.930 2727.490 204.110 2728.670 ;
        RECT 202.930 2549.090 204.110 2550.270 ;
        RECT 202.930 2547.490 204.110 2548.670 ;
        RECT 202.930 2369.090 204.110 2370.270 ;
        RECT 202.930 2367.490 204.110 2368.670 ;
        RECT 202.930 2189.090 204.110 2190.270 ;
        RECT 202.930 2187.490 204.110 2188.670 ;
        RECT 202.930 2009.090 204.110 2010.270 ;
        RECT 202.930 2007.490 204.110 2008.670 ;
        RECT 202.930 1829.090 204.110 1830.270 ;
        RECT 202.930 1827.490 204.110 1828.670 ;
        RECT 202.930 1649.090 204.110 1650.270 ;
        RECT 202.930 1647.490 204.110 1648.670 ;
        RECT 202.930 1469.090 204.110 1470.270 ;
        RECT 202.930 1467.490 204.110 1468.670 ;
        RECT 202.930 1289.090 204.110 1290.270 ;
        RECT 202.930 1287.490 204.110 1288.670 ;
        RECT 202.930 1109.090 204.110 1110.270 ;
        RECT 202.930 1107.490 204.110 1108.670 ;
        RECT 202.930 929.090 204.110 930.270 ;
        RECT 202.930 927.490 204.110 928.670 ;
        RECT 202.930 749.090 204.110 750.270 ;
        RECT 202.930 747.490 204.110 748.670 ;
        RECT 202.930 569.090 204.110 570.270 ;
        RECT 202.930 567.490 204.110 568.670 ;
        RECT 202.930 389.090 204.110 390.270 ;
        RECT 202.930 387.490 204.110 388.670 ;
        RECT 202.930 209.090 204.110 210.270 ;
        RECT 202.930 207.490 204.110 208.670 ;
        RECT 202.930 29.090 204.110 30.270 ;
        RECT 202.930 27.490 204.110 28.670 ;
        RECT 202.930 -12.110 204.110 -10.930 ;
        RECT 202.930 -13.710 204.110 -12.530 ;
        RECT 382.930 3532.210 384.110 3533.390 ;
        RECT 382.930 3530.610 384.110 3531.790 ;
        RECT 382.930 3449.090 384.110 3450.270 ;
        RECT 382.930 3447.490 384.110 3448.670 ;
        RECT 382.930 3269.090 384.110 3270.270 ;
        RECT 382.930 3267.490 384.110 3268.670 ;
        RECT 382.930 3089.090 384.110 3090.270 ;
        RECT 382.930 3087.490 384.110 3088.670 ;
        RECT 382.930 2909.090 384.110 2910.270 ;
        RECT 382.930 2907.490 384.110 2908.670 ;
        RECT 382.930 2729.090 384.110 2730.270 ;
        RECT 382.930 2727.490 384.110 2728.670 ;
        RECT 382.930 2549.090 384.110 2550.270 ;
        RECT 382.930 2547.490 384.110 2548.670 ;
        RECT 382.930 2369.090 384.110 2370.270 ;
        RECT 382.930 2367.490 384.110 2368.670 ;
        RECT 382.930 2189.090 384.110 2190.270 ;
        RECT 382.930 2187.490 384.110 2188.670 ;
        RECT 382.930 2009.090 384.110 2010.270 ;
        RECT 382.930 2007.490 384.110 2008.670 ;
        RECT 382.930 1829.090 384.110 1830.270 ;
        RECT 382.930 1827.490 384.110 1828.670 ;
        RECT 382.930 1649.090 384.110 1650.270 ;
        RECT 382.930 1647.490 384.110 1648.670 ;
        RECT 382.930 1469.090 384.110 1470.270 ;
        RECT 382.930 1467.490 384.110 1468.670 ;
        RECT 382.930 1289.090 384.110 1290.270 ;
        RECT 382.930 1287.490 384.110 1288.670 ;
        RECT 382.930 1109.090 384.110 1110.270 ;
        RECT 382.930 1107.490 384.110 1108.670 ;
        RECT 382.930 929.090 384.110 930.270 ;
        RECT 382.930 927.490 384.110 928.670 ;
        RECT 382.930 749.090 384.110 750.270 ;
        RECT 382.930 747.490 384.110 748.670 ;
        RECT 382.930 569.090 384.110 570.270 ;
        RECT 382.930 567.490 384.110 568.670 ;
        RECT 382.930 389.090 384.110 390.270 ;
        RECT 382.930 387.490 384.110 388.670 ;
        RECT 382.930 209.090 384.110 210.270 ;
        RECT 382.930 207.490 384.110 208.670 ;
        RECT 382.930 29.090 384.110 30.270 ;
        RECT 382.930 27.490 384.110 28.670 ;
        RECT 382.930 -12.110 384.110 -10.930 ;
        RECT 382.930 -13.710 384.110 -12.530 ;
        RECT 562.930 3532.210 564.110 3533.390 ;
        RECT 562.930 3530.610 564.110 3531.790 ;
        RECT 562.930 3449.090 564.110 3450.270 ;
        RECT 562.930 3447.490 564.110 3448.670 ;
        RECT 562.930 3269.090 564.110 3270.270 ;
        RECT 562.930 3267.490 564.110 3268.670 ;
        RECT 562.930 3089.090 564.110 3090.270 ;
        RECT 562.930 3087.490 564.110 3088.670 ;
        RECT 562.930 2909.090 564.110 2910.270 ;
        RECT 562.930 2907.490 564.110 2908.670 ;
        RECT 562.930 2729.090 564.110 2730.270 ;
        RECT 562.930 2727.490 564.110 2728.670 ;
        RECT 562.930 2549.090 564.110 2550.270 ;
        RECT 562.930 2547.490 564.110 2548.670 ;
        RECT 562.930 2369.090 564.110 2370.270 ;
        RECT 562.930 2367.490 564.110 2368.670 ;
        RECT 562.930 2189.090 564.110 2190.270 ;
        RECT 562.930 2187.490 564.110 2188.670 ;
        RECT 562.930 2009.090 564.110 2010.270 ;
        RECT 562.930 2007.490 564.110 2008.670 ;
        RECT 562.930 1829.090 564.110 1830.270 ;
        RECT 562.930 1827.490 564.110 1828.670 ;
        RECT 562.930 1649.090 564.110 1650.270 ;
        RECT 562.930 1647.490 564.110 1648.670 ;
        RECT 562.930 1469.090 564.110 1470.270 ;
        RECT 562.930 1467.490 564.110 1468.670 ;
        RECT 562.930 1289.090 564.110 1290.270 ;
        RECT 562.930 1287.490 564.110 1288.670 ;
        RECT 562.930 1109.090 564.110 1110.270 ;
        RECT 562.930 1107.490 564.110 1108.670 ;
        RECT 562.930 929.090 564.110 930.270 ;
        RECT 562.930 927.490 564.110 928.670 ;
        RECT 562.930 749.090 564.110 750.270 ;
        RECT 562.930 747.490 564.110 748.670 ;
        RECT 562.930 569.090 564.110 570.270 ;
        RECT 562.930 567.490 564.110 568.670 ;
        RECT 562.930 389.090 564.110 390.270 ;
        RECT 562.930 387.490 564.110 388.670 ;
        RECT 562.930 209.090 564.110 210.270 ;
        RECT 562.930 207.490 564.110 208.670 ;
        RECT 562.930 29.090 564.110 30.270 ;
        RECT 562.930 27.490 564.110 28.670 ;
        RECT 562.930 -12.110 564.110 -10.930 ;
        RECT 562.930 -13.710 564.110 -12.530 ;
        RECT 742.930 3532.210 744.110 3533.390 ;
        RECT 742.930 3530.610 744.110 3531.790 ;
        RECT 742.930 3449.090 744.110 3450.270 ;
        RECT 742.930 3447.490 744.110 3448.670 ;
        RECT 742.930 3269.090 744.110 3270.270 ;
        RECT 742.930 3267.490 744.110 3268.670 ;
        RECT 742.930 3089.090 744.110 3090.270 ;
        RECT 742.930 3087.490 744.110 3088.670 ;
        RECT 742.930 2909.090 744.110 2910.270 ;
        RECT 742.930 2907.490 744.110 2908.670 ;
        RECT 742.930 2729.090 744.110 2730.270 ;
        RECT 742.930 2727.490 744.110 2728.670 ;
        RECT 742.930 2549.090 744.110 2550.270 ;
        RECT 742.930 2547.490 744.110 2548.670 ;
        RECT 742.930 2369.090 744.110 2370.270 ;
        RECT 742.930 2367.490 744.110 2368.670 ;
        RECT 742.930 2189.090 744.110 2190.270 ;
        RECT 742.930 2187.490 744.110 2188.670 ;
        RECT 742.930 2009.090 744.110 2010.270 ;
        RECT 742.930 2007.490 744.110 2008.670 ;
        RECT 742.930 1829.090 744.110 1830.270 ;
        RECT 742.930 1827.490 744.110 1828.670 ;
        RECT 742.930 1649.090 744.110 1650.270 ;
        RECT 742.930 1647.490 744.110 1648.670 ;
        RECT 742.930 1469.090 744.110 1470.270 ;
        RECT 742.930 1467.490 744.110 1468.670 ;
        RECT 742.930 1289.090 744.110 1290.270 ;
        RECT 742.930 1287.490 744.110 1288.670 ;
        RECT 742.930 1109.090 744.110 1110.270 ;
        RECT 742.930 1107.490 744.110 1108.670 ;
        RECT 742.930 929.090 744.110 930.270 ;
        RECT 742.930 927.490 744.110 928.670 ;
        RECT 742.930 749.090 744.110 750.270 ;
        RECT 742.930 747.490 744.110 748.670 ;
        RECT 742.930 569.090 744.110 570.270 ;
        RECT 742.930 567.490 744.110 568.670 ;
        RECT 742.930 389.090 744.110 390.270 ;
        RECT 742.930 387.490 744.110 388.670 ;
        RECT 742.930 209.090 744.110 210.270 ;
        RECT 742.930 207.490 744.110 208.670 ;
        RECT 742.930 29.090 744.110 30.270 ;
        RECT 742.930 27.490 744.110 28.670 ;
        RECT 742.930 -12.110 744.110 -10.930 ;
        RECT 742.930 -13.710 744.110 -12.530 ;
        RECT 922.930 3532.210 924.110 3533.390 ;
        RECT 922.930 3530.610 924.110 3531.790 ;
        RECT 922.930 3449.090 924.110 3450.270 ;
        RECT 922.930 3447.490 924.110 3448.670 ;
        RECT 922.930 3269.090 924.110 3270.270 ;
        RECT 922.930 3267.490 924.110 3268.670 ;
        RECT 922.930 3089.090 924.110 3090.270 ;
        RECT 922.930 3087.490 924.110 3088.670 ;
        RECT 922.930 2909.090 924.110 2910.270 ;
        RECT 922.930 2907.490 924.110 2908.670 ;
        RECT 922.930 2729.090 924.110 2730.270 ;
        RECT 922.930 2727.490 924.110 2728.670 ;
        RECT 922.930 2549.090 924.110 2550.270 ;
        RECT 922.930 2547.490 924.110 2548.670 ;
        RECT 922.930 2369.090 924.110 2370.270 ;
        RECT 922.930 2367.490 924.110 2368.670 ;
        RECT 922.930 2189.090 924.110 2190.270 ;
        RECT 922.930 2187.490 924.110 2188.670 ;
        RECT 922.930 2009.090 924.110 2010.270 ;
        RECT 922.930 2007.490 924.110 2008.670 ;
        RECT 922.930 1829.090 924.110 1830.270 ;
        RECT 922.930 1827.490 924.110 1828.670 ;
        RECT 922.930 1649.090 924.110 1650.270 ;
        RECT 922.930 1647.490 924.110 1648.670 ;
        RECT 922.930 1469.090 924.110 1470.270 ;
        RECT 922.930 1467.490 924.110 1468.670 ;
        RECT 922.930 1289.090 924.110 1290.270 ;
        RECT 922.930 1287.490 924.110 1288.670 ;
        RECT 922.930 1109.090 924.110 1110.270 ;
        RECT 922.930 1107.490 924.110 1108.670 ;
        RECT 922.930 929.090 924.110 930.270 ;
        RECT 922.930 927.490 924.110 928.670 ;
        RECT 922.930 749.090 924.110 750.270 ;
        RECT 922.930 747.490 924.110 748.670 ;
        RECT 922.930 569.090 924.110 570.270 ;
        RECT 922.930 567.490 924.110 568.670 ;
        RECT 922.930 389.090 924.110 390.270 ;
        RECT 922.930 387.490 924.110 388.670 ;
        RECT 922.930 209.090 924.110 210.270 ;
        RECT 922.930 207.490 924.110 208.670 ;
        RECT 922.930 29.090 924.110 30.270 ;
        RECT 922.930 27.490 924.110 28.670 ;
        RECT 922.930 -12.110 924.110 -10.930 ;
        RECT 922.930 -13.710 924.110 -12.530 ;
        RECT 1102.930 3532.210 1104.110 3533.390 ;
        RECT 1102.930 3530.610 1104.110 3531.790 ;
        RECT 1102.930 3449.090 1104.110 3450.270 ;
        RECT 1102.930 3447.490 1104.110 3448.670 ;
        RECT 1102.930 3269.090 1104.110 3270.270 ;
        RECT 1102.930 3267.490 1104.110 3268.670 ;
        RECT 1102.930 3089.090 1104.110 3090.270 ;
        RECT 1102.930 3087.490 1104.110 3088.670 ;
        RECT 1102.930 2909.090 1104.110 2910.270 ;
        RECT 1102.930 2907.490 1104.110 2908.670 ;
        RECT 1102.930 2729.090 1104.110 2730.270 ;
        RECT 1102.930 2727.490 1104.110 2728.670 ;
        RECT 1102.930 2549.090 1104.110 2550.270 ;
        RECT 1102.930 2547.490 1104.110 2548.670 ;
        RECT 1102.930 2369.090 1104.110 2370.270 ;
        RECT 1102.930 2367.490 1104.110 2368.670 ;
        RECT 1102.930 2189.090 1104.110 2190.270 ;
        RECT 1102.930 2187.490 1104.110 2188.670 ;
        RECT 1102.930 2009.090 1104.110 2010.270 ;
        RECT 1102.930 2007.490 1104.110 2008.670 ;
        RECT 1102.930 1829.090 1104.110 1830.270 ;
        RECT 1102.930 1827.490 1104.110 1828.670 ;
        RECT 1102.930 1649.090 1104.110 1650.270 ;
        RECT 1102.930 1647.490 1104.110 1648.670 ;
        RECT 1102.930 1469.090 1104.110 1470.270 ;
        RECT 1102.930 1467.490 1104.110 1468.670 ;
        RECT 1102.930 1289.090 1104.110 1290.270 ;
        RECT 1102.930 1287.490 1104.110 1288.670 ;
        RECT 1102.930 1109.090 1104.110 1110.270 ;
        RECT 1102.930 1107.490 1104.110 1108.670 ;
        RECT 1102.930 929.090 1104.110 930.270 ;
        RECT 1102.930 927.490 1104.110 928.670 ;
        RECT 1102.930 749.090 1104.110 750.270 ;
        RECT 1102.930 747.490 1104.110 748.670 ;
        RECT 1102.930 569.090 1104.110 570.270 ;
        RECT 1102.930 567.490 1104.110 568.670 ;
        RECT 1102.930 389.090 1104.110 390.270 ;
        RECT 1102.930 387.490 1104.110 388.670 ;
        RECT 1102.930 209.090 1104.110 210.270 ;
        RECT 1102.930 207.490 1104.110 208.670 ;
        RECT 1102.930 29.090 1104.110 30.270 ;
        RECT 1102.930 27.490 1104.110 28.670 ;
        RECT 1102.930 -12.110 1104.110 -10.930 ;
        RECT 1102.930 -13.710 1104.110 -12.530 ;
        RECT 1282.930 3532.210 1284.110 3533.390 ;
        RECT 1282.930 3530.610 1284.110 3531.790 ;
        RECT 1282.930 3449.090 1284.110 3450.270 ;
        RECT 1282.930 3447.490 1284.110 3448.670 ;
        RECT 1282.930 3269.090 1284.110 3270.270 ;
        RECT 1282.930 3267.490 1284.110 3268.670 ;
        RECT 1282.930 3089.090 1284.110 3090.270 ;
        RECT 1282.930 3087.490 1284.110 3088.670 ;
        RECT 1282.930 2909.090 1284.110 2910.270 ;
        RECT 1282.930 2907.490 1284.110 2908.670 ;
        RECT 1282.930 2729.090 1284.110 2730.270 ;
        RECT 1282.930 2727.490 1284.110 2728.670 ;
        RECT 1282.930 2549.090 1284.110 2550.270 ;
        RECT 1282.930 2547.490 1284.110 2548.670 ;
        RECT 1282.930 2369.090 1284.110 2370.270 ;
        RECT 1282.930 2367.490 1284.110 2368.670 ;
        RECT 1282.930 2189.090 1284.110 2190.270 ;
        RECT 1282.930 2187.490 1284.110 2188.670 ;
        RECT 1282.930 2009.090 1284.110 2010.270 ;
        RECT 1282.930 2007.490 1284.110 2008.670 ;
        RECT 1282.930 1829.090 1284.110 1830.270 ;
        RECT 1282.930 1827.490 1284.110 1828.670 ;
        RECT 1282.930 1649.090 1284.110 1650.270 ;
        RECT 1282.930 1647.490 1284.110 1648.670 ;
        RECT 1282.930 1469.090 1284.110 1470.270 ;
        RECT 1282.930 1467.490 1284.110 1468.670 ;
        RECT 1282.930 1289.090 1284.110 1290.270 ;
        RECT 1282.930 1287.490 1284.110 1288.670 ;
        RECT 1282.930 1109.090 1284.110 1110.270 ;
        RECT 1282.930 1107.490 1284.110 1108.670 ;
        RECT 1282.930 929.090 1284.110 930.270 ;
        RECT 1282.930 927.490 1284.110 928.670 ;
        RECT 1282.930 749.090 1284.110 750.270 ;
        RECT 1282.930 747.490 1284.110 748.670 ;
        RECT 1282.930 569.090 1284.110 570.270 ;
        RECT 1282.930 567.490 1284.110 568.670 ;
        RECT 1282.930 389.090 1284.110 390.270 ;
        RECT 1282.930 387.490 1284.110 388.670 ;
        RECT 1282.930 209.090 1284.110 210.270 ;
        RECT 1282.930 207.490 1284.110 208.670 ;
        RECT 1282.930 29.090 1284.110 30.270 ;
        RECT 1282.930 27.490 1284.110 28.670 ;
        RECT 1282.930 -12.110 1284.110 -10.930 ;
        RECT 1282.930 -13.710 1284.110 -12.530 ;
        RECT 1462.930 3532.210 1464.110 3533.390 ;
        RECT 1462.930 3530.610 1464.110 3531.790 ;
        RECT 1462.930 3449.090 1464.110 3450.270 ;
        RECT 1462.930 3447.490 1464.110 3448.670 ;
        RECT 1462.930 3269.090 1464.110 3270.270 ;
        RECT 1462.930 3267.490 1464.110 3268.670 ;
        RECT 1462.930 3089.090 1464.110 3090.270 ;
        RECT 1462.930 3087.490 1464.110 3088.670 ;
        RECT 1462.930 2909.090 1464.110 2910.270 ;
        RECT 1462.930 2907.490 1464.110 2908.670 ;
        RECT 1462.930 2729.090 1464.110 2730.270 ;
        RECT 1462.930 2727.490 1464.110 2728.670 ;
        RECT 1462.930 2549.090 1464.110 2550.270 ;
        RECT 1462.930 2547.490 1464.110 2548.670 ;
        RECT 1462.930 2369.090 1464.110 2370.270 ;
        RECT 1462.930 2367.490 1464.110 2368.670 ;
        RECT 1462.930 2189.090 1464.110 2190.270 ;
        RECT 1462.930 2187.490 1464.110 2188.670 ;
        RECT 1462.930 2009.090 1464.110 2010.270 ;
        RECT 1462.930 2007.490 1464.110 2008.670 ;
        RECT 1462.930 1829.090 1464.110 1830.270 ;
        RECT 1462.930 1827.490 1464.110 1828.670 ;
        RECT 1462.930 1649.090 1464.110 1650.270 ;
        RECT 1462.930 1647.490 1464.110 1648.670 ;
        RECT 1462.930 1469.090 1464.110 1470.270 ;
        RECT 1462.930 1467.490 1464.110 1468.670 ;
        RECT 1462.930 1289.090 1464.110 1290.270 ;
        RECT 1462.930 1287.490 1464.110 1288.670 ;
        RECT 1462.930 1109.090 1464.110 1110.270 ;
        RECT 1462.930 1107.490 1464.110 1108.670 ;
        RECT 1462.930 929.090 1464.110 930.270 ;
        RECT 1462.930 927.490 1464.110 928.670 ;
        RECT 1462.930 749.090 1464.110 750.270 ;
        RECT 1462.930 747.490 1464.110 748.670 ;
        RECT 1462.930 569.090 1464.110 570.270 ;
        RECT 1462.930 567.490 1464.110 568.670 ;
        RECT 1462.930 389.090 1464.110 390.270 ;
        RECT 1462.930 387.490 1464.110 388.670 ;
        RECT 1462.930 209.090 1464.110 210.270 ;
        RECT 1462.930 207.490 1464.110 208.670 ;
        RECT 1462.930 29.090 1464.110 30.270 ;
        RECT 1462.930 27.490 1464.110 28.670 ;
        RECT 1462.930 -12.110 1464.110 -10.930 ;
        RECT 1462.930 -13.710 1464.110 -12.530 ;
        RECT 1642.930 3532.210 1644.110 3533.390 ;
        RECT 1642.930 3530.610 1644.110 3531.790 ;
        RECT 1642.930 3449.090 1644.110 3450.270 ;
        RECT 1642.930 3447.490 1644.110 3448.670 ;
        RECT 1642.930 3269.090 1644.110 3270.270 ;
        RECT 1642.930 3267.490 1644.110 3268.670 ;
        RECT 1642.930 3089.090 1644.110 3090.270 ;
        RECT 1642.930 3087.490 1644.110 3088.670 ;
        RECT 1642.930 2909.090 1644.110 2910.270 ;
        RECT 1642.930 2907.490 1644.110 2908.670 ;
        RECT 1642.930 2729.090 1644.110 2730.270 ;
        RECT 1642.930 2727.490 1644.110 2728.670 ;
        RECT 1642.930 2549.090 1644.110 2550.270 ;
        RECT 1642.930 2547.490 1644.110 2548.670 ;
        RECT 1642.930 2369.090 1644.110 2370.270 ;
        RECT 1642.930 2367.490 1644.110 2368.670 ;
        RECT 1642.930 2189.090 1644.110 2190.270 ;
        RECT 1642.930 2187.490 1644.110 2188.670 ;
        RECT 1642.930 2009.090 1644.110 2010.270 ;
        RECT 1642.930 2007.490 1644.110 2008.670 ;
        RECT 1642.930 1829.090 1644.110 1830.270 ;
        RECT 1642.930 1827.490 1644.110 1828.670 ;
        RECT 1642.930 1649.090 1644.110 1650.270 ;
        RECT 1642.930 1647.490 1644.110 1648.670 ;
        RECT 1642.930 1469.090 1644.110 1470.270 ;
        RECT 1642.930 1467.490 1644.110 1468.670 ;
        RECT 1642.930 1289.090 1644.110 1290.270 ;
        RECT 1642.930 1287.490 1644.110 1288.670 ;
        RECT 1642.930 1109.090 1644.110 1110.270 ;
        RECT 1642.930 1107.490 1644.110 1108.670 ;
        RECT 1642.930 929.090 1644.110 930.270 ;
        RECT 1642.930 927.490 1644.110 928.670 ;
        RECT 1642.930 749.090 1644.110 750.270 ;
        RECT 1642.930 747.490 1644.110 748.670 ;
        RECT 1642.930 569.090 1644.110 570.270 ;
        RECT 1642.930 567.490 1644.110 568.670 ;
        RECT 1642.930 389.090 1644.110 390.270 ;
        RECT 1642.930 387.490 1644.110 388.670 ;
        RECT 1642.930 209.090 1644.110 210.270 ;
        RECT 1642.930 207.490 1644.110 208.670 ;
        RECT 1642.930 29.090 1644.110 30.270 ;
        RECT 1642.930 27.490 1644.110 28.670 ;
        RECT 1642.930 -12.110 1644.110 -10.930 ;
        RECT 1642.930 -13.710 1644.110 -12.530 ;
        RECT 1822.930 3532.210 1824.110 3533.390 ;
        RECT 1822.930 3530.610 1824.110 3531.790 ;
        RECT 1822.930 3449.090 1824.110 3450.270 ;
        RECT 1822.930 3447.490 1824.110 3448.670 ;
        RECT 1822.930 3269.090 1824.110 3270.270 ;
        RECT 1822.930 3267.490 1824.110 3268.670 ;
        RECT 1822.930 3089.090 1824.110 3090.270 ;
        RECT 1822.930 3087.490 1824.110 3088.670 ;
        RECT 1822.930 2909.090 1824.110 2910.270 ;
        RECT 1822.930 2907.490 1824.110 2908.670 ;
        RECT 1822.930 2729.090 1824.110 2730.270 ;
        RECT 1822.930 2727.490 1824.110 2728.670 ;
        RECT 1822.930 2549.090 1824.110 2550.270 ;
        RECT 1822.930 2547.490 1824.110 2548.670 ;
        RECT 1822.930 2369.090 1824.110 2370.270 ;
        RECT 1822.930 2367.490 1824.110 2368.670 ;
        RECT 1822.930 2189.090 1824.110 2190.270 ;
        RECT 1822.930 2187.490 1824.110 2188.670 ;
        RECT 1822.930 2009.090 1824.110 2010.270 ;
        RECT 1822.930 2007.490 1824.110 2008.670 ;
        RECT 1822.930 1829.090 1824.110 1830.270 ;
        RECT 1822.930 1827.490 1824.110 1828.670 ;
        RECT 1822.930 1649.090 1824.110 1650.270 ;
        RECT 1822.930 1647.490 1824.110 1648.670 ;
        RECT 1822.930 1469.090 1824.110 1470.270 ;
        RECT 1822.930 1467.490 1824.110 1468.670 ;
        RECT 1822.930 1289.090 1824.110 1290.270 ;
        RECT 1822.930 1287.490 1824.110 1288.670 ;
        RECT 1822.930 1109.090 1824.110 1110.270 ;
        RECT 1822.930 1107.490 1824.110 1108.670 ;
        RECT 1822.930 929.090 1824.110 930.270 ;
        RECT 1822.930 927.490 1824.110 928.670 ;
        RECT 1822.930 749.090 1824.110 750.270 ;
        RECT 1822.930 747.490 1824.110 748.670 ;
        RECT 1822.930 569.090 1824.110 570.270 ;
        RECT 1822.930 567.490 1824.110 568.670 ;
        RECT 1822.930 389.090 1824.110 390.270 ;
        RECT 1822.930 387.490 1824.110 388.670 ;
        RECT 1822.930 209.090 1824.110 210.270 ;
        RECT 1822.930 207.490 1824.110 208.670 ;
        RECT 1822.930 29.090 1824.110 30.270 ;
        RECT 1822.930 27.490 1824.110 28.670 ;
        RECT 1822.930 -12.110 1824.110 -10.930 ;
        RECT 1822.930 -13.710 1824.110 -12.530 ;
        RECT 2002.930 3532.210 2004.110 3533.390 ;
        RECT 2002.930 3530.610 2004.110 3531.790 ;
        RECT 2002.930 3449.090 2004.110 3450.270 ;
        RECT 2002.930 3447.490 2004.110 3448.670 ;
        RECT 2002.930 3269.090 2004.110 3270.270 ;
        RECT 2002.930 3267.490 2004.110 3268.670 ;
        RECT 2002.930 3089.090 2004.110 3090.270 ;
        RECT 2002.930 3087.490 2004.110 3088.670 ;
        RECT 2002.930 2909.090 2004.110 2910.270 ;
        RECT 2002.930 2907.490 2004.110 2908.670 ;
        RECT 2002.930 2729.090 2004.110 2730.270 ;
        RECT 2002.930 2727.490 2004.110 2728.670 ;
        RECT 2002.930 2549.090 2004.110 2550.270 ;
        RECT 2002.930 2547.490 2004.110 2548.670 ;
        RECT 2002.930 2369.090 2004.110 2370.270 ;
        RECT 2002.930 2367.490 2004.110 2368.670 ;
        RECT 2002.930 2189.090 2004.110 2190.270 ;
        RECT 2002.930 2187.490 2004.110 2188.670 ;
        RECT 2002.930 2009.090 2004.110 2010.270 ;
        RECT 2002.930 2007.490 2004.110 2008.670 ;
        RECT 2002.930 1829.090 2004.110 1830.270 ;
        RECT 2002.930 1827.490 2004.110 1828.670 ;
        RECT 2002.930 1649.090 2004.110 1650.270 ;
        RECT 2002.930 1647.490 2004.110 1648.670 ;
        RECT 2002.930 1469.090 2004.110 1470.270 ;
        RECT 2002.930 1467.490 2004.110 1468.670 ;
        RECT 2002.930 1289.090 2004.110 1290.270 ;
        RECT 2002.930 1287.490 2004.110 1288.670 ;
        RECT 2002.930 1109.090 2004.110 1110.270 ;
        RECT 2002.930 1107.490 2004.110 1108.670 ;
        RECT 2002.930 929.090 2004.110 930.270 ;
        RECT 2002.930 927.490 2004.110 928.670 ;
        RECT 2002.930 749.090 2004.110 750.270 ;
        RECT 2002.930 747.490 2004.110 748.670 ;
        RECT 2002.930 569.090 2004.110 570.270 ;
        RECT 2002.930 567.490 2004.110 568.670 ;
        RECT 2002.930 389.090 2004.110 390.270 ;
        RECT 2002.930 387.490 2004.110 388.670 ;
        RECT 2002.930 209.090 2004.110 210.270 ;
        RECT 2002.930 207.490 2004.110 208.670 ;
        RECT 2002.930 29.090 2004.110 30.270 ;
        RECT 2002.930 27.490 2004.110 28.670 ;
        RECT 2002.930 -12.110 2004.110 -10.930 ;
        RECT 2002.930 -13.710 2004.110 -12.530 ;
        RECT 2182.930 3532.210 2184.110 3533.390 ;
        RECT 2182.930 3530.610 2184.110 3531.790 ;
        RECT 2182.930 3449.090 2184.110 3450.270 ;
        RECT 2182.930 3447.490 2184.110 3448.670 ;
        RECT 2182.930 3269.090 2184.110 3270.270 ;
        RECT 2182.930 3267.490 2184.110 3268.670 ;
        RECT 2182.930 3089.090 2184.110 3090.270 ;
        RECT 2182.930 3087.490 2184.110 3088.670 ;
        RECT 2182.930 2909.090 2184.110 2910.270 ;
        RECT 2182.930 2907.490 2184.110 2908.670 ;
        RECT 2182.930 2729.090 2184.110 2730.270 ;
        RECT 2182.930 2727.490 2184.110 2728.670 ;
        RECT 2182.930 2549.090 2184.110 2550.270 ;
        RECT 2182.930 2547.490 2184.110 2548.670 ;
        RECT 2182.930 2369.090 2184.110 2370.270 ;
        RECT 2182.930 2367.490 2184.110 2368.670 ;
        RECT 2182.930 2189.090 2184.110 2190.270 ;
        RECT 2182.930 2187.490 2184.110 2188.670 ;
        RECT 2182.930 2009.090 2184.110 2010.270 ;
        RECT 2182.930 2007.490 2184.110 2008.670 ;
        RECT 2182.930 1829.090 2184.110 1830.270 ;
        RECT 2182.930 1827.490 2184.110 1828.670 ;
        RECT 2182.930 1649.090 2184.110 1650.270 ;
        RECT 2182.930 1647.490 2184.110 1648.670 ;
        RECT 2182.930 1469.090 2184.110 1470.270 ;
        RECT 2182.930 1467.490 2184.110 1468.670 ;
        RECT 2182.930 1289.090 2184.110 1290.270 ;
        RECT 2182.930 1287.490 2184.110 1288.670 ;
        RECT 2182.930 1109.090 2184.110 1110.270 ;
        RECT 2182.930 1107.490 2184.110 1108.670 ;
        RECT 2182.930 929.090 2184.110 930.270 ;
        RECT 2182.930 927.490 2184.110 928.670 ;
        RECT 2182.930 749.090 2184.110 750.270 ;
        RECT 2182.930 747.490 2184.110 748.670 ;
        RECT 2182.930 569.090 2184.110 570.270 ;
        RECT 2182.930 567.490 2184.110 568.670 ;
        RECT 2182.930 389.090 2184.110 390.270 ;
        RECT 2182.930 387.490 2184.110 388.670 ;
        RECT 2182.930 209.090 2184.110 210.270 ;
        RECT 2182.930 207.490 2184.110 208.670 ;
        RECT 2182.930 29.090 2184.110 30.270 ;
        RECT 2182.930 27.490 2184.110 28.670 ;
        RECT 2182.930 -12.110 2184.110 -10.930 ;
        RECT 2182.930 -13.710 2184.110 -12.530 ;
        RECT 2362.930 3532.210 2364.110 3533.390 ;
        RECT 2362.930 3530.610 2364.110 3531.790 ;
        RECT 2362.930 3449.090 2364.110 3450.270 ;
        RECT 2362.930 3447.490 2364.110 3448.670 ;
        RECT 2362.930 3269.090 2364.110 3270.270 ;
        RECT 2362.930 3267.490 2364.110 3268.670 ;
        RECT 2362.930 3089.090 2364.110 3090.270 ;
        RECT 2362.930 3087.490 2364.110 3088.670 ;
        RECT 2362.930 2909.090 2364.110 2910.270 ;
        RECT 2362.930 2907.490 2364.110 2908.670 ;
        RECT 2362.930 2729.090 2364.110 2730.270 ;
        RECT 2362.930 2727.490 2364.110 2728.670 ;
        RECT 2362.930 2549.090 2364.110 2550.270 ;
        RECT 2362.930 2547.490 2364.110 2548.670 ;
        RECT 2362.930 2369.090 2364.110 2370.270 ;
        RECT 2362.930 2367.490 2364.110 2368.670 ;
        RECT 2362.930 2189.090 2364.110 2190.270 ;
        RECT 2362.930 2187.490 2364.110 2188.670 ;
        RECT 2362.930 2009.090 2364.110 2010.270 ;
        RECT 2362.930 2007.490 2364.110 2008.670 ;
        RECT 2362.930 1829.090 2364.110 1830.270 ;
        RECT 2362.930 1827.490 2364.110 1828.670 ;
        RECT 2362.930 1649.090 2364.110 1650.270 ;
        RECT 2362.930 1647.490 2364.110 1648.670 ;
        RECT 2362.930 1469.090 2364.110 1470.270 ;
        RECT 2362.930 1467.490 2364.110 1468.670 ;
        RECT 2362.930 1289.090 2364.110 1290.270 ;
        RECT 2362.930 1287.490 2364.110 1288.670 ;
        RECT 2362.930 1109.090 2364.110 1110.270 ;
        RECT 2362.930 1107.490 2364.110 1108.670 ;
        RECT 2362.930 929.090 2364.110 930.270 ;
        RECT 2362.930 927.490 2364.110 928.670 ;
        RECT 2362.930 749.090 2364.110 750.270 ;
        RECT 2362.930 747.490 2364.110 748.670 ;
        RECT 2362.930 569.090 2364.110 570.270 ;
        RECT 2362.930 567.490 2364.110 568.670 ;
        RECT 2362.930 389.090 2364.110 390.270 ;
        RECT 2362.930 387.490 2364.110 388.670 ;
        RECT 2362.930 209.090 2364.110 210.270 ;
        RECT 2362.930 207.490 2364.110 208.670 ;
        RECT 2362.930 29.090 2364.110 30.270 ;
        RECT 2362.930 27.490 2364.110 28.670 ;
        RECT 2362.930 -12.110 2364.110 -10.930 ;
        RECT 2362.930 -13.710 2364.110 -12.530 ;
        RECT 2542.930 3532.210 2544.110 3533.390 ;
        RECT 2542.930 3530.610 2544.110 3531.790 ;
        RECT 2542.930 3449.090 2544.110 3450.270 ;
        RECT 2542.930 3447.490 2544.110 3448.670 ;
        RECT 2542.930 3269.090 2544.110 3270.270 ;
        RECT 2542.930 3267.490 2544.110 3268.670 ;
        RECT 2542.930 3089.090 2544.110 3090.270 ;
        RECT 2542.930 3087.490 2544.110 3088.670 ;
        RECT 2542.930 2909.090 2544.110 2910.270 ;
        RECT 2542.930 2907.490 2544.110 2908.670 ;
        RECT 2542.930 2729.090 2544.110 2730.270 ;
        RECT 2542.930 2727.490 2544.110 2728.670 ;
        RECT 2542.930 2549.090 2544.110 2550.270 ;
        RECT 2542.930 2547.490 2544.110 2548.670 ;
        RECT 2542.930 2369.090 2544.110 2370.270 ;
        RECT 2542.930 2367.490 2544.110 2368.670 ;
        RECT 2542.930 2189.090 2544.110 2190.270 ;
        RECT 2542.930 2187.490 2544.110 2188.670 ;
        RECT 2542.930 2009.090 2544.110 2010.270 ;
        RECT 2542.930 2007.490 2544.110 2008.670 ;
        RECT 2542.930 1829.090 2544.110 1830.270 ;
        RECT 2542.930 1827.490 2544.110 1828.670 ;
        RECT 2542.930 1649.090 2544.110 1650.270 ;
        RECT 2542.930 1647.490 2544.110 1648.670 ;
        RECT 2542.930 1469.090 2544.110 1470.270 ;
        RECT 2542.930 1467.490 2544.110 1468.670 ;
        RECT 2542.930 1289.090 2544.110 1290.270 ;
        RECT 2542.930 1287.490 2544.110 1288.670 ;
        RECT 2542.930 1109.090 2544.110 1110.270 ;
        RECT 2542.930 1107.490 2544.110 1108.670 ;
        RECT 2542.930 929.090 2544.110 930.270 ;
        RECT 2542.930 927.490 2544.110 928.670 ;
        RECT 2542.930 749.090 2544.110 750.270 ;
        RECT 2542.930 747.490 2544.110 748.670 ;
        RECT 2542.930 569.090 2544.110 570.270 ;
        RECT 2542.930 567.490 2544.110 568.670 ;
        RECT 2542.930 389.090 2544.110 390.270 ;
        RECT 2542.930 387.490 2544.110 388.670 ;
        RECT 2542.930 209.090 2544.110 210.270 ;
        RECT 2542.930 207.490 2544.110 208.670 ;
        RECT 2542.930 29.090 2544.110 30.270 ;
        RECT 2542.930 27.490 2544.110 28.670 ;
        RECT 2542.930 -12.110 2544.110 -10.930 ;
        RECT 2542.930 -13.710 2544.110 -12.530 ;
        RECT 2722.930 3532.210 2724.110 3533.390 ;
        RECT 2722.930 3530.610 2724.110 3531.790 ;
        RECT 2722.930 3449.090 2724.110 3450.270 ;
        RECT 2722.930 3447.490 2724.110 3448.670 ;
        RECT 2722.930 3269.090 2724.110 3270.270 ;
        RECT 2722.930 3267.490 2724.110 3268.670 ;
        RECT 2722.930 3089.090 2724.110 3090.270 ;
        RECT 2722.930 3087.490 2724.110 3088.670 ;
        RECT 2722.930 2909.090 2724.110 2910.270 ;
        RECT 2722.930 2907.490 2724.110 2908.670 ;
        RECT 2722.930 2729.090 2724.110 2730.270 ;
        RECT 2722.930 2727.490 2724.110 2728.670 ;
        RECT 2722.930 2549.090 2724.110 2550.270 ;
        RECT 2722.930 2547.490 2724.110 2548.670 ;
        RECT 2722.930 2369.090 2724.110 2370.270 ;
        RECT 2722.930 2367.490 2724.110 2368.670 ;
        RECT 2722.930 2189.090 2724.110 2190.270 ;
        RECT 2722.930 2187.490 2724.110 2188.670 ;
        RECT 2722.930 2009.090 2724.110 2010.270 ;
        RECT 2722.930 2007.490 2724.110 2008.670 ;
        RECT 2722.930 1829.090 2724.110 1830.270 ;
        RECT 2722.930 1827.490 2724.110 1828.670 ;
        RECT 2722.930 1649.090 2724.110 1650.270 ;
        RECT 2722.930 1647.490 2724.110 1648.670 ;
        RECT 2722.930 1469.090 2724.110 1470.270 ;
        RECT 2722.930 1467.490 2724.110 1468.670 ;
        RECT 2722.930 1289.090 2724.110 1290.270 ;
        RECT 2722.930 1287.490 2724.110 1288.670 ;
        RECT 2722.930 1109.090 2724.110 1110.270 ;
        RECT 2722.930 1107.490 2724.110 1108.670 ;
        RECT 2722.930 929.090 2724.110 930.270 ;
        RECT 2722.930 927.490 2724.110 928.670 ;
        RECT 2722.930 749.090 2724.110 750.270 ;
        RECT 2722.930 747.490 2724.110 748.670 ;
        RECT 2722.930 569.090 2724.110 570.270 ;
        RECT 2722.930 567.490 2724.110 568.670 ;
        RECT 2722.930 389.090 2724.110 390.270 ;
        RECT 2722.930 387.490 2724.110 388.670 ;
        RECT 2722.930 209.090 2724.110 210.270 ;
        RECT 2722.930 207.490 2724.110 208.670 ;
        RECT 2722.930 29.090 2724.110 30.270 ;
        RECT 2722.930 27.490 2724.110 28.670 ;
        RECT 2722.930 -12.110 2724.110 -10.930 ;
        RECT 2722.930 -13.710 2724.110 -12.530 ;
        RECT 2902.930 3532.210 2904.110 3533.390 ;
        RECT 2902.930 3530.610 2904.110 3531.790 ;
        RECT 2902.930 3449.090 2904.110 3450.270 ;
        RECT 2902.930 3447.490 2904.110 3448.670 ;
        RECT 2902.930 3269.090 2904.110 3270.270 ;
        RECT 2902.930 3267.490 2904.110 3268.670 ;
        RECT 2902.930 3089.090 2904.110 3090.270 ;
        RECT 2902.930 3087.490 2904.110 3088.670 ;
        RECT 2902.930 2909.090 2904.110 2910.270 ;
        RECT 2902.930 2907.490 2904.110 2908.670 ;
        RECT 2902.930 2729.090 2904.110 2730.270 ;
        RECT 2902.930 2727.490 2904.110 2728.670 ;
        RECT 2902.930 2549.090 2904.110 2550.270 ;
        RECT 2902.930 2547.490 2904.110 2548.670 ;
        RECT 2902.930 2369.090 2904.110 2370.270 ;
        RECT 2902.930 2367.490 2904.110 2368.670 ;
        RECT 2902.930 2189.090 2904.110 2190.270 ;
        RECT 2902.930 2187.490 2904.110 2188.670 ;
        RECT 2902.930 2009.090 2904.110 2010.270 ;
        RECT 2902.930 2007.490 2904.110 2008.670 ;
        RECT 2902.930 1829.090 2904.110 1830.270 ;
        RECT 2902.930 1827.490 2904.110 1828.670 ;
        RECT 2902.930 1649.090 2904.110 1650.270 ;
        RECT 2902.930 1647.490 2904.110 1648.670 ;
        RECT 2902.930 1469.090 2904.110 1470.270 ;
        RECT 2902.930 1467.490 2904.110 1468.670 ;
        RECT 2902.930 1289.090 2904.110 1290.270 ;
        RECT 2902.930 1287.490 2904.110 1288.670 ;
        RECT 2902.930 1109.090 2904.110 1110.270 ;
        RECT 2902.930 1107.490 2904.110 1108.670 ;
        RECT 2902.930 929.090 2904.110 930.270 ;
        RECT 2902.930 927.490 2904.110 928.670 ;
        RECT 2902.930 749.090 2904.110 750.270 ;
        RECT 2902.930 747.490 2904.110 748.670 ;
        RECT 2902.930 569.090 2904.110 570.270 ;
        RECT 2902.930 567.490 2904.110 568.670 ;
        RECT 2902.930 389.090 2904.110 390.270 ;
        RECT 2902.930 387.490 2904.110 388.670 ;
        RECT 2902.930 209.090 2904.110 210.270 ;
        RECT 2902.930 207.490 2904.110 208.670 ;
        RECT 2902.930 29.090 2904.110 30.270 ;
        RECT 2902.930 27.490 2904.110 28.670 ;
        RECT 2902.930 -12.110 2904.110 -10.930 ;
        RECT 2902.930 -13.710 2904.110 -12.530 ;
        RECT 2936.710 3532.210 2937.890 3533.390 ;
        RECT 2936.710 3530.610 2937.890 3531.790 ;
        RECT 2936.710 3449.090 2937.890 3450.270 ;
        RECT 2936.710 3447.490 2937.890 3448.670 ;
        RECT 2936.710 3269.090 2937.890 3270.270 ;
        RECT 2936.710 3267.490 2937.890 3268.670 ;
        RECT 2936.710 3089.090 2937.890 3090.270 ;
        RECT 2936.710 3087.490 2937.890 3088.670 ;
        RECT 2936.710 2909.090 2937.890 2910.270 ;
        RECT 2936.710 2907.490 2937.890 2908.670 ;
        RECT 2936.710 2729.090 2937.890 2730.270 ;
        RECT 2936.710 2727.490 2937.890 2728.670 ;
        RECT 2936.710 2549.090 2937.890 2550.270 ;
        RECT 2936.710 2547.490 2937.890 2548.670 ;
        RECT 2936.710 2369.090 2937.890 2370.270 ;
        RECT 2936.710 2367.490 2937.890 2368.670 ;
        RECT 2936.710 2189.090 2937.890 2190.270 ;
        RECT 2936.710 2187.490 2937.890 2188.670 ;
        RECT 2936.710 2009.090 2937.890 2010.270 ;
        RECT 2936.710 2007.490 2937.890 2008.670 ;
        RECT 2936.710 1829.090 2937.890 1830.270 ;
        RECT 2936.710 1827.490 2937.890 1828.670 ;
        RECT 2936.710 1649.090 2937.890 1650.270 ;
        RECT 2936.710 1647.490 2937.890 1648.670 ;
        RECT 2936.710 1469.090 2937.890 1470.270 ;
        RECT 2936.710 1467.490 2937.890 1468.670 ;
        RECT 2936.710 1289.090 2937.890 1290.270 ;
        RECT 2936.710 1287.490 2937.890 1288.670 ;
        RECT 2936.710 1109.090 2937.890 1110.270 ;
        RECT 2936.710 1107.490 2937.890 1108.670 ;
        RECT 2936.710 929.090 2937.890 930.270 ;
        RECT 2936.710 927.490 2937.890 928.670 ;
        RECT 2936.710 749.090 2937.890 750.270 ;
        RECT 2936.710 747.490 2937.890 748.670 ;
        RECT 2936.710 569.090 2937.890 570.270 ;
        RECT 2936.710 567.490 2937.890 568.670 ;
        RECT 2936.710 389.090 2937.890 390.270 ;
        RECT 2936.710 387.490 2937.890 388.670 ;
        RECT 2936.710 209.090 2937.890 210.270 ;
        RECT 2936.710 207.490 2937.890 208.670 ;
        RECT 2936.710 29.090 2937.890 30.270 ;
        RECT 2936.710 27.490 2937.890 28.670 ;
        RECT 2936.710 -12.110 2937.890 -10.930 ;
        RECT 2936.710 -13.710 2937.890 -12.530 ;
      LAYER met5 ;
        RECT -19.180 3533.500 -16.180 3533.510 ;
        RECT 22.020 3533.500 25.020 3533.510 ;
        RECT 202.020 3533.500 205.020 3533.510 ;
        RECT 382.020 3533.500 385.020 3533.510 ;
        RECT 562.020 3533.500 565.020 3533.510 ;
        RECT 742.020 3533.500 745.020 3533.510 ;
        RECT 922.020 3533.500 925.020 3533.510 ;
        RECT 1102.020 3533.500 1105.020 3533.510 ;
        RECT 1282.020 3533.500 1285.020 3533.510 ;
        RECT 1462.020 3533.500 1465.020 3533.510 ;
        RECT 1642.020 3533.500 1645.020 3533.510 ;
        RECT 1822.020 3533.500 1825.020 3533.510 ;
        RECT 2002.020 3533.500 2005.020 3533.510 ;
        RECT 2182.020 3533.500 2185.020 3533.510 ;
        RECT 2362.020 3533.500 2365.020 3533.510 ;
        RECT 2542.020 3533.500 2545.020 3533.510 ;
        RECT 2722.020 3533.500 2725.020 3533.510 ;
        RECT 2902.020 3533.500 2905.020 3533.510 ;
        RECT 2935.800 3533.500 2938.800 3533.510 ;
        RECT -19.180 3530.500 2938.800 3533.500 ;
        RECT -19.180 3530.490 -16.180 3530.500 ;
        RECT 22.020 3530.490 25.020 3530.500 ;
        RECT 202.020 3530.490 205.020 3530.500 ;
        RECT 382.020 3530.490 385.020 3530.500 ;
        RECT 562.020 3530.490 565.020 3530.500 ;
        RECT 742.020 3530.490 745.020 3530.500 ;
        RECT 922.020 3530.490 925.020 3530.500 ;
        RECT 1102.020 3530.490 1105.020 3530.500 ;
        RECT 1282.020 3530.490 1285.020 3530.500 ;
        RECT 1462.020 3530.490 1465.020 3530.500 ;
        RECT 1642.020 3530.490 1645.020 3530.500 ;
        RECT 1822.020 3530.490 1825.020 3530.500 ;
        RECT 2002.020 3530.490 2005.020 3530.500 ;
        RECT 2182.020 3530.490 2185.020 3530.500 ;
        RECT 2362.020 3530.490 2365.020 3530.500 ;
        RECT 2542.020 3530.490 2545.020 3530.500 ;
        RECT 2722.020 3530.490 2725.020 3530.500 ;
        RECT 2902.020 3530.490 2905.020 3530.500 ;
        RECT 2935.800 3530.490 2938.800 3530.500 ;
        RECT -19.180 3450.380 -16.180 3450.390 ;
        RECT 22.020 3450.380 25.020 3450.390 ;
        RECT 202.020 3450.380 205.020 3450.390 ;
        RECT 382.020 3450.380 385.020 3450.390 ;
        RECT 562.020 3450.380 565.020 3450.390 ;
        RECT 742.020 3450.380 745.020 3450.390 ;
        RECT 922.020 3450.380 925.020 3450.390 ;
        RECT 1102.020 3450.380 1105.020 3450.390 ;
        RECT 1282.020 3450.380 1285.020 3450.390 ;
        RECT 1462.020 3450.380 1465.020 3450.390 ;
        RECT 1642.020 3450.380 1645.020 3450.390 ;
        RECT 1822.020 3450.380 1825.020 3450.390 ;
        RECT 2002.020 3450.380 2005.020 3450.390 ;
        RECT 2182.020 3450.380 2185.020 3450.390 ;
        RECT 2362.020 3450.380 2365.020 3450.390 ;
        RECT 2542.020 3450.380 2545.020 3450.390 ;
        RECT 2722.020 3450.380 2725.020 3450.390 ;
        RECT 2902.020 3450.380 2905.020 3450.390 ;
        RECT 2935.800 3450.380 2938.800 3450.390 ;
        RECT -23.780 3447.380 2943.400 3450.380 ;
        RECT -19.180 3447.370 -16.180 3447.380 ;
        RECT 22.020 3447.370 25.020 3447.380 ;
        RECT 202.020 3447.370 205.020 3447.380 ;
        RECT 382.020 3447.370 385.020 3447.380 ;
        RECT 562.020 3447.370 565.020 3447.380 ;
        RECT 742.020 3447.370 745.020 3447.380 ;
        RECT 922.020 3447.370 925.020 3447.380 ;
        RECT 1102.020 3447.370 1105.020 3447.380 ;
        RECT 1282.020 3447.370 1285.020 3447.380 ;
        RECT 1462.020 3447.370 1465.020 3447.380 ;
        RECT 1642.020 3447.370 1645.020 3447.380 ;
        RECT 1822.020 3447.370 1825.020 3447.380 ;
        RECT 2002.020 3447.370 2005.020 3447.380 ;
        RECT 2182.020 3447.370 2185.020 3447.380 ;
        RECT 2362.020 3447.370 2365.020 3447.380 ;
        RECT 2542.020 3447.370 2545.020 3447.380 ;
        RECT 2722.020 3447.370 2725.020 3447.380 ;
        RECT 2902.020 3447.370 2905.020 3447.380 ;
        RECT 2935.800 3447.370 2938.800 3447.380 ;
        RECT -19.180 3270.380 -16.180 3270.390 ;
        RECT 22.020 3270.380 25.020 3270.390 ;
        RECT 202.020 3270.380 205.020 3270.390 ;
        RECT 382.020 3270.380 385.020 3270.390 ;
        RECT 562.020 3270.380 565.020 3270.390 ;
        RECT 742.020 3270.380 745.020 3270.390 ;
        RECT 922.020 3270.380 925.020 3270.390 ;
        RECT 1102.020 3270.380 1105.020 3270.390 ;
        RECT 1282.020 3270.380 1285.020 3270.390 ;
        RECT 1462.020 3270.380 1465.020 3270.390 ;
        RECT 1642.020 3270.380 1645.020 3270.390 ;
        RECT 1822.020 3270.380 1825.020 3270.390 ;
        RECT 2002.020 3270.380 2005.020 3270.390 ;
        RECT 2182.020 3270.380 2185.020 3270.390 ;
        RECT 2362.020 3270.380 2365.020 3270.390 ;
        RECT 2542.020 3270.380 2545.020 3270.390 ;
        RECT 2722.020 3270.380 2725.020 3270.390 ;
        RECT 2902.020 3270.380 2905.020 3270.390 ;
        RECT 2935.800 3270.380 2938.800 3270.390 ;
        RECT -23.780 3267.380 2943.400 3270.380 ;
        RECT -19.180 3267.370 -16.180 3267.380 ;
        RECT 22.020 3267.370 25.020 3267.380 ;
        RECT 202.020 3267.370 205.020 3267.380 ;
        RECT 382.020 3267.370 385.020 3267.380 ;
        RECT 562.020 3267.370 565.020 3267.380 ;
        RECT 742.020 3267.370 745.020 3267.380 ;
        RECT 922.020 3267.370 925.020 3267.380 ;
        RECT 1102.020 3267.370 1105.020 3267.380 ;
        RECT 1282.020 3267.370 1285.020 3267.380 ;
        RECT 1462.020 3267.370 1465.020 3267.380 ;
        RECT 1642.020 3267.370 1645.020 3267.380 ;
        RECT 1822.020 3267.370 1825.020 3267.380 ;
        RECT 2002.020 3267.370 2005.020 3267.380 ;
        RECT 2182.020 3267.370 2185.020 3267.380 ;
        RECT 2362.020 3267.370 2365.020 3267.380 ;
        RECT 2542.020 3267.370 2545.020 3267.380 ;
        RECT 2722.020 3267.370 2725.020 3267.380 ;
        RECT 2902.020 3267.370 2905.020 3267.380 ;
        RECT 2935.800 3267.370 2938.800 3267.380 ;
        RECT -19.180 3090.380 -16.180 3090.390 ;
        RECT 22.020 3090.380 25.020 3090.390 ;
        RECT 202.020 3090.380 205.020 3090.390 ;
        RECT 382.020 3090.380 385.020 3090.390 ;
        RECT 562.020 3090.380 565.020 3090.390 ;
        RECT 742.020 3090.380 745.020 3090.390 ;
        RECT 922.020 3090.380 925.020 3090.390 ;
        RECT 1102.020 3090.380 1105.020 3090.390 ;
        RECT 1282.020 3090.380 1285.020 3090.390 ;
        RECT 1462.020 3090.380 1465.020 3090.390 ;
        RECT 1642.020 3090.380 1645.020 3090.390 ;
        RECT 1822.020 3090.380 1825.020 3090.390 ;
        RECT 2002.020 3090.380 2005.020 3090.390 ;
        RECT 2182.020 3090.380 2185.020 3090.390 ;
        RECT 2362.020 3090.380 2365.020 3090.390 ;
        RECT 2542.020 3090.380 2545.020 3090.390 ;
        RECT 2722.020 3090.380 2725.020 3090.390 ;
        RECT 2902.020 3090.380 2905.020 3090.390 ;
        RECT 2935.800 3090.380 2938.800 3090.390 ;
        RECT -23.780 3087.380 2943.400 3090.380 ;
        RECT -19.180 3087.370 -16.180 3087.380 ;
        RECT 22.020 3087.370 25.020 3087.380 ;
        RECT 202.020 3087.370 205.020 3087.380 ;
        RECT 382.020 3087.370 385.020 3087.380 ;
        RECT 562.020 3087.370 565.020 3087.380 ;
        RECT 742.020 3087.370 745.020 3087.380 ;
        RECT 922.020 3087.370 925.020 3087.380 ;
        RECT 1102.020 3087.370 1105.020 3087.380 ;
        RECT 1282.020 3087.370 1285.020 3087.380 ;
        RECT 1462.020 3087.370 1465.020 3087.380 ;
        RECT 1642.020 3087.370 1645.020 3087.380 ;
        RECT 1822.020 3087.370 1825.020 3087.380 ;
        RECT 2002.020 3087.370 2005.020 3087.380 ;
        RECT 2182.020 3087.370 2185.020 3087.380 ;
        RECT 2362.020 3087.370 2365.020 3087.380 ;
        RECT 2542.020 3087.370 2545.020 3087.380 ;
        RECT 2722.020 3087.370 2725.020 3087.380 ;
        RECT 2902.020 3087.370 2905.020 3087.380 ;
        RECT 2935.800 3087.370 2938.800 3087.380 ;
        RECT -19.180 2910.380 -16.180 2910.390 ;
        RECT 22.020 2910.380 25.020 2910.390 ;
        RECT 202.020 2910.380 205.020 2910.390 ;
        RECT 382.020 2910.380 385.020 2910.390 ;
        RECT 562.020 2910.380 565.020 2910.390 ;
        RECT 742.020 2910.380 745.020 2910.390 ;
        RECT 922.020 2910.380 925.020 2910.390 ;
        RECT 1102.020 2910.380 1105.020 2910.390 ;
        RECT 1282.020 2910.380 1285.020 2910.390 ;
        RECT 1462.020 2910.380 1465.020 2910.390 ;
        RECT 1642.020 2910.380 1645.020 2910.390 ;
        RECT 1822.020 2910.380 1825.020 2910.390 ;
        RECT 2002.020 2910.380 2005.020 2910.390 ;
        RECT 2182.020 2910.380 2185.020 2910.390 ;
        RECT 2362.020 2910.380 2365.020 2910.390 ;
        RECT 2542.020 2910.380 2545.020 2910.390 ;
        RECT 2722.020 2910.380 2725.020 2910.390 ;
        RECT 2902.020 2910.380 2905.020 2910.390 ;
        RECT 2935.800 2910.380 2938.800 2910.390 ;
        RECT -23.780 2907.380 2943.400 2910.380 ;
        RECT -19.180 2907.370 -16.180 2907.380 ;
        RECT 22.020 2907.370 25.020 2907.380 ;
        RECT 202.020 2907.370 205.020 2907.380 ;
        RECT 382.020 2907.370 385.020 2907.380 ;
        RECT 562.020 2907.370 565.020 2907.380 ;
        RECT 742.020 2907.370 745.020 2907.380 ;
        RECT 922.020 2907.370 925.020 2907.380 ;
        RECT 1102.020 2907.370 1105.020 2907.380 ;
        RECT 1282.020 2907.370 1285.020 2907.380 ;
        RECT 1462.020 2907.370 1465.020 2907.380 ;
        RECT 1642.020 2907.370 1645.020 2907.380 ;
        RECT 1822.020 2907.370 1825.020 2907.380 ;
        RECT 2002.020 2907.370 2005.020 2907.380 ;
        RECT 2182.020 2907.370 2185.020 2907.380 ;
        RECT 2362.020 2907.370 2365.020 2907.380 ;
        RECT 2542.020 2907.370 2545.020 2907.380 ;
        RECT 2722.020 2907.370 2725.020 2907.380 ;
        RECT 2902.020 2907.370 2905.020 2907.380 ;
        RECT 2935.800 2907.370 2938.800 2907.380 ;
        RECT -19.180 2730.380 -16.180 2730.390 ;
        RECT 22.020 2730.380 25.020 2730.390 ;
        RECT 202.020 2730.380 205.020 2730.390 ;
        RECT 382.020 2730.380 385.020 2730.390 ;
        RECT 562.020 2730.380 565.020 2730.390 ;
        RECT 742.020 2730.380 745.020 2730.390 ;
        RECT 922.020 2730.380 925.020 2730.390 ;
        RECT 1102.020 2730.380 1105.020 2730.390 ;
        RECT 1282.020 2730.380 1285.020 2730.390 ;
        RECT 1462.020 2730.380 1465.020 2730.390 ;
        RECT 1642.020 2730.380 1645.020 2730.390 ;
        RECT 1822.020 2730.380 1825.020 2730.390 ;
        RECT 2002.020 2730.380 2005.020 2730.390 ;
        RECT 2182.020 2730.380 2185.020 2730.390 ;
        RECT 2362.020 2730.380 2365.020 2730.390 ;
        RECT 2542.020 2730.380 2545.020 2730.390 ;
        RECT 2722.020 2730.380 2725.020 2730.390 ;
        RECT 2902.020 2730.380 2905.020 2730.390 ;
        RECT 2935.800 2730.380 2938.800 2730.390 ;
        RECT -23.780 2727.380 2943.400 2730.380 ;
        RECT -19.180 2727.370 -16.180 2727.380 ;
        RECT 22.020 2727.370 25.020 2727.380 ;
        RECT 202.020 2727.370 205.020 2727.380 ;
        RECT 382.020 2727.370 385.020 2727.380 ;
        RECT 562.020 2727.370 565.020 2727.380 ;
        RECT 742.020 2727.370 745.020 2727.380 ;
        RECT 922.020 2727.370 925.020 2727.380 ;
        RECT 1102.020 2727.370 1105.020 2727.380 ;
        RECT 1282.020 2727.370 1285.020 2727.380 ;
        RECT 1462.020 2727.370 1465.020 2727.380 ;
        RECT 1642.020 2727.370 1645.020 2727.380 ;
        RECT 1822.020 2727.370 1825.020 2727.380 ;
        RECT 2002.020 2727.370 2005.020 2727.380 ;
        RECT 2182.020 2727.370 2185.020 2727.380 ;
        RECT 2362.020 2727.370 2365.020 2727.380 ;
        RECT 2542.020 2727.370 2545.020 2727.380 ;
        RECT 2722.020 2727.370 2725.020 2727.380 ;
        RECT 2902.020 2727.370 2905.020 2727.380 ;
        RECT 2935.800 2727.370 2938.800 2727.380 ;
        RECT -19.180 2550.380 -16.180 2550.390 ;
        RECT 22.020 2550.380 25.020 2550.390 ;
        RECT 202.020 2550.380 205.020 2550.390 ;
        RECT 382.020 2550.380 385.020 2550.390 ;
        RECT 562.020 2550.380 565.020 2550.390 ;
        RECT 742.020 2550.380 745.020 2550.390 ;
        RECT 922.020 2550.380 925.020 2550.390 ;
        RECT 1102.020 2550.380 1105.020 2550.390 ;
        RECT 1282.020 2550.380 1285.020 2550.390 ;
        RECT 1462.020 2550.380 1465.020 2550.390 ;
        RECT 1642.020 2550.380 1645.020 2550.390 ;
        RECT 1822.020 2550.380 1825.020 2550.390 ;
        RECT 2002.020 2550.380 2005.020 2550.390 ;
        RECT 2182.020 2550.380 2185.020 2550.390 ;
        RECT 2362.020 2550.380 2365.020 2550.390 ;
        RECT 2542.020 2550.380 2545.020 2550.390 ;
        RECT 2722.020 2550.380 2725.020 2550.390 ;
        RECT 2902.020 2550.380 2905.020 2550.390 ;
        RECT 2935.800 2550.380 2938.800 2550.390 ;
        RECT -23.780 2547.380 2943.400 2550.380 ;
        RECT -19.180 2547.370 -16.180 2547.380 ;
        RECT 22.020 2547.370 25.020 2547.380 ;
        RECT 202.020 2547.370 205.020 2547.380 ;
        RECT 382.020 2547.370 385.020 2547.380 ;
        RECT 562.020 2547.370 565.020 2547.380 ;
        RECT 742.020 2547.370 745.020 2547.380 ;
        RECT 922.020 2547.370 925.020 2547.380 ;
        RECT 1102.020 2547.370 1105.020 2547.380 ;
        RECT 1282.020 2547.370 1285.020 2547.380 ;
        RECT 1462.020 2547.370 1465.020 2547.380 ;
        RECT 1642.020 2547.370 1645.020 2547.380 ;
        RECT 1822.020 2547.370 1825.020 2547.380 ;
        RECT 2002.020 2547.370 2005.020 2547.380 ;
        RECT 2182.020 2547.370 2185.020 2547.380 ;
        RECT 2362.020 2547.370 2365.020 2547.380 ;
        RECT 2542.020 2547.370 2545.020 2547.380 ;
        RECT 2722.020 2547.370 2725.020 2547.380 ;
        RECT 2902.020 2547.370 2905.020 2547.380 ;
        RECT 2935.800 2547.370 2938.800 2547.380 ;
        RECT -19.180 2370.380 -16.180 2370.390 ;
        RECT 22.020 2370.380 25.020 2370.390 ;
        RECT 202.020 2370.380 205.020 2370.390 ;
        RECT 382.020 2370.380 385.020 2370.390 ;
        RECT 562.020 2370.380 565.020 2370.390 ;
        RECT 742.020 2370.380 745.020 2370.390 ;
        RECT 922.020 2370.380 925.020 2370.390 ;
        RECT 1102.020 2370.380 1105.020 2370.390 ;
        RECT 1282.020 2370.380 1285.020 2370.390 ;
        RECT 1462.020 2370.380 1465.020 2370.390 ;
        RECT 1642.020 2370.380 1645.020 2370.390 ;
        RECT 1822.020 2370.380 1825.020 2370.390 ;
        RECT 2002.020 2370.380 2005.020 2370.390 ;
        RECT 2182.020 2370.380 2185.020 2370.390 ;
        RECT 2362.020 2370.380 2365.020 2370.390 ;
        RECT 2542.020 2370.380 2545.020 2370.390 ;
        RECT 2722.020 2370.380 2725.020 2370.390 ;
        RECT 2902.020 2370.380 2905.020 2370.390 ;
        RECT 2935.800 2370.380 2938.800 2370.390 ;
        RECT -23.780 2367.380 2943.400 2370.380 ;
        RECT -19.180 2367.370 -16.180 2367.380 ;
        RECT 22.020 2367.370 25.020 2367.380 ;
        RECT 202.020 2367.370 205.020 2367.380 ;
        RECT 382.020 2367.370 385.020 2367.380 ;
        RECT 562.020 2367.370 565.020 2367.380 ;
        RECT 742.020 2367.370 745.020 2367.380 ;
        RECT 922.020 2367.370 925.020 2367.380 ;
        RECT 1102.020 2367.370 1105.020 2367.380 ;
        RECT 1282.020 2367.370 1285.020 2367.380 ;
        RECT 1462.020 2367.370 1465.020 2367.380 ;
        RECT 1642.020 2367.370 1645.020 2367.380 ;
        RECT 1822.020 2367.370 1825.020 2367.380 ;
        RECT 2002.020 2367.370 2005.020 2367.380 ;
        RECT 2182.020 2367.370 2185.020 2367.380 ;
        RECT 2362.020 2367.370 2365.020 2367.380 ;
        RECT 2542.020 2367.370 2545.020 2367.380 ;
        RECT 2722.020 2367.370 2725.020 2367.380 ;
        RECT 2902.020 2367.370 2905.020 2367.380 ;
        RECT 2935.800 2367.370 2938.800 2367.380 ;
        RECT -19.180 2190.380 -16.180 2190.390 ;
        RECT 22.020 2190.380 25.020 2190.390 ;
        RECT 202.020 2190.380 205.020 2190.390 ;
        RECT 382.020 2190.380 385.020 2190.390 ;
        RECT 562.020 2190.380 565.020 2190.390 ;
        RECT 742.020 2190.380 745.020 2190.390 ;
        RECT 922.020 2190.380 925.020 2190.390 ;
        RECT 1102.020 2190.380 1105.020 2190.390 ;
        RECT 1282.020 2190.380 1285.020 2190.390 ;
        RECT 1462.020 2190.380 1465.020 2190.390 ;
        RECT 1642.020 2190.380 1645.020 2190.390 ;
        RECT 1822.020 2190.380 1825.020 2190.390 ;
        RECT 2002.020 2190.380 2005.020 2190.390 ;
        RECT 2182.020 2190.380 2185.020 2190.390 ;
        RECT 2362.020 2190.380 2365.020 2190.390 ;
        RECT 2542.020 2190.380 2545.020 2190.390 ;
        RECT 2722.020 2190.380 2725.020 2190.390 ;
        RECT 2902.020 2190.380 2905.020 2190.390 ;
        RECT 2935.800 2190.380 2938.800 2190.390 ;
        RECT -23.780 2187.380 2943.400 2190.380 ;
        RECT -19.180 2187.370 -16.180 2187.380 ;
        RECT 22.020 2187.370 25.020 2187.380 ;
        RECT 202.020 2187.370 205.020 2187.380 ;
        RECT 382.020 2187.370 385.020 2187.380 ;
        RECT 562.020 2187.370 565.020 2187.380 ;
        RECT 742.020 2187.370 745.020 2187.380 ;
        RECT 922.020 2187.370 925.020 2187.380 ;
        RECT 1102.020 2187.370 1105.020 2187.380 ;
        RECT 1282.020 2187.370 1285.020 2187.380 ;
        RECT 1462.020 2187.370 1465.020 2187.380 ;
        RECT 1642.020 2187.370 1645.020 2187.380 ;
        RECT 1822.020 2187.370 1825.020 2187.380 ;
        RECT 2002.020 2187.370 2005.020 2187.380 ;
        RECT 2182.020 2187.370 2185.020 2187.380 ;
        RECT 2362.020 2187.370 2365.020 2187.380 ;
        RECT 2542.020 2187.370 2545.020 2187.380 ;
        RECT 2722.020 2187.370 2725.020 2187.380 ;
        RECT 2902.020 2187.370 2905.020 2187.380 ;
        RECT 2935.800 2187.370 2938.800 2187.380 ;
        RECT -19.180 2010.380 -16.180 2010.390 ;
        RECT 22.020 2010.380 25.020 2010.390 ;
        RECT 202.020 2010.380 205.020 2010.390 ;
        RECT 382.020 2010.380 385.020 2010.390 ;
        RECT 562.020 2010.380 565.020 2010.390 ;
        RECT 742.020 2010.380 745.020 2010.390 ;
        RECT 922.020 2010.380 925.020 2010.390 ;
        RECT 1102.020 2010.380 1105.020 2010.390 ;
        RECT 1282.020 2010.380 1285.020 2010.390 ;
        RECT 1462.020 2010.380 1465.020 2010.390 ;
        RECT 1642.020 2010.380 1645.020 2010.390 ;
        RECT 1822.020 2010.380 1825.020 2010.390 ;
        RECT 2002.020 2010.380 2005.020 2010.390 ;
        RECT 2182.020 2010.380 2185.020 2010.390 ;
        RECT 2362.020 2010.380 2365.020 2010.390 ;
        RECT 2542.020 2010.380 2545.020 2010.390 ;
        RECT 2722.020 2010.380 2725.020 2010.390 ;
        RECT 2902.020 2010.380 2905.020 2010.390 ;
        RECT 2935.800 2010.380 2938.800 2010.390 ;
        RECT -23.780 2007.380 2943.400 2010.380 ;
        RECT -19.180 2007.370 -16.180 2007.380 ;
        RECT 22.020 2007.370 25.020 2007.380 ;
        RECT 202.020 2007.370 205.020 2007.380 ;
        RECT 382.020 2007.370 385.020 2007.380 ;
        RECT 562.020 2007.370 565.020 2007.380 ;
        RECT 742.020 2007.370 745.020 2007.380 ;
        RECT 922.020 2007.370 925.020 2007.380 ;
        RECT 1102.020 2007.370 1105.020 2007.380 ;
        RECT 1282.020 2007.370 1285.020 2007.380 ;
        RECT 1462.020 2007.370 1465.020 2007.380 ;
        RECT 1642.020 2007.370 1645.020 2007.380 ;
        RECT 1822.020 2007.370 1825.020 2007.380 ;
        RECT 2002.020 2007.370 2005.020 2007.380 ;
        RECT 2182.020 2007.370 2185.020 2007.380 ;
        RECT 2362.020 2007.370 2365.020 2007.380 ;
        RECT 2542.020 2007.370 2545.020 2007.380 ;
        RECT 2722.020 2007.370 2725.020 2007.380 ;
        RECT 2902.020 2007.370 2905.020 2007.380 ;
        RECT 2935.800 2007.370 2938.800 2007.380 ;
        RECT -19.180 1830.380 -16.180 1830.390 ;
        RECT 22.020 1830.380 25.020 1830.390 ;
        RECT 202.020 1830.380 205.020 1830.390 ;
        RECT 382.020 1830.380 385.020 1830.390 ;
        RECT 562.020 1830.380 565.020 1830.390 ;
        RECT 742.020 1830.380 745.020 1830.390 ;
        RECT 922.020 1830.380 925.020 1830.390 ;
        RECT 1102.020 1830.380 1105.020 1830.390 ;
        RECT 1282.020 1830.380 1285.020 1830.390 ;
        RECT 1462.020 1830.380 1465.020 1830.390 ;
        RECT 1642.020 1830.380 1645.020 1830.390 ;
        RECT 1822.020 1830.380 1825.020 1830.390 ;
        RECT 2002.020 1830.380 2005.020 1830.390 ;
        RECT 2182.020 1830.380 2185.020 1830.390 ;
        RECT 2362.020 1830.380 2365.020 1830.390 ;
        RECT 2542.020 1830.380 2545.020 1830.390 ;
        RECT 2722.020 1830.380 2725.020 1830.390 ;
        RECT 2902.020 1830.380 2905.020 1830.390 ;
        RECT 2935.800 1830.380 2938.800 1830.390 ;
        RECT -23.780 1827.380 2943.400 1830.380 ;
        RECT -19.180 1827.370 -16.180 1827.380 ;
        RECT 22.020 1827.370 25.020 1827.380 ;
        RECT 202.020 1827.370 205.020 1827.380 ;
        RECT 382.020 1827.370 385.020 1827.380 ;
        RECT 562.020 1827.370 565.020 1827.380 ;
        RECT 742.020 1827.370 745.020 1827.380 ;
        RECT 922.020 1827.370 925.020 1827.380 ;
        RECT 1102.020 1827.370 1105.020 1827.380 ;
        RECT 1282.020 1827.370 1285.020 1827.380 ;
        RECT 1462.020 1827.370 1465.020 1827.380 ;
        RECT 1642.020 1827.370 1645.020 1827.380 ;
        RECT 1822.020 1827.370 1825.020 1827.380 ;
        RECT 2002.020 1827.370 2005.020 1827.380 ;
        RECT 2182.020 1827.370 2185.020 1827.380 ;
        RECT 2362.020 1827.370 2365.020 1827.380 ;
        RECT 2542.020 1827.370 2545.020 1827.380 ;
        RECT 2722.020 1827.370 2725.020 1827.380 ;
        RECT 2902.020 1827.370 2905.020 1827.380 ;
        RECT 2935.800 1827.370 2938.800 1827.380 ;
        RECT -19.180 1650.380 -16.180 1650.390 ;
        RECT 22.020 1650.380 25.020 1650.390 ;
        RECT 202.020 1650.380 205.020 1650.390 ;
        RECT 382.020 1650.380 385.020 1650.390 ;
        RECT 562.020 1650.380 565.020 1650.390 ;
        RECT 742.020 1650.380 745.020 1650.390 ;
        RECT 922.020 1650.380 925.020 1650.390 ;
        RECT 1102.020 1650.380 1105.020 1650.390 ;
        RECT 1282.020 1650.380 1285.020 1650.390 ;
        RECT 1462.020 1650.380 1465.020 1650.390 ;
        RECT 1642.020 1650.380 1645.020 1650.390 ;
        RECT 1822.020 1650.380 1825.020 1650.390 ;
        RECT 2002.020 1650.380 2005.020 1650.390 ;
        RECT 2182.020 1650.380 2185.020 1650.390 ;
        RECT 2362.020 1650.380 2365.020 1650.390 ;
        RECT 2542.020 1650.380 2545.020 1650.390 ;
        RECT 2722.020 1650.380 2725.020 1650.390 ;
        RECT 2902.020 1650.380 2905.020 1650.390 ;
        RECT 2935.800 1650.380 2938.800 1650.390 ;
        RECT -23.780 1647.380 2943.400 1650.380 ;
        RECT -19.180 1647.370 -16.180 1647.380 ;
        RECT 22.020 1647.370 25.020 1647.380 ;
        RECT 202.020 1647.370 205.020 1647.380 ;
        RECT 382.020 1647.370 385.020 1647.380 ;
        RECT 562.020 1647.370 565.020 1647.380 ;
        RECT 742.020 1647.370 745.020 1647.380 ;
        RECT 922.020 1647.370 925.020 1647.380 ;
        RECT 1102.020 1647.370 1105.020 1647.380 ;
        RECT 1282.020 1647.370 1285.020 1647.380 ;
        RECT 1462.020 1647.370 1465.020 1647.380 ;
        RECT 1642.020 1647.370 1645.020 1647.380 ;
        RECT 1822.020 1647.370 1825.020 1647.380 ;
        RECT 2002.020 1647.370 2005.020 1647.380 ;
        RECT 2182.020 1647.370 2185.020 1647.380 ;
        RECT 2362.020 1647.370 2365.020 1647.380 ;
        RECT 2542.020 1647.370 2545.020 1647.380 ;
        RECT 2722.020 1647.370 2725.020 1647.380 ;
        RECT 2902.020 1647.370 2905.020 1647.380 ;
        RECT 2935.800 1647.370 2938.800 1647.380 ;
        RECT -19.180 1470.380 -16.180 1470.390 ;
        RECT 22.020 1470.380 25.020 1470.390 ;
        RECT 202.020 1470.380 205.020 1470.390 ;
        RECT 382.020 1470.380 385.020 1470.390 ;
        RECT 562.020 1470.380 565.020 1470.390 ;
        RECT 742.020 1470.380 745.020 1470.390 ;
        RECT 922.020 1470.380 925.020 1470.390 ;
        RECT 1102.020 1470.380 1105.020 1470.390 ;
        RECT 1282.020 1470.380 1285.020 1470.390 ;
        RECT 1462.020 1470.380 1465.020 1470.390 ;
        RECT 1642.020 1470.380 1645.020 1470.390 ;
        RECT 1822.020 1470.380 1825.020 1470.390 ;
        RECT 2002.020 1470.380 2005.020 1470.390 ;
        RECT 2182.020 1470.380 2185.020 1470.390 ;
        RECT 2362.020 1470.380 2365.020 1470.390 ;
        RECT 2542.020 1470.380 2545.020 1470.390 ;
        RECT 2722.020 1470.380 2725.020 1470.390 ;
        RECT 2902.020 1470.380 2905.020 1470.390 ;
        RECT 2935.800 1470.380 2938.800 1470.390 ;
        RECT -23.780 1467.380 2943.400 1470.380 ;
        RECT -19.180 1467.370 -16.180 1467.380 ;
        RECT 22.020 1467.370 25.020 1467.380 ;
        RECT 202.020 1467.370 205.020 1467.380 ;
        RECT 382.020 1467.370 385.020 1467.380 ;
        RECT 562.020 1467.370 565.020 1467.380 ;
        RECT 742.020 1467.370 745.020 1467.380 ;
        RECT 922.020 1467.370 925.020 1467.380 ;
        RECT 1102.020 1467.370 1105.020 1467.380 ;
        RECT 1282.020 1467.370 1285.020 1467.380 ;
        RECT 1462.020 1467.370 1465.020 1467.380 ;
        RECT 1642.020 1467.370 1645.020 1467.380 ;
        RECT 1822.020 1467.370 1825.020 1467.380 ;
        RECT 2002.020 1467.370 2005.020 1467.380 ;
        RECT 2182.020 1467.370 2185.020 1467.380 ;
        RECT 2362.020 1467.370 2365.020 1467.380 ;
        RECT 2542.020 1467.370 2545.020 1467.380 ;
        RECT 2722.020 1467.370 2725.020 1467.380 ;
        RECT 2902.020 1467.370 2905.020 1467.380 ;
        RECT 2935.800 1467.370 2938.800 1467.380 ;
        RECT -19.180 1290.380 -16.180 1290.390 ;
        RECT 22.020 1290.380 25.020 1290.390 ;
        RECT 202.020 1290.380 205.020 1290.390 ;
        RECT 382.020 1290.380 385.020 1290.390 ;
        RECT 562.020 1290.380 565.020 1290.390 ;
        RECT 742.020 1290.380 745.020 1290.390 ;
        RECT 922.020 1290.380 925.020 1290.390 ;
        RECT 1102.020 1290.380 1105.020 1290.390 ;
        RECT 1282.020 1290.380 1285.020 1290.390 ;
        RECT 1462.020 1290.380 1465.020 1290.390 ;
        RECT 1642.020 1290.380 1645.020 1290.390 ;
        RECT 1822.020 1290.380 1825.020 1290.390 ;
        RECT 2002.020 1290.380 2005.020 1290.390 ;
        RECT 2182.020 1290.380 2185.020 1290.390 ;
        RECT 2362.020 1290.380 2365.020 1290.390 ;
        RECT 2542.020 1290.380 2545.020 1290.390 ;
        RECT 2722.020 1290.380 2725.020 1290.390 ;
        RECT 2902.020 1290.380 2905.020 1290.390 ;
        RECT 2935.800 1290.380 2938.800 1290.390 ;
        RECT -23.780 1287.380 2943.400 1290.380 ;
        RECT -19.180 1287.370 -16.180 1287.380 ;
        RECT 22.020 1287.370 25.020 1287.380 ;
        RECT 202.020 1287.370 205.020 1287.380 ;
        RECT 382.020 1287.370 385.020 1287.380 ;
        RECT 562.020 1287.370 565.020 1287.380 ;
        RECT 742.020 1287.370 745.020 1287.380 ;
        RECT 922.020 1287.370 925.020 1287.380 ;
        RECT 1102.020 1287.370 1105.020 1287.380 ;
        RECT 1282.020 1287.370 1285.020 1287.380 ;
        RECT 1462.020 1287.370 1465.020 1287.380 ;
        RECT 1642.020 1287.370 1645.020 1287.380 ;
        RECT 1822.020 1287.370 1825.020 1287.380 ;
        RECT 2002.020 1287.370 2005.020 1287.380 ;
        RECT 2182.020 1287.370 2185.020 1287.380 ;
        RECT 2362.020 1287.370 2365.020 1287.380 ;
        RECT 2542.020 1287.370 2545.020 1287.380 ;
        RECT 2722.020 1287.370 2725.020 1287.380 ;
        RECT 2902.020 1287.370 2905.020 1287.380 ;
        RECT 2935.800 1287.370 2938.800 1287.380 ;
        RECT -19.180 1110.380 -16.180 1110.390 ;
        RECT 22.020 1110.380 25.020 1110.390 ;
        RECT 202.020 1110.380 205.020 1110.390 ;
        RECT 382.020 1110.380 385.020 1110.390 ;
        RECT 562.020 1110.380 565.020 1110.390 ;
        RECT 742.020 1110.380 745.020 1110.390 ;
        RECT 922.020 1110.380 925.020 1110.390 ;
        RECT 1102.020 1110.380 1105.020 1110.390 ;
        RECT 1282.020 1110.380 1285.020 1110.390 ;
        RECT 1462.020 1110.380 1465.020 1110.390 ;
        RECT 1642.020 1110.380 1645.020 1110.390 ;
        RECT 1822.020 1110.380 1825.020 1110.390 ;
        RECT 2002.020 1110.380 2005.020 1110.390 ;
        RECT 2182.020 1110.380 2185.020 1110.390 ;
        RECT 2362.020 1110.380 2365.020 1110.390 ;
        RECT 2542.020 1110.380 2545.020 1110.390 ;
        RECT 2722.020 1110.380 2725.020 1110.390 ;
        RECT 2902.020 1110.380 2905.020 1110.390 ;
        RECT 2935.800 1110.380 2938.800 1110.390 ;
        RECT -23.780 1107.380 2943.400 1110.380 ;
        RECT -19.180 1107.370 -16.180 1107.380 ;
        RECT 22.020 1107.370 25.020 1107.380 ;
        RECT 202.020 1107.370 205.020 1107.380 ;
        RECT 382.020 1107.370 385.020 1107.380 ;
        RECT 562.020 1107.370 565.020 1107.380 ;
        RECT 742.020 1107.370 745.020 1107.380 ;
        RECT 922.020 1107.370 925.020 1107.380 ;
        RECT 1102.020 1107.370 1105.020 1107.380 ;
        RECT 1282.020 1107.370 1285.020 1107.380 ;
        RECT 1462.020 1107.370 1465.020 1107.380 ;
        RECT 1642.020 1107.370 1645.020 1107.380 ;
        RECT 1822.020 1107.370 1825.020 1107.380 ;
        RECT 2002.020 1107.370 2005.020 1107.380 ;
        RECT 2182.020 1107.370 2185.020 1107.380 ;
        RECT 2362.020 1107.370 2365.020 1107.380 ;
        RECT 2542.020 1107.370 2545.020 1107.380 ;
        RECT 2722.020 1107.370 2725.020 1107.380 ;
        RECT 2902.020 1107.370 2905.020 1107.380 ;
        RECT 2935.800 1107.370 2938.800 1107.380 ;
        RECT -19.180 930.380 -16.180 930.390 ;
        RECT 22.020 930.380 25.020 930.390 ;
        RECT 202.020 930.380 205.020 930.390 ;
        RECT 382.020 930.380 385.020 930.390 ;
        RECT 562.020 930.380 565.020 930.390 ;
        RECT 742.020 930.380 745.020 930.390 ;
        RECT 922.020 930.380 925.020 930.390 ;
        RECT 1102.020 930.380 1105.020 930.390 ;
        RECT 1282.020 930.380 1285.020 930.390 ;
        RECT 1462.020 930.380 1465.020 930.390 ;
        RECT 1642.020 930.380 1645.020 930.390 ;
        RECT 1822.020 930.380 1825.020 930.390 ;
        RECT 2002.020 930.380 2005.020 930.390 ;
        RECT 2182.020 930.380 2185.020 930.390 ;
        RECT 2362.020 930.380 2365.020 930.390 ;
        RECT 2542.020 930.380 2545.020 930.390 ;
        RECT 2722.020 930.380 2725.020 930.390 ;
        RECT 2902.020 930.380 2905.020 930.390 ;
        RECT 2935.800 930.380 2938.800 930.390 ;
        RECT -23.780 927.380 2943.400 930.380 ;
        RECT -19.180 927.370 -16.180 927.380 ;
        RECT 22.020 927.370 25.020 927.380 ;
        RECT 202.020 927.370 205.020 927.380 ;
        RECT 382.020 927.370 385.020 927.380 ;
        RECT 562.020 927.370 565.020 927.380 ;
        RECT 742.020 927.370 745.020 927.380 ;
        RECT 922.020 927.370 925.020 927.380 ;
        RECT 1102.020 927.370 1105.020 927.380 ;
        RECT 1282.020 927.370 1285.020 927.380 ;
        RECT 1462.020 927.370 1465.020 927.380 ;
        RECT 1642.020 927.370 1645.020 927.380 ;
        RECT 1822.020 927.370 1825.020 927.380 ;
        RECT 2002.020 927.370 2005.020 927.380 ;
        RECT 2182.020 927.370 2185.020 927.380 ;
        RECT 2362.020 927.370 2365.020 927.380 ;
        RECT 2542.020 927.370 2545.020 927.380 ;
        RECT 2722.020 927.370 2725.020 927.380 ;
        RECT 2902.020 927.370 2905.020 927.380 ;
        RECT 2935.800 927.370 2938.800 927.380 ;
        RECT -19.180 750.380 -16.180 750.390 ;
        RECT 22.020 750.380 25.020 750.390 ;
        RECT 202.020 750.380 205.020 750.390 ;
        RECT 382.020 750.380 385.020 750.390 ;
        RECT 562.020 750.380 565.020 750.390 ;
        RECT 742.020 750.380 745.020 750.390 ;
        RECT 922.020 750.380 925.020 750.390 ;
        RECT 1102.020 750.380 1105.020 750.390 ;
        RECT 1282.020 750.380 1285.020 750.390 ;
        RECT 1462.020 750.380 1465.020 750.390 ;
        RECT 1642.020 750.380 1645.020 750.390 ;
        RECT 1822.020 750.380 1825.020 750.390 ;
        RECT 2002.020 750.380 2005.020 750.390 ;
        RECT 2182.020 750.380 2185.020 750.390 ;
        RECT 2362.020 750.380 2365.020 750.390 ;
        RECT 2542.020 750.380 2545.020 750.390 ;
        RECT 2722.020 750.380 2725.020 750.390 ;
        RECT 2902.020 750.380 2905.020 750.390 ;
        RECT 2935.800 750.380 2938.800 750.390 ;
        RECT -23.780 747.380 2943.400 750.380 ;
        RECT -19.180 747.370 -16.180 747.380 ;
        RECT 22.020 747.370 25.020 747.380 ;
        RECT 202.020 747.370 205.020 747.380 ;
        RECT 382.020 747.370 385.020 747.380 ;
        RECT 562.020 747.370 565.020 747.380 ;
        RECT 742.020 747.370 745.020 747.380 ;
        RECT 922.020 747.370 925.020 747.380 ;
        RECT 1102.020 747.370 1105.020 747.380 ;
        RECT 1282.020 747.370 1285.020 747.380 ;
        RECT 1462.020 747.370 1465.020 747.380 ;
        RECT 1642.020 747.370 1645.020 747.380 ;
        RECT 1822.020 747.370 1825.020 747.380 ;
        RECT 2002.020 747.370 2005.020 747.380 ;
        RECT 2182.020 747.370 2185.020 747.380 ;
        RECT 2362.020 747.370 2365.020 747.380 ;
        RECT 2542.020 747.370 2545.020 747.380 ;
        RECT 2722.020 747.370 2725.020 747.380 ;
        RECT 2902.020 747.370 2905.020 747.380 ;
        RECT 2935.800 747.370 2938.800 747.380 ;
        RECT -19.180 570.380 -16.180 570.390 ;
        RECT 22.020 570.380 25.020 570.390 ;
        RECT 202.020 570.380 205.020 570.390 ;
        RECT 382.020 570.380 385.020 570.390 ;
        RECT 562.020 570.380 565.020 570.390 ;
        RECT 742.020 570.380 745.020 570.390 ;
        RECT 922.020 570.380 925.020 570.390 ;
        RECT 1102.020 570.380 1105.020 570.390 ;
        RECT 1282.020 570.380 1285.020 570.390 ;
        RECT 1462.020 570.380 1465.020 570.390 ;
        RECT 1642.020 570.380 1645.020 570.390 ;
        RECT 1822.020 570.380 1825.020 570.390 ;
        RECT 2002.020 570.380 2005.020 570.390 ;
        RECT 2182.020 570.380 2185.020 570.390 ;
        RECT 2362.020 570.380 2365.020 570.390 ;
        RECT 2542.020 570.380 2545.020 570.390 ;
        RECT 2722.020 570.380 2725.020 570.390 ;
        RECT 2902.020 570.380 2905.020 570.390 ;
        RECT 2935.800 570.380 2938.800 570.390 ;
        RECT -23.780 567.380 2943.400 570.380 ;
        RECT -19.180 567.370 -16.180 567.380 ;
        RECT 22.020 567.370 25.020 567.380 ;
        RECT 202.020 567.370 205.020 567.380 ;
        RECT 382.020 567.370 385.020 567.380 ;
        RECT 562.020 567.370 565.020 567.380 ;
        RECT 742.020 567.370 745.020 567.380 ;
        RECT 922.020 567.370 925.020 567.380 ;
        RECT 1102.020 567.370 1105.020 567.380 ;
        RECT 1282.020 567.370 1285.020 567.380 ;
        RECT 1462.020 567.370 1465.020 567.380 ;
        RECT 1642.020 567.370 1645.020 567.380 ;
        RECT 1822.020 567.370 1825.020 567.380 ;
        RECT 2002.020 567.370 2005.020 567.380 ;
        RECT 2182.020 567.370 2185.020 567.380 ;
        RECT 2362.020 567.370 2365.020 567.380 ;
        RECT 2542.020 567.370 2545.020 567.380 ;
        RECT 2722.020 567.370 2725.020 567.380 ;
        RECT 2902.020 567.370 2905.020 567.380 ;
        RECT 2935.800 567.370 2938.800 567.380 ;
        RECT -19.180 390.380 -16.180 390.390 ;
        RECT 22.020 390.380 25.020 390.390 ;
        RECT 202.020 390.380 205.020 390.390 ;
        RECT 382.020 390.380 385.020 390.390 ;
        RECT 562.020 390.380 565.020 390.390 ;
        RECT 742.020 390.380 745.020 390.390 ;
        RECT 922.020 390.380 925.020 390.390 ;
        RECT 1102.020 390.380 1105.020 390.390 ;
        RECT 1282.020 390.380 1285.020 390.390 ;
        RECT 1462.020 390.380 1465.020 390.390 ;
        RECT 1642.020 390.380 1645.020 390.390 ;
        RECT 1822.020 390.380 1825.020 390.390 ;
        RECT 2002.020 390.380 2005.020 390.390 ;
        RECT 2182.020 390.380 2185.020 390.390 ;
        RECT 2362.020 390.380 2365.020 390.390 ;
        RECT 2542.020 390.380 2545.020 390.390 ;
        RECT 2722.020 390.380 2725.020 390.390 ;
        RECT 2902.020 390.380 2905.020 390.390 ;
        RECT 2935.800 390.380 2938.800 390.390 ;
        RECT -23.780 387.380 2943.400 390.380 ;
        RECT -19.180 387.370 -16.180 387.380 ;
        RECT 22.020 387.370 25.020 387.380 ;
        RECT 202.020 387.370 205.020 387.380 ;
        RECT 382.020 387.370 385.020 387.380 ;
        RECT 562.020 387.370 565.020 387.380 ;
        RECT 742.020 387.370 745.020 387.380 ;
        RECT 922.020 387.370 925.020 387.380 ;
        RECT 1102.020 387.370 1105.020 387.380 ;
        RECT 1282.020 387.370 1285.020 387.380 ;
        RECT 1462.020 387.370 1465.020 387.380 ;
        RECT 1642.020 387.370 1645.020 387.380 ;
        RECT 1822.020 387.370 1825.020 387.380 ;
        RECT 2002.020 387.370 2005.020 387.380 ;
        RECT 2182.020 387.370 2185.020 387.380 ;
        RECT 2362.020 387.370 2365.020 387.380 ;
        RECT 2542.020 387.370 2545.020 387.380 ;
        RECT 2722.020 387.370 2725.020 387.380 ;
        RECT 2902.020 387.370 2905.020 387.380 ;
        RECT 2935.800 387.370 2938.800 387.380 ;
        RECT -19.180 210.380 -16.180 210.390 ;
        RECT 22.020 210.380 25.020 210.390 ;
        RECT 202.020 210.380 205.020 210.390 ;
        RECT 382.020 210.380 385.020 210.390 ;
        RECT 562.020 210.380 565.020 210.390 ;
        RECT 742.020 210.380 745.020 210.390 ;
        RECT 922.020 210.380 925.020 210.390 ;
        RECT 1102.020 210.380 1105.020 210.390 ;
        RECT 1282.020 210.380 1285.020 210.390 ;
        RECT 1462.020 210.380 1465.020 210.390 ;
        RECT 1642.020 210.380 1645.020 210.390 ;
        RECT 1822.020 210.380 1825.020 210.390 ;
        RECT 2002.020 210.380 2005.020 210.390 ;
        RECT 2182.020 210.380 2185.020 210.390 ;
        RECT 2362.020 210.380 2365.020 210.390 ;
        RECT 2542.020 210.380 2545.020 210.390 ;
        RECT 2722.020 210.380 2725.020 210.390 ;
        RECT 2902.020 210.380 2905.020 210.390 ;
        RECT 2935.800 210.380 2938.800 210.390 ;
        RECT -23.780 207.380 2943.400 210.380 ;
        RECT -19.180 207.370 -16.180 207.380 ;
        RECT 22.020 207.370 25.020 207.380 ;
        RECT 202.020 207.370 205.020 207.380 ;
        RECT 382.020 207.370 385.020 207.380 ;
        RECT 562.020 207.370 565.020 207.380 ;
        RECT 742.020 207.370 745.020 207.380 ;
        RECT 922.020 207.370 925.020 207.380 ;
        RECT 1102.020 207.370 1105.020 207.380 ;
        RECT 1282.020 207.370 1285.020 207.380 ;
        RECT 1462.020 207.370 1465.020 207.380 ;
        RECT 1642.020 207.370 1645.020 207.380 ;
        RECT 1822.020 207.370 1825.020 207.380 ;
        RECT 2002.020 207.370 2005.020 207.380 ;
        RECT 2182.020 207.370 2185.020 207.380 ;
        RECT 2362.020 207.370 2365.020 207.380 ;
        RECT 2542.020 207.370 2545.020 207.380 ;
        RECT 2722.020 207.370 2725.020 207.380 ;
        RECT 2902.020 207.370 2905.020 207.380 ;
        RECT 2935.800 207.370 2938.800 207.380 ;
        RECT -19.180 30.380 -16.180 30.390 ;
        RECT 22.020 30.380 25.020 30.390 ;
        RECT 202.020 30.380 205.020 30.390 ;
        RECT 382.020 30.380 385.020 30.390 ;
        RECT 562.020 30.380 565.020 30.390 ;
        RECT 742.020 30.380 745.020 30.390 ;
        RECT 922.020 30.380 925.020 30.390 ;
        RECT 1102.020 30.380 1105.020 30.390 ;
        RECT 1282.020 30.380 1285.020 30.390 ;
        RECT 1462.020 30.380 1465.020 30.390 ;
        RECT 1642.020 30.380 1645.020 30.390 ;
        RECT 1822.020 30.380 1825.020 30.390 ;
        RECT 2002.020 30.380 2005.020 30.390 ;
        RECT 2182.020 30.380 2185.020 30.390 ;
        RECT 2362.020 30.380 2365.020 30.390 ;
        RECT 2542.020 30.380 2545.020 30.390 ;
        RECT 2722.020 30.380 2725.020 30.390 ;
        RECT 2902.020 30.380 2905.020 30.390 ;
        RECT 2935.800 30.380 2938.800 30.390 ;
        RECT -23.780 27.380 2943.400 30.380 ;
        RECT -19.180 27.370 -16.180 27.380 ;
        RECT 22.020 27.370 25.020 27.380 ;
        RECT 202.020 27.370 205.020 27.380 ;
        RECT 382.020 27.370 385.020 27.380 ;
        RECT 562.020 27.370 565.020 27.380 ;
        RECT 742.020 27.370 745.020 27.380 ;
        RECT 922.020 27.370 925.020 27.380 ;
        RECT 1102.020 27.370 1105.020 27.380 ;
        RECT 1282.020 27.370 1285.020 27.380 ;
        RECT 1462.020 27.370 1465.020 27.380 ;
        RECT 1642.020 27.370 1645.020 27.380 ;
        RECT 1822.020 27.370 1825.020 27.380 ;
        RECT 2002.020 27.370 2005.020 27.380 ;
        RECT 2182.020 27.370 2185.020 27.380 ;
        RECT 2362.020 27.370 2365.020 27.380 ;
        RECT 2542.020 27.370 2545.020 27.380 ;
        RECT 2722.020 27.370 2725.020 27.380 ;
        RECT 2902.020 27.370 2905.020 27.380 ;
        RECT 2935.800 27.370 2938.800 27.380 ;
        RECT -19.180 -10.820 -16.180 -10.810 ;
        RECT 22.020 -10.820 25.020 -10.810 ;
        RECT 202.020 -10.820 205.020 -10.810 ;
        RECT 382.020 -10.820 385.020 -10.810 ;
        RECT 562.020 -10.820 565.020 -10.810 ;
        RECT 742.020 -10.820 745.020 -10.810 ;
        RECT 922.020 -10.820 925.020 -10.810 ;
        RECT 1102.020 -10.820 1105.020 -10.810 ;
        RECT 1282.020 -10.820 1285.020 -10.810 ;
        RECT 1462.020 -10.820 1465.020 -10.810 ;
        RECT 1642.020 -10.820 1645.020 -10.810 ;
        RECT 1822.020 -10.820 1825.020 -10.810 ;
        RECT 2002.020 -10.820 2005.020 -10.810 ;
        RECT 2182.020 -10.820 2185.020 -10.810 ;
        RECT 2362.020 -10.820 2365.020 -10.810 ;
        RECT 2542.020 -10.820 2545.020 -10.810 ;
        RECT 2722.020 -10.820 2725.020 -10.810 ;
        RECT 2902.020 -10.820 2905.020 -10.810 ;
        RECT 2935.800 -10.820 2938.800 -10.810 ;
        RECT -19.180 -13.820 2938.800 -10.820 ;
        RECT -19.180 -13.830 -16.180 -13.820 ;
        RECT 22.020 -13.830 25.020 -13.820 ;
        RECT 202.020 -13.830 205.020 -13.820 ;
        RECT 382.020 -13.830 385.020 -13.820 ;
        RECT 562.020 -13.830 565.020 -13.820 ;
        RECT 742.020 -13.830 745.020 -13.820 ;
        RECT 922.020 -13.830 925.020 -13.820 ;
        RECT 1102.020 -13.830 1105.020 -13.820 ;
        RECT 1282.020 -13.830 1285.020 -13.820 ;
        RECT 1462.020 -13.830 1465.020 -13.820 ;
        RECT 1642.020 -13.830 1645.020 -13.820 ;
        RECT 1822.020 -13.830 1825.020 -13.820 ;
        RECT 2002.020 -13.830 2005.020 -13.820 ;
        RECT 2182.020 -13.830 2185.020 -13.820 ;
        RECT 2362.020 -13.830 2365.020 -13.820 ;
        RECT 2542.020 -13.830 2545.020 -13.820 ;
        RECT 2722.020 -13.830 2725.020 -13.820 ;
        RECT 2902.020 -13.830 2905.020 -13.820 ;
        RECT 2935.800 -13.830 2938.800 -13.820 ;
    END
  END vccd2
  PIN vssd2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -23.780 -18.420 -20.780 3538.100 ;
        RECT 112.020 -18.420 115.020 3538.100 ;
        RECT 292.020 -18.420 295.020 3538.100 ;
        RECT 472.020 -18.420 475.020 3538.100 ;
        RECT 652.020 -18.420 655.020 3538.100 ;
        RECT 832.020 -18.420 835.020 3538.100 ;
        RECT 1012.020 -18.420 1015.020 3538.100 ;
        RECT 1192.020 -18.420 1195.020 3538.100 ;
        RECT 1372.020 -18.420 1375.020 3538.100 ;
        RECT 1552.020 -18.420 1555.020 3538.100 ;
        RECT 1732.020 -18.420 1735.020 3538.100 ;
        RECT 1912.020 -18.420 1915.020 3538.100 ;
        RECT 2092.020 -18.420 2095.020 3538.100 ;
        RECT 2272.020 -18.420 2275.020 3538.100 ;
        RECT 2452.020 -18.420 2455.020 3538.100 ;
        RECT 2632.020 -18.420 2635.020 3538.100 ;
        RECT 2812.020 -18.420 2815.020 3538.100 ;
        RECT 2940.400 -18.420 2943.400 3538.100 ;
      LAYER via4 ;
        RECT -22.870 3536.810 -21.690 3537.990 ;
        RECT -22.870 3535.210 -21.690 3536.390 ;
        RECT -22.870 3359.090 -21.690 3360.270 ;
        RECT -22.870 3357.490 -21.690 3358.670 ;
        RECT -22.870 3179.090 -21.690 3180.270 ;
        RECT -22.870 3177.490 -21.690 3178.670 ;
        RECT -22.870 2999.090 -21.690 3000.270 ;
        RECT -22.870 2997.490 -21.690 2998.670 ;
        RECT -22.870 2819.090 -21.690 2820.270 ;
        RECT -22.870 2817.490 -21.690 2818.670 ;
        RECT -22.870 2639.090 -21.690 2640.270 ;
        RECT -22.870 2637.490 -21.690 2638.670 ;
        RECT -22.870 2459.090 -21.690 2460.270 ;
        RECT -22.870 2457.490 -21.690 2458.670 ;
        RECT -22.870 2279.090 -21.690 2280.270 ;
        RECT -22.870 2277.490 -21.690 2278.670 ;
        RECT -22.870 2099.090 -21.690 2100.270 ;
        RECT -22.870 2097.490 -21.690 2098.670 ;
        RECT -22.870 1919.090 -21.690 1920.270 ;
        RECT -22.870 1917.490 -21.690 1918.670 ;
        RECT -22.870 1739.090 -21.690 1740.270 ;
        RECT -22.870 1737.490 -21.690 1738.670 ;
        RECT -22.870 1559.090 -21.690 1560.270 ;
        RECT -22.870 1557.490 -21.690 1558.670 ;
        RECT -22.870 1379.090 -21.690 1380.270 ;
        RECT -22.870 1377.490 -21.690 1378.670 ;
        RECT -22.870 1199.090 -21.690 1200.270 ;
        RECT -22.870 1197.490 -21.690 1198.670 ;
        RECT -22.870 1019.090 -21.690 1020.270 ;
        RECT -22.870 1017.490 -21.690 1018.670 ;
        RECT -22.870 839.090 -21.690 840.270 ;
        RECT -22.870 837.490 -21.690 838.670 ;
        RECT -22.870 659.090 -21.690 660.270 ;
        RECT -22.870 657.490 -21.690 658.670 ;
        RECT -22.870 479.090 -21.690 480.270 ;
        RECT -22.870 477.490 -21.690 478.670 ;
        RECT -22.870 299.090 -21.690 300.270 ;
        RECT -22.870 297.490 -21.690 298.670 ;
        RECT -22.870 119.090 -21.690 120.270 ;
        RECT -22.870 117.490 -21.690 118.670 ;
        RECT -22.870 -16.710 -21.690 -15.530 ;
        RECT -22.870 -18.310 -21.690 -17.130 ;
        RECT 112.930 3536.810 114.110 3537.990 ;
        RECT 112.930 3535.210 114.110 3536.390 ;
        RECT 112.930 3359.090 114.110 3360.270 ;
        RECT 112.930 3357.490 114.110 3358.670 ;
        RECT 112.930 3179.090 114.110 3180.270 ;
        RECT 112.930 3177.490 114.110 3178.670 ;
        RECT 112.930 2999.090 114.110 3000.270 ;
        RECT 112.930 2997.490 114.110 2998.670 ;
        RECT 112.930 2819.090 114.110 2820.270 ;
        RECT 112.930 2817.490 114.110 2818.670 ;
        RECT 112.930 2639.090 114.110 2640.270 ;
        RECT 112.930 2637.490 114.110 2638.670 ;
        RECT 112.930 2459.090 114.110 2460.270 ;
        RECT 112.930 2457.490 114.110 2458.670 ;
        RECT 112.930 2279.090 114.110 2280.270 ;
        RECT 112.930 2277.490 114.110 2278.670 ;
        RECT 112.930 2099.090 114.110 2100.270 ;
        RECT 112.930 2097.490 114.110 2098.670 ;
        RECT 112.930 1919.090 114.110 1920.270 ;
        RECT 112.930 1917.490 114.110 1918.670 ;
        RECT 112.930 1739.090 114.110 1740.270 ;
        RECT 112.930 1737.490 114.110 1738.670 ;
        RECT 112.930 1559.090 114.110 1560.270 ;
        RECT 112.930 1557.490 114.110 1558.670 ;
        RECT 112.930 1379.090 114.110 1380.270 ;
        RECT 112.930 1377.490 114.110 1378.670 ;
        RECT 112.930 1199.090 114.110 1200.270 ;
        RECT 112.930 1197.490 114.110 1198.670 ;
        RECT 112.930 1019.090 114.110 1020.270 ;
        RECT 112.930 1017.490 114.110 1018.670 ;
        RECT 112.930 839.090 114.110 840.270 ;
        RECT 112.930 837.490 114.110 838.670 ;
        RECT 112.930 659.090 114.110 660.270 ;
        RECT 112.930 657.490 114.110 658.670 ;
        RECT 112.930 479.090 114.110 480.270 ;
        RECT 112.930 477.490 114.110 478.670 ;
        RECT 112.930 299.090 114.110 300.270 ;
        RECT 112.930 297.490 114.110 298.670 ;
        RECT 112.930 119.090 114.110 120.270 ;
        RECT 112.930 117.490 114.110 118.670 ;
        RECT 112.930 -16.710 114.110 -15.530 ;
        RECT 112.930 -18.310 114.110 -17.130 ;
        RECT 292.930 3536.810 294.110 3537.990 ;
        RECT 292.930 3535.210 294.110 3536.390 ;
        RECT 292.930 3359.090 294.110 3360.270 ;
        RECT 292.930 3357.490 294.110 3358.670 ;
        RECT 292.930 3179.090 294.110 3180.270 ;
        RECT 292.930 3177.490 294.110 3178.670 ;
        RECT 292.930 2999.090 294.110 3000.270 ;
        RECT 292.930 2997.490 294.110 2998.670 ;
        RECT 292.930 2819.090 294.110 2820.270 ;
        RECT 292.930 2817.490 294.110 2818.670 ;
        RECT 292.930 2639.090 294.110 2640.270 ;
        RECT 292.930 2637.490 294.110 2638.670 ;
        RECT 292.930 2459.090 294.110 2460.270 ;
        RECT 292.930 2457.490 294.110 2458.670 ;
        RECT 292.930 2279.090 294.110 2280.270 ;
        RECT 292.930 2277.490 294.110 2278.670 ;
        RECT 292.930 2099.090 294.110 2100.270 ;
        RECT 292.930 2097.490 294.110 2098.670 ;
        RECT 292.930 1919.090 294.110 1920.270 ;
        RECT 292.930 1917.490 294.110 1918.670 ;
        RECT 292.930 1739.090 294.110 1740.270 ;
        RECT 292.930 1737.490 294.110 1738.670 ;
        RECT 292.930 1559.090 294.110 1560.270 ;
        RECT 292.930 1557.490 294.110 1558.670 ;
        RECT 292.930 1379.090 294.110 1380.270 ;
        RECT 292.930 1377.490 294.110 1378.670 ;
        RECT 292.930 1199.090 294.110 1200.270 ;
        RECT 292.930 1197.490 294.110 1198.670 ;
        RECT 292.930 1019.090 294.110 1020.270 ;
        RECT 292.930 1017.490 294.110 1018.670 ;
        RECT 292.930 839.090 294.110 840.270 ;
        RECT 292.930 837.490 294.110 838.670 ;
        RECT 292.930 659.090 294.110 660.270 ;
        RECT 292.930 657.490 294.110 658.670 ;
        RECT 292.930 479.090 294.110 480.270 ;
        RECT 292.930 477.490 294.110 478.670 ;
        RECT 292.930 299.090 294.110 300.270 ;
        RECT 292.930 297.490 294.110 298.670 ;
        RECT 292.930 119.090 294.110 120.270 ;
        RECT 292.930 117.490 294.110 118.670 ;
        RECT 292.930 -16.710 294.110 -15.530 ;
        RECT 292.930 -18.310 294.110 -17.130 ;
        RECT 472.930 3536.810 474.110 3537.990 ;
        RECT 472.930 3535.210 474.110 3536.390 ;
        RECT 472.930 3359.090 474.110 3360.270 ;
        RECT 472.930 3357.490 474.110 3358.670 ;
        RECT 472.930 3179.090 474.110 3180.270 ;
        RECT 472.930 3177.490 474.110 3178.670 ;
        RECT 472.930 2999.090 474.110 3000.270 ;
        RECT 472.930 2997.490 474.110 2998.670 ;
        RECT 472.930 2819.090 474.110 2820.270 ;
        RECT 472.930 2817.490 474.110 2818.670 ;
        RECT 472.930 2639.090 474.110 2640.270 ;
        RECT 472.930 2637.490 474.110 2638.670 ;
        RECT 472.930 2459.090 474.110 2460.270 ;
        RECT 472.930 2457.490 474.110 2458.670 ;
        RECT 472.930 2279.090 474.110 2280.270 ;
        RECT 472.930 2277.490 474.110 2278.670 ;
        RECT 472.930 2099.090 474.110 2100.270 ;
        RECT 472.930 2097.490 474.110 2098.670 ;
        RECT 472.930 1919.090 474.110 1920.270 ;
        RECT 472.930 1917.490 474.110 1918.670 ;
        RECT 472.930 1739.090 474.110 1740.270 ;
        RECT 472.930 1737.490 474.110 1738.670 ;
        RECT 472.930 1559.090 474.110 1560.270 ;
        RECT 472.930 1557.490 474.110 1558.670 ;
        RECT 472.930 1379.090 474.110 1380.270 ;
        RECT 472.930 1377.490 474.110 1378.670 ;
        RECT 472.930 1199.090 474.110 1200.270 ;
        RECT 472.930 1197.490 474.110 1198.670 ;
        RECT 472.930 1019.090 474.110 1020.270 ;
        RECT 472.930 1017.490 474.110 1018.670 ;
        RECT 472.930 839.090 474.110 840.270 ;
        RECT 472.930 837.490 474.110 838.670 ;
        RECT 472.930 659.090 474.110 660.270 ;
        RECT 472.930 657.490 474.110 658.670 ;
        RECT 472.930 479.090 474.110 480.270 ;
        RECT 472.930 477.490 474.110 478.670 ;
        RECT 472.930 299.090 474.110 300.270 ;
        RECT 472.930 297.490 474.110 298.670 ;
        RECT 472.930 119.090 474.110 120.270 ;
        RECT 472.930 117.490 474.110 118.670 ;
        RECT 472.930 -16.710 474.110 -15.530 ;
        RECT 472.930 -18.310 474.110 -17.130 ;
        RECT 652.930 3536.810 654.110 3537.990 ;
        RECT 652.930 3535.210 654.110 3536.390 ;
        RECT 652.930 3359.090 654.110 3360.270 ;
        RECT 652.930 3357.490 654.110 3358.670 ;
        RECT 652.930 3179.090 654.110 3180.270 ;
        RECT 652.930 3177.490 654.110 3178.670 ;
        RECT 652.930 2999.090 654.110 3000.270 ;
        RECT 652.930 2997.490 654.110 2998.670 ;
        RECT 652.930 2819.090 654.110 2820.270 ;
        RECT 652.930 2817.490 654.110 2818.670 ;
        RECT 652.930 2639.090 654.110 2640.270 ;
        RECT 652.930 2637.490 654.110 2638.670 ;
        RECT 652.930 2459.090 654.110 2460.270 ;
        RECT 652.930 2457.490 654.110 2458.670 ;
        RECT 652.930 2279.090 654.110 2280.270 ;
        RECT 652.930 2277.490 654.110 2278.670 ;
        RECT 652.930 2099.090 654.110 2100.270 ;
        RECT 652.930 2097.490 654.110 2098.670 ;
        RECT 652.930 1919.090 654.110 1920.270 ;
        RECT 652.930 1917.490 654.110 1918.670 ;
        RECT 652.930 1739.090 654.110 1740.270 ;
        RECT 652.930 1737.490 654.110 1738.670 ;
        RECT 652.930 1559.090 654.110 1560.270 ;
        RECT 652.930 1557.490 654.110 1558.670 ;
        RECT 652.930 1379.090 654.110 1380.270 ;
        RECT 652.930 1377.490 654.110 1378.670 ;
        RECT 652.930 1199.090 654.110 1200.270 ;
        RECT 652.930 1197.490 654.110 1198.670 ;
        RECT 652.930 1019.090 654.110 1020.270 ;
        RECT 652.930 1017.490 654.110 1018.670 ;
        RECT 652.930 839.090 654.110 840.270 ;
        RECT 652.930 837.490 654.110 838.670 ;
        RECT 652.930 659.090 654.110 660.270 ;
        RECT 652.930 657.490 654.110 658.670 ;
        RECT 652.930 479.090 654.110 480.270 ;
        RECT 652.930 477.490 654.110 478.670 ;
        RECT 652.930 299.090 654.110 300.270 ;
        RECT 652.930 297.490 654.110 298.670 ;
        RECT 652.930 119.090 654.110 120.270 ;
        RECT 652.930 117.490 654.110 118.670 ;
        RECT 652.930 -16.710 654.110 -15.530 ;
        RECT 652.930 -18.310 654.110 -17.130 ;
        RECT 832.930 3536.810 834.110 3537.990 ;
        RECT 832.930 3535.210 834.110 3536.390 ;
        RECT 832.930 3359.090 834.110 3360.270 ;
        RECT 832.930 3357.490 834.110 3358.670 ;
        RECT 832.930 3179.090 834.110 3180.270 ;
        RECT 832.930 3177.490 834.110 3178.670 ;
        RECT 832.930 2999.090 834.110 3000.270 ;
        RECT 832.930 2997.490 834.110 2998.670 ;
        RECT 832.930 2819.090 834.110 2820.270 ;
        RECT 832.930 2817.490 834.110 2818.670 ;
        RECT 832.930 2639.090 834.110 2640.270 ;
        RECT 832.930 2637.490 834.110 2638.670 ;
        RECT 832.930 2459.090 834.110 2460.270 ;
        RECT 832.930 2457.490 834.110 2458.670 ;
        RECT 832.930 2279.090 834.110 2280.270 ;
        RECT 832.930 2277.490 834.110 2278.670 ;
        RECT 832.930 2099.090 834.110 2100.270 ;
        RECT 832.930 2097.490 834.110 2098.670 ;
        RECT 832.930 1919.090 834.110 1920.270 ;
        RECT 832.930 1917.490 834.110 1918.670 ;
        RECT 832.930 1739.090 834.110 1740.270 ;
        RECT 832.930 1737.490 834.110 1738.670 ;
        RECT 832.930 1559.090 834.110 1560.270 ;
        RECT 832.930 1557.490 834.110 1558.670 ;
        RECT 832.930 1379.090 834.110 1380.270 ;
        RECT 832.930 1377.490 834.110 1378.670 ;
        RECT 832.930 1199.090 834.110 1200.270 ;
        RECT 832.930 1197.490 834.110 1198.670 ;
        RECT 832.930 1019.090 834.110 1020.270 ;
        RECT 832.930 1017.490 834.110 1018.670 ;
        RECT 832.930 839.090 834.110 840.270 ;
        RECT 832.930 837.490 834.110 838.670 ;
        RECT 832.930 659.090 834.110 660.270 ;
        RECT 832.930 657.490 834.110 658.670 ;
        RECT 832.930 479.090 834.110 480.270 ;
        RECT 832.930 477.490 834.110 478.670 ;
        RECT 832.930 299.090 834.110 300.270 ;
        RECT 832.930 297.490 834.110 298.670 ;
        RECT 832.930 119.090 834.110 120.270 ;
        RECT 832.930 117.490 834.110 118.670 ;
        RECT 832.930 -16.710 834.110 -15.530 ;
        RECT 832.930 -18.310 834.110 -17.130 ;
        RECT 1012.930 3536.810 1014.110 3537.990 ;
        RECT 1012.930 3535.210 1014.110 3536.390 ;
        RECT 1012.930 3359.090 1014.110 3360.270 ;
        RECT 1012.930 3357.490 1014.110 3358.670 ;
        RECT 1012.930 3179.090 1014.110 3180.270 ;
        RECT 1012.930 3177.490 1014.110 3178.670 ;
        RECT 1012.930 2999.090 1014.110 3000.270 ;
        RECT 1012.930 2997.490 1014.110 2998.670 ;
        RECT 1012.930 2819.090 1014.110 2820.270 ;
        RECT 1012.930 2817.490 1014.110 2818.670 ;
        RECT 1012.930 2639.090 1014.110 2640.270 ;
        RECT 1012.930 2637.490 1014.110 2638.670 ;
        RECT 1012.930 2459.090 1014.110 2460.270 ;
        RECT 1012.930 2457.490 1014.110 2458.670 ;
        RECT 1012.930 2279.090 1014.110 2280.270 ;
        RECT 1012.930 2277.490 1014.110 2278.670 ;
        RECT 1012.930 2099.090 1014.110 2100.270 ;
        RECT 1012.930 2097.490 1014.110 2098.670 ;
        RECT 1012.930 1919.090 1014.110 1920.270 ;
        RECT 1012.930 1917.490 1014.110 1918.670 ;
        RECT 1012.930 1739.090 1014.110 1740.270 ;
        RECT 1012.930 1737.490 1014.110 1738.670 ;
        RECT 1012.930 1559.090 1014.110 1560.270 ;
        RECT 1012.930 1557.490 1014.110 1558.670 ;
        RECT 1012.930 1379.090 1014.110 1380.270 ;
        RECT 1012.930 1377.490 1014.110 1378.670 ;
        RECT 1012.930 1199.090 1014.110 1200.270 ;
        RECT 1012.930 1197.490 1014.110 1198.670 ;
        RECT 1012.930 1019.090 1014.110 1020.270 ;
        RECT 1012.930 1017.490 1014.110 1018.670 ;
        RECT 1012.930 839.090 1014.110 840.270 ;
        RECT 1012.930 837.490 1014.110 838.670 ;
        RECT 1012.930 659.090 1014.110 660.270 ;
        RECT 1012.930 657.490 1014.110 658.670 ;
        RECT 1012.930 479.090 1014.110 480.270 ;
        RECT 1012.930 477.490 1014.110 478.670 ;
        RECT 1012.930 299.090 1014.110 300.270 ;
        RECT 1012.930 297.490 1014.110 298.670 ;
        RECT 1012.930 119.090 1014.110 120.270 ;
        RECT 1012.930 117.490 1014.110 118.670 ;
        RECT 1012.930 -16.710 1014.110 -15.530 ;
        RECT 1012.930 -18.310 1014.110 -17.130 ;
        RECT 1192.930 3536.810 1194.110 3537.990 ;
        RECT 1192.930 3535.210 1194.110 3536.390 ;
        RECT 1192.930 3359.090 1194.110 3360.270 ;
        RECT 1192.930 3357.490 1194.110 3358.670 ;
        RECT 1192.930 3179.090 1194.110 3180.270 ;
        RECT 1192.930 3177.490 1194.110 3178.670 ;
        RECT 1192.930 2999.090 1194.110 3000.270 ;
        RECT 1192.930 2997.490 1194.110 2998.670 ;
        RECT 1192.930 2819.090 1194.110 2820.270 ;
        RECT 1192.930 2817.490 1194.110 2818.670 ;
        RECT 1192.930 2639.090 1194.110 2640.270 ;
        RECT 1192.930 2637.490 1194.110 2638.670 ;
        RECT 1192.930 2459.090 1194.110 2460.270 ;
        RECT 1192.930 2457.490 1194.110 2458.670 ;
        RECT 1192.930 2279.090 1194.110 2280.270 ;
        RECT 1192.930 2277.490 1194.110 2278.670 ;
        RECT 1192.930 2099.090 1194.110 2100.270 ;
        RECT 1192.930 2097.490 1194.110 2098.670 ;
        RECT 1192.930 1919.090 1194.110 1920.270 ;
        RECT 1192.930 1917.490 1194.110 1918.670 ;
        RECT 1192.930 1739.090 1194.110 1740.270 ;
        RECT 1192.930 1737.490 1194.110 1738.670 ;
        RECT 1192.930 1559.090 1194.110 1560.270 ;
        RECT 1192.930 1557.490 1194.110 1558.670 ;
        RECT 1192.930 1379.090 1194.110 1380.270 ;
        RECT 1192.930 1377.490 1194.110 1378.670 ;
        RECT 1192.930 1199.090 1194.110 1200.270 ;
        RECT 1192.930 1197.490 1194.110 1198.670 ;
        RECT 1192.930 1019.090 1194.110 1020.270 ;
        RECT 1192.930 1017.490 1194.110 1018.670 ;
        RECT 1192.930 839.090 1194.110 840.270 ;
        RECT 1192.930 837.490 1194.110 838.670 ;
        RECT 1192.930 659.090 1194.110 660.270 ;
        RECT 1192.930 657.490 1194.110 658.670 ;
        RECT 1192.930 479.090 1194.110 480.270 ;
        RECT 1192.930 477.490 1194.110 478.670 ;
        RECT 1192.930 299.090 1194.110 300.270 ;
        RECT 1192.930 297.490 1194.110 298.670 ;
        RECT 1192.930 119.090 1194.110 120.270 ;
        RECT 1192.930 117.490 1194.110 118.670 ;
        RECT 1192.930 -16.710 1194.110 -15.530 ;
        RECT 1192.930 -18.310 1194.110 -17.130 ;
        RECT 1372.930 3536.810 1374.110 3537.990 ;
        RECT 1372.930 3535.210 1374.110 3536.390 ;
        RECT 1372.930 3359.090 1374.110 3360.270 ;
        RECT 1372.930 3357.490 1374.110 3358.670 ;
        RECT 1372.930 3179.090 1374.110 3180.270 ;
        RECT 1372.930 3177.490 1374.110 3178.670 ;
        RECT 1372.930 2999.090 1374.110 3000.270 ;
        RECT 1372.930 2997.490 1374.110 2998.670 ;
        RECT 1372.930 2819.090 1374.110 2820.270 ;
        RECT 1372.930 2817.490 1374.110 2818.670 ;
        RECT 1372.930 2639.090 1374.110 2640.270 ;
        RECT 1372.930 2637.490 1374.110 2638.670 ;
        RECT 1372.930 2459.090 1374.110 2460.270 ;
        RECT 1372.930 2457.490 1374.110 2458.670 ;
        RECT 1372.930 2279.090 1374.110 2280.270 ;
        RECT 1372.930 2277.490 1374.110 2278.670 ;
        RECT 1372.930 2099.090 1374.110 2100.270 ;
        RECT 1372.930 2097.490 1374.110 2098.670 ;
        RECT 1372.930 1919.090 1374.110 1920.270 ;
        RECT 1372.930 1917.490 1374.110 1918.670 ;
        RECT 1372.930 1739.090 1374.110 1740.270 ;
        RECT 1372.930 1737.490 1374.110 1738.670 ;
        RECT 1372.930 1559.090 1374.110 1560.270 ;
        RECT 1372.930 1557.490 1374.110 1558.670 ;
        RECT 1372.930 1379.090 1374.110 1380.270 ;
        RECT 1372.930 1377.490 1374.110 1378.670 ;
        RECT 1372.930 1199.090 1374.110 1200.270 ;
        RECT 1372.930 1197.490 1374.110 1198.670 ;
        RECT 1372.930 1019.090 1374.110 1020.270 ;
        RECT 1372.930 1017.490 1374.110 1018.670 ;
        RECT 1372.930 839.090 1374.110 840.270 ;
        RECT 1372.930 837.490 1374.110 838.670 ;
        RECT 1372.930 659.090 1374.110 660.270 ;
        RECT 1372.930 657.490 1374.110 658.670 ;
        RECT 1372.930 479.090 1374.110 480.270 ;
        RECT 1372.930 477.490 1374.110 478.670 ;
        RECT 1372.930 299.090 1374.110 300.270 ;
        RECT 1372.930 297.490 1374.110 298.670 ;
        RECT 1372.930 119.090 1374.110 120.270 ;
        RECT 1372.930 117.490 1374.110 118.670 ;
        RECT 1372.930 -16.710 1374.110 -15.530 ;
        RECT 1372.930 -18.310 1374.110 -17.130 ;
        RECT 1552.930 3536.810 1554.110 3537.990 ;
        RECT 1552.930 3535.210 1554.110 3536.390 ;
        RECT 1552.930 3359.090 1554.110 3360.270 ;
        RECT 1552.930 3357.490 1554.110 3358.670 ;
        RECT 1552.930 3179.090 1554.110 3180.270 ;
        RECT 1552.930 3177.490 1554.110 3178.670 ;
        RECT 1552.930 2999.090 1554.110 3000.270 ;
        RECT 1552.930 2997.490 1554.110 2998.670 ;
        RECT 1552.930 2819.090 1554.110 2820.270 ;
        RECT 1552.930 2817.490 1554.110 2818.670 ;
        RECT 1552.930 2639.090 1554.110 2640.270 ;
        RECT 1552.930 2637.490 1554.110 2638.670 ;
        RECT 1552.930 2459.090 1554.110 2460.270 ;
        RECT 1552.930 2457.490 1554.110 2458.670 ;
        RECT 1552.930 2279.090 1554.110 2280.270 ;
        RECT 1552.930 2277.490 1554.110 2278.670 ;
        RECT 1552.930 2099.090 1554.110 2100.270 ;
        RECT 1552.930 2097.490 1554.110 2098.670 ;
        RECT 1552.930 1919.090 1554.110 1920.270 ;
        RECT 1552.930 1917.490 1554.110 1918.670 ;
        RECT 1552.930 1739.090 1554.110 1740.270 ;
        RECT 1552.930 1737.490 1554.110 1738.670 ;
        RECT 1552.930 1559.090 1554.110 1560.270 ;
        RECT 1552.930 1557.490 1554.110 1558.670 ;
        RECT 1552.930 1379.090 1554.110 1380.270 ;
        RECT 1552.930 1377.490 1554.110 1378.670 ;
        RECT 1552.930 1199.090 1554.110 1200.270 ;
        RECT 1552.930 1197.490 1554.110 1198.670 ;
        RECT 1552.930 1019.090 1554.110 1020.270 ;
        RECT 1552.930 1017.490 1554.110 1018.670 ;
        RECT 1552.930 839.090 1554.110 840.270 ;
        RECT 1552.930 837.490 1554.110 838.670 ;
        RECT 1552.930 659.090 1554.110 660.270 ;
        RECT 1552.930 657.490 1554.110 658.670 ;
        RECT 1552.930 479.090 1554.110 480.270 ;
        RECT 1552.930 477.490 1554.110 478.670 ;
        RECT 1552.930 299.090 1554.110 300.270 ;
        RECT 1552.930 297.490 1554.110 298.670 ;
        RECT 1552.930 119.090 1554.110 120.270 ;
        RECT 1552.930 117.490 1554.110 118.670 ;
        RECT 1552.930 -16.710 1554.110 -15.530 ;
        RECT 1552.930 -18.310 1554.110 -17.130 ;
        RECT 1732.930 3536.810 1734.110 3537.990 ;
        RECT 1732.930 3535.210 1734.110 3536.390 ;
        RECT 1732.930 3359.090 1734.110 3360.270 ;
        RECT 1732.930 3357.490 1734.110 3358.670 ;
        RECT 1732.930 3179.090 1734.110 3180.270 ;
        RECT 1732.930 3177.490 1734.110 3178.670 ;
        RECT 1732.930 2999.090 1734.110 3000.270 ;
        RECT 1732.930 2997.490 1734.110 2998.670 ;
        RECT 1732.930 2819.090 1734.110 2820.270 ;
        RECT 1732.930 2817.490 1734.110 2818.670 ;
        RECT 1732.930 2639.090 1734.110 2640.270 ;
        RECT 1732.930 2637.490 1734.110 2638.670 ;
        RECT 1732.930 2459.090 1734.110 2460.270 ;
        RECT 1732.930 2457.490 1734.110 2458.670 ;
        RECT 1732.930 2279.090 1734.110 2280.270 ;
        RECT 1732.930 2277.490 1734.110 2278.670 ;
        RECT 1732.930 2099.090 1734.110 2100.270 ;
        RECT 1732.930 2097.490 1734.110 2098.670 ;
        RECT 1732.930 1919.090 1734.110 1920.270 ;
        RECT 1732.930 1917.490 1734.110 1918.670 ;
        RECT 1732.930 1739.090 1734.110 1740.270 ;
        RECT 1732.930 1737.490 1734.110 1738.670 ;
        RECT 1732.930 1559.090 1734.110 1560.270 ;
        RECT 1732.930 1557.490 1734.110 1558.670 ;
        RECT 1732.930 1379.090 1734.110 1380.270 ;
        RECT 1732.930 1377.490 1734.110 1378.670 ;
        RECT 1732.930 1199.090 1734.110 1200.270 ;
        RECT 1732.930 1197.490 1734.110 1198.670 ;
        RECT 1732.930 1019.090 1734.110 1020.270 ;
        RECT 1732.930 1017.490 1734.110 1018.670 ;
        RECT 1732.930 839.090 1734.110 840.270 ;
        RECT 1732.930 837.490 1734.110 838.670 ;
        RECT 1732.930 659.090 1734.110 660.270 ;
        RECT 1732.930 657.490 1734.110 658.670 ;
        RECT 1732.930 479.090 1734.110 480.270 ;
        RECT 1732.930 477.490 1734.110 478.670 ;
        RECT 1732.930 299.090 1734.110 300.270 ;
        RECT 1732.930 297.490 1734.110 298.670 ;
        RECT 1732.930 119.090 1734.110 120.270 ;
        RECT 1732.930 117.490 1734.110 118.670 ;
        RECT 1732.930 -16.710 1734.110 -15.530 ;
        RECT 1732.930 -18.310 1734.110 -17.130 ;
        RECT 1912.930 3536.810 1914.110 3537.990 ;
        RECT 1912.930 3535.210 1914.110 3536.390 ;
        RECT 1912.930 3359.090 1914.110 3360.270 ;
        RECT 1912.930 3357.490 1914.110 3358.670 ;
        RECT 1912.930 3179.090 1914.110 3180.270 ;
        RECT 1912.930 3177.490 1914.110 3178.670 ;
        RECT 1912.930 2999.090 1914.110 3000.270 ;
        RECT 1912.930 2997.490 1914.110 2998.670 ;
        RECT 1912.930 2819.090 1914.110 2820.270 ;
        RECT 1912.930 2817.490 1914.110 2818.670 ;
        RECT 1912.930 2639.090 1914.110 2640.270 ;
        RECT 1912.930 2637.490 1914.110 2638.670 ;
        RECT 1912.930 2459.090 1914.110 2460.270 ;
        RECT 1912.930 2457.490 1914.110 2458.670 ;
        RECT 1912.930 2279.090 1914.110 2280.270 ;
        RECT 1912.930 2277.490 1914.110 2278.670 ;
        RECT 1912.930 2099.090 1914.110 2100.270 ;
        RECT 1912.930 2097.490 1914.110 2098.670 ;
        RECT 1912.930 1919.090 1914.110 1920.270 ;
        RECT 1912.930 1917.490 1914.110 1918.670 ;
        RECT 1912.930 1739.090 1914.110 1740.270 ;
        RECT 1912.930 1737.490 1914.110 1738.670 ;
        RECT 1912.930 1559.090 1914.110 1560.270 ;
        RECT 1912.930 1557.490 1914.110 1558.670 ;
        RECT 1912.930 1379.090 1914.110 1380.270 ;
        RECT 1912.930 1377.490 1914.110 1378.670 ;
        RECT 1912.930 1199.090 1914.110 1200.270 ;
        RECT 1912.930 1197.490 1914.110 1198.670 ;
        RECT 1912.930 1019.090 1914.110 1020.270 ;
        RECT 1912.930 1017.490 1914.110 1018.670 ;
        RECT 1912.930 839.090 1914.110 840.270 ;
        RECT 1912.930 837.490 1914.110 838.670 ;
        RECT 1912.930 659.090 1914.110 660.270 ;
        RECT 1912.930 657.490 1914.110 658.670 ;
        RECT 1912.930 479.090 1914.110 480.270 ;
        RECT 1912.930 477.490 1914.110 478.670 ;
        RECT 1912.930 299.090 1914.110 300.270 ;
        RECT 1912.930 297.490 1914.110 298.670 ;
        RECT 1912.930 119.090 1914.110 120.270 ;
        RECT 1912.930 117.490 1914.110 118.670 ;
        RECT 1912.930 -16.710 1914.110 -15.530 ;
        RECT 1912.930 -18.310 1914.110 -17.130 ;
        RECT 2092.930 3536.810 2094.110 3537.990 ;
        RECT 2092.930 3535.210 2094.110 3536.390 ;
        RECT 2092.930 3359.090 2094.110 3360.270 ;
        RECT 2092.930 3357.490 2094.110 3358.670 ;
        RECT 2092.930 3179.090 2094.110 3180.270 ;
        RECT 2092.930 3177.490 2094.110 3178.670 ;
        RECT 2092.930 2999.090 2094.110 3000.270 ;
        RECT 2092.930 2997.490 2094.110 2998.670 ;
        RECT 2092.930 2819.090 2094.110 2820.270 ;
        RECT 2092.930 2817.490 2094.110 2818.670 ;
        RECT 2092.930 2639.090 2094.110 2640.270 ;
        RECT 2092.930 2637.490 2094.110 2638.670 ;
        RECT 2092.930 2459.090 2094.110 2460.270 ;
        RECT 2092.930 2457.490 2094.110 2458.670 ;
        RECT 2092.930 2279.090 2094.110 2280.270 ;
        RECT 2092.930 2277.490 2094.110 2278.670 ;
        RECT 2092.930 2099.090 2094.110 2100.270 ;
        RECT 2092.930 2097.490 2094.110 2098.670 ;
        RECT 2092.930 1919.090 2094.110 1920.270 ;
        RECT 2092.930 1917.490 2094.110 1918.670 ;
        RECT 2092.930 1739.090 2094.110 1740.270 ;
        RECT 2092.930 1737.490 2094.110 1738.670 ;
        RECT 2092.930 1559.090 2094.110 1560.270 ;
        RECT 2092.930 1557.490 2094.110 1558.670 ;
        RECT 2092.930 1379.090 2094.110 1380.270 ;
        RECT 2092.930 1377.490 2094.110 1378.670 ;
        RECT 2092.930 1199.090 2094.110 1200.270 ;
        RECT 2092.930 1197.490 2094.110 1198.670 ;
        RECT 2092.930 1019.090 2094.110 1020.270 ;
        RECT 2092.930 1017.490 2094.110 1018.670 ;
        RECT 2092.930 839.090 2094.110 840.270 ;
        RECT 2092.930 837.490 2094.110 838.670 ;
        RECT 2092.930 659.090 2094.110 660.270 ;
        RECT 2092.930 657.490 2094.110 658.670 ;
        RECT 2092.930 479.090 2094.110 480.270 ;
        RECT 2092.930 477.490 2094.110 478.670 ;
        RECT 2092.930 299.090 2094.110 300.270 ;
        RECT 2092.930 297.490 2094.110 298.670 ;
        RECT 2092.930 119.090 2094.110 120.270 ;
        RECT 2092.930 117.490 2094.110 118.670 ;
        RECT 2092.930 -16.710 2094.110 -15.530 ;
        RECT 2092.930 -18.310 2094.110 -17.130 ;
        RECT 2272.930 3536.810 2274.110 3537.990 ;
        RECT 2272.930 3535.210 2274.110 3536.390 ;
        RECT 2272.930 3359.090 2274.110 3360.270 ;
        RECT 2272.930 3357.490 2274.110 3358.670 ;
        RECT 2272.930 3179.090 2274.110 3180.270 ;
        RECT 2272.930 3177.490 2274.110 3178.670 ;
        RECT 2272.930 2999.090 2274.110 3000.270 ;
        RECT 2272.930 2997.490 2274.110 2998.670 ;
        RECT 2272.930 2819.090 2274.110 2820.270 ;
        RECT 2272.930 2817.490 2274.110 2818.670 ;
        RECT 2272.930 2639.090 2274.110 2640.270 ;
        RECT 2272.930 2637.490 2274.110 2638.670 ;
        RECT 2272.930 2459.090 2274.110 2460.270 ;
        RECT 2272.930 2457.490 2274.110 2458.670 ;
        RECT 2272.930 2279.090 2274.110 2280.270 ;
        RECT 2272.930 2277.490 2274.110 2278.670 ;
        RECT 2272.930 2099.090 2274.110 2100.270 ;
        RECT 2272.930 2097.490 2274.110 2098.670 ;
        RECT 2272.930 1919.090 2274.110 1920.270 ;
        RECT 2272.930 1917.490 2274.110 1918.670 ;
        RECT 2272.930 1739.090 2274.110 1740.270 ;
        RECT 2272.930 1737.490 2274.110 1738.670 ;
        RECT 2272.930 1559.090 2274.110 1560.270 ;
        RECT 2272.930 1557.490 2274.110 1558.670 ;
        RECT 2272.930 1379.090 2274.110 1380.270 ;
        RECT 2272.930 1377.490 2274.110 1378.670 ;
        RECT 2272.930 1199.090 2274.110 1200.270 ;
        RECT 2272.930 1197.490 2274.110 1198.670 ;
        RECT 2272.930 1019.090 2274.110 1020.270 ;
        RECT 2272.930 1017.490 2274.110 1018.670 ;
        RECT 2272.930 839.090 2274.110 840.270 ;
        RECT 2272.930 837.490 2274.110 838.670 ;
        RECT 2272.930 659.090 2274.110 660.270 ;
        RECT 2272.930 657.490 2274.110 658.670 ;
        RECT 2272.930 479.090 2274.110 480.270 ;
        RECT 2272.930 477.490 2274.110 478.670 ;
        RECT 2272.930 299.090 2274.110 300.270 ;
        RECT 2272.930 297.490 2274.110 298.670 ;
        RECT 2272.930 119.090 2274.110 120.270 ;
        RECT 2272.930 117.490 2274.110 118.670 ;
        RECT 2272.930 -16.710 2274.110 -15.530 ;
        RECT 2272.930 -18.310 2274.110 -17.130 ;
        RECT 2452.930 3536.810 2454.110 3537.990 ;
        RECT 2452.930 3535.210 2454.110 3536.390 ;
        RECT 2452.930 3359.090 2454.110 3360.270 ;
        RECT 2452.930 3357.490 2454.110 3358.670 ;
        RECT 2452.930 3179.090 2454.110 3180.270 ;
        RECT 2452.930 3177.490 2454.110 3178.670 ;
        RECT 2452.930 2999.090 2454.110 3000.270 ;
        RECT 2452.930 2997.490 2454.110 2998.670 ;
        RECT 2452.930 2819.090 2454.110 2820.270 ;
        RECT 2452.930 2817.490 2454.110 2818.670 ;
        RECT 2452.930 2639.090 2454.110 2640.270 ;
        RECT 2452.930 2637.490 2454.110 2638.670 ;
        RECT 2452.930 2459.090 2454.110 2460.270 ;
        RECT 2452.930 2457.490 2454.110 2458.670 ;
        RECT 2452.930 2279.090 2454.110 2280.270 ;
        RECT 2452.930 2277.490 2454.110 2278.670 ;
        RECT 2452.930 2099.090 2454.110 2100.270 ;
        RECT 2452.930 2097.490 2454.110 2098.670 ;
        RECT 2452.930 1919.090 2454.110 1920.270 ;
        RECT 2452.930 1917.490 2454.110 1918.670 ;
        RECT 2452.930 1739.090 2454.110 1740.270 ;
        RECT 2452.930 1737.490 2454.110 1738.670 ;
        RECT 2452.930 1559.090 2454.110 1560.270 ;
        RECT 2452.930 1557.490 2454.110 1558.670 ;
        RECT 2452.930 1379.090 2454.110 1380.270 ;
        RECT 2452.930 1377.490 2454.110 1378.670 ;
        RECT 2452.930 1199.090 2454.110 1200.270 ;
        RECT 2452.930 1197.490 2454.110 1198.670 ;
        RECT 2452.930 1019.090 2454.110 1020.270 ;
        RECT 2452.930 1017.490 2454.110 1018.670 ;
        RECT 2452.930 839.090 2454.110 840.270 ;
        RECT 2452.930 837.490 2454.110 838.670 ;
        RECT 2452.930 659.090 2454.110 660.270 ;
        RECT 2452.930 657.490 2454.110 658.670 ;
        RECT 2452.930 479.090 2454.110 480.270 ;
        RECT 2452.930 477.490 2454.110 478.670 ;
        RECT 2452.930 299.090 2454.110 300.270 ;
        RECT 2452.930 297.490 2454.110 298.670 ;
        RECT 2452.930 119.090 2454.110 120.270 ;
        RECT 2452.930 117.490 2454.110 118.670 ;
        RECT 2452.930 -16.710 2454.110 -15.530 ;
        RECT 2452.930 -18.310 2454.110 -17.130 ;
        RECT 2632.930 3536.810 2634.110 3537.990 ;
        RECT 2632.930 3535.210 2634.110 3536.390 ;
        RECT 2632.930 3359.090 2634.110 3360.270 ;
        RECT 2632.930 3357.490 2634.110 3358.670 ;
        RECT 2632.930 3179.090 2634.110 3180.270 ;
        RECT 2632.930 3177.490 2634.110 3178.670 ;
        RECT 2632.930 2999.090 2634.110 3000.270 ;
        RECT 2632.930 2997.490 2634.110 2998.670 ;
        RECT 2632.930 2819.090 2634.110 2820.270 ;
        RECT 2632.930 2817.490 2634.110 2818.670 ;
        RECT 2632.930 2639.090 2634.110 2640.270 ;
        RECT 2632.930 2637.490 2634.110 2638.670 ;
        RECT 2632.930 2459.090 2634.110 2460.270 ;
        RECT 2632.930 2457.490 2634.110 2458.670 ;
        RECT 2632.930 2279.090 2634.110 2280.270 ;
        RECT 2632.930 2277.490 2634.110 2278.670 ;
        RECT 2632.930 2099.090 2634.110 2100.270 ;
        RECT 2632.930 2097.490 2634.110 2098.670 ;
        RECT 2632.930 1919.090 2634.110 1920.270 ;
        RECT 2632.930 1917.490 2634.110 1918.670 ;
        RECT 2632.930 1739.090 2634.110 1740.270 ;
        RECT 2632.930 1737.490 2634.110 1738.670 ;
        RECT 2632.930 1559.090 2634.110 1560.270 ;
        RECT 2632.930 1557.490 2634.110 1558.670 ;
        RECT 2632.930 1379.090 2634.110 1380.270 ;
        RECT 2632.930 1377.490 2634.110 1378.670 ;
        RECT 2632.930 1199.090 2634.110 1200.270 ;
        RECT 2632.930 1197.490 2634.110 1198.670 ;
        RECT 2632.930 1019.090 2634.110 1020.270 ;
        RECT 2632.930 1017.490 2634.110 1018.670 ;
        RECT 2632.930 839.090 2634.110 840.270 ;
        RECT 2632.930 837.490 2634.110 838.670 ;
        RECT 2632.930 659.090 2634.110 660.270 ;
        RECT 2632.930 657.490 2634.110 658.670 ;
        RECT 2632.930 479.090 2634.110 480.270 ;
        RECT 2632.930 477.490 2634.110 478.670 ;
        RECT 2632.930 299.090 2634.110 300.270 ;
        RECT 2632.930 297.490 2634.110 298.670 ;
        RECT 2632.930 119.090 2634.110 120.270 ;
        RECT 2632.930 117.490 2634.110 118.670 ;
        RECT 2632.930 -16.710 2634.110 -15.530 ;
        RECT 2632.930 -18.310 2634.110 -17.130 ;
        RECT 2812.930 3536.810 2814.110 3537.990 ;
        RECT 2812.930 3535.210 2814.110 3536.390 ;
        RECT 2812.930 3359.090 2814.110 3360.270 ;
        RECT 2812.930 3357.490 2814.110 3358.670 ;
        RECT 2812.930 3179.090 2814.110 3180.270 ;
        RECT 2812.930 3177.490 2814.110 3178.670 ;
        RECT 2812.930 2999.090 2814.110 3000.270 ;
        RECT 2812.930 2997.490 2814.110 2998.670 ;
        RECT 2812.930 2819.090 2814.110 2820.270 ;
        RECT 2812.930 2817.490 2814.110 2818.670 ;
        RECT 2812.930 2639.090 2814.110 2640.270 ;
        RECT 2812.930 2637.490 2814.110 2638.670 ;
        RECT 2812.930 2459.090 2814.110 2460.270 ;
        RECT 2812.930 2457.490 2814.110 2458.670 ;
        RECT 2812.930 2279.090 2814.110 2280.270 ;
        RECT 2812.930 2277.490 2814.110 2278.670 ;
        RECT 2812.930 2099.090 2814.110 2100.270 ;
        RECT 2812.930 2097.490 2814.110 2098.670 ;
        RECT 2812.930 1919.090 2814.110 1920.270 ;
        RECT 2812.930 1917.490 2814.110 1918.670 ;
        RECT 2812.930 1739.090 2814.110 1740.270 ;
        RECT 2812.930 1737.490 2814.110 1738.670 ;
        RECT 2812.930 1559.090 2814.110 1560.270 ;
        RECT 2812.930 1557.490 2814.110 1558.670 ;
        RECT 2812.930 1379.090 2814.110 1380.270 ;
        RECT 2812.930 1377.490 2814.110 1378.670 ;
        RECT 2812.930 1199.090 2814.110 1200.270 ;
        RECT 2812.930 1197.490 2814.110 1198.670 ;
        RECT 2812.930 1019.090 2814.110 1020.270 ;
        RECT 2812.930 1017.490 2814.110 1018.670 ;
        RECT 2812.930 839.090 2814.110 840.270 ;
        RECT 2812.930 837.490 2814.110 838.670 ;
        RECT 2812.930 659.090 2814.110 660.270 ;
        RECT 2812.930 657.490 2814.110 658.670 ;
        RECT 2812.930 479.090 2814.110 480.270 ;
        RECT 2812.930 477.490 2814.110 478.670 ;
        RECT 2812.930 299.090 2814.110 300.270 ;
        RECT 2812.930 297.490 2814.110 298.670 ;
        RECT 2812.930 119.090 2814.110 120.270 ;
        RECT 2812.930 117.490 2814.110 118.670 ;
        RECT 2812.930 -16.710 2814.110 -15.530 ;
        RECT 2812.930 -18.310 2814.110 -17.130 ;
        RECT 2941.310 3536.810 2942.490 3537.990 ;
        RECT 2941.310 3535.210 2942.490 3536.390 ;
        RECT 2941.310 3359.090 2942.490 3360.270 ;
        RECT 2941.310 3357.490 2942.490 3358.670 ;
        RECT 2941.310 3179.090 2942.490 3180.270 ;
        RECT 2941.310 3177.490 2942.490 3178.670 ;
        RECT 2941.310 2999.090 2942.490 3000.270 ;
        RECT 2941.310 2997.490 2942.490 2998.670 ;
        RECT 2941.310 2819.090 2942.490 2820.270 ;
        RECT 2941.310 2817.490 2942.490 2818.670 ;
        RECT 2941.310 2639.090 2942.490 2640.270 ;
        RECT 2941.310 2637.490 2942.490 2638.670 ;
        RECT 2941.310 2459.090 2942.490 2460.270 ;
        RECT 2941.310 2457.490 2942.490 2458.670 ;
        RECT 2941.310 2279.090 2942.490 2280.270 ;
        RECT 2941.310 2277.490 2942.490 2278.670 ;
        RECT 2941.310 2099.090 2942.490 2100.270 ;
        RECT 2941.310 2097.490 2942.490 2098.670 ;
        RECT 2941.310 1919.090 2942.490 1920.270 ;
        RECT 2941.310 1917.490 2942.490 1918.670 ;
        RECT 2941.310 1739.090 2942.490 1740.270 ;
        RECT 2941.310 1737.490 2942.490 1738.670 ;
        RECT 2941.310 1559.090 2942.490 1560.270 ;
        RECT 2941.310 1557.490 2942.490 1558.670 ;
        RECT 2941.310 1379.090 2942.490 1380.270 ;
        RECT 2941.310 1377.490 2942.490 1378.670 ;
        RECT 2941.310 1199.090 2942.490 1200.270 ;
        RECT 2941.310 1197.490 2942.490 1198.670 ;
        RECT 2941.310 1019.090 2942.490 1020.270 ;
        RECT 2941.310 1017.490 2942.490 1018.670 ;
        RECT 2941.310 839.090 2942.490 840.270 ;
        RECT 2941.310 837.490 2942.490 838.670 ;
        RECT 2941.310 659.090 2942.490 660.270 ;
        RECT 2941.310 657.490 2942.490 658.670 ;
        RECT 2941.310 479.090 2942.490 480.270 ;
        RECT 2941.310 477.490 2942.490 478.670 ;
        RECT 2941.310 299.090 2942.490 300.270 ;
        RECT 2941.310 297.490 2942.490 298.670 ;
        RECT 2941.310 119.090 2942.490 120.270 ;
        RECT 2941.310 117.490 2942.490 118.670 ;
        RECT 2941.310 -16.710 2942.490 -15.530 ;
        RECT 2941.310 -18.310 2942.490 -17.130 ;
      LAYER met5 ;
        RECT -23.780 3538.100 -20.780 3538.110 ;
        RECT 112.020 3538.100 115.020 3538.110 ;
        RECT 292.020 3538.100 295.020 3538.110 ;
        RECT 472.020 3538.100 475.020 3538.110 ;
        RECT 652.020 3538.100 655.020 3538.110 ;
        RECT 832.020 3538.100 835.020 3538.110 ;
        RECT 1012.020 3538.100 1015.020 3538.110 ;
        RECT 1192.020 3538.100 1195.020 3538.110 ;
        RECT 1372.020 3538.100 1375.020 3538.110 ;
        RECT 1552.020 3538.100 1555.020 3538.110 ;
        RECT 1732.020 3538.100 1735.020 3538.110 ;
        RECT 1912.020 3538.100 1915.020 3538.110 ;
        RECT 2092.020 3538.100 2095.020 3538.110 ;
        RECT 2272.020 3538.100 2275.020 3538.110 ;
        RECT 2452.020 3538.100 2455.020 3538.110 ;
        RECT 2632.020 3538.100 2635.020 3538.110 ;
        RECT 2812.020 3538.100 2815.020 3538.110 ;
        RECT 2940.400 3538.100 2943.400 3538.110 ;
        RECT -23.780 3535.100 2943.400 3538.100 ;
        RECT -23.780 3535.090 -20.780 3535.100 ;
        RECT 112.020 3535.090 115.020 3535.100 ;
        RECT 292.020 3535.090 295.020 3535.100 ;
        RECT 472.020 3535.090 475.020 3535.100 ;
        RECT 652.020 3535.090 655.020 3535.100 ;
        RECT 832.020 3535.090 835.020 3535.100 ;
        RECT 1012.020 3535.090 1015.020 3535.100 ;
        RECT 1192.020 3535.090 1195.020 3535.100 ;
        RECT 1372.020 3535.090 1375.020 3535.100 ;
        RECT 1552.020 3535.090 1555.020 3535.100 ;
        RECT 1732.020 3535.090 1735.020 3535.100 ;
        RECT 1912.020 3535.090 1915.020 3535.100 ;
        RECT 2092.020 3535.090 2095.020 3535.100 ;
        RECT 2272.020 3535.090 2275.020 3535.100 ;
        RECT 2452.020 3535.090 2455.020 3535.100 ;
        RECT 2632.020 3535.090 2635.020 3535.100 ;
        RECT 2812.020 3535.090 2815.020 3535.100 ;
        RECT 2940.400 3535.090 2943.400 3535.100 ;
        RECT -23.780 3360.380 -20.780 3360.390 ;
        RECT 112.020 3360.380 115.020 3360.390 ;
        RECT 292.020 3360.380 295.020 3360.390 ;
        RECT 472.020 3360.380 475.020 3360.390 ;
        RECT 652.020 3360.380 655.020 3360.390 ;
        RECT 832.020 3360.380 835.020 3360.390 ;
        RECT 1012.020 3360.380 1015.020 3360.390 ;
        RECT 1192.020 3360.380 1195.020 3360.390 ;
        RECT 1372.020 3360.380 1375.020 3360.390 ;
        RECT 1552.020 3360.380 1555.020 3360.390 ;
        RECT 1732.020 3360.380 1735.020 3360.390 ;
        RECT 1912.020 3360.380 1915.020 3360.390 ;
        RECT 2092.020 3360.380 2095.020 3360.390 ;
        RECT 2272.020 3360.380 2275.020 3360.390 ;
        RECT 2452.020 3360.380 2455.020 3360.390 ;
        RECT 2632.020 3360.380 2635.020 3360.390 ;
        RECT 2812.020 3360.380 2815.020 3360.390 ;
        RECT 2940.400 3360.380 2943.400 3360.390 ;
        RECT -23.780 3357.380 2943.400 3360.380 ;
        RECT -23.780 3357.370 -20.780 3357.380 ;
        RECT 112.020 3357.370 115.020 3357.380 ;
        RECT 292.020 3357.370 295.020 3357.380 ;
        RECT 472.020 3357.370 475.020 3357.380 ;
        RECT 652.020 3357.370 655.020 3357.380 ;
        RECT 832.020 3357.370 835.020 3357.380 ;
        RECT 1012.020 3357.370 1015.020 3357.380 ;
        RECT 1192.020 3357.370 1195.020 3357.380 ;
        RECT 1372.020 3357.370 1375.020 3357.380 ;
        RECT 1552.020 3357.370 1555.020 3357.380 ;
        RECT 1732.020 3357.370 1735.020 3357.380 ;
        RECT 1912.020 3357.370 1915.020 3357.380 ;
        RECT 2092.020 3357.370 2095.020 3357.380 ;
        RECT 2272.020 3357.370 2275.020 3357.380 ;
        RECT 2452.020 3357.370 2455.020 3357.380 ;
        RECT 2632.020 3357.370 2635.020 3357.380 ;
        RECT 2812.020 3357.370 2815.020 3357.380 ;
        RECT 2940.400 3357.370 2943.400 3357.380 ;
        RECT -23.780 3180.380 -20.780 3180.390 ;
        RECT 112.020 3180.380 115.020 3180.390 ;
        RECT 292.020 3180.380 295.020 3180.390 ;
        RECT 472.020 3180.380 475.020 3180.390 ;
        RECT 652.020 3180.380 655.020 3180.390 ;
        RECT 832.020 3180.380 835.020 3180.390 ;
        RECT 1012.020 3180.380 1015.020 3180.390 ;
        RECT 1192.020 3180.380 1195.020 3180.390 ;
        RECT 1372.020 3180.380 1375.020 3180.390 ;
        RECT 1552.020 3180.380 1555.020 3180.390 ;
        RECT 1732.020 3180.380 1735.020 3180.390 ;
        RECT 1912.020 3180.380 1915.020 3180.390 ;
        RECT 2092.020 3180.380 2095.020 3180.390 ;
        RECT 2272.020 3180.380 2275.020 3180.390 ;
        RECT 2452.020 3180.380 2455.020 3180.390 ;
        RECT 2632.020 3180.380 2635.020 3180.390 ;
        RECT 2812.020 3180.380 2815.020 3180.390 ;
        RECT 2940.400 3180.380 2943.400 3180.390 ;
        RECT -23.780 3177.380 2943.400 3180.380 ;
        RECT -23.780 3177.370 -20.780 3177.380 ;
        RECT 112.020 3177.370 115.020 3177.380 ;
        RECT 292.020 3177.370 295.020 3177.380 ;
        RECT 472.020 3177.370 475.020 3177.380 ;
        RECT 652.020 3177.370 655.020 3177.380 ;
        RECT 832.020 3177.370 835.020 3177.380 ;
        RECT 1012.020 3177.370 1015.020 3177.380 ;
        RECT 1192.020 3177.370 1195.020 3177.380 ;
        RECT 1372.020 3177.370 1375.020 3177.380 ;
        RECT 1552.020 3177.370 1555.020 3177.380 ;
        RECT 1732.020 3177.370 1735.020 3177.380 ;
        RECT 1912.020 3177.370 1915.020 3177.380 ;
        RECT 2092.020 3177.370 2095.020 3177.380 ;
        RECT 2272.020 3177.370 2275.020 3177.380 ;
        RECT 2452.020 3177.370 2455.020 3177.380 ;
        RECT 2632.020 3177.370 2635.020 3177.380 ;
        RECT 2812.020 3177.370 2815.020 3177.380 ;
        RECT 2940.400 3177.370 2943.400 3177.380 ;
        RECT -23.780 3000.380 -20.780 3000.390 ;
        RECT 112.020 3000.380 115.020 3000.390 ;
        RECT 292.020 3000.380 295.020 3000.390 ;
        RECT 472.020 3000.380 475.020 3000.390 ;
        RECT 652.020 3000.380 655.020 3000.390 ;
        RECT 832.020 3000.380 835.020 3000.390 ;
        RECT 1012.020 3000.380 1015.020 3000.390 ;
        RECT 1192.020 3000.380 1195.020 3000.390 ;
        RECT 1372.020 3000.380 1375.020 3000.390 ;
        RECT 1552.020 3000.380 1555.020 3000.390 ;
        RECT 1732.020 3000.380 1735.020 3000.390 ;
        RECT 1912.020 3000.380 1915.020 3000.390 ;
        RECT 2092.020 3000.380 2095.020 3000.390 ;
        RECT 2272.020 3000.380 2275.020 3000.390 ;
        RECT 2452.020 3000.380 2455.020 3000.390 ;
        RECT 2632.020 3000.380 2635.020 3000.390 ;
        RECT 2812.020 3000.380 2815.020 3000.390 ;
        RECT 2940.400 3000.380 2943.400 3000.390 ;
        RECT -23.780 2997.380 2943.400 3000.380 ;
        RECT -23.780 2997.370 -20.780 2997.380 ;
        RECT 112.020 2997.370 115.020 2997.380 ;
        RECT 292.020 2997.370 295.020 2997.380 ;
        RECT 472.020 2997.370 475.020 2997.380 ;
        RECT 652.020 2997.370 655.020 2997.380 ;
        RECT 832.020 2997.370 835.020 2997.380 ;
        RECT 1012.020 2997.370 1015.020 2997.380 ;
        RECT 1192.020 2997.370 1195.020 2997.380 ;
        RECT 1372.020 2997.370 1375.020 2997.380 ;
        RECT 1552.020 2997.370 1555.020 2997.380 ;
        RECT 1732.020 2997.370 1735.020 2997.380 ;
        RECT 1912.020 2997.370 1915.020 2997.380 ;
        RECT 2092.020 2997.370 2095.020 2997.380 ;
        RECT 2272.020 2997.370 2275.020 2997.380 ;
        RECT 2452.020 2997.370 2455.020 2997.380 ;
        RECT 2632.020 2997.370 2635.020 2997.380 ;
        RECT 2812.020 2997.370 2815.020 2997.380 ;
        RECT 2940.400 2997.370 2943.400 2997.380 ;
        RECT -23.780 2820.380 -20.780 2820.390 ;
        RECT 112.020 2820.380 115.020 2820.390 ;
        RECT 292.020 2820.380 295.020 2820.390 ;
        RECT 472.020 2820.380 475.020 2820.390 ;
        RECT 652.020 2820.380 655.020 2820.390 ;
        RECT 832.020 2820.380 835.020 2820.390 ;
        RECT 1012.020 2820.380 1015.020 2820.390 ;
        RECT 1192.020 2820.380 1195.020 2820.390 ;
        RECT 1372.020 2820.380 1375.020 2820.390 ;
        RECT 1552.020 2820.380 1555.020 2820.390 ;
        RECT 1732.020 2820.380 1735.020 2820.390 ;
        RECT 1912.020 2820.380 1915.020 2820.390 ;
        RECT 2092.020 2820.380 2095.020 2820.390 ;
        RECT 2272.020 2820.380 2275.020 2820.390 ;
        RECT 2452.020 2820.380 2455.020 2820.390 ;
        RECT 2632.020 2820.380 2635.020 2820.390 ;
        RECT 2812.020 2820.380 2815.020 2820.390 ;
        RECT 2940.400 2820.380 2943.400 2820.390 ;
        RECT -23.780 2817.380 2943.400 2820.380 ;
        RECT -23.780 2817.370 -20.780 2817.380 ;
        RECT 112.020 2817.370 115.020 2817.380 ;
        RECT 292.020 2817.370 295.020 2817.380 ;
        RECT 472.020 2817.370 475.020 2817.380 ;
        RECT 652.020 2817.370 655.020 2817.380 ;
        RECT 832.020 2817.370 835.020 2817.380 ;
        RECT 1012.020 2817.370 1015.020 2817.380 ;
        RECT 1192.020 2817.370 1195.020 2817.380 ;
        RECT 1372.020 2817.370 1375.020 2817.380 ;
        RECT 1552.020 2817.370 1555.020 2817.380 ;
        RECT 1732.020 2817.370 1735.020 2817.380 ;
        RECT 1912.020 2817.370 1915.020 2817.380 ;
        RECT 2092.020 2817.370 2095.020 2817.380 ;
        RECT 2272.020 2817.370 2275.020 2817.380 ;
        RECT 2452.020 2817.370 2455.020 2817.380 ;
        RECT 2632.020 2817.370 2635.020 2817.380 ;
        RECT 2812.020 2817.370 2815.020 2817.380 ;
        RECT 2940.400 2817.370 2943.400 2817.380 ;
        RECT -23.780 2640.380 -20.780 2640.390 ;
        RECT 112.020 2640.380 115.020 2640.390 ;
        RECT 292.020 2640.380 295.020 2640.390 ;
        RECT 472.020 2640.380 475.020 2640.390 ;
        RECT 652.020 2640.380 655.020 2640.390 ;
        RECT 832.020 2640.380 835.020 2640.390 ;
        RECT 1012.020 2640.380 1015.020 2640.390 ;
        RECT 1192.020 2640.380 1195.020 2640.390 ;
        RECT 1372.020 2640.380 1375.020 2640.390 ;
        RECT 1552.020 2640.380 1555.020 2640.390 ;
        RECT 1732.020 2640.380 1735.020 2640.390 ;
        RECT 1912.020 2640.380 1915.020 2640.390 ;
        RECT 2092.020 2640.380 2095.020 2640.390 ;
        RECT 2272.020 2640.380 2275.020 2640.390 ;
        RECT 2452.020 2640.380 2455.020 2640.390 ;
        RECT 2632.020 2640.380 2635.020 2640.390 ;
        RECT 2812.020 2640.380 2815.020 2640.390 ;
        RECT 2940.400 2640.380 2943.400 2640.390 ;
        RECT -23.780 2637.380 2943.400 2640.380 ;
        RECT -23.780 2637.370 -20.780 2637.380 ;
        RECT 112.020 2637.370 115.020 2637.380 ;
        RECT 292.020 2637.370 295.020 2637.380 ;
        RECT 472.020 2637.370 475.020 2637.380 ;
        RECT 652.020 2637.370 655.020 2637.380 ;
        RECT 832.020 2637.370 835.020 2637.380 ;
        RECT 1012.020 2637.370 1015.020 2637.380 ;
        RECT 1192.020 2637.370 1195.020 2637.380 ;
        RECT 1372.020 2637.370 1375.020 2637.380 ;
        RECT 1552.020 2637.370 1555.020 2637.380 ;
        RECT 1732.020 2637.370 1735.020 2637.380 ;
        RECT 1912.020 2637.370 1915.020 2637.380 ;
        RECT 2092.020 2637.370 2095.020 2637.380 ;
        RECT 2272.020 2637.370 2275.020 2637.380 ;
        RECT 2452.020 2637.370 2455.020 2637.380 ;
        RECT 2632.020 2637.370 2635.020 2637.380 ;
        RECT 2812.020 2637.370 2815.020 2637.380 ;
        RECT 2940.400 2637.370 2943.400 2637.380 ;
        RECT -23.780 2460.380 -20.780 2460.390 ;
        RECT 112.020 2460.380 115.020 2460.390 ;
        RECT 292.020 2460.380 295.020 2460.390 ;
        RECT 472.020 2460.380 475.020 2460.390 ;
        RECT 652.020 2460.380 655.020 2460.390 ;
        RECT 832.020 2460.380 835.020 2460.390 ;
        RECT 1012.020 2460.380 1015.020 2460.390 ;
        RECT 1192.020 2460.380 1195.020 2460.390 ;
        RECT 1372.020 2460.380 1375.020 2460.390 ;
        RECT 1552.020 2460.380 1555.020 2460.390 ;
        RECT 1732.020 2460.380 1735.020 2460.390 ;
        RECT 1912.020 2460.380 1915.020 2460.390 ;
        RECT 2092.020 2460.380 2095.020 2460.390 ;
        RECT 2272.020 2460.380 2275.020 2460.390 ;
        RECT 2452.020 2460.380 2455.020 2460.390 ;
        RECT 2632.020 2460.380 2635.020 2460.390 ;
        RECT 2812.020 2460.380 2815.020 2460.390 ;
        RECT 2940.400 2460.380 2943.400 2460.390 ;
        RECT -23.780 2457.380 2943.400 2460.380 ;
        RECT -23.780 2457.370 -20.780 2457.380 ;
        RECT 112.020 2457.370 115.020 2457.380 ;
        RECT 292.020 2457.370 295.020 2457.380 ;
        RECT 472.020 2457.370 475.020 2457.380 ;
        RECT 652.020 2457.370 655.020 2457.380 ;
        RECT 832.020 2457.370 835.020 2457.380 ;
        RECT 1012.020 2457.370 1015.020 2457.380 ;
        RECT 1192.020 2457.370 1195.020 2457.380 ;
        RECT 1372.020 2457.370 1375.020 2457.380 ;
        RECT 1552.020 2457.370 1555.020 2457.380 ;
        RECT 1732.020 2457.370 1735.020 2457.380 ;
        RECT 1912.020 2457.370 1915.020 2457.380 ;
        RECT 2092.020 2457.370 2095.020 2457.380 ;
        RECT 2272.020 2457.370 2275.020 2457.380 ;
        RECT 2452.020 2457.370 2455.020 2457.380 ;
        RECT 2632.020 2457.370 2635.020 2457.380 ;
        RECT 2812.020 2457.370 2815.020 2457.380 ;
        RECT 2940.400 2457.370 2943.400 2457.380 ;
        RECT -23.780 2280.380 -20.780 2280.390 ;
        RECT 112.020 2280.380 115.020 2280.390 ;
        RECT 292.020 2280.380 295.020 2280.390 ;
        RECT 472.020 2280.380 475.020 2280.390 ;
        RECT 652.020 2280.380 655.020 2280.390 ;
        RECT 832.020 2280.380 835.020 2280.390 ;
        RECT 1012.020 2280.380 1015.020 2280.390 ;
        RECT 1192.020 2280.380 1195.020 2280.390 ;
        RECT 1372.020 2280.380 1375.020 2280.390 ;
        RECT 1552.020 2280.380 1555.020 2280.390 ;
        RECT 1732.020 2280.380 1735.020 2280.390 ;
        RECT 1912.020 2280.380 1915.020 2280.390 ;
        RECT 2092.020 2280.380 2095.020 2280.390 ;
        RECT 2272.020 2280.380 2275.020 2280.390 ;
        RECT 2452.020 2280.380 2455.020 2280.390 ;
        RECT 2632.020 2280.380 2635.020 2280.390 ;
        RECT 2812.020 2280.380 2815.020 2280.390 ;
        RECT 2940.400 2280.380 2943.400 2280.390 ;
        RECT -23.780 2277.380 2943.400 2280.380 ;
        RECT -23.780 2277.370 -20.780 2277.380 ;
        RECT 112.020 2277.370 115.020 2277.380 ;
        RECT 292.020 2277.370 295.020 2277.380 ;
        RECT 472.020 2277.370 475.020 2277.380 ;
        RECT 652.020 2277.370 655.020 2277.380 ;
        RECT 832.020 2277.370 835.020 2277.380 ;
        RECT 1012.020 2277.370 1015.020 2277.380 ;
        RECT 1192.020 2277.370 1195.020 2277.380 ;
        RECT 1372.020 2277.370 1375.020 2277.380 ;
        RECT 1552.020 2277.370 1555.020 2277.380 ;
        RECT 1732.020 2277.370 1735.020 2277.380 ;
        RECT 1912.020 2277.370 1915.020 2277.380 ;
        RECT 2092.020 2277.370 2095.020 2277.380 ;
        RECT 2272.020 2277.370 2275.020 2277.380 ;
        RECT 2452.020 2277.370 2455.020 2277.380 ;
        RECT 2632.020 2277.370 2635.020 2277.380 ;
        RECT 2812.020 2277.370 2815.020 2277.380 ;
        RECT 2940.400 2277.370 2943.400 2277.380 ;
        RECT -23.780 2100.380 -20.780 2100.390 ;
        RECT 112.020 2100.380 115.020 2100.390 ;
        RECT 292.020 2100.380 295.020 2100.390 ;
        RECT 472.020 2100.380 475.020 2100.390 ;
        RECT 652.020 2100.380 655.020 2100.390 ;
        RECT 832.020 2100.380 835.020 2100.390 ;
        RECT 1012.020 2100.380 1015.020 2100.390 ;
        RECT 1192.020 2100.380 1195.020 2100.390 ;
        RECT 1372.020 2100.380 1375.020 2100.390 ;
        RECT 1552.020 2100.380 1555.020 2100.390 ;
        RECT 1732.020 2100.380 1735.020 2100.390 ;
        RECT 1912.020 2100.380 1915.020 2100.390 ;
        RECT 2092.020 2100.380 2095.020 2100.390 ;
        RECT 2272.020 2100.380 2275.020 2100.390 ;
        RECT 2452.020 2100.380 2455.020 2100.390 ;
        RECT 2632.020 2100.380 2635.020 2100.390 ;
        RECT 2812.020 2100.380 2815.020 2100.390 ;
        RECT 2940.400 2100.380 2943.400 2100.390 ;
        RECT -23.780 2097.380 2943.400 2100.380 ;
        RECT -23.780 2097.370 -20.780 2097.380 ;
        RECT 112.020 2097.370 115.020 2097.380 ;
        RECT 292.020 2097.370 295.020 2097.380 ;
        RECT 472.020 2097.370 475.020 2097.380 ;
        RECT 652.020 2097.370 655.020 2097.380 ;
        RECT 832.020 2097.370 835.020 2097.380 ;
        RECT 1012.020 2097.370 1015.020 2097.380 ;
        RECT 1192.020 2097.370 1195.020 2097.380 ;
        RECT 1372.020 2097.370 1375.020 2097.380 ;
        RECT 1552.020 2097.370 1555.020 2097.380 ;
        RECT 1732.020 2097.370 1735.020 2097.380 ;
        RECT 1912.020 2097.370 1915.020 2097.380 ;
        RECT 2092.020 2097.370 2095.020 2097.380 ;
        RECT 2272.020 2097.370 2275.020 2097.380 ;
        RECT 2452.020 2097.370 2455.020 2097.380 ;
        RECT 2632.020 2097.370 2635.020 2097.380 ;
        RECT 2812.020 2097.370 2815.020 2097.380 ;
        RECT 2940.400 2097.370 2943.400 2097.380 ;
        RECT -23.780 1920.380 -20.780 1920.390 ;
        RECT 112.020 1920.380 115.020 1920.390 ;
        RECT 292.020 1920.380 295.020 1920.390 ;
        RECT 472.020 1920.380 475.020 1920.390 ;
        RECT 652.020 1920.380 655.020 1920.390 ;
        RECT 832.020 1920.380 835.020 1920.390 ;
        RECT 1012.020 1920.380 1015.020 1920.390 ;
        RECT 1192.020 1920.380 1195.020 1920.390 ;
        RECT 1372.020 1920.380 1375.020 1920.390 ;
        RECT 1552.020 1920.380 1555.020 1920.390 ;
        RECT 1732.020 1920.380 1735.020 1920.390 ;
        RECT 1912.020 1920.380 1915.020 1920.390 ;
        RECT 2092.020 1920.380 2095.020 1920.390 ;
        RECT 2272.020 1920.380 2275.020 1920.390 ;
        RECT 2452.020 1920.380 2455.020 1920.390 ;
        RECT 2632.020 1920.380 2635.020 1920.390 ;
        RECT 2812.020 1920.380 2815.020 1920.390 ;
        RECT 2940.400 1920.380 2943.400 1920.390 ;
        RECT -23.780 1917.380 2943.400 1920.380 ;
        RECT -23.780 1917.370 -20.780 1917.380 ;
        RECT 112.020 1917.370 115.020 1917.380 ;
        RECT 292.020 1917.370 295.020 1917.380 ;
        RECT 472.020 1917.370 475.020 1917.380 ;
        RECT 652.020 1917.370 655.020 1917.380 ;
        RECT 832.020 1917.370 835.020 1917.380 ;
        RECT 1012.020 1917.370 1015.020 1917.380 ;
        RECT 1192.020 1917.370 1195.020 1917.380 ;
        RECT 1372.020 1917.370 1375.020 1917.380 ;
        RECT 1552.020 1917.370 1555.020 1917.380 ;
        RECT 1732.020 1917.370 1735.020 1917.380 ;
        RECT 1912.020 1917.370 1915.020 1917.380 ;
        RECT 2092.020 1917.370 2095.020 1917.380 ;
        RECT 2272.020 1917.370 2275.020 1917.380 ;
        RECT 2452.020 1917.370 2455.020 1917.380 ;
        RECT 2632.020 1917.370 2635.020 1917.380 ;
        RECT 2812.020 1917.370 2815.020 1917.380 ;
        RECT 2940.400 1917.370 2943.400 1917.380 ;
        RECT -23.780 1740.380 -20.780 1740.390 ;
        RECT 112.020 1740.380 115.020 1740.390 ;
        RECT 292.020 1740.380 295.020 1740.390 ;
        RECT 472.020 1740.380 475.020 1740.390 ;
        RECT 652.020 1740.380 655.020 1740.390 ;
        RECT 832.020 1740.380 835.020 1740.390 ;
        RECT 1012.020 1740.380 1015.020 1740.390 ;
        RECT 1192.020 1740.380 1195.020 1740.390 ;
        RECT 1372.020 1740.380 1375.020 1740.390 ;
        RECT 1552.020 1740.380 1555.020 1740.390 ;
        RECT 1732.020 1740.380 1735.020 1740.390 ;
        RECT 1912.020 1740.380 1915.020 1740.390 ;
        RECT 2092.020 1740.380 2095.020 1740.390 ;
        RECT 2272.020 1740.380 2275.020 1740.390 ;
        RECT 2452.020 1740.380 2455.020 1740.390 ;
        RECT 2632.020 1740.380 2635.020 1740.390 ;
        RECT 2812.020 1740.380 2815.020 1740.390 ;
        RECT 2940.400 1740.380 2943.400 1740.390 ;
        RECT -23.780 1737.380 2943.400 1740.380 ;
        RECT -23.780 1737.370 -20.780 1737.380 ;
        RECT 112.020 1737.370 115.020 1737.380 ;
        RECT 292.020 1737.370 295.020 1737.380 ;
        RECT 472.020 1737.370 475.020 1737.380 ;
        RECT 652.020 1737.370 655.020 1737.380 ;
        RECT 832.020 1737.370 835.020 1737.380 ;
        RECT 1012.020 1737.370 1015.020 1737.380 ;
        RECT 1192.020 1737.370 1195.020 1737.380 ;
        RECT 1372.020 1737.370 1375.020 1737.380 ;
        RECT 1552.020 1737.370 1555.020 1737.380 ;
        RECT 1732.020 1737.370 1735.020 1737.380 ;
        RECT 1912.020 1737.370 1915.020 1737.380 ;
        RECT 2092.020 1737.370 2095.020 1737.380 ;
        RECT 2272.020 1737.370 2275.020 1737.380 ;
        RECT 2452.020 1737.370 2455.020 1737.380 ;
        RECT 2632.020 1737.370 2635.020 1737.380 ;
        RECT 2812.020 1737.370 2815.020 1737.380 ;
        RECT 2940.400 1737.370 2943.400 1737.380 ;
        RECT -23.780 1560.380 -20.780 1560.390 ;
        RECT 112.020 1560.380 115.020 1560.390 ;
        RECT 292.020 1560.380 295.020 1560.390 ;
        RECT 472.020 1560.380 475.020 1560.390 ;
        RECT 652.020 1560.380 655.020 1560.390 ;
        RECT 832.020 1560.380 835.020 1560.390 ;
        RECT 1012.020 1560.380 1015.020 1560.390 ;
        RECT 1192.020 1560.380 1195.020 1560.390 ;
        RECT 1372.020 1560.380 1375.020 1560.390 ;
        RECT 1552.020 1560.380 1555.020 1560.390 ;
        RECT 1732.020 1560.380 1735.020 1560.390 ;
        RECT 1912.020 1560.380 1915.020 1560.390 ;
        RECT 2092.020 1560.380 2095.020 1560.390 ;
        RECT 2272.020 1560.380 2275.020 1560.390 ;
        RECT 2452.020 1560.380 2455.020 1560.390 ;
        RECT 2632.020 1560.380 2635.020 1560.390 ;
        RECT 2812.020 1560.380 2815.020 1560.390 ;
        RECT 2940.400 1560.380 2943.400 1560.390 ;
        RECT -23.780 1557.380 2943.400 1560.380 ;
        RECT -23.780 1557.370 -20.780 1557.380 ;
        RECT 112.020 1557.370 115.020 1557.380 ;
        RECT 292.020 1557.370 295.020 1557.380 ;
        RECT 472.020 1557.370 475.020 1557.380 ;
        RECT 652.020 1557.370 655.020 1557.380 ;
        RECT 832.020 1557.370 835.020 1557.380 ;
        RECT 1012.020 1557.370 1015.020 1557.380 ;
        RECT 1192.020 1557.370 1195.020 1557.380 ;
        RECT 1372.020 1557.370 1375.020 1557.380 ;
        RECT 1552.020 1557.370 1555.020 1557.380 ;
        RECT 1732.020 1557.370 1735.020 1557.380 ;
        RECT 1912.020 1557.370 1915.020 1557.380 ;
        RECT 2092.020 1557.370 2095.020 1557.380 ;
        RECT 2272.020 1557.370 2275.020 1557.380 ;
        RECT 2452.020 1557.370 2455.020 1557.380 ;
        RECT 2632.020 1557.370 2635.020 1557.380 ;
        RECT 2812.020 1557.370 2815.020 1557.380 ;
        RECT 2940.400 1557.370 2943.400 1557.380 ;
        RECT -23.780 1380.380 -20.780 1380.390 ;
        RECT 112.020 1380.380 115.020 1380.390 ;
        RECT 292.020 1380.380 295.020 1380.390 ;
        RECT 472.020 1380.380 475.020 1380.390 ;
        RECT 652.020 1380.380 655.020 1380.390 ;
        RECT 832.020 1380.380 835.020 1380.390 ;
        RECT 1012.020 1380.380 1015.020 1380.390 ;
        RECT 1192.020 1380.380 1195.020 1380.390 ;
        RECT 1372.020 1380.380 1375.020 1380.390 ;
        RECT 1552.020 1380.380 1555.020 1380.390 ;
        RECT 1732.020 1380.380 1735.020 1380.390 ;
        RECT 1912.020 1380.380 1915.020 1380.390 ;
        RECT 2092.020 1380.380 2095.020 1380.390 ;
        RECT 2272.020 1380.380 2275.020 1380.390 ;
        RECT 2452.020 1380.380 2455.020 1380.390 ;
        RECT 2632.020 1380.380 2635.020 1380.390 ;
        RECT 2812.020 1380.380 2815.020 1380.390 ;
        RECT 2940.400 1380.380 2943.400 1380.390 ;
        RECT -23.780 1377.380 2943.400 1380.380 ;
        RECT -23.780 1377.370 -20.780 1377.380 ;
        RECT 112.020 1377.370 115.020 1377.380 ;
        RECT 292.020 1377.370 295.020 1377.380 ;
        RECT 472.020 1377.370 475.020 1377.380 ;
        RECT 652.020 1377.370 655.020 1377.380 ;
        RECT 832.020 1377.370 835.020 1377.380 ;
        RECT 1012.020 1377.370 1015.020 1377.380 ;
        RECT 1192.020 1377.370 1195.020 1377.380 ;
        RECT 1372.020 1377.370 1375.020 1377.380 ;
        RECT 1552.020 1377.370 1555.020 1377.380 ;
        RECT 1732.020 1377.370 1735.020 1377.380 ;
        RECT 1912.020 1377.370 1915.020 1377.380 ;
        RECT 2092.020 1377.370 2095.020 1377.380 ;
        RECT 2272.020 1377.370 2275.020 1377.380 ;
        RECT 2452.020 1377.370 2455.020 1377.380 ;
        RECT 2632.020 1377.370 2635.020 1377.380 ;
        RECT 2812.020 1377.370 2815.020 1377.380 ;
        RECT 2940.400 1377.370 2943.400 1377.380 ;
        RECT -23.780 1200.380 -20.780 1200.390 ;
        RECT 112.020 1200.380 115.020 1200.390 ;
        RECT 292.020 1200.380 295.020 1200.390 ;
        RECT 472.020 1200.380 475.020 1200.390 ;
        RECT 652.020 1200.380 655.020 1200.390 ;
        RECT 832.020 1200.380 835.020 1200.390 ;
        RECT 1012.020 1200.380 1015.020 1200.390 ;
        RECT 1192.020 1200.380 1195.020 1200.390 ;
        RECT 1372.020 1200.380 1375.020 1200.390 ;
        RECT 1552.020 1200.380 1555.020 1200.390 ;
        RECT 1732.020 1200.380 1735.020 1200.390 ;
        RECT 1912.020 1200.380 1915.020 1200.390 ;
        RECT 2092.020 1200.380 2095.020 1200.390 ;
        RECT 2272.020 1200.380 2275.020 1200.390 ;
        RECT 2452.020 1200.380 2455.020 1200.390 ;
        RECT 2632.020 1200.380 2635.020 1200.390 ;
        RECT 2812.020 1200.380 2815.020 1200.390 ;
        RECT 2940.400 1200.380 2943.400 1200.390 ;
        RECT -23.780 1197.380 2943.400 1200.380 ;
        RECT -23.780 1197.370 -20.780 1197.380 ;
        RECT 112.020 1197.370 115.020 1197.380 ;
        RECT 292.020 1197.370 295.020 1197.380 ;
        RECT 472.020 1197.370 475.020 1197.380 ;
        RECT 652.020 1197.370 655.020 1197.380 ;
        RECT 832.020 1197.370 835.020 1197.380 ;
        RECT 1012.020 1197.370 1015.020 1197.380 ;
        RECT 1192.020 1197.370 1195.020 1197.380 ;
        RECT 1372.020 1197.370 1375.020 1197.380 ;
        RECT 1552.020 1197.370 1555.020 1197.380 ;
        RECT 1732.020 1197.370 1735.020 1197.380 ;
        RECT 1912.020 1197.370 1915.020 1197.380 ;
        RECT 2092.020 1197.370 2095.020 1197.380 ;
        RECT 2272.020 1197.370 2275.020 1197.380 ;
        RECT 2452.020 1197.370 2455.020 1197.380 ;
        RECT 2632.020 1197.370 2635.020 1197.380 ;
        RECT 2812.020 1197.370 2815.020 1197.380 ;
        RECT 2940.400 1197.370 2943.400 1197.380 ;
        RECT -23.780 1020.380 -20.780 1020.390 ;
        RECT 112.020 1020.380 115.020 1020.390 ;
        RECT 292.020 1020.380 295.020 1020.390 ;
        RECT 472.020 1020.380 475.020 1020.390 ;
        RECT 652.020 1020.380 655.020 1020.390 ;
        RECT 832.020 1020.380 835.020 1020.390 ;
        RECT 1012.020 1020.380 1015.020 1020.390 ;
        RECT 1192.020 1020.380 1195.020 1020.390 ;
        RECT 1372.020 1020.380 1375.020 1020.390 ;
        RECT 1552.020 1020.380 1555.020 1020.390 ;
        RECT 1732.020 1020.380 1735.020 1020.390 ;
        RECT 1912.020 1020.380 1915.020 1020.390 ;
        RECT 2092.020 1020.380 2095.020 1020.390 ;
        RECT 2272.020 1020.380 2275.020 1020.390 ;
        RECT 2452.020 1020.380 2455.020 1020.390 ;
        RECT 2632.020 1020.380 2635.020 1020.390 ;
        RECT 2812.020 1020.380 2815.020 1020.390 ;
        RECT 2940.400 1020.380 2943.400 1020.390 ;
        RECT -23.780 1017.380 2943.400 1020.380 ;
        RECT -23.780 1017.370 -20.780 1017.380 ;
        RECT 112.020 1017.370 115.020 1017.380 ;
        RECT 292.020 1017.370 295.020 1017.380 ;
        RECT 472.020 1017.370 475.020 1017.380 ;
        RECT 652.020 1017.370 655.020 1017.380 ;
        RECT 832.020 1017.370 835.020 1017.380 ;
        RECT 1012.020 1017.370 1015.020 1017.380 ;
        RECT 1192.020 1017.370 1195.020 1017.380 ;
        RECT 1372.020 1017.370 1375.020 1017.380 ;
        RECT 1552.020 1017.370 1555.020 1017.380 ;
        RECT 1732.020 1017.370 1735.020 1017.380 ;
        RECT 1912.020 1017.370 1915.020 1017.380 ;
        RECT 2092.020 1017.370 2095.020 1017.380 ;
        RECT 2272.020 1017.370 2275.020 1017.380 ;
        RECT 2452.020 1017.370 2455.020 1017.380 ;
        RECT 2632.020 1017.370 2635.020 1017.380 ;
        RECT 2812.020 1017.370 2815.020 1017.380 ;
        RECT 2940.400 1017.370 2943.400 1017.380 ;
        RECT -23.780 840.380 -20.780 840.390 ;
        RECT 112.020 840.380 115.020 840.390 ;
        RECT 292.020 840.380 295.020 840.390 ;
        RECT 472.020 840.380 475.020 840.390 ;
        RECT 652.020 840.380 655.020 840.390 ;
        RECT 832.020 840.380 835.020 840.390 ;
        RECT 1012.020 840.380 1015.020 840.390 ;
        RECT 1192.020 840.380 1195.020 840.390 ;
        RECT 1372.020 840.380 1375.020 840.390 ;
        RECT 1552.020 840.380 1555.020 840.390 ;
        RECT 1732.020 840.380 1735.020 840.390 ;
        RECT 1912.020 840.380 1915.020 840.390 ;
        RECT 2092.020 840.380 2095.020 840.390 ;
        RECT 2272.020 840.380 2275.020 840.390 ;
        RECT 2452.020 840.380 2455.020 840.390 ;
        RECT 2632.020 840.380 2635.020 840.390 ;
        RECT 2812.020 840.380 2815.020 840.390 ;
        RECT 2940.400 840.380 2943.400 840.390 ;
        RECT -23.780 837.380 2943.400 840.380 ;
        RECT -23.780 837.370 -20.780 837.380 ;
        RECT 112.020 837.370 115.020 837.380 ;
        RECT 292.020 837.370 295.020 837.380 ;
        RECT 472.020 837.370 475.020 837.380 ;
        RECT 652.020 837.370 655.020 837.380 ;
        RECT 832.020 837.370 835.020 837.380 ;
        RECT 1012.020 837.370 1015.020 837.380 ;
        RECT 1192.020 837.370 1195.020 837.380 ;
        RECT 1372.020 837.370 1375.020 837.380 ;
        RECT 1552.020 837.370 1555.020 837.380 ;
        RECT 1732.020 837.370 1735.020 837.380 ;
        RECT 1912.020 837.370 1915.020 837.380 ;
        RECT 2092.020 837.370 2095.020 837.380 ;
        RECT 2272.020 837.370 2275.020 837.380 ;
        RECT 2452.020 837.370 2455.020 837.380 ;
        RECT 2632.020 837.370 2635.020 837.380 ;
        RECT 2812.020 837.370 2815.020 837.380 ;
        RECT 2940.400 837.370 2943.400 837.380 ;
        RECT -23.780 660.380 -20.780 660.390 ;
        RECT 112.020 660.380 115.020 660.390 ;
        RECT 292.020 660.380 295.020 660.390 ;
        RECT 472.020 660.380 475.020 660.390 ;
        RECT 652.020 660.380 655.020 660.390 ;
        RECT 832.020 660.380 835.020 660.390 ;
        RECT 1012.020 660.380 1015.020 660.390 ;
        RECT 1192.020 660.380 1195.020 660.390 ;
        RECT 1372.020 660.380 1375.020 660.390 ;
        RECT 1552.020 660.380 1555.020 660.390 ;
        RECT 1732.020 660.380 1735.020 660.390 ;
        RECT 1912.020 660.380 1915.020 660.390 ;
        RECT 2092.020 660.380 2095.020 660.390 ;
        RECT 2272.020 660.380 2275.020 660.390 ;
        RECT 2452.020 660.380 2455.020 660.390 ;
        RECT 2632.020 660.380 2635.020 660.390 ;
        RECT 2812.020 660.380 2815.020 660.390 ;
        RECT 2940.400 660.380 2943.400 660.390 ;
        RECT -23.780 657.380 2943.400 660.380 ;
        RECT -23.780 657.370 -20.780 657.380 ;
        RECT 112.020 657.370 115.020 657.380 ;
        RECT 292.020 657.370 295.020 657.380 ;
        RECT 472.020 657.370 475.020 657.380 ;
        RECT 652.020 657.370 655.020 657.380 ;
        RECT 832.020 657.370 835.020 657.380 ;
        RECT 1012.020 657.370 1015.020 657.380 ;
        RECT 1192.020 657.370 1195.020 657.380 ;
        RECT 1372.020 657.370 1375.020 657.380 ;
        RECT 1552.020 657.370 1555.020 657.380 ;
        RECT 1732.020 657.370 1735.020 657.380 ;
        RECT 1912.020 657.370 1915.020 657.380 ;
        RECT 2092.020 657.370 2095.020 657.380 ;
        RECT 2272.020 657.370 2275.020 657.380 ;
        RECT 2452.020 657.370 2455.020 657.380 ;
        RECT 2632.020 657.370 2635.020 657.380 ;
        RECT 2812.020 657.370 2815.020 657.380 ;
        RECT 2940.400 657.370 2943.400 657.380 ;
        RECT -23.780 480.380 -20.780 480.390 ;
        RECT 112.020 480.380 115.020 480.390 ;
        RECT 292.020 480.380 295.020 480.390 ;
        RECT 472.020 480.380 475.020 480.390 ;
        RECT 652.020 480.380 655.020 480.390 ;
        RECT 832.020 480.380 835.020 480.390 ;
        RECT 1012.020 480.380 1015.020 480.390 ;
        RECT 1192.020 480.380 1195.020 480.390 ;
        RECT 1372.020 480.380 1375.020 480.390 ;
        RECT 1552.020 480.380 1555.020 480.390 ;
        RECT 1732.020 480.380 1735.020 480.390 ;
        RECT 1912.020 480.380 1915.020 480.390 ;
        RECT 2092.020 480.380 2095.020 480.390 ;
        RECT 2272.020 480.380 2275.020 480.390 ;
        RECT 2452.020 480.380 2455.020 480.390 ;
        RECT 2632.020 480.380 2635.020 480.390 ;
        RECT 2812.020 480.380 2815.020 480.390 ;
        RECT 2940.400 480.380 2943.400 480.390 ;
        RECT -23.780 477.380 2943.400 480.380 ;
        RECT -23.780 477.370 -20.780 477.380 ;
        RECT 112.020 477.370 115.020 477.380 ;
        RECT 292.020 477.370 295.020 477.380 ;
        RECT 472.020 477.370 475.020 477.380 ;
        RECT 652.020 477.370 655.020 477.380 ;
        RECT 832.020 477.370 835.020 477.380 ;
        RECT 1012.020 477.370 1015.020 477.380 ;
        RECT 1192.020 477.370 1195.020 477.380 ;
        RECT 1372.020 477.370 1375.020 477.380 ;
        RECT 1552.020 477.370 1555.020 477.380 ;
        RECT 1732.020 477.370 1735.020 477.380 ;
        RECT 1912.020 477.370 1915.020 477.380 ;
        RECT 2092.020 477.370 2095.020 477.380 ;
        RECT 2272.020 477.370 2275.020 477.380 ;
        RECT 2452.020 477.370 2455.020 477.380 ;
        RECT 2632.020 477.370 2635.020 477.380 ;
        RECT 2812.020 477.370 2815.020 477.380 ;
        RECT 2940.400 477.370 2943.400 477.380 ;
        RECT -23.780 300.380 -20.780 300.390 ;
        RECT 112.020 300.380 115.020 300.390 ;
        RECT 292.020 300.380 295.020 300.390 ;
        RECT 472.020 300.380 475.020 300.390 ;
        RECT 652.020 300.380 655.020 300.390 ;
        RECT 832.020 300.380 835.020 300.390 ;
        RECT 1012.020 300.380 1015.020 300.390 ;
        RECT 1192.020 300.380 1195.020 300.390 ;
        RECT 1372.020 300.380 1375.020 300.390 ;
        RECT 1552.020 300.380 1555.020 300.390 ;
        RECT 1732.020 300.380 1735.020 300.390 ;
        RECT 1912.020 300.380 1915.020 300.390 ;
        RECT 2092.020 300.380 2095.020 300.390 ;
        RECT 2272.020 300.380 2275.020 300.390 ;
        RECT 2452.020 300.380 2455.020 300.390 ;
        RECT 2632.020 300.380 2635.020 300.390 ;
        RECT 2812.020 300.380 2815.020 300.390 ;
        RECT 2940.400 300.380 2943.400 300.390 ;
        RECT -23.780 297.380 2943.400 300.380 ;
        RECT -23.780 297.370 -20.780 297.380 ;
        RECT 112.020 297.370 115.020 297.380 ;
        RECT 292.020 297.370 295.020 297.380 ;
        RECT 472.020 297.370 475.020 297.380 ;
        RECT 652.020 297.370 655.020 297.380 ;
        RECT 832.020 297.370 835.020 297.380 ;
        RECT 1012.020 297.370 1015.020 297.380 ;
        RECT 1192.020 297.370 1195.020 297.380 ;
        RECT 1372.020 297.370 1375.020 297.380 ;
        RECT 1552.020 297.370 1555.020 297.380 ;
        RECT 1732.020 297.370 1735.020 297.380 ;
        RECT 1912.020 297.370 1915.020 297.380 ;
        RECT 2092.020 297.370 2095.020 297.380 ;
        RECT 2272.020 297.370 2275.020 297.380 ;
        RECT 2452.020 297.370 2455.020 297.380 ;
        RECT 2632.020 297.370 2635.020 297.380 ;
        RECT 2812.020 297.370 2815.020 297.380 ;
        RECT 2940.400 297.370 2943.400 297.380 ;
        RECT -23.780 120.380 -20.780 120.390 ;
        RECT 112.020 120.380 115.020 120.390 ;
        RECT 292.020 120.380 295.020 120.390 ;
        RECT 472.020 120.380 475.020 120.390 ;
        RECT 652.020 120.380 655.020 120.390 ;
        RECT 832.020 120.380 835.020 120.390 ;
        RECT 1012.020 120.380 1015.020 120.390 ;
        RECT 1192.020 120.380 1195.020 120.390 ;
        RECT 1372.020 120.380 1375.020 120.390 ;
        RECT 1552.020 120.380 1555.020 120.390 ;
        RECT 1732.020 120.380 1735.020 120.390 ;
        RECT 1912.020 120.380 1915.020 120.390 ;
        RECT 2092.020 120.380 2095.020 120.390 ;
        RECT 2272.020 120.380 2275.020 120.390 ;
        RECT 2452.020 120.380 2455.020 120.390 ;
        RECT 2632.020 120.380 2635.020 120.390 ;
        RECT 2812.020 120.380 2815.020 120.390 ;
        RECT 2940.400 120.380 2943.400 120.390 ;
        RECT -23.780 117.380 2943.400 120.380 ;
        RECT -23.780 117.370 -20.780 117.380 ;
        RECT 112.020 117.370 115.020 117.380 ;
        RECT 292.020 117.370 295.020 117.380 ;
        RECT 472.020 117.370 475.020 117.380 ;
        RECT 652.020 117.370 655.020 117.380 ;
        RECT 832.020 117.370 835.020 117.380 ;
        RECT 1012.020 117.370 1015.020 117.380 ;
        RECT 1192.020 117.370 1195.020 117.380 ;
        RECT 1372.020 117.370 1375.020 117.380 ;
        RECT 1552.020 117.370 1555.020 117.380 ;
        RECT 1732.020 117.370 1735.020 117.380 ;
        RECT 1912.020 117.370 1915.020 117.380 ;
        RECT 2092.020 117.370 2095.020 117.380 ;
        RECT 2272.020 117.370 2275.020 117.380 ;
        RECT 2452.020 117.370 2455.020 117.380 ;
        RECT 2632.020 117.370 2635.020 117.380 ;
        RECT 2812.020 117.370 2815.020 117.380 ;
        RECT 2940.400 117.370 2943.400 117.380 ;
        RECT -23.780 -15.420 -20.780 -15.410 ;
        RECT 112.020 -15.420 115.020 -15.410 ;
        RECT 292.020 -15.420 295.020 -15.410 ;
        RECT 472.020 -15.420 475.020 -15.410 ;
        RECT 652.020 -15.420 655.020 -15.410 ;
        RECT 832.020 -15.420 835.020 -15.410 ;
        RECT 1012.020 -15.420 1015.020 -15.410 ;
        RECT 1192.020 -15.420 1195.020 -15.410 ;
        RECT 1372.020 -15.420 1375.020 -15.410 ;
        RECT 1552.020 -15.420 1555.020 -15.410 ;
        RECT 1732.020 -15.420 1735.020 -15.410 ;
        RECT 1912.020 -15.420 1915.020 -15.410 ;
        RECT 2092.020 -15.420 2095.020 -15.410 ;
        RECT 2272.020 -15.420 2275.020 -15.410 ;
        RECT 2452.020 -15.420 2455.020 -15.410 ;
        RECT 2632.020 -15.420 2635.020 -15.410 ;
        RECT 2812.020 -15.420 2815.020 -15.410 ;
        RECT 2940.400 -15.420 2943.400 -15.410 ;
        RECT -23.780 -18.420 2943.400 -15.420 ;
        RECT -23.780 -18.430 -20.780 -18.420 ;
        RECT 112.020 -18.430 115.020 -18.420 ;
        RECT 292.020 -18.430 295.020 -18.420 ;
        RECT 472.020 -18.430 475.020 -18.420 ;
        RECT 652.020 -18.430 655.020 -18.420 ;
        RECT 832.020 -18.430 835.020 -18.420 ;
        RECT 1012.020 -18.430 1015.020 -18.420 ;
        RECT 1192.020 -18.430 1195.020 -18.420 ;
        RECT 1372.020 -18.430 1375.020 -18.420 ;
        RECT 1552.020 -18.430 1555.020 -18.420 ;
        RECT 1732.020 -18.430 1735.020 -18.420 ;
        RECT 1912.020 -18.430 1915.020 -18.420 ;
        RECT 2092.020 -18.430 2095.020 -18.420 ;
        RECT 2272.020 -18.430 2275.020 -18.420 ;
        RECT 2452.020 -18.430 2455.020 -18.420 ;
        RECT 2632.020 -18.430 2635.020 -18.420 ;
        RECT 2812.020 -18.430 2815.020 -18.420 ;
        RECT 2940.400 -18.430 2943.400 -18.420 ;
    END
  END vssd2
  PIN vdda1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -28.380 -23.020 -25.380 3542.700 ;
        RECT 40.020 -27.620 43.020 3547.300 ;
        RECT 220.020 -27.620 223.020 3547.300 ;
        RECT 400.020 -27.620 403.020 3547.300 ;
        RECT 580.020 -27.620 583.020 3547.300 ;
        RECT 760.020 -27.620 763.020 3547.300 ;
        RECT 940.020 -27.620 943.020 3547.300 ;
        RECT 1120.020 -27.620 1123.020 3547.300 ;
        RECT 1300.020 -27.620 1303.020 3547.300 ;
        RECT 1480.020 -27.620 1483.020 3547.300 ;
        RECT 1660.020 -27.620 1663.020 3547.300 ;
        RECT 1840.020 -27.620 1843.020 3547.300 ;
        RECT 2020.020 -27.620 2023.020 3547.300 ;
        RECT 2200.020 -27.620 2203.020 3547.300 ;
        RECT 2380.020 -27.620 2383.020 3547.300 ;
        RECT 2560.020 -27.620 2563.020 3547.300 ;
        RECT 2740.020 -27.620 2743.020 3547.300 ;
        RECT 2945.000 -23.020 2948.000 3542.700 ;
      LAYER via4 ;
        RECT -27.470 3541.410 -26.290 3542.590 ;
        RECT -27.470 3539.810 -26.290 3540.990 ;
        RECT -27.470 3467.090 -26.290 3468.270 ;
        RECT -27.470 3465.490 -26.290 3466.670 ;
        RECT -27.470 3287.090 -26.290 3288.270 ;
        RECT -27.470 3285.490 -26.290 3286.670 ;
        RECT -27.470 3107.090 -26.290 3108.270 ;
        RECT -27.470 3105.490 -26.290 3106.670 ;
        RECT -27.470 2927.090 -26.290 2928.270 ;
        RECT -27.470 2925.490 -26.290 2926.670 ;
        RECT -27.470 2747.090 -26.290 2748.270 ;
        RECT -27.470 2745.490 -26.290 2746.670 ;
        RECT -27.470 2567.090 -26.290 2568.270 ;
        RECT -27.470 2565.490 -26.290 2566.670 ;
        RECT -27.470 2387.090 -26.290 2388.270 ;
        RECT -27.470 2385.490 -26.290 2386.670 ;
        RECT -27.470 2207.090 -26.290 2208.270 ;
        RECT -27.470 2205.490 -26.290 2206.670 ;
        RECT -27.470 2027.090 -26.290 2028.270 ;
        RECT -27.470 2025.490 -26.290 2026.670 ;
        RECT -27.470 1847.090 -26.290 1848.270 ;
        RECT -27.470 1845.490 -26.290 1846.670 ;
        RECT -27.470 1667.090 -26.290 1668.270 ;
        RECT -27.470 1665.490 -26.290 1666.670 ;
        RECT -27.470 1487.090 -26.290 1488.270 ;
        RECT -27.470 1485.490 -26.290 1486.670 ;
        RECT -27.470 1307.090 -26.290 1308.270 ;
        RECT -27.470 1305.490 -26.290 1306.670 ;
        RECT -27.470 1127.090 -26.290 1128.270 ;
        RECT -27.470 1125.490 -26.290 1126.670 ;
        RECT -27.470 947.090 -26.290 948.270 ;
        RECT -27.470 945.490 -26.290 946.670 ;
        RECT -27.470 767.090 -26.290 768.270 ;
        RECT -27.470 765.490 -26.290 766.670 ;
        RECT -27.470 587.090 -26.290 588.270 ;
        RECT -27.470 585.490 -26.290 586.670 ;
        RECT -27.470 407.090 -26.290 408.270 ;
        RECT -27.470 405.490 -26.290 406.670 ;
        RECT -27.470 227.090 -26.290 228.270 ;
        RECT -27.470 225.490 -26.290 226.670 ;
        RECT -27.470 47.090 -26.290 48.270 ;
        RECT -27.470 45.490 -26.290 46.670 ;
        RECT -27.470 -21.310 -26.290 -20.130 ;
        RECT -27.470 -22.910 -26.290 -21.730 ;
        RECT 40.930 3541.410 42.110 3542.590 ;
        RECT 40.930 3539.810 42.110 3540.990 ;
        RECT 40.930 3467.090 42.110 3468.270 ;
        RECT 40.930 3465.490 42.110 3466.670 ;
        RECT 40.930 3287.090 42.110 3288.270 ;
        RECT 40.930 3285.490 42.110 3286.670 ;
        RECT 40.930 3107.090 42.110 3108.270 ;
        RECT 40.930 3105.490 42.110 3106.670 ;
        RECT 40.930 2927.090 42.110 2928.270 ;
        RECT 40.930 2925.490 42.110 2926.670 ;
        RECT 40.930 2747.090 42.110 2748.270 ;
        RECT 40.930 2745.490 42.110 2746.670 ;
        RECT 40.930 2567.090 42.110 2568.270 ;
        RECT 40.930 2565.490 42.110 2566.670 ;
        RECT 40.930 2387.090 42.110 2388.270 ;
        RECT 40.930 2385.490 42.110 2386.670 ;
        RECT 40.930 2207.090 42.110 2208.270 ;
        RECT 40.930 2205.490 42.110 2206.670 ;
        RECT 40.930 2027.090 42.110 2028.270 ;
        RECT 40.930 2025.490 42.110 2026.670 ;
        RECT 40.930 1847.090 42.110 1848.270 ;
        RECT 40.930 1845.490 42.110 1846.670 ;
        RECT 40.930 1667.090 42.110 1668.270 ;
        RECT 40.930 1665.490 42.110 1666.670 ;
        RECT 40.930 1487.090 42.110 1488.270 ;
        RECT 40.930 1485.490 42.110 1486.670 ;
        RECT 40.930 1307.090 42.110 1308.270 ;
        RECT 40.930 1305.490 42.110 1306.670 ;
        RECT 40.930 1127.090 42.110 1128.270 ;
        RECT 40.930 1125.490 42.110 1126.670 ;
        RECT 40.930 947.090 42.110 948.270 ;
        RECT 40.930 945.490 42.110 946.670 ;
        RECT 40.930 767.090 42.110 768.270 ;
        RECT 40.930 765.490 42.110 766.670 ;
        RECT 40.930 587.090 42.110 588.270 ;
        RECT 40.930 585.490 42.110 586.670 ;
        RECT 40.930 407.090 42.110 408.270 ;
        RECT 40.930 405.490 42.110 406.670 ;
        RECT 40.930 227.090 42.110 228.270 ;
        RECT 40.930 225.490 42.110 226.670 ;
        RECT 40.930 47.090 42.110 48.270 ;
        RECT 40.930 45.490 42.110 46.670 ;
        RECT 40.930 -21.310 42.110 -20.130 ;
        RECT 40.930 -22.910 42.110 -21.730 ;
        RECT 220.930 3541.410 222.110 3542.590 ;
        RECT 220.930 3539.810 222.110 3540.990 ;
        RECT 220.930 3467.090 222.110 3468.270 ;
        RECT 220.930 3465.490 222.110 3466.670 ;
        RECT 220.930 3287.090 222.110 3288.270 ;
        RECT 220.930 3285.490 222.110 3286.670 ;
        RECT 220.930 3107.090 222.110 3108.270 ;
        RECT 220.930 3105.490 222.110 3106.670 ;
        RECT 220.930 2927.090 222.110 2928.270 ;
        RECT 220.930 2925.490 222.110 2926.670 ;
        RECT 220.930 2747.090 222.110 2748.270 ;
        RECT 220.930 2745.490 222.110 2746.670 ;
        RECT 220.930 2567.090 222.110 2568.270 ;
        RECT 220.930 2565.490 222.110 2566.670 ;
        RECT 220.930 2387.090 222.110 2388.270 ;
        RECT 220.930 2385.490 222.110 2386.670 ;
        RECT 220.930 2207.090 222.110 2208.270 ;
        RECT 220.930 2205.490 222.110 2206.670 ;
        RECT 220.930 2027.090 222.110 2028.270 ;
        RECT 220.930 2025.490 222.110 2026.670 ;
        RECT 220.930 1847.090 222.110 1848.270 ;
        RECT 220.930 1845.490 222.110 1846.670 ;
        RECT 220.930 1667.090 222.110 1668.270 ;
        RECT 220.930 1665.490 222.110 1666.670 ;
        RECT 220.930 1487.090 222.110 1488.270 ;
        RECT 220.930 1485.490 222.110 1486.670 ;
        RECT 220.930 1307.090 222.110 1308.270 ;
        RECT 220.930 1305.490 222.110 1306.670 ;
        RECT 220.930 1127.090 222.110 1128.270 ;
        RECT 220.930 1125.490 222.110 1126.670 ;
        RECT 220.930 947.090 222.110 948.270 ;
        RECT 220.930 945.490 222.110 946.670 ;
        RECT 220.930 767.090 222.110 768.270 ;
        RECT 220.930 765.490 222.110 766.670 ;
        RECT 220.930 587.090 222.110 588.270 ;
        RECT 220.930 585.490 222.110 586.670 ;
        RECT 220.930 407.090 222.110 408.270 ;
        RECT 220.930 405.490 222.110 406.670 ;
        RECT 220.930 227.090 222.110 228.270 ;
        RECT 220.930 225.490 222.110 226.670 ;
        RECT 220.930 47.090 222.110 48.270 ;
        RECT 220.930 45.490 222.110 46.670 ;
        RECT 220.930 -21.310 222.110 -20.130 ;
        RECT 220.930 -22.910 222.110 -21.730 ;
        RECT 400.930 3541.410 402.110 3542.590 ;
        RECT 400.930 3539.810 402.110 3540.990 ;
        RECT 400.930 3467.090 402.110 3468.270 ;
        RECT 400.930 3465.490 402.110 3466.670 ;
        RECT 400.930 3287.090 402.110 3288.270 ;
        RECT 400.930 3285.490 402.110 3286.670 ;
        RECT 400.930 3107.090 402.110 3108.270 ;
        RECT 400.930 3105.490 402.110 3106.670 ;
        RECT 400.930 2927.090 402.110 2928.270 ;
        RECT 400.930 2925.490 402.110 2926.670 ;
        RECT 400.930 2747.090 402.110 2748.270 ;
        RECT 400.930 2745.490 402.110 2746.670 ;
        RECT 400.930 2567.090 402.110 2568.270 ;
        RECT 400.930 2565.490 402.110 2566.670 ;
        RECT 400.930 2387.090 402.110 2388.270 ;
        RECT 400.930 2385.490 402.110 2386.670 ;
        RECT 400.930 2207.090 402.110 2208.270 ;
        RECT 400.930 2205.490 402.110 2206.670 ;
        RECT 400.930 2027.090 402.110 2028.270 ;
        RECT 400.930 2025.490 402.110 2026.670 ;
        RECT 400.930 1847.090 402.110 1848.270 ;
        RECT 400.930 1845.490 402.110 1846.670 ;
        RECT 400.930 1667.090 402.110 1668.270 ;
        RECT 400.930 1665.490 402.110 1666.670 ;
        RECT 400.930 1487.090 402.110 1488.270 ;
        RECT 400.930 1485.490 402.110 1486.670 ;
        RECT 400.930 1307.090 402.110 1308.270 ;
        RECT 400.930 1305.490 402.110 1306.670 ;
        RECT 400.930 1127.090 402.110 1128.270 ;
        RECT 400.930 1125.490 402.110 1126.670 ;
        RECT 400.930 947.090 402.110 948.270 ;
        RECT 400.930 945.490 402.110 946.670 ;
        RECT 400.930 767.090 402.110 768.270 ;
        RECT 400.930 765.490 402.110 766.670 ;
        RECT 400.930 587.090 402.110 588.270 ;
        RECT 400.930 585.490 402.110 586.670 ;
        RECT 400.930 407.090 402.110 408.270 ;
        RECT 400.930 405.490 402.110 406.670 ;
        RECT 400.930 227.090 402.110 228.270 ;
        RECT 400.930 225.490 402.110 226.670 ;
        RECT 400.930 47.090 402.110 48.270 ;
        RECT 400.930 45.490 402.110 46.670 ;
        RECT 400.930 -21.310 402.110 -20.130 ;
        RECT 400.930 -22.910 402.110 -21.730 ;
        RECT 580.930 3541.410 582.110 3542.590 ;
        RECT 580.930 3539.810 582.110 3540.990 ;
        RECT 580.930 3467.090 582.110 3468.270 ;
        RECT 580.930 3465.490 582.110 3466.670 ;
        RECT 580.930 3287.090 582.110 3288.270 ;
        RECT 580.930 3285.490 582.110 3286.670 ;
        RECT 580.930 3107.090 582.110 3108.270 ;
        RECT 580.930 3105.490 582.110 3106.670 ;
        RECT 580.930 2927.090 582.110 2928.270 ;
        RECT 580.930 2925.490 582.110 2926.670 ;
        RECT 580.930 2747.090 582.110 2748.270 ;
        RECT 580.930 2745.490 582.110 2746.670 ;
        RECT 580.930 2567.090 582.110 2568.270 ;
        RECT 580.930 2565.490 582.110 2566.670 ;
        RECT 580.930 2387.090 582.110 2388.270 ;
        RECT 580.930 2385.490 582.110 2386.670 ;
        RECT 580.930 2207.090 582.110 2208.270 ;
        RECT 580.930 2205.490 582.110 2206.670 ;
        RECT 580.930 2027.090 582.110 2028.270 ;
        RECT 580.930 2025.490 582.110 2026.670 ;
        RECT 580.930 1847.090 582.110 1848.270 ;
        RECT 580.930 1845.490 582.110 1846.670 ;
        RECT 580.930 1667.090 582.110 1668.270 ;
        RECT 580.930 1665.490 582.110 1666.670 ;
        RECT 580.930 1487.090 582.110 1488.270 ;
        RECT 580.930 1485.490 582.110 1486.670 ;
        RECT 580.930 1307.090 582.110 1308.270 ;
        RECT 580.930 1305.490 582.110 1306.670 ;
        RECT 580.930 1127.090 582.110 1128.270 ;
        RECT 580.930 1125.490 582.110 1126.670 ;
        RECT 580.930 947.090 582.110 948.270 ;
        RECT 580.930 945.490 582.110 946.670 ;
        RECT 580.930 767.090 582.110 768.270 ;
        RECT 580.930 765.490 582.110 766.670 ;
        RECT 580.930 587.090 582.110 588.270 ;
        RECT 580.930 585.490 582.110 586.670 ;
        RECT 580.930 407.090 582.110 408.270 ;
        RECT 580.930 405.490 582.110 406.670 ;
        RECT 580.930 227.090 582.110 228.270 ;
        RECT 580.930 225.490 582.110 226.670 ;
        RECT 580.930 47.090 582.110 48.270 ;
        RECT 580.930 45.490 582.110 46.670 ;
        RECT 580.930 -21.310 582.110 -20.130 ;
        RECT 580.930 -22.910 582.110 -21.730 ;
        RECT 760.930 3541.410 762.110 3542.590 ;
        RECT 760.930 3539.810 762.110 3540.990 ;
        RECT 760.930 3467.090 762.110 3468.270 ;
        RECT 760.930 3465.490 762.110 3466.670 ;
        RECT 760.930 3287.090 762.110 3288.270 ;
        RECT 760.930 3285.490 762.110 3286.670 ;
        RECT 760.930 3107.090 762.110 3108.270 ;
        RECT 760.930 3105.490 762.110 3106.670 ;
        RECT 760.930 2927.090 762.110 2928.270 ;
        RECT 760.930 2925.490 762.110 2926.670 ;
        RECT 760.930 2747.090 762.110 2748.270 ;
        RECT 760.930 2745.490 762.110 2746.670 ;
        RECT 760.930 2567.090 762.110 2568.270 ;
        RECT 760.930 2565.490 762.110 2566.670 ;
        RECT 760.930 2387.090 762.110 2388.270 ;
        RECT 760.930 2385.490 762.110 2386.670 ;
        RECT 760.930 2207.090 762.110 2208.270 ;
        RECT 760.930 2205.490 762.110 2206.670 ;
        RECT 760.930 2027.090 762.110 2028.270 ;
        RECT 760.930 2025.490 762.110 2026.670 ;
        RECT 760.930 1847.090 762.110 1848.270 ;
        RECT 760.930 1845.490 762.110 1846.670 ;
        RECT 760.930 1667.090 762.110 1668.270 ;
        RECT 760.930 1665.490 762.110 1666.670 ;
        RECT 760.930 1487.090 762.110 1488.270 ;
        RECT 760.930 1485.490 762.110 1486.670 ;
        RECT 760.930 1307.090 762.110 1308.270 ;
        RECT 760.930 1305.490 762.110 1306.670 ;
        RECT 760.930 1127.090 762.110 1128.270 ;
        RECT 760.930 1125.490 762.110 1126.670 ;
        RECT 760.930 947.090 762.110 948.270 ;
        RECT 760.930 945.490 762.110 946.670 ;
        RECT 760.930 767.090 762.110 768.270 ;
        RECT 760.930 765.490 762.110 766.670 ;
        RECT 760.930 587.090 762.110 588.270 ;
        RECT 760.930 585.490 762.110 586.670 ;
        RECT 760.930 407.090 762.110 408.270 ;
        RECT 760.930 405.490 762.110 406.670 ;
        RECT 760.930 227.090 762.110 228.270 ;
        RECT 760.930 225.490 762.110 226.670 ;
        RECT 760.930 47.090 762.110 48.270 ;
        RECT 760.930 45.490 762.110 46.670 ;
        RECT 760.930 -21.310 762.110 -20.130 ;
        RECT 760.930 -22.910 762.110 -21.730 ;
        RECT 940.930 3541.410 942.110 3542.590 ;
        RECT 940.930 3539.810 942.110 3540.990 ;
        RECT 940.930 3467.090 942.110 3468.270 ;
        RECT 940.930 3465.490 942.110 3466.670 ;
        RECT 940.930 3287.090 942.110 3288.270 ;
        RECT 940.930 3285.490 942.110 3286.670 ;
        RECT 940.930 3107.090 942.110 3108.270 ;
        RECT 940.930 3105.490 942.110 3106.670 ;
        RECT 940.930 2927.090 942.110 2928.270 ;
        RECT 940.930 2925.490 942.110 2926.670 ;
        RECT 940.930 2747.090 942.110 2748.270 ;
        RECT 940.930 2745.490 942.110 2746.670 ;
        RECT 940.930 2567.090 942.110 2568.270 ;
        RECT 940.930 2565.490 942.110 2566.670 ;
        RECT 940.930 2387.090 942.110 2388.270 ;
        RECT 940.930 2385.490 942.110 2386.670 ;
        RECT 940.930 2207.090 942.110 2208.270 ;
        RECT 940.930 2205.490 942.110 2206.670 ;
        RECT 940.930 2027.090 942.110 2028.270 ;
        RECT 940.930 2025.490 942.110 2026.670 ;
        RECT 940.930 1847.090 942.110 1848.270 ;
        RECT 940.930 1845.490 942.110 1846.670 ;
        RECT 940.930 1667.090 942.110 1668.270 ;
        RECT 940.930 1665.490 942.110 1666.670 ;
        RECT 940.930 1487.090 942.110 1488.270 ;
        RECT 940.930 1485.490 942.110 1486.670 ;
        RECT 940.930 1307.090 942.110 1308.270 ;
        RECT 940.930 1305.490 942.110 1306.670 ;
        RECT 940.930 1127.090 942.110 1128.270 ;
        RECT 940.930 1125.490 942.110 1126.670 ;
        RECT 940.930 947.090 942.110 948.270 ;
        RECT 940.930 945.490 942.110 946.670 ;
        RECT 940.930 767.090 942.110 768.270 ;
        RECT 940.930 765.490 942.110 766.670 ;
        RECT 940.930 587.090 942.110 588.270 ;
        RECT 940.930 585.490 942.110 586.670 ;
        RECT 940.930 407.090 942.110 408.270 ;
        RECT 940.930 405.490 942.110 406.670 ;
        RECT 940.930 227.090 942.110 228.270 ;
        RECT 940.930 225.490 942.110 226.670 ;
        RECT 940.930 47.090 942.110 48.270 ;
        RECT 940.930 45.490 942.110 46.670 ;
        RECT 940.930 -21.310 942.110 -20.130 ;
        RECT 940.930 -22.910 942.110 -21.730 ;
        RECT 1120.930 3541.410 1122.110 3542.590 ;
        RECT 1120.930 3539.810 1122.110 3540.990 ;
        RECT 1120.930 3467.090 1122.110 3468.270 ;
        RECT 1120.930 3465.490 1122.110 3466.670 ;
        RECT 1120.930 3287.090 1122.110 3288.270 ;
        RECT 1120.930 3285.490 1122.110 3286.670 ;
        RECT 1120.930 3107.090 1122.110 3108.270 ;
        RECT 1120.930 3105.490 1122.110 3106.670 ;
        RECT 1120.930 2927.090 1122.110 2928.270 ;
        RECT 1120.930 2925.490 1122.110 2926.670 ;
        RECT 1120.930 2747.090 1122.110 2748.270 ;
        RECT 1120.930 2745.490 1122.110 2746.670 ;
        RECT 1120.930 2567.090 1122.110 2568.270 ;
        RECT 1120.930 2565.490 1122.110 2566.670 ;
        RECT 1120.930 2387.090 1122.110 2388.270 ;
        RECT 1120.930 2385.490 1122.110 2386.670 ;
        RECT 1120.930 2207.090 1122.110 2208.270 ;
        RECT 1120.930 2205.490 1122.110 2206.670 ;
        RECT 1120.930 2027.090 1122.110 2028.270 ;
        RECT 1120.930 2025.490 1122.110 2026.670 ;
        RECT 1120.930 1847.090 1122.110 1848.270 ;
        RECT 1120.930 1845.490 1122.110 1846.670 ;
        RECT 1120.930 1667.090 1122.110 1668.270 ;
        RECT 1120.930 1665.490 1122.110 1666.670 ;
        RECT 1120.930 1487.090 1122.110 1488.270 ;
        RECT 1120.930 1485.490 1122.110 1486.670 ;
        RECT 1120.930 1307.090 1122.110 1308.270 ;
        RECT 1120.930 1305.490 1122.110 1306.670 ;
        RECT 1120.930 1127.090 1122.110 1128.270 ;
        RECT 1120.930 1125.490 1122.110 1126.670 ;
        RECT 1120.930 947.090 1122.110 948.270 ;
        RECT 1120.930 945.490 1122.110 946.670 ;
        RECT 1120.930 767.090 1122.110 768.270 ;
        RECT 1120.930 765.490 1122.110 766.670 ;
        RECT 1120.930 587.090 1122.110 588.270 ;
        RECT 1120.930 585.490 1122.110 586.670 ;
        RECT 1120.930 407.090 1122.110 408.270 ;
        RECT 1120.930 405.490 1122.110 406.670 ;
        RECT 1120.930 227.090 1122.110 228.270 ;
        RECT 1120.930 225.490 1122.110 226.670 ;
        RECT 1120.930 47.090 1122.110 48.270 ;
        RECT 1120.930 45.490 1122.110 46.670 ;
        RECT 1120.930 -21.310 1122.110 -20.130 ;
        RECT 1120.930 -22.910 1122.110 -21.730 ;
        RECT 1300.930 3541.410 1302.110 3542.590 ;
        RECT 1300.930 3539.810 1302.110 3540.990 ;
        RECT 1300.930 3467.090 1302.110 3468.270 ;
        RECT 1300.930 3465.490 1302.110 3466.670 ;
        RECT 1300.930 3287.090 1302.110 3288.270 ;
        RECT 1300.930 3285.490 1302.110 3286.670 ;
        RECT 1300.930 3107.090 1302.110 3108.270 ;
        RECT 1300.930 3105.490 1302.110 3106.670 ;
        RECT 1300.930 2927.090 1302.110 2928.270 ;
        RECT 1300.930 2925.490 1302.110 2926.670 ;
        RECT 1300.930 2747.090 1302.110 2748.270 ;
        RECT 1300.930 2745.490 1302.110 2746.670 ;
        RECT 1300.930 2567.090 1302.110 2568.270 ;
        RECT 1300.930 2565.490 1302.110 2566.670 ;
        RECT 1300.930 2387.090 1302.110 2388.270 ;
        RECT 1300.930 2385.490 1302.110 2386.670 ;
        RECT 1300.930 2207.090 1302.110 2208.270 ;
        RECT 1300.930 2205.490 1302.110 2206.670 ;
        RECT 1300.930 2027.090 1302.110 2028.270 ;
        RECT 1300.930 2025.490 1302.110 2026.670 ;
        RECT 1300.930 1847.090 1302.110 1848.270 ;
        RECT 1300.930 1845.490 1302.110 1846.670 ;
        RECT 1300.930 1667.090 1302.110 1668.270 ;
        RECT 1300.930 1665.490 1302.110 1666.670 ;
        RECT 1300.930 1487.090 1302.110 1488.270 ;
        RECT 1300.930 1485.490 1302.110 1486.670 ;
        RECT 1300.930 1307.090 1302.110 1308.270 ;
        RECT 1300.930 1305.490 1302.110 1306.670 ;
        RECT 1300.930 1127.090 1302.110 1128.270 ;
        RECT 1300.930 1125.490 1302.110 1126.670 ;
        RECT 1300.930 947.090 1302.110 948.270 ;
        RECT 1300.930 945.490 1302.110 946.670 ;
        RECT 1300.930 767.090 1302.110 768.270 ;
        RECT 1300.930 765.490 1302.110 766.670 ;
        RECT 1300.930 587.090 1302.110 588.270 ;
        RECT 1300.930 585.490 1302.110 586.670 ;
        RECT 1300.930 407.090 1302.110 408.270 ;
        RECT 1300.930 405.490 1302.110 406.670 ;
        RECT 1300.930 227.090 1302.110 228.270 ;
        RECT 1300.930 225.490 1302.110 226.670 ;
        RECT 1300.930 47.090 1302.110 48.270 ;
        RECT 1300.930 45.490 1302.110 46.670 ;
        RECT 1300.930 -21.310 1302.110 -20.130 ;
        RECT 1300.930 -22.910 1302.110 -21.730 ;
        RECT 1480.930 3541.410 1482.110 3542.590 ;
        RECT 1480.930 3539.810 1482.110 3540.990 ;
        RECT 1480.930 3467.090 1482.110 3468.270 ;
        RECT 1480.930 3465.490 1482.110 3466.670 ;
        RECT 1480.930 3287.090 1482.110 3288.270 ;
        RECT 1480.930 3285.490 1482.110 3286.670 ;
        RECT 1480.930 3107.090 1482.110 3108.270 ;
        RECT 1480.930 3105.490 1482.110 3106.670 ;
        RECT 1480.930 2927.090 1482.110 2928.270 ;
        RECT 1480.930 2925.490 1482.110 2926.670 ;
        RECT 1480.930 2747.090 1482.110 2748.270 ;
        RECT 1480.930 2745.490 1482.110 2746.670 ;
        RECT 1480.930 2567.090 1482.110 2568.270 ;
        RECT 1480.930 2565.490 1482.110 2566.670 ;
        RECT 1480.930 2387.090 1482.110 2388.270 ;
        RECT 1480.930 2385.490 1482.110 2386.670 ;
        RECT 1480.930 2207.090 1482.110 2208.270 ;
        RECT 1480.930 2205.490 1482.110 2206.670 ;
        RECT 1480.930 2027.090 1482.110 2028.270 ;
        RECT 1480.930 2025.490 1482.110 2026.670 ;
        RECT 1480.930 1847.090 1482.110 1848.270 ;
        RECT 1480.930 1845.490 1482.110 1846.670 ;
        RECT 1480.930 1667.090 1482.110 1668.270 ;
        RECT 1480.930 1665.490 1482.110 1666.670 ;
        RECT 1480.930 1487.090 1482.110 1488.270 ;
        RECT 1480.930 1485.490 1482.110 1486.670 ;
        RECT 1480.930 1307.090 1482.110 1308.270 ;
        RECT 1480.930 1305.490 1482.110 1306.670 ;
        RECT 1480.930 1127.090 1482.110 1128.270 ;
        RECT 1480.930 1125.490 1482.110 1126.670 ;
        RECT 1480.930 947.090 1482.110 948.270 ;
        RECT 1480.930 945.490 1482.110 946.670 ;
        RECT 1480.930 767.090 1482.110 768.270 ;
        RECT 1480.930 765.490 1482.110 766.670 ;
        RECT 1480.930 587.090 1482.110 588.270 ;
        RECT 1480.930 585.490 1482.110 586.670 ;
        RECT 1480.930 407.090 1482.110 408.270 ;
        RECT 1480.930 405.490 1482.110 406.670 ;
        RECT 1480.930 227.090 1482.110 228.270 ;
        RECT 1480.930 225.490 1482.110 226.670 ;
        RECT 1480.930 47.090 1482.110 48.270 ;
        RECT 1480.930 45.490 1482.110 46.670 ;
        RECT 1480.930 -21.310 1482.110 -20.130 ;
        RECT 1480.930 -22.910 1482.110 -21.730 ;
        RECT 1660.930 3541.410 1662.110 3542.590 ;
        RECT 1660.930 3539.810 1662.110 3540.990 ;
        RECT 1660.930 3467.090 1662.110 3468.270 ;
        RECT 1660.930 3465.490 1662.110 3466.670 ;
        RECT 1660.930 3287.090 1662.110 3288.270 ;
        RECT 1660.930 3285.490 1662.110 3286.670 ;
        RECT 1660.930 3107.090 1662.110 3108.270 ;
        RECT 1660.930 3105.490 1662.110 3106.670 ;
        RECT 1660.930 2927.090 1662.110 2928.270 ;
        RECT 1660.930 2925.490 1662.110 2926.670 ;
        RECT 1660.930 2747.090 1662.110 2748.270 ;
        RECT 1660.930 2745.490 1662.110 2746.670 ;
        RECT 1660.930 2567.090 1662.110 2568.270 ;
        RECT 1660.930 2565.490 1662.110 2566.670 ;
        RECT 1660.930 2387.090 1662.110 2388.270 ;
        RECT 1660.930 2385.490 1662.110 2386.670 ;
        RECT 1660.930 2207.090 1662.110 2208.270 ;
        RECT 1660.930 2205.490 1662.110 2206.670 ;
        RECT 1660.930 2027.090 1662.110 2028.270 ;
        RECT 1660.930 2025.490 1662.110 2026.670 ;
        RECT 1660.930 1847.090 1662.110 1848.270 ;
        RECT 1660.930 1845.490 1662.110 1846.670 ;
        RECT 1660.930 1667.090 1662.110 1668.270 ;
        RECT 1660.930 1665.490 1662.110 1666.670 ;
        RECT 1660.930 1487.090 1662.110 1488.270 ;
        RECT 1660.930 1485.490 1662.110 1486.670 ;
        RECT 1660.930 1307.090 1662.110 1308.270 ;
        RECT 1660.930 1305.490 1662.110 1306.670 ;
        RECT 1660.930 1127.090 1662.110 1128.270 ;
        RECT 1660.930 1125.490 1662.110 1126.670 ;
        RECT 1660.930 947.090 1662.110 948.270 ;
        RECT 1660.930 945.490 1662.110 946.670 ;
        RECT 1660.930 767.090 1662.110 768.270 ;
        RECT 1660.930 765.490 1662.110 766.670 ;
        RECT 1660.930 587.090 1662.110 588.270 ;
        RECT 1660.930 585.490 1662.110 586.670 ;
        RECT 1660.930 407.090 1662.110 408.270 ;
        RECT 1660.930 405.490 1662.110 406.670 ;
        RECT 1660.930 227.090 1662.110 228.270 ;
        RECT 1660.930 225.490 1662.110 226.670 ;
        RECT 1660.930 47.090 1662.110 48.270 ;
        RECT 1660.930 45.490 1662.110 46.670 ;
        RECT 1660.930 -21.310 1662.110 -20.130 ;
        RECT 1660.930 -22.910 1662.110 -21.730 ;
        RECT 1840.930 3541.410 1842.110 3542.590 ;
        RECT 1840.930 3539.810 1842.110 3540.990 ;
        RECT 1840.930 3467.090 1842.110 3468.270 ;
        RECT 1840.930 3465.490 1842.110 3466.670 ;
        RECT 1840.930 3287.090 1842.110 3288.270 ;
        RECT 1840.930 3285.490 1842.110 3286.670 ;
        RECT 1840.930 3107.090 1842.110 3108.270 ;
        RECT 1840.930 3105.490 1842.110 3106.670 ;
        RECT 1840.930 2927.090 1842.110 2928.270 ;
        RECT 1840.930 2925.490 1842.110 2926.670 ;
        RECT 1840.930 2747.090 1842.110 2748.270 ;
        RECT 1840.930 2745.490 1842.110 2746.670 ;
        RECT 1840.930 2567.090 1842.110 2568.270 ;
        RECT 1840.930 2565.490 1842.110 2566.670 ;
        RECT 1840.930 2387.090 1842.110 2388.270 ;
        RECT 1840.930 2385.490 1842.110 2386.670 ;
        RECT 1840.930 2207.090 1842.110 2208.270 ;
        RECT 1840.930 2205.490 1842.110 2206.670 ;
        RECT 1840.930 2027.090 1842.110 2028.270 ;
        RECT 1840.930 2025.490 1842.110 2026.670 ;
        RECT 1840.930 1847.090 1842.110 1848.270 ;
        RECT 1840.930 1845.490 1842.110 1846.670 ;
        RECT 1840.930 1667.090 1842.110 1668.270 ;
        RECT 1840.930 1665.490 1842.110 1666.670 ;
        RECT 1840.930 1487.090 1842.110 1488.270 ;
        RECT 1840.930 1485.490 1842.110 1486.670 ;
        RECT 1840.930 1307.090 1842.110 1308.270 ;
        RECT 1840.930 1305.490 1842.110 1306.670 ;
        RECT 1840.930 1127.090 1842.110 1128.270 ;
        RECT 1840.930 1125.490 1842.110 1126.670 ;
        RECT 1840.930 947.090 1842.110 948.270 ;
        RECT 1840.930 945.490 1842.110 946.670 ;
        RECT 1840.930 767.090 1842.110 768.270 ;
        RECT 1840.930 765.490 1842.110 766.670 ;
        RECT 1840.930 587.090 1842.110 588.270 ;
        RECT 1840.930 585.490 1842.110 586.670 ;
        RECT 1840.930 407.090 1842.110 408.270 ;
        RECT 1840.930 405.490 1842.110 406.670 ;
        RECT 1840.930 227.090 1842.110 228.270 ;
        RECT 1840.930 225.490 1842.110 226.670 ;
        RECT 1840.930 47.090 1842.110 48.270 ;
        RECT 1840.930 45.490 1842.110 46.670 ;
        RECT 1840.930 -21.310 1842.110 -20.130 ;
        RECT 1840.930 -22.910 1842.110 -21.730 ;
        RECT 2020.930 3541.410 2022.110 3542.590 ;
        RECT 2020.930 3539.810 2022.110 3540.990 ;
        RECT 2020.930 3467.090 2022.110 3468.270 ;
        RECT 2020.930 3465.490 2022.110 3466.670 ;
        RECT 2020.930 3287.090 2022.110 3288.270 ;
        RECT 2020.930 3285.490 2022.110 3286.670 ;
        RECT 2020.930 3107.090 2022.110 3108.270 ;
        RECT 2020.930 3105.490 2022.110 3106.670 ;
        RECT 2020.930 2927.090 2022.110 2928.270 ;
        RECT 2020.930 2925.490 2022.110 2926.670 ;
        RECT 2020.930 2747.090 2022.110 2748.270 ;
        RECT 2020.930 2745.490 2022.110 2746.670 ;
        RECT 2020.930 2567.090 2022.110 2568.270 ;
        RECT 2020.930 2565.490 2022.110 2566.670 ;
        RECT 2020.930 2387.090 2022.110 2388.270 ;
        RECT 2020.930 2385.490 2022.110 2386.670 ;
        RECT 2020.930 2207.090 2022.110 2208.270 ;
        RECT 2020.930 2205.490 2022.110 2206.670 ;
        RECT 2020.930 2027.090 2022.110 2028.270 ;
        RECT 2020.930 2025.490 2022.110 2026.670 ;
        RECT 2020.930 1847.090 2022.110 1848.270 ;
        RECT 2020.930 1845.490 2022.110 1846.670 ;
        RECT 2020.930 1667.090 2022.110 1668.270 ;
        RECT 2020.930 1665.490 2022.110 1666.670 ;
        RECT 2020.930 1487.090 2022.110 1488.270 ;
        RECT 2020.930 1485.490 2022.110 1486.670 ;
        RECT 2020.930 1307.090 2022.110 1308.270 ;
        RECT 2020.930 1305.490 2022.110 1306.670 ;
        RECT 2020.930 1127.090 2022.110 1128.270 ;
        RECT 2020.930 1125.490 2022.110 1126.670 ;
        RECT 2020.930 947.090 2022.110 948.270 ;
        RECT 2020.930 945.490 2022.110 946.670 ;
        RECT 2020.930 767.090 2022.110 768.270 ;
        RECT 2020.930 765.490 2022.110 766.670 ;
        RECT 2020.930 587.090 2022.110 588.270 ;
        RECT 2020.930 585.490 2022.110 586.670 ;
        RECT 2020.930 407.090 2022.110 408.270 ;
        RECT 2020.930 405.490 2022.110 406.670 ;
        RECT 2020.930 227.090 2022.110 228.270 ;
        RECT 2020.930 225.490 2022.110 226.670 ;
        RECT 2020.930 47.090 2022.110 48.270 ;
        RECT 2020.930 45.490 2022.110 46.670 ;
        RECT 2020.930 -21.310 2022.110 -20.130 ;
        RECT 2020.930 -22.910 2022.110 -21.730 ;
        RECT 2200.930 3541.410 2202.110 3542.590 ;
        RECT 2200.930 3539.810 2202.110 3540.990 ;
        RECT 2200.930 3467.090 2202.110 3468.270 ;
        RECT 2200.930 3465.490 2202.110 3466.670 ;
        RECT 2200.930 3287.090 2202.110 3288.270 ;
        RECT 2200.930 3285.490 2202.110 3286.670 ;
        RECT 2200.930 3107.090 2202.110 3108.270 ;
        RECT 2200.930 3105.490 2202.110 3106.670 ;
        RECT 2200.930 2927.090 2202.110 2928.270 ;
        RECT 2200.930 2925.490 2202.110 2926.670 ;
        RECT 2200.930 2747.090 2202.110 2748.270 ;
        RECT 2200.930 2745.490 2202.110 2746.670 ;
        RECT 2200.930 2567.090 2202.110 2568.270 ;
        RECT 2200.930 2565.490 2202.110 2566.670 ;
        RECT 2200.930 2387.090 2202.110 2388.270 ;
        RECT 2200.930 2385.490 2202.110 2386.670 ;
        RECT 2200.930 2207.090 2202.110 2208.270 ;
        RECT 2200.930 2205.490 2202.110 2206.670 ;
        RECT 2200.930 2027.090 2202.110 2028.270 ;
        RECT 2200.930 2025.490 2202.110 2026.670 ;
        RECT 2200.930 1847.090 2202.110 1848.270 ;
        RECT 2200.930 1845.490 2202.110 1846.670 ;
        RECT 2200.930 1667.090 2202.110 1668.270 ;
        RECT 2200.930 1665.490 2202.110 1666.670 ;
        RECT 2200.930 1487.090 2202.110 1488.270 ;
        RECT 2200.930 1485.490 2202.110 1486.670 ;
        RECT 2200.930 1307.090 2202.110 1308.270 ;
        RECT 2200.930 1305.490 2202.110 1306.670 ;
        RECT 2200.930 1127.090 2202.110 1128.270 ;
        RECT 2200.930 1125.490 2202.110 1126.670 ;
        RECT 2200.930 947.090 2202.110 948.270 ;
        RECT 2200.930 945.490 2202.110 946.670 ;
        RECT 2200.930 767.090 2202.110 768.270 ;
        RECT 2200.930 765.490 2202.110 766.670 ;
        RECT 2200.930 587.090 2202.110 588.270 ;
        RECT 2200.930 585.490 2202.110 586.670 ;
        RECT 2200.930 407.090 2202.110 408.270 ;
        RECT 2200.930 405.490 2202.110 406.670 ;
        RECT 2200.930 227.090 2202.110 228.270 ;
        RECT 2200.930 225.490 2202.110 226.670 ;
        RECT 2200.930 47.090 2202.110 48.270 ;
        RECT 2200.930 45.490 2202.110 46.670 ;
        RECT 2200.930 -21.310 2202.110 -20.130 ;
        RECT 2200.930 -22.910 2202.110 -21.730 ;
        RECT 2380.930 3541.410 2382.110 3542.590 ;
        RECT 2380.930 3539.810 2382.110 3540.990 ;
        RECT 2380.930 3467.090 2382.110 3468.270 ;
        RECT 2380.930 3465.490 2382.110 3466.670 ;
        RECT 2380.930 3287.090 2382.110 3288.270 ;
        RECT 2380.930 3285.490 2382.110 3286.670 ;
        RECT 2380.930 3107.090 2382.110 3108.270 ;
        RECT 2380.930 3105.490 2382.110 3106.670 ;
        RECT 2380.930 2927.090 2382.110 2928.270 ;
        RECT 2380.930 2925.490 2382.110 2926.670 ;
        RECT 2380.930 2747.090 2382.110 2748.270 ;
        RECT 2380.930 2745.490 2382.110 2746.670 ;
        RECT 2380.930 2567.090 2382.110 2568.270 ;
        RECT 2380.930 2565.490 2382.110 2566.670 ;
        RECT 2380.930 2387.090 2382.110 2388.270 ;
        RECT 2380.930 2385.490 2382.110 2386.670 ;
        RECT 2380.930 2207.090 2382.110 2208.270 ;
        RECT 2380.930 2205.490 2382.110 2206.670 ;
        RECT 2380.930 2027.090 2382.110 2028.270 ;
        RECT 2380.930 2025.490 2382.110 2026.670 ;
        RECT 2380.930 1847.090 2382.110 1848.270 ;
        RECT 2380.930 1845.490 2382.110 1846.670 ;
        RECT 2380.930 1667.090 2382.110 1668.270 ;
        RECT 2380.930 1665.490 2382.110 1666.670 ;
        RECT 2380.930 1487.090 2382.110 1488.270 ;
        RECT 2380.930 1485.490 2382.110 1486.670 ;
        RECT 2380.930 1307.090 2382.110 1308.270 ;
        RECT 2380.930 1305.490 2382.110 1306.670 ;
        RECT 2380.930 1127.090 2382.110 1128.270 ;
        RECT 2380.930 1125.490 2382.110 1126.670 ;
        RECT 2380.930 947.090 2382.110 948.270 ;
        RECT 2380.930 945.490 2382.110 946.670 ;
        RECT 2380.930 767.090 2382.110 768.270 ;
        RECT 2380.930 765.490 2382.110 766.670 ;
        RECT 2380.930 587.090 2382.110 588.270 ;
        RECT 2380.930 585.490 2382.110 586.670 ;
        RECT 2380.930 407.090 2382.110 408.270 ;
        RECT 2380.930 405.490 2382.110 406.670 ;
        RECT 2380.930 227.090 2382.110 228.270 ;
        RECT 2380.930 225.490 2382.110 226.670 ;
        RECT 2380.930 47.090 2382.110 48.270 ;
        RECT 2380.930 45.490 2382.110 46.670 ;
        RECT 2380.930 -21.310 2382.110 -20.130 ;
        RECT 2380.930 -22.910 2382.110 -21.730 ;
        RECT 2560.930 3541.410 2562.110 3542.590 ;
        RECT 2560.930 3539.810 2562.110 3540.990 ;
        RECT 2560.930 3467.090 2562.110 3468.270 ;
        RECT 2560.930 3465.490 2562.110 3466.670 ;
        RECT 2560.930 3287.090 2562.110 3288.270 ;
        RECT 2560.930 3285.490 2562.110 3286.670 ;
        RECT 2560.930 3107.090 2562.110 3108.270 ;
        RECT 2560.930 3105.490 2562.110 3106.670 ;
        RECT 2560.930 2927.090 2562.110 2928.270 ;
        RECT 2560.930 2925.490 2562.110 2926.670 ;
        RECT 2560.930 2747.090 2562.110 2748.270 ;
        RECT 2560.930 2745.490 2562.110 2746.670 ;
        RECT 2560.930 2567.090 2562.110 2568.270 ;
        RECT 2560.930 2565.490 2562.110 2566.670 ;
        RECT 2560.930 2387.090 2562.110 2388.270 ;
        RECT 2560.930 2385.490 2562.110 2386.670 ;
        RECT 2560.930 2207.090 2562.110 2208.270 ;
        RECT 2560.930 2205.490 2562.110 2206.670 ;
        RECT 2560.930 2027.090 2562.110 2028.270 ;
        RECT 2560.930 2025.490 2562.110 2026.670 ;
        RECT 2560.930 1847.090 2562.110 1848.270 ;
        RECT 2560.930 1845.490 2562.110 1846.670 ;
        RECT 2560.930 1667.090 2562.110 1668.270 ;
        RECT 2560.930 1665.490 2562.110 1666.670 ;
        RECT 2560.930 1487.090 2562.110 1488.270 ;
        RECT 2560.930 1485.490 2562.110 1486.670 ;
        RECT 2560.930 1307.090 2562.110 1308.270 ;
        RECT 2560.930 1305.490 2562.110 1306.670 ;
        RECT 2560.930 1127.090 2562.110 1128.270 ;
        RECT 2560.930 1125.490 2562.110 1126.670 ;
        RECT 2560.930 947.090 2562.110 948.270 ;
        RECT 2560.930 945.490 2562.110 946.670 ;
        RECT 2560.930 767.090 2562.110 768.270 ;
        RECT 2560.930 765.490 2562.110 766.670 ;
        RECT 2560.930 587.090 2562.110 588.270 ;
        RECT 2560.930 585.490 2562.110 586.670 ;
        RECT 2560.930 407.090 2562.110 408.270 ;
        RECT 2560.930 405.490 2562.110 406.670 ;
        RECT 2560.930 227.090 2562.110 228.270 ;
        RECT 2560.930 225.490 2562.110 226.670 ;
        RECT 2560.930 47.090 2562.110 48.270 ;
        RECT 2560.930 45.490 2562.110 46.670 ;
        RECT 2560.930 -21.310 2562.110 -20.130 ;
        RECT 2560.930 -22.910 2562.110 -21.730 ;
        RECT 2740.930 3541.410 2742.110 3542.590 ;
        RECT 2740.930 3539.810 2742.110 3540.990 ;
        RECT 2740.930 3467.090 2742.110 3468.270 ;
        RECT 2740.930 3465.490 2742.110 3466.670 ;
        RECT 2740.930 3287.090 2742.110 3288.270 ;
        RECT 2740.930 3285.490 2742.110 3286.670 ;
        RECT 2740.930 3107.090 2742.110 3108.270 ;
        RECT 2740.930 3105.490 2742.110 3106.670 ;
        RECT 2740.930 2927.090 2742.110 2928.270 ;
        RECT 2740.930 2925.490 2742.110 2926.670 ;
        RECT 2740.930 2747.090 2742.110 2748.270 ;
        RECT 2740.930 2745.490 2742.110 2746.670 ;
        RECT 2740.930 2567.090 2742.110 2568.270 ;
        RECT 2740.930 2565.490 2742.110 2566.670 ;
        RECT 2740.930 2387.090 2742.110 2388.270 ;
        RECT 2740.930 2385.490 2742.110 2386.670 ;
        RECT 2740.930 2207.090 2742.110 2208.270 ;
        RECT 2740.930 2205.490 2742.110 2206.670 ;
        RECT 2740.930 2027.090 2742.110 2028.270 ;
        RECT 2740.930 2025.490 2742.110 2026.670 ;
        RECT 2740.930 1847.090 2742.110 1848.270 ;
        RECT 2740.930 1845.490 2742.110 1846.670 ;
        RECT 2740.930 1667.090 2742.110 1668.270 ;
        RECT 2740.930 1665.490 2742.110 1666.670 ;
        RECT 2740.930 1487.090 2742.110 1488.270 ;
        RECT 2740.930 1485.490 2742.110 1486.670 ;
        RECT 2740.930 1307.090 2742.110 1308.270 ;
        RECT 2740.930 1305.490 2742.110 1306.670 ;
        RECT 2740.930 1127.090 2742.110 1128.270 ;
        RECT 2740.930 1125.490 2742.110 1126.670 ;
        RECT 2740.930 947.090 2742.110 948.270 ;
        RECT 2740.930 945.490 2742.110 946.670 ;
        RECT 2740.930 767.090 2742.110 768.270 ;
        RECT 2740.930 765.490 2742.110 766.670 ;
        RECT 2740.930 587.090 2742.110 588.270 ;
        RECT 2740.930 585.490 2742.110 586.670 ;
        RECT 2740.930 407.090 2742.110 408.270 ;
        RECT 2740.930 405.490 2742.110 406.670 ;
        RECT 2740.930 227.090 2742.110 228.270 ;
        RECT 2740.930 225.490 2742.110 226.670 ;
        RECT 2740.930 47.090 2742.110 48.270 ;
        RECT 2740.930 45.490 2742.110 46.670 ;
        RECT 2740.930 -21.310 2742.110 -20.130 ;
        RECT 2740.930 -22.910 2742.110 -21.730 ;
        RECT 2945.910 3541.410 2947.090 3542.590 ;
        RECT 2945.910 3539.810 2947.090 3540.990 ;
        RECT 2945.910 3467.090 2947.090 3468.270 ;
        RECT 2945.910 3465.490 2947.090 3466.670 ;
        RECT 2945.910 3287.090 2947.090 3288.270 ;
        RECT 2945.910 3285.490 2947.090 3286.670 ;
        RECT 2945.910 3107.090 2947.090 3108.270 ;
        RECT 2945.910 3105.490 2947.090 3106.670 ;
        RECT 2945.910 2927.090 2947.090 2928.270 ;
        RECT 2945.910 2925.490 2947.090 2926.670 ;
        RECT 2945.910 2747.090 2947.090 2748.270 ;
        RECT 2945.910 2745.490 2947.090 2746.670 ;
        RECT 2945.910 2567.090 2947.090 2568.270 ;
        RECT 2945.910 2565.490 2947.090 2566.670 ;
        RECT 2945.910 2387.090 2947.090 2388.270 ;
        RECT 2945.910 2385.490 2947.090 2386.670 ;
        RECT 2945.910 2207.090 2947.090 2208.270 ;
        RECT 2945.910 2205.490 2947.090 2206.670 ;
        RECT 2945.910 2027.090 2947.090 2028.270 ;
        RECT 2945.910 2025.490 2947.090 2026.670 ;
        RECT 2945.910 1847.090 2947.090 1848.270 ;
        RECT 2945.910 1845.490 2947.090 1846.670 ;
        RECT 2945.910 1667.090 2947.090 1668.270 ;
        RECT 2945.910 1665.490 2947.090 1666.670 ;
        RECT 2945.910 1487.090 2947.090 1488.270 ;
        RECT 2945.910 1485.490 2947.090 1486.670 ;
        RECT 2945.910 1307.090 2947.090 1308.270 ;
        RECT 2945.910 1305.490 2947.090 1306.670 ;
        RECT 2945.910 1127.090 2947.090 1128.270 ;
        RECT 2945.910 1125.490 2947.090 1126.670 ;
        RECT 2945.910 947.090 2947.090 948.270 ;
        RECT 2945.910 945.490 2947.090 946.670 ;
        RECT 2945.910 767.090 2947.090 768.270 ;
        RECT 2945.910 765.490 2947.090 766.670 ;
        RECT 2945.910 587.090 2947.090 588.270 ;
        RECT 2945.910 585.490 2947.090 586.670 ;
        RECT 2945.910 407.090 2947.090 408.270 ;
        RECT 2945.910 405.490 2947.090 406.670 ;
        RECT 2945.910 227.090 2947.090 228.270 ;
        RECT 2945.910 225.490 2947.090 226.670 ;
        RECT 2945.910 47.090 2947.090 48.270 ;
        RECT 2945.910 45.490 2947.090 46.670 ;
        RECT 2945.910 -21.310 2947.090 -20.130 ;
        RECT 2945.910 -22.910 2947.090 -21.730 ;
      LAYER met5 ;
        RECT -28.380 3542.700 -25.380 3542.710 ;
        RECT 40.020 3542.700 43.020 3542.710 ;
        RECT 220.020 3542.700 223.020 3542.710 ;
        RECT 400.020 3542.700 403.020 3542.710 ;
        RECT 580.020 3542.700 583.020 3542.710 ;
        RECT 760.020 3542.700 763.020 3542.710 ;
        RECT 940.020 3542.700 943.020 3542.710 ;
        RECT 1120.020 3542.700 1123.020 3542.710 ;
        RECT 1300.020 3542.700 1303.020 3542.710 ;
        RECT 1480.020 3542.700 1483.020 3542.710 ;
        RECT 1660.020 3542.700 1663.020 3542.710 ;
        RECT 1840.020 3542.700 1843.020 3542.710 ;
        RECT 2020.020 3542.700 2023.020 3542.710 ;
        RECT 2200.020 3542.700 2203.020 3542.710 ;
        RECT 2380.020 3542.700 2383.020 3542.710 ;
        RECT 2560.020 3542.700 2563.020 3542.710 ;
        RECT 2740.020 3542.700 2743.020 3542.710 ;
        RECT 2945.000 3542.700 2948.000 3542.710 ;
        RECT -28.380 3539.700 2948.000 3542.700 ;
        RECT -28.380 3539.690 -25.380 3539.700 ;
        RECT 40.020 3539.690 43.020 3539.700 ;
        RECT 220.020 3539.690 223.020 3539.700 ;
        RECT 400.020 3539.690 403.020 3539.700 ;
        RECT 580.020 3539.690 583.020 3539.700 ;
        RECT 760.020 3539.690 763.020 3539.700 ;
        RECT 940.020 3539.690 943.020 3539.700 ;
        RECT 1120.020 3539.690 1123.020 3539.700 ;
        RECT 1300.020 3539.690 1303.020 3539.700 ;
        RECT 1480.020 3539.690 1483.020 3539.700 ;
        RECT 1660.020 3539.690 1663.020 3539.700 ;
        RECT 1840.020 3539.690 1843.020 3539.700 ;
        RECT 2020.020 3539.690 2023.020 3539.700 ;
        RECT 2200.020 3539.690 2203.020 3539.700 ;
        RECT 2380.020 3539.690 2383.020 3539.700 ;
        RECT 2560.020 3539.690 2563.020 3539.700 ;
        RECT 2740.020 3539.690 2743.020 3539.700 ;
        RECT 2945.000 3539.690 2948.000 3539.700 ;
        RECT -28.380 3468.380 -25.380 3468.390 ;
        RECT 40.020 3468.380 43.020 3468.390 ;
        RECT 220.020 3468.380 223.020 3468.390 ;
        RECT 400.020 3468.380 403.020 3468.390 ;
        RECT 580.020 3468.380 583.020 3468.390 ;
        RECT 760.020 3468.380 763.020 3468.390 ;
        RECT 940.020 3468.380 943.020 3468.390 ;
        RECT 1120.020 3468.380 1123.020 3468.390 ;
        RECT 1300.020 3468.380 1303.020 3468.390 ;
        RECT 1480.020 3468.380 1483.020 3468.390 ;
        RECT 1660.020 3468.380 1663.020 3468.390 ;
        RECT 1840.020 3468.380 1843.020 3468.390 ;
        RECT 2020.020 3468.380 2023.020 3468.390 ;
        RECT 2200.020 3468.380 2203.020 3468.390 ;
        RECT 2380.020 3468.380 2383.020 3468.390 ;
        RECT 2560.020 3468.380 2563.020 3468.390 ;
        RECT 2740.020 3468.380 2743.020 3468.390 ;
        RECT 2945.000 3468.380 2948.000 3468.390 ;
        RECT -32.980 3465.380 2952.600 3468.380 ;
        RECT -28.380 3465.370 -25.380 3465.380 ;
        RECT 40.020 3465.370 43.020 3465.380 ;
        RECT 220.020 3465.370 223.020 3465.380 ;
        RECT 400.020 3465.370 403.020 3465.380 ;
        RECT 580.020 3465.370 583.020 3465.380 ;
        RECT 760.020 3465.370 763.020 3465.380 ;
        RECT 940.020 3465.370 943.020 3465.380 ;
        RECT 1120.020 3465.370 1123.020 3465.380 ;
        RECT 1300.020 3465.370 1303.020 3465.380 ;
        RECT 1480.020 3465.370 1483.020 3465.380 ;
        RECT 1660.020 3465.370 1663.020 3465.380 ;
        RECT 1840.020 3465.370 1843.020 3465.380 ;
        RECT 2020.020 3465.370 2023.020 3465.380 ;
        RECT 2200.020 3465.370 2203.020 3465.380 ;
        RECT 2380.020 3465.370 2383.020 3465.380 ;
        RECT 2560.020 3465.370 2563.020 3465.380 ;
        RECT 2740.020 3465.370 2743.020 3465.380 ;
        RECT 2945.000 3465.370 2948.000 3465.380 ;
        RECT -28.380 3288.380 -25.380 3288.390 ;
        RECT 40.020 3288.380 43.020 3288.390 ;
        RECT 220.020 3288.380 223.020 3288.390 ;
        RECT 400.020 3288.380 403.020 3288.390 ;
        RECT 580.020 3288.380 583.020 3288.390 ;
        RECT 760.020 3288.380 763.020 3288.390 ;
        RECT 940.020 3288.380 943.020 3288.390 ;
        RECT 1120.020 3288.380 1123.020 3288.390 ;
        RECT 1300.020 3288.380 1303.020 3288.390 ;
        RECT 1480.020 3288.380 1483.020 3288.390 ;
        RECT 1660.020 3288.380 1663.020 3288.390 ;
        RECT 1840.020 3288.380 1843.020 3288.390 ;
        RECT 2020.020 3288.380 2023.020 3288.390 ;
        RECT 2200.020 3288.380 2203.020 3288.390 ;
        RECT 2380.020 3288.380 2383.020 3288.390 ;
        RECT 2560.020 3288.380 2563.020 3288.390 ;
        RECT 2740.020 3288.380 2743.020 3288.390 ;
        RECT 2945.000 3288.380 2948.000 3288.390 ;
        RECT -32.980 3285.380 2952.600 3288.380 ;
        RECT -28.380 3285.370 -25.380 3285.380 ;
        RECT 40.020 3285.370 43.020 3285.380 ;
        RECT 220.020 3285.370 223.020 3285.380 ;
        RECT 400.020 3285.370 403.020 3285.380 ;
        RECT 580.020 3285.370 583.020 3285.380 ;
        RECT 760.020 3285.370 763.020 3285.380 ;
        RECT 940.020 3285.370 943.020 3285.380 ;
        RECT 1120.020 3285.370 1123.020 3285.380 ;
        RECT 1300.020 3285.370 1303.020 3285.380 ;
        RECT 1480.020 3285.370 1483.020 3285.380 ;
        RECT 1660.020 3285.370 1663.020 3285.380 ;
        RECT 1840.020 3285.370 1843.020 3285.380 ;
        RECT 2020.020 3285.370 2023.020 3285.380 ;
        RECT 2200.020 3285.370 2203.020 3285.380 ;
        RECT 2380.020 3285.370 2383.020 3285.380 ;
        RECT 2560.020 3285.370 2563.020 3285.380 ;
        RECT 2740.020 3285.370 2743.020 3285.380 ;
        RECT 2945.000 3285.370 2948.000 3285.380 ;
        RECT -28.380 3108.380 -25.380 3108.390 ;
        RECT 40.020 3108.380 43.020 3108.390 ;
        RECT 220.020 3108.380 223.020 3108.390 ;
        RECT 400.020 3108.380 403.020 3108.390 ;
        RECT 580.020 3108.380 583.020 3108.390 ;
        RECT 760.020 3108.380 763.020 3108.390 ;
        RECT 940.020 3108.380 943.020 3108.390 ;
        RECT 1120.020 3108.380 1123.020 3108.390 ;
        RECT 1300.020 3108.380 1303.020 3108.390 ;
        RECT 1480.020 3108.380 1483.020 3108.390 ;
        RECT 1660.020 3108.380 1663.020 3108.390 ;
        RECT 1840.020 3108.380 1843.020 3108.390 ;
        RECT 2020.020 3108.380 2023.020 3108.390 ;
        RECT 2200.020 3108.380 2203.020 3108.390 ;
        RECT 2380.020 3108.380 2383.020 3108.390 ;
        RECT 2560.020 3108.380 2563.020 3108.390 ;
        RECT 2740.020 3108.380 2743.020 3108.390 ;
        RECT 2945.000 3108.380 2948.000 3108.390 ;
        RECT -32.980 3105.380 2952.600 3108.380 ;
        RECT -28.380 3105.370 -25.380 3105.380 ;
        RECT 40.020 3105.370 43.020 3105.380 ;
        RECT 220.020 3105.370 223.020 3105.380 ;
        RECT 400.020 3105.370 403.020 3105.380 ;
        RECT 580.020 3105.370 583.020 3105.380 ;
        RECT 760.020 3105.370 763.020 3105.380 ;
        RECT 940.020 3105.370 943.020 3105.380 ;
        RECT 1120.020 3105.370 1123.020 3105.380 ;
        RECT 1300.020 3105.370 1303.020 3105.380 ;
        RECT 1480.020 3105.370 1483.020 3105.380 ;
        RECT 1660.020 3105.370 1663.020 3105.380 ;
        RECT 1840.020 3105.370 1843.020 3105.380 ;
        RECT 2020.020 3105.370 2023.020 3105.380 ;
        RECT 2200.020 3105.370 2203.020 3105.380 ;
        RECT 2380.020 3105.370 2383.020 3105.380 ;
        RECT 2560.020 3105.370 2563.020 3105.380 ;
        RECT 2740.020 3105.370 2743.020 3105.380 ;
        RECT 2945.000 3105.370 2948.000 3105.380 ;
        RECT -28.380 2928.380 -25.380 2928.390 ;
        RECT 40.020 2928.380 43.020 2928.390 ;
        RECT 220.020 2928.380 223.020 2928.390 ;
        RECT 400.020 2928.380 403.020 2928.390 ;
        RECT 580.020 2928.380 583.020 2928.390 ;
        RECT 760.020 2928.380 763.020 2928.390 ;
        RECT 940.020 2928.380 943.020 2928.390 ;
        RECT 1120.020 2928.380 1123.020 2928.390 ;
        RECT 1300.020 2928.380 1303.020 2928.390 ;
        RECT 1480.020 2928.380 1483.020 2928.390 ;
        RECT 1660.020 2928.380 1663.020 2928.390 ;
        RECT 1840.020 2928.380 1843.020 2928.390 ;
        RECT 2020.020 2928.380 2023.020 2928.390 ;
        RECT 2200.020 2928.380 2203.020 2928.390 ;
        RECT 2380.020 2928.380 2383.020 2928.390 ;
        RECT 2560.020 2928.380 2563.020 2928.390 ;
        RECT 2740.020 2928.380 2743.020 2928.390 ;
        RECT 2945.000 2928.380 2948.000 2928.390 ;
        RECT -32.980 2925.380 2952.600 2928.380 ;
        RECT -28.380 2925.370 -25.380 2925.380 ;
        RECT 40.020 2925.370 43.020 2925.380 ;
        RECT 220.020 2925.370 223.020 2925.380 ;
        RECT 400.020 2925.370 403.020 2925.380 ;
        RECT 580.020 2925.370 583.020 2925.380 ;
        RECT 760.020 2925.370 763.020 2925.380 ;
        RECT 940.020 2925.370 943.020 2925.380 ;
        RECT 1120.020 2925.370 1123.020 2925.380 ;
        RECT 1300.020 2925.370 1303.020 2925.380 ;
        RECT 1480.020 2925.370 1483.020 2925.380 ;
        RECT 1660.020 2925.370 1663.020 2925.380 ;
        RECT 1840.020 2925.370 1843.020 2925.380 ;
        RECT 2020.020 2925.370 2023.020 2925.380 ;
        RECT 2200.020 2925.370 2203.020 2925.380 ;
        RECT 2380.020 2925.370 2383.020 2925.380 ;
        RECT 2560.020 2925.370 2563.020 2925.380 ;
        RECT 2740.020 2925.370 2743.020 2925.380 ;
        RECT 2945.000 2925.370 2948.000 2925.380 ;
        RECT -28.380 2748.380 -25.380 2748.390 ;
        RECT 40.020 2748.380 43.020 2748.390 ;
        RECT 220.020 2748.380 223.020 2748.390 ;
        RECT 400.020 2748.380 403.020 2748.390 ;
        RECT 580.020 2748.380 583.020 2748.390 ;
        RECT 760.020 2748.380 763.020 2748.390 ;
        RECT 940.020 2748.380 943.020 2748.390 ;
        RECT 1120.020 2748.380 1123.020 2748.390 ;
        RECT 1300.020 2748.380 1303.020 2748.390 ;
        RECT 1480.020 2748.380 1483.020 2748.390 ;
        RECT 1660.020 2748.380 1663.020 2748.390 ;
        RECT 1840.020 2748.380 1843.020 2748.390 ;
        RECT 2020.020 2748.380 2023.020 2748.390 ;
        RECT 2200.020 2748.380 2203.020 2748.390 ;
        RECT 2380.020 2748.380 2383.020 2748.390 ;
        RECT 2560.020 2748.380 2563.020 2748.390 ;
        RECT 2740.020 2748.380 2743.020 2748.390 ;
        RECT 2945.000 2748.380 2948.000 2748.390 ;
        RECT -32.980 2745.380 2952.600 2748.380 ;
        RECT -28.380 2745.370 -25.380 2745.380 ;
        RECT 40.020 2745.370 43.020 2745.380 ;
        RECT 220.020 2745.370 223.020 2745.380 ;
        RECT 400.020 2745.370 403.020 2745.380 ;
        RECT 580.020 2745.370 583.020 2745.380 ;
        RECT 760.020 2745.370 763.020 2745.380 ;
        RECT 940.020 2745.370 943.020 2745.380 ;
        RECT 1120.020 2745.370 1123.020 2745.380 ;
        RECT 1300.020 2745.370 1303.020 2745.380 ;
        RECT 1480.020 2745.370 1483.020 2745.380 ;
        RECT 1660.020 2745.370 1663.020 2745.380 ;
        RECT 1840.020 2745.370 1843.020 2745.380 ;
        RECT 2020.020 2745.370 2023.020 2745.380 ;
        RECT 2200.020 2745.370 2203.020 2745.380 ;
        RECT 2380.020 2745.370 2383.020 2745.380 ;
        RECT 2560.020 2745.370 2563.020 2745.380 ;
        RECT 2740.020 2745.370 2743.020 2745.380 ;
        RECT 2945.000 2745.370 2948.000 2745.380 ;
        RECT -28.380 2568.380 -25.380 2568.390 ;
        RECT 40.020 2568.380 43.020 2568.390 ;
        RECT 220.020 2568.380 223.020 2568.390 ;
        RECT 400.020 2568.380 403.020 2568.390 ;
        RECT 580.020 2568.380 583.020 2568.390 ;
        RECT 760.020 2568.380 763.020 2568.390 ;
        RECT 940.020 2568.380 943.020 2568.390 ;
        RECT 1120.020 2568.380 1123.020 2568.390 ;
        RECT 1300.020 2568.380 1303.020 2568.390 ;
        RECT 1480.020 2568.380 1483.020 2568.390 ;
        RECT 1660.020 2568.380 1663.020 2568.390 ;
        RECT 1840.020 2568.380 1843.020 2568.390 ;
        RECT 2020.020 2568.380 2023.020 2568.390 ;
        RECT 2200.020 2568.380 2203.020 2568.390 ;
        RECT 2380.020 2568.380 2383.020 2568.390 ;
        RECT 2560.020 2568.380 2563.020 2568.390 ;
        RECT 2740.020 2568.380 2743.020 2568.390 ;
        RECT 2945.000 2568.380 2948.000 2568.390 ;
        RECT -32.980 2565.380 2952.600 2568.380 ;
        RECT -28.380 2565.370 -25.380 2565.380 ;
        RECT 40.020 2565.370 43.020 2565.380 ;
        RECT 220.020 2565.370 223.020 2565.380 ;
        RECT 400.020 2565.370 403.020 2565.380 ;
        RECT 580.020 2565.370 583.020 2565.380 ;
        RECT 760.020 2565.370 763.020 2565.380 ;
        RECT 940.020 2565.370 943.020 2565.380 ;
        RECT 1120.020 2565.370 1123.020 2565.380 ;
        RECT 1300.020 2565.370 1303.020 2565.380 ;
        RECT 1480.020 2565.370 1483.020 2565.380 ;
        RECT 1660.020 2565.370 1663.020 2565.380 ;
        RECT 1840.020 2565.370 1843.020 2565.380 ;
        RECT 2020.020 2565.370 2023.020 2565.380 ;
        RECT 2200.020 2565.370 2203.020 2565.380 ;
        RECT 2380.020 2565.370 2383.020 2565.380 ;
        RECT 2560.020 2565.370 2563.020 2565.380 ;
        RECT 2740.020 2565.370 2743.020 2565.380 ;
        RECT 2945.000 2565.370 2948.000 2565.380 ;
        RECT -28.380 2388.380 -25.380 2388.390 ;
        RECT 40.020 2388.380 43.020 2388.390 ;
        RECT 220.020 2388.380 223.020 2388.390 ;
        RECT 400.020 2388.380 403.020 2388.390 ;
        RECT 580.020 2388.380 583.020 2388.390 ;
        RECT 760.020 2388.380 763.020 2388.390 ;
        RECT 940.020 2388.380 943.020 2388.390 ;
        RECT 1120.020 2388.380 1123.020 2388.390 ;
        RECT 1300.020 2388.380 1303.020 2388.390 ;
        RECT 1480.020 2388.380 1483.020 2388.390 ;
        RECT 1660.020 2388.380 1663.020 2388.390 ;
        RECT 1840.020 2388.380 1843.020 2388.390 ;
        RECT 2020.020 2388.380 2023.020 2388.390 ;
        RECT 2200.020 2388.380 2203.020 2388.390 ;
        RECT 2380.020 2388.380 2383.020 2388.390 ;
        RECT 2560.020 2388.380 2563.020 2388.390 ;
        RECT 2740.020 2388.380 2743.020 2388.390 ;
        RECT 2945.000 2388.380 2948.000 2388.390 ;
        RECT -32.980 2385.380 2952.600 2388.380 ;
        RECT -28.380 2385.370 -25.380 2385.380 ;
        RECT 40.020 2385.370 43.020 2385.380 ;
        RECT 220.020 2385.370 223.020 2385.380 ;
        RECT 400.020 2385.370 403.020 2385.380 ;
        RECT 580.020 2385.370 583.020 2385.380 ;
        RECT 760.020 2385.370 763.020 2385.380 ;
        RECT 940.020 2385.370 943.020 2385.380 ;
        RECT 1120.020 2385.370 1123.020 2385.380 ;
        RECT 1300.020 2385.370 1303.020 2385.380 ;
        RECT 1480.020 2385.370 1483.020 2385.380 ;
        RECT 1660.020 2385.370 1663.020 2385.380 ;
        RECT 1840.020 2385.370 1843.020 2385.380 ;
        RECT 2020.020 2385.370 2023.020 2385.380 ;
        RECT 2200.020 2385.370 2203.020 2385.380 ;
        RECT 2380.020 2385.370 2383.020 2385.380 ;
        RECT 2560.020 2385.370 2563.020 2385.380 ;
        RECT 2740.020 2385.370 2743.020 2385.380 ;
        RECT 2945.000 2385.370 2948.000 2385.380 ;
        RECT -28.380 2208.380 -25.380 2208.390 ;
        RECT 40.020 2208.380 43.020 2208.390 ;
        RECT 220.020 2208.380 223.020 2208.390 ;
        RECT 400.020 2208.380 403.020 2208.390 ;
        RECT 580.020 2208.380 583.020 2208.390 ;
        RECT 760.020 2208.380 763.020 2208.390 ;
        RECT 940.020 2208.380 943.020 2208.390 ;
        RECT 1120.020 2208.380 1123.020 2208.390 ;
        RECT 1300.020 2208.380 1303.020 2208.390 ;
        RECT 1480.020 2208.380 1483.020 2208.390 ;
        RECT 1660.020 2208.380 1663.020 2208.390 ;
        RECT 1840.020 2208.380 1843.020 2208.390 ;
        RECT 2020.020 2208.380 2023.020 2208.390 ;
        RECT 2200.020 2208.380 2203.020 2208.390 ;
        RECT 2380.020 2208.380 2383.020 2208.390 ;
        RECT 2560.020 2208.380 2563.020 2208.390 ;
        RECT 2740.020 2208.380 2743.020 2208.390 ;
        RECT 2945.000 2208.380 2948.000 2208.390 ;
        RECT -32.980 2205.380 2952.600 2208.380 ;
        RECT -28.380 2205.370 -25.380 2205.380 ;
        RECT 40.020 2205.370 43.020 2205.380 ;
        RECT 220.020 2205.370 223.020 2205.380 ;
        RECT 400.020 2205.370 403.020 2205.380 ;
        RECT 580.020 2205.370 583.020 2205.380 ;
        RECT 760.020 2205.370 763.020 2205.380 ;
        RECT 940.020 2205.370 943.020 2205.380 ;
        RECT 1120.020 2205.370 1123.020 2205.380 ;
        RECT 1300.020 2205.370 1303.020 2205.380 ;
        RECT 1480.020 2205.370 1483.020 2205.380 ;
        RECT 1660.020 2205.370 1663.020 2205.380 ;
        RECT 1840.020 2205.370 1843.020 2205.380 ;
        RECT 2020.020 2205.370 2023.020 2205.380 ;
        RECT 2200.020 2205.370 2203.020 2205.380 ;
        RECT 2380.020 2205.370 2383.020 2205.380 ;
        RECT 2560.020 2205.370 2563.020 2205.380 ;
        RECT 2740.020 2205.370 2743.020 2205.380 ;
        RECT 2945.000 2205.370 2948.000 2205.380 ;
        RECT -28.380 2028.380 -25.380 2028.390 ;
        RECT 40.020 2028.380 43.020 2028.390 ;
        RECT 220.020 2028.380 223.020 2028.390 ;
        RECT 400.020 2028.380 403.020 2028.390 ;
        RECT 580.020 2028.380 583.020 2028.390 ;
        RECT 760.020 2028.380 763.020 2028.390 ;
        RECT 940.020 2028.380 943.020 2028.390 ;
        RECT 1120.020 2028.380 1123.020 2028.390 ;
        RECT 1300.020 2028.380 1303.020 2028.390 ;
        RECT 1480.020 2028.380 1483.020 2028.390 ;
        RECT 1660.020 2028.380 1663.020 2028.390 ;
        RECT 1840.020 2028.380 1843.020 2028.390 ;
        RECT 2020.020 2028.380 2023.020 2028.390 ;
        RECT 2200.020 2028.380 2203.020 2028.390 ;
        RECT 2380.020 2028.380 2383.020 2028.390 ;
        RECT 2560.020 2028.380 2563.020 2028.390 ;
        RECT 2740.020 2028.380 2743.020 2028.390 ;
        RECT 2945.000 2028.380 2948.000 2028.390 ;
        RECT -32.980 2025.380 2952.600 2028.380 ;
        RECT -28.380 2025.370 -25.380 2025.380 ;
        RECT 40.020 2025.370 43.020 2025.380 ;
        RECT 220.020 2025.370 223.020 2025.380 ;
        RECT 400.020 2025.370 403.020 2025.380 ;
        RECT 580.020 2025.370 583.020 2025.380 ;
        RECT 760.020 2025.370 763.020 2025.380 ;
        RECT 940.020 2025.370 943.020 2025.380 ;
        RECT 1120.020 2025.370 1123.020 2025.380 ;
        RECT 1300.020 2025.370 1303.020 2025.380 ;
        RECT 1480.020 2025.370 1483.020 2025.380 ;
        RECT 1660.020 2025.370 1663.020 2025.380 ;
        RECT 1840.020 2025.370 1843.020 2025.380 ;
        RECT 2020.020 2025.370 2023.020 2025.380 ;
        RECT 2200.020 2025.370 2203.020 2025.380 ;
        RECT 2380.020 2025.370 2383.020 2025.380 ;
        RECT 2560.020 2025.370 2563.020 2025.380 ;
        RECT 2740.020 2025.370 2743.020 2025.380 ;
        RECT 2945.000 2025.370 2948.000 2025.380 ;
        RECT -28.380 1848.380 -25.380 1848.390 ;
        RECT 40.020 1848.380 43.020 1848.390 ;
        RECT 220.020 1848.380 223.020 1848.390 ;
        RECT 400.020 1848.380 403.020 1848.390 ;
        RECT 580.020 1848.380 583.020 1848.390 ;
        RECT 760.020 1848.380 763.020 1848.390 ;
        RECT 940.020 1848.380 943.020 1848.390 ;
        RECT 1120.020 1848.380 1123.020 1848.390 ;
        RECT 1300.020 1848.380 1303.020 1848.390 ;
        RECT 1480.020 1848.380 1483.020 1848.390 ;
        RECT 1660.020 1848.380 1663.020 1848.390 ;
        RECT 1840.020 1848.380 1843.020 1848.390 ;
        RECT 2020.020 1848.380 2023.020 1848.390 ;
        RECT 2200.020 1848.380 2203.020 1848.390 ;
        RECT 2380.020 1848.380 2383.020 1848.390 ;
        RECT 2560.020 1848.380 2563.020 1848.390 ;
        RECT 2740.020 1848.380 2743.020 1848.390 ;
        RECT 2945.000 1848.380 2948.000 1848.390 ;
        RECT -32.980 1845.380 2952.600 1848.380 ;
        RECT -28.380 1845.370 -25.380 1845.380 ;
        RECT 40.020 1845.370 43.020 1845.380 ;
        RECT 220.020 1845.370 223.020 1845.380 ;
        RECT 400.020 1845.370 403.020 1845.380 ;
        RECT 580.020 1845.370 583.020 1845.380 ;
        RECT 760.020 1845.370 763.020 1845.380 ;
        RECT 940.020 1845.370 943.020 1845.380 ;
        RECT 1120.020 1845.370 1123.020 1845.380 ;
        RECT 1300.020 1845.370 1303.020 1845.380 ;
        RECT 1480.020 1845.370 1483.020 1845.380 ;
        RECT 1660.020 1845.370 1663.020 1845.380 ;
        RECT 1840.020 1845.370 1843.020 1845.380 ;
        RECT 2020.020 1845.370 2023.020 1845.380 ;
        RECT 2200.020 1845.370 2203.020 1845.380 ;
        RECT 2380.020 1845.370 2383.020 1845.380 ;
        RECT 2560.020 1845.370 2563.020 1845.380 ;
        RECT 2740.020 1845.370 2743.020 1845.380 ;
        RECT 2945.000 1845.370 2948.000 1845.380 ;
        RECT -28.380 1668.380 -25.380 1668.390 ;
        RECT 40.020 1668.380 43.020 1668.390 ;
        RECT 220.020 1668.380 223.020 1668.390 ;
        RECT 400.020 1668.380 403.020 1668.390 ;
        RECT 580.020 1668.380 583.020 1668.390 ;
        RECT 760.020 1668.380 763.020 1668.390 ;
        RECT 940.020 1668.380 943.020 1668.390 ;
        RECT 1120.020 1668.380 1123.020 1668.390 ;
        RECT 1300.020 1668.380 1303.020 1668.390 ;
        RECT 1480.020 1668.380 1483.020 1668.390 ;
        RECT 1660.020 1668.380 1663.020 1668.390 ;
        RECT 1840.020 1668.380 1843.020 1668.390 ;
        RECT 2020.020 1668.380 2023.020 1668.390 ;
        RECT 2200.020 1668.380 2203.020 1668.390 ;
        RECT 2380.020 1668.380 2383.020 1668.390 ;
        RECT 2560.020 1668.380 2563.020 1668.390 ;
        RECT 2740.020 1668.380 2743.020 1668.390 ;
        RECT 2945.000 1668.380 2948.000 1668.390 ;
        RECT -32.980 1665.380 2952.600 1668.380 ;
        RECT -28.380 1665.370 -25.380 1665.380 ;
        RECT 40.020 1665.370 43.020 1665.380 ;
        RECT 220.020 1665.370 223.020 1665.380 ;
        RECT 400.020 1665.370 403.020 1665.380 ;
        RECT 580.020 1665.370 583.020 1665.380 ;
        RECT 760.020 1665.370 763.020 1665.380 ;
        RECT 940.020 1665.370 943.020 1665.380 ;
        RECT 1120.020 1665.370 1123.020 1665.380 ;
        RECT 1300.020 1665.370 1303.020 1665.380 ;
        RECT 1480.020 1665.370 1483.020 1665.380 ;
        RECT 1660.020 1665.370 1663.020 1665.380 ;
        RECT 1840.020 1665.370 1843.020 1665.380 ;
        RECT 2020.020 1665.370 2023.020 1665.380 ;
        RECT 2200.020 1665.370 2203.020 1665.380 ;
        RECT 2380.020 1665.370 2383.020 1665.380 ;
        RECT 2560.020 1665.370 2563.020 1665.380 ;
        RECT 2740.020 1665.370 2743.020 1665.380 ;
        RECT 2945.000 1665.370 2948.000 1665.380 ;
        RECT -28.380 1488.380 -25.380 1488.390 ;
        RECT 40.020 1488.380 43.020 1488.390 ;
        RECT 220.020 1488.380 223.020 1488.390 ;
        RECT 400.020 1488.380 403.020 1488.390 ;
        RECT 580.020 1488.380 583.020 1488.390 ;
        RECT 760.020 1488.380 763.020 1488.390 ;
        RECT 940.020 1488.380 943.020 1488.390 ;
        RECT 1120.020 1488.380 1123.020 1488.390 ;
        RECT 1300.020 1488.380 1303.020 1488.390 ;
        RECT 1480.020 1488.380 1483.020 1488.390 ;
        RECT 1660.020 1488.380 1663.020 1488.390 ;
        RECT 1840.020 1488.380 1843.020 1488.390 ;
        RECT 2020.020 1488.380 2023.020 1488.390 ;
        RECT 2200.020 1488.380 2203.020 1488.390 ;
        RECT 2380.020 1488.380 2383.020 1488.390 ;
        RECT 2560.020 1488.380 2563.020 1488.390 ;
        RECT 2740.020 1488.380 2743.020 1488.390 ;
        RECT 2945.000 1488.380 2948.000 1488.390 ;
        RECT -32.980 1485.380 2952.600 1488.380 ;
        RECT -28.380 1485.370 -25.380 1485.380 ;
        RECT 40.020 1485.370 43.020 1485.380 ;
        RECT 220.020 1485.370 223.020 1485.380 ;
        RECT 400.020 1485.370 403.020 1485.380 ;
        RECT 580.020 1485.370 583.020 1485.380 ;
        RECT 760.020 1485.370 763.020 1485.380 ;
        RECT 940.020 1485.370 943.020 1485.380 ;
        RECT 1120.020 1485.370 1123.020 1485.380 ;
        RECT 1300.020 1485.370 1303.020 1485.380 ;
        RECT 1480.020 1485.370 1483.020 1485.380 ;
        RECT 1660.020 1485.370 1663.020 1485.380 ;
        RECT 1840.020 1485.370 1843.020 1485.380 ;
        RECT 2020.020 1485.370 2023.020 1485.380 ;
        RECT 2200.020 1485.370 2203.020 1485.380 ;
        RECT 2380.020 1485.370 2383.020 1485.380 ;
        RECT 2560.020 1485.370 2563.020 1485.380 ;
        RECT 2740.020 1485.370 2743.020 1485.380 ;
        RECT 2945.000 1485.370 2948.000 1485.380 ;
        RECT -28.380 1308.380 -25.380 1308.390 ;
        RECT 40.020 1308.380 43.020 1308.390 ;
        RECT 220.020 1308.380 223.020 1308.390 ;
        RECT 400.020 1308.380 403.020 1308.390 ;
        RECT 580.020 1308.380 583.020 1308.390 ;
        RECT 760.020 1308.380 763.020 1308.390 ;
        RECT 940.020 1308.380 943.020 1308.390 ;
        RECT 1120.020 1308.380 1123.020 1308.390 ;
        RECT 1300.020 1308.380 1303.020 1308.390 ;
        RECT 1480.020 1308.380 1483.020 1308.390 ;
        RECT 1660.020 1308.380 1663.020 1308.390 ;
        RECT 1840.020 1308.380 1843.020 1308.390 ;
        RECT 2020.020 1308.380 2023.020 1308.390 ;
        RECT 2200.020 1308.380 2203.020 1308.390 ;
        RECT 2380.020 1308.380 2383.020 1308.390 ;
        RECT 2560.020 1308.380 2563.020 1308.390 ;
        RECT 2740.020 1308.380 2743.020 1308.390 ;
        RECT 2945.000 1308.380 2948.000 1308.390 ;
        RECT -32.980 1305.380 2952.600 1308.380 ;
        RECT -28.380 1305.370 -25.380 1305.380 ;
        RECT 40.020 1305.370 43.020 1305.380 ;
        RECT 220.020 1305.370 223.020 1305.380 ;
        RECT 400.020 1305.370 403.020 1305.380 ;
        RECT 580.020 1305.370 583.020 1305.380 ;
        RECT 760.020 1305.370 763.020 1305.380 ;
        RECT 940.020 1305.370 943.020 1305.380 ;
        RECT 1120.020 1305.370 1123.020 1305.380 ;
        RECT 1300.020 1305.370 1303.020 1305.380 ;
        RECT 1480.020 1305.370 1483.020 1305.380 ;
        RECT 1660.020 1305.370 1663.020 1305.380 ;
        RECT 1840.020 1305.370 1843.020 1305.380 ;
        RECT 2020.020 1305.370 2023.020 1305.380 ;
        RECT 2200.020 1305.370 2203.020 1305.380 ;
        RECT 2380.020 1305.370 2383.020 1305.380 ;
        RECT 2560.020 1305.370 2563.020 1305.380 ;
        RECT 2740.020 1305.370 2743.020 1305.380 ;
        RECT 2945.000 1305.370 2948.000 1305.380 ;
        RECT -28.380 1128.380 -25.380 1128.390 ;
        RECT 40.020 1128.380 43.020 1128.390 ;
        RECT 220.020 1128.380 223.020 1128.390 ;
        RECT 400.020 1128.380 403.020 1128.390 ;
        RECT 580.020 1128.380 583.020 1128.390 ;
        RECT 760.020 1128.380 763.020 1128.390 ;
        RECT 940.020 1128.380 943.020 1128.390 ;
        RECT 1120.020 1128.380 1123.020 1128.390 ;
        RECT 1300.020 1128.380 1303.020 1128.390 ;
        RECT 1480.020 1128.380 1483.020 1128.390 ;
        RECT 1660.020 1128.380 1663.020 1128.390 ;
        RECT 1840.020 1128.380 1843.020 1128.390 ;
        RECT 2020.020 1128.380 2023.020 1128.390 ;
        RECT 2200.020 1128.380 2203.020 1128.390 ;
        RECT 2380.020 1128.380 2383.020 1128.390 ;
        RECT 2560.020 1128.380 2563.020 1128.390 ;
        RECT 2740.020 1128.380 2743.020 1128.390 ;
        RECT 2945.000 1128.380 2948.000 1128.390 ;
        RECT -32.980 1125.380 2952.600 1128.380 ;
        RECT -28.380 1125.370 -25.380 1125.380 ;
        RECT 40.020 1125.370 43.020 1125.380 ;
        RECT 220.020 1125.370 223.020 1125.380 ;
        RECT 400.020 1125.370 403.020 1125.380 ;
        RECT 580.020 1125.370 583.020 1125.380 ;
        RECT 760.020 1125.370 763.020 1125.380 ;
        RECT 940.020 1125.370 943.020 1125.380 ;
        RECT 1120.020 1125.370 1123.020 1125.380 ;
        RECT 1300.020 1125.370 1303.020 1125.380 ;
        RECT 1480.020 1125.370 1483.020 1125.380 ;
        RECT 1660.020 1125.370 1663.020 1125.380 ;
        RECT 1840.020 1125.370 1843.020 1125.380 ;
        RECT 2020.020 1125.370 2023.020 1125.380 ;
        RECT 2200.020 1125.370 2203.020 1125.380 ;
        RECT 2380.020 1125.370 2383.020 1125.380 ;
        RECT 2560.020 1125.370 2563.020 1125.380 ;
        RECT 2740.020 1125.370 2743.020 1125.380 ;
        RECT 2945.000 1125.370 2948.000 1125.380 ;
        RECT -28.380 948.380 -25.380 948.390 ;
        RECT 40.020 948.380 43.020 948.390 ;
        RECT 220.020 948.380 223.020 948.390 ;
        RECT 400.020 948.380 403.020 948.390 ;
        RECT 580.020 948.380 583.020 948.390 ;
        RECT 760.020 948.380 763.020 948.390 ;
        RECT 940.020 948.380 943.020 948.390 ;
        RECT 1120.020 948.380 1123.020 948.390 ;
        RECT 1300.020 948.380 1303.020 948.390 ;
        RECT 1480.020 948.380 1483.020 948.390 ;
        RECT 1660.020 948.380 1663.020 948.390 ;
        RECT 1840.020 948.380 1843.020 948.390 ;
        RECT 2020.020 948.380 2023.020 948.390 ;
        RECT 2200.020 948.380 2203.020 948.390 ;
        RECT 2380.020 948.380 2383.020 948.390 ;
        RECT 2560.020 948.380 2563.020 948.390 ;
        RECT 2740.020 948.380 2743.020 948.390 ;
        RECT 2945.000 948.380 2948.000 948.390 ;
        RECT -32.980 945.380 2952.600 948.380 ;
        RECT -28.380 945.370 -25.380 945.380 ;
        RECT 40.020 945.370 43.020 945.380 ;
        RECT 220.020 945.370 223.020 945.380 ;
        RECT 400.020 945.370 403.020 945.380 ;
        RECT 580.020 945.370 583.020 945.380 ;
        RECT 760.020 945.370 763.020 945.380 ;
        RECT 940.020 945.370 943.020 945.380 ;
        RECT 1120.020 945.370 1123.020 945.380 ;
        RECT 1300.020 945.370 1303.020 945.380 ;
        RECT 1480.020 945.370 1483.020 945.380 ;
        RECT 1660.020 945.370 1663.020 945.380 ;
        RECT 1840.020 945.370 1843.020 945.380 ;
        RECT 2020.020 945.370 2023.020 945.380 ;
        RECT 2200.020 945.370 2203.020 945.380 ;
        RECT 2380.020 945.370 2383.020 945.380 ;
        RECT 2560.020 945.370 2563.020 945.380 ;
        RECT 2740.020 945.370 2743.020 945.380 ;
        RECT 2945.000 945.370 2948.000 945.380 ;
        RECT -28.380 768.380 -25.380 768.390 ;
        RECT 40.020 768.380 43.020 768.390 ;
        RECT 220.020 768.380 223.020 768.390 ;
        RECT 400.020 768.380 403.020 768.390 ;
        RECT 580.020 768.380 583.020 768.390 ;
        RECT 760.020 768.380 763.020 768.390 ;
        RECT 940.020 768.380 943.020 768.390 ;
        RECT 1120.020 768.380 1123.020 768.390 ;
        RECT 1300.020 768.380 1303.020 768.390 ;
        RECT 1480.020 768.380 1483.020 768.390 ;
        RECT 1660.020 768.380 1663.020 768.390 ;
        RECT 1840.020 768.380 1843.020 768.390 ;
        RECT 2020.020 768.380 2023.020 768.390 ;
        RECT 2200.020 768.380 2203.020 768.390 ;
        RECT 2380.020 768.380 2383.020 768.390 ;
        RECT 2560.020 768.380 2563.020 768.390 ;
        RECT 2740.020 768.380 2743.020 768.390 ;
        RECT 2945.000 768.380 2948.000 768.390 ;
        RECT -32.980 765.380 2952.600 768.380 ;
        RECT -28.380 765.370 -25.380 765.380 ;
        RECT 40.020 765.370 43.020 765.380 ;
        RECT 220.020 765.370 223.020 765.380 ;
        RECT 400.020 765.370 403.020 765.380 ;
        RECT 580.020 765.370 583.020 765.380 ;
        RECT 760.020 765.370 763.020 765.380 ;
        RECT 940.020 765.370 943.020 765.380 ;
        RECT 1120.020 765.370 1123.020 765.380 ;
        RECT 1300.020 765.370 1303.020 765.380 ;
        RECT 1480.020 765.370 1483.020 765.380 ;
        RECT 1660.020 765.370 1663.020 765.380 ;
        RECT 1840.020 765.370 1843.020 765.380 ;
        RECT 2020.020 765.370 2023.020 765.380 ;
        RECT 2200.020 765.370 2203.020 765.380 ;
        RECT 2380.020 765.370 2383.020 765.380 ;
        RECT 2560.020 765.370 2563.020 765.380 ;
        RECT 2740.020 765.370 2743.020 765.380 ;
        RECT 2945.000 765.370 2948.000 765.380 ;
        RECT -28.380 588.380 -25.380 588.390 ;
        RECT 40.020 588.380 43.020 588.390 ;
        RECT 220.020 588.380 223.020 588.390 ;
        RECT 400.020 588.380 403.020 588.390 ;
        RECT 580.020 588.380 583.020 588.390 ;
        RECT 760.020 588.380 763.020 588.390 ;
        RECT 940.020 588.380 943.020 588.390 ;
        RECT 1120.020 588.380 1123.020 588.390 ;
        RECT 1300.020 588.380 1303.020 588.390 ;
        RECT 1480.020 588.380 1483.020 588.390 ;
        RECT 1660.020 588.380 1663.020 588.390 ;
        RECT 1840.020 588.380 1843.020 588.390 ;
        RECT 2020.020 588.380 2023.020 588.390 ;
        RECT 2200.020 588.380 2203.020 588.390 ;
        RECT 2380.020 588.380 2383.020 588.390 ;
        RECT 2560.020 588.380 2563.020 588.390 ;
        RECT 2740.020 588.380 2743.020 588.390 ;
        RECT 2945.000 588.380 2948.000 588.390 ;
        RECT -32.980 585.380 2952.600 588.380 ;
        RECT -28.380 585.370 -25.380 585.380 ;
        RECT 40.020 585.370 43.020 585.380 ;
        RECT 220.020 585.370 223.020 585.380 ;
        RECT 400.020 585.370 403.020 585.380 ;
        RECT 580.020 585.370 583.020 585.380 ;
        RECT 760.020 585.370 763.020 585.380 ;
        RECT 940.020 585.370 943.020 585.380 ;
        RECT 1120.020 585.370 1123.020 585.380 ;
        RECT 1300.020 585.370 1303.020 585.380 ;
        RECT 1480.020 585.370 1483.020 585.380 ;
        RECT 1660.020 585.370 1663.020 585.380 ;
        RECT 1840.020 585.370 1843.020 585.380 ;
        RECT 2020.020 585.370 2023.020 585.380 ;
        RECT 2200.020 585.370 2203.020 585.380 ;
        RECT 2380.020 585.370 2383.020 585.380 ;
        RECT 2560.020 585.370 2563.020 585.380 ;
        RECT 2740.020 585.370 2743.020 585.380 ;
        RECT 2945.000 585.370 2948.000 585.380 ;
        RECT -28.380 408.380 -25.380 408.390 ;
        RECT 40.020 408.380 43.020 408.390 ;
        RECT 220.020 408.380 223.020 408.390 ;
        RECT 400.020 408.380 403.020 408.390 ;
        RECT 580.020 408.380 583.020 408.390 ;
        RECT 760.020 408.380 763.020 408.390 ;
        RECT 940.020 408.380 943.020 408.390 ;
        RECT 1120.020 408.380 1123.020 408.390 ;
        RECT 1300.020 408.380 1303.020 408.390 ;
        RECT 1480.020 408.380 1483.020 408.390 ;
        RECT 1660.020 408.380 1663.020 408.390 ;
        RECT 1840.020 408.380 1843.020 408.390 ;
        RECT 2020.020 408.380 2023.020 408.390 ;
        RECT 2200.020 408.380 2203.020 408.390 ;
        RECT 2380.020 408.380 2383.020 408.390 ;
        RECT 2560.020 408.380 2563.020 408.390 ;
        RECT 2740.020 408.380 2743.020 408.390 ;
        RECT 2945.000 408.380 2948.000 408.390 ;
        RECT -32.980 405.380 2952.600 408.380 ;
        RECT -28.380 405.370 -25.380 405.380 ;
        RECT 40.020 405.370 43.020 405.380 ;
        RECT 220.020 405.370 223.020 405.380 ;
        RECT 400.020 405.370 403.020 405.380 ;
        RECT 580.020 405.370 583.020 405.380 ;
        RECT 760.020 405.370 763.020 405.380 ;
        RECT 940.020 405.370 943.020 405.380 ;
        RECT 1120.020 405.370 1123.020 405.380 ;
        RECT 1300.020 405.370 1303.020 405.380 ;
        RECT 1480.020 405.370 1483.020 405.380 ;
        RECT 1660.020 405.370 1663.020 405.380 ;
        RECT 1840.020 405.370 1843.020 405.380 ;
        RECT 2020.020 405.370 2023.020 405.380 ;
        RECT 2200.020 405.370 2203.020 405.380 ;
        RECT 2380.020 405.370 2383.020 405.380 ;
        RECT 2560.020 405.370 2563.020 405.380 ;
        RECT 2740.020 405.370 2743.020 405.380 ;
        RECT 2945.000 405.370 2948.000 405.380 ;
        RECT -28.380 228.380 -25.380 228.390 ;
        RECT 40.020 228.380 43.020 228.390 ;
        RECT 220.020 228.380 223.020 228.390 ;
        RECT 400.020 228.380 403.020 228.390 ;
        RECT 580.020 228.380 583.020 228.390 ;
        RECT 760.020 228.380 763.020 228.390 ;
        RECT 940.020 228.380 943.020 228.390 ;
        RECT 1120.020 228.380 1123.020 228.390 ;
        RECT 1300.020 228.380 1303.020 228.390 ;
        RECT 1480.020 228.380 1483.020 228.390 ;
        RECT 1660.020 228.380 1663.020 228.390 ;
        RECT 1840.020 228.380 1843.020 228.390 ;
        RECT 2020.020 228.380 2023.020 228.390 ;
        RECT 2200.020 228.380 2203.020 228.390 ;
        RECT 2380.020 228.380 2383.020 228.390 ;
        RECT 2560.020 228.380 2563.020 228.390 ;
        RECT 2740.020 228.380 2743.020 228.390 ;
        RECT 2945.000 228.380 2948.000 228.390 ;
        RECT -32.980 225.380 2952.600 228.380 ;
        RECT -28.380 225.370 -25.380 225.380 ;
        RECT 40.020 225.370 43.020 225.380 ;
        RECT 220.020 225.370 223.020 225.380 ;
        RECT 400.020 225.370 403.020 225.380 ;
        RECT 580.020 225.370 583.020 225.380 ;
        RECT 760.020 225.370 763.020 225.380 ;
        RECT 940.020 225.370 943.020 225.380 ;
        RECT 1120.020 225.370 1123.020 225.380 ;
        RECT 1300.020 225.370 1303.020 225.380 ;
        RECT 1480.020 225.370 1483.020 225.380 ;
        RECT 1660.020 225.370 1663.020 225.380 ;
        RECT 1840.020 225.370 1843.020 225.380 ;
        RECT 2020.020 225.370 2023.020 225.380 ;
        RECT 2200.020 225.370 2203.020 225.380 ;
        RECT 2380.020 225.370 2383.020 225.380 ;
        RECT 2560.020 225.370 2563.020 225.380 ;
        RECT 2740.020 225.370 2743.020 225.380 ;
        RECT 2945.000 225.370 2948.000 225.380 ;
        RECT -28.380 48.380 -25.380 48.390 ;
        RECT 40.020 48.380 43.020 48.390 ;
        RECT 220.020 48.380 223.020 48.390 ;
        RECT 400.020 48.380 403.020 48.390 ;
        RECT 580.020 48.380 583.020 48.390 ;
        RECT 760.020 48.380 763.020 48.390 ;
        RECT 940.020 48.380 943.020 48.390 ;
        RECT 1120.020 48.380 1123.020 48.390 ;
        RECT 1300.020 48.380 1303.020 48.390 ;
        RECT 1480.020 48.380 1483.020 48.390 ;
        RECT 1660.020 48.380 1663.020 48.390 ;
        RECT 1840.020 48.380 1843.020 48.390 ;
        RECT 2020.020 48.380 2023.020 48.390 ;
        RECT 2200.020 48.380 2203.020 48.390 ;
        RECT 2380.020 48.380 2383.020 48.390 ;
        RECT 2560.020 48.380 2563.020 48.390 ;
        RECT 2740.020 48.380 2743.020 48.390 ;
        RECT 2945.000 48.380 2948.000 48.390 ;
        RECT -32.980 45.380 2952.600 48.380 ;
        RECT -28.380 45.370 -25.380 45.380 ;
        RECT 40.020 45.370 43.020 45.380 ;
        RECT 220.020 45.370 223.020 45.380 ;
        RECT 400.020 45.370 403.020 45.380 ;
        RECT 580.020 45.370 583.020 45.380 ;
        RECT 760.020 45.370 763.020 45.380 ;
        RECT 940.020 45.370 943.020 45.380 ;
        RECT 1120.020 45.370 1123.020 45.380 ;
        RECT 1300.020 45.370 1303.020 45.380 ;
        RECT 1480.020 45.370 1483.020 45.380 ;
        RECT 1660.020 45.370 1663.020 45.380 ;
        RECT 1840.020 45.370 1843.020 45.380 ;
        RECT 2020.020 45.370 2023.020 45.380 ;
        RECT 2200.020 45.370 2203.020 45.380 ;
        RECT 2380.020 45.370 2383.020 45.380 ;
        RECT 2560.020 45.370 2563.020 45.380 ;
        RECT 2740.020 45.370 2743.020 45.380 ;
        RECT 2945.000 45.370 2948.000 45.380 ;
        RECT -28.380 -20.020 -25.380 -20.010 ;
        RECT 40.020 -20.020 43.020 -20.010 ;
        RECT 220.020 -20.020 223.020 -20.010 ;
        RECT 400.020 -20.020 403.020 -20.010 ;
        RECT 580.020 -20.020 583.020 -20.010 ;
        RECT 760.020 -20.020 763.020 -20.010 ;
        RECT 940.020 -20.020 943.020 -20.010 ;
        RECT 1120.020 -20.020 1123.020 -20.010 ;
        RECT 1300.020 -20.020 1303.020 -20.010 ;
        RECT 1480.020 -20.020 1483.020 -20.010 ;
        RECT 1660.020 -20.020 1663.020 -20.010 ;
        RECT 1840.020 -20.020 1843.020 -20.010 ;
        RECT 2020.020 -20.020 2023.020 -20.010 ;
        RECT 2200.020 -20.020 2203.020 -20.010 ;
        RECT 2380.020 -20.020 2383.020 -20.010 ;
        RECT 2560.020 -20.020 2563.020 -20.010 ;
        RECT 2740.020 -20.020 2743.020 -20.010 ;
        RECT 2945.000 -20.020 2948.000 -20.010 ;
        RECT -28.380 -23.020 2948.000 -20.020 ;
        RECT -28.380 -23.030 -25.380 -23.020 ;
        RECT 40.020 -23.030 43.020 -23.020 ;
        RECT 220.020 -23.030 223.020 -23.020 ;
        RECT 400.020 -23.030 403.020 -23.020 ;
        RECT 580.020 -23.030 583.020 -23.020 ;
        RECT 760.020 -23.030 763.020 -23.020 ;
        RECT 940.020 -23.030 943.020 -23.020 ;
        RECT 1120.020 -23.030 1123.020 -23.020 ;
        RECT 1300.020 -23.030 1303.020 -23.020 ;
        RECT 1480.020 -23.030 1483.020 -23.020 ;
        RECT 1660.020 -23.030 1663.020 -23.020 ;
        RECT 1840.020 -23.030 1843.020 -23.020 ;
        RECT 2020.020 -23.030 2023.020 -23.020 ;
        RECT 2200.020 -23.030 2203.020 -23.020 ;
        RECT 2380.020 -23.030 2383.020 -23.020 ;
        RECT 2560.020 -23.030 2563.020 -23.020 ;
        RECT 2740.020 -23.030 2743.020 -23.020 ;
        RECT 2945.000 -23.030 2948.000 -23.020 ;
    END
  END vdda1
  PIN vssa1
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -32.980 -27.620 -29.980 3547.300 ;
        RECT 130.020 -27.620 133.020 3547.300 ;
        RECT 310.020 -27.620 313.020 3547.300 ;
        RECT 490.020 -27.620 493.020 3547.300 ;
        RECT 670.020 -27.620 673.020 3547.300 ;
        RECT 850.020 -27.620 853.020 3547.300 ;
        RECT 1030.020 -27.620 1033.020 3547.300 ;
        RECT 1210.020 -27.620 1213.020 3547.300 ;
        RECT 1390.020 -27.620 1393.020 3547.300 ;
        RECT 1570.020 -27.620 1573.020 3547.300 ;
        RECT 1750.020 -27.620 1753.020 3547.300 ;
        RECT 1930.020 -27.620 1933.020 3547.300 ;
        RECT 2110.020 -27.620 2113.020 3547.300 ;
        RECT 2290.020 -27.620 2293.020 3547.300 ;
        RECT 2470.020 -27.620 2473.020 3547.300 ;
        RECT 2650.020 -27.620 2653.020 3547.300 ;
        RECT 2830.020 -27.620 2833.020 3547.300 ;
        RECT 2949.600 -27.620 2952.600 3547.300 ;
      LAYER via4 ;
        RECT -32.070 3546.010 -30.890 3547.190 ;
        RECT -32.070 3544.410 -30.890 3545.590 ;
        RECT -32.070 3377.090 -30.890 3378.270 ;
        RECT -32.070 3375.490 -30.890 3376.670 ;
        RECT -32.070 3197.090 -30.890 3198.270 ;
        RECT -32.070 3195.490 -30.890 3196.670 ;
        RECT -32.070 3017.090 -30.890 3018.270 ;
        RECT -32.070 3015.490 -30.890 3016.670 ;
        RECT -32.070 2837.090 -30.890 2838.270 ;
        RECT -32.070 2835.490 -30.890 2836.670 ;
        RECT -32.070 2657.090 -30.890 2658.270 ;
        RECT -32.070 2655.490 -30.890 2656.670 ;
        RECT -32.070 2477.090 -30.890 2478.270 ;
        RECT -32.070 2475.490 -30.890 2476.670 ;
        RECT -32.070 2297.090 -30.890 2298.270 ;
        RECT -32.070 2295.490 -30.890 2296.670 ;
        RECT -32.070 2117.090 -30.890 2118.270 ;
        RECT -32.070 2115.490 -30.890 2116.670 ;
        RECT -32.070 1937.090 -30.890 1938.270 ;
        RECT -32.070 1935.490 -30.890 1936.670 ;
        RECT -32.070 1757.090 -30.890 1758.270 ;
        RECT -32.070 1755.490 -30.890 1756.670 ;
        RECT -32.070 1577.090 -30.890 1578.270 ;
        RECT -32.070 1575.490 -30.890 1576.670 ;
        RECT -32.070 1397.090 -30.890 1398.270 ;
        RECT -32.070 1395.490 -30.890 1396.670 ;
        RECT -32.070 1217.090 -30.890 1218.270 ;
        RECT -32.070 1215.490 -30.890 1216.670 ;
        RECT -32.070 1037.090 -30.890 1038.270 ;
        RECT -32.070 1035.490 -30.890 1036.670 ;
        RECT -32.070 857.090 -30.890 858.270 ;
        RECT -32.070 855.490 -30.890 856.670 ;
        RECT -32.070 677.090 -30.890 678.270 ;
        RECT -32.070 675.490 -30.890 676.670 ;
        RECT -32.070 497.090 -30.890 498.270 ;
        RECT -32.070 495.490 -30.890 496.670 ;
        RECT -32.070 317.090 -30.890 318.270 ;
        RECT -32.070 315.490 -30.890 316.670 ;
        RECT -32.070 137.090 -30.890 138.270 ;
        RECT -32.070 135.490 -30.890 136.670 ;
        RECT -32.070 -25.910 -30.890 -24.730 ;
        RECT -32.070 -27.510 -30.890 -26.330 ;
        RECT 130.930 3546.010 132.110 3547.190 ;
        RECT 130.930 3544.410 132.110 3545.590 ;
        RECT 130.930 3377.090 132.110 3378.270 ;
        RECT 130.930 3375.490 132.110 3376.670 ;
        RECT 130.930 3197.090 132.110 3198.270 ;
        RECT 130.930 3195.490 132.110 3196.670 ;
        RECT 130.930 3017.090 132.110 3018.270 ;
        RECT 130.930 3015.490 132.110 3016.670 ;
        RECT 130.930 2837.090 132.110 2838.270 ;
        RECT 130.930 2835.490 132.110 2836.670 ;
        RECT 130.930 2657.090 132.110 2658.270 ;
        RECT 130.930 2655.490 132.110 2656.670 ;
        RECT 130.930 2477.090 132.110 2478.270 ;
        RECT 130.930 2475.490 132.110 2476.670 ;
        RECT 130.930 2297.090 132.110 2298.270 ;
        RECT 130.930 2295.490 132.110 2296.670 ;
        RECT 130.930 2117.090 132.110 2118.270 ;
        RECT 130.930 2115.490 132.110 2116.670 ;
        RECT 130.930 1937.090 132.110 1938.270 ;
        RECT 130.930 1935.490 132.110 1936.670 ;
        RECT 130.930 1757.090 132.110 1758.270 ;
        RECT 130.930 1755.490 132.110 1756.670 ;
        RECT 130.930 1577.090 132.110 1578.270 ;
        RECT 130.930 1575.490 132.110 1576.670 ;
        RECT 130.930 1397.090 132.110 1398.270 ;
        RECT 130.930 1395.490 132.110 1396.670 ;
        RECT 130.930 1217.090 132.110 1218.270 ;
        RECT 130.930 1215.490 132.110 1216.670 ;
        RECT 130.930 1037.090 132.110 1038.270 ;
        RECT 130.930 1035.490 132.110 1036.670 ;
        RECT 130.930 857.090 132.110 858.270 ;
        RECT 130.930 855.490 132.110 856.670 ;
        RECT 130.930 677.090 132.110 678.270 ;
        RECT 130.930 675.490 132.110 676.670 ;
        RECT 130.930 497.090 132.110 498.270 ;
        RECT 130.930 495.490 132.110 496.670 ;
        RECT 130.930 317.090 132.110 318.270 ;
        RECT 130.930 315.490 132.110 316.670 ;
        RECT 130.930 137.090 132.110 138.270 ;
        RECT 130.930 135.490 132.110 136.670 ;
        RECT 130.930 -25.910 132.110 -24.730 ;
        RECT 130.930 -27.510 132.110 -26.330 ;
        RECT 310.930 3546.010 312.110 3547.190 ;
        RECT 310.930 3544.410 312.110 3545.590 ;
        RECT 310.930 3377.090 312.110 3378.270 ;
        RECT 310.930 3375.490 312.110 3376.670 ;
        RECT 310.930 3197.090 312.110 3198.270 ;
        RECT 310.930 3195.490 312.110 3196.670 ;
        RECT 310.930 3017.090 312.110 3018.270 ;
        RECT 310.930 3015.490 312.110 3016.670 ;
        RECT 310.930 2837.090 312.110 2838.270 ;
        RECT 310.930 2835.490 312.110 2836.670 ;
        RECT 310.930 2657.090 312.110 2658.270 ;
        RECT 310.930 2655.490 312.110 2656.670 ;
        RECT 310.930 2477.090 312.110 2478.270 ;
        RECT 310.930 2475.490 312.110 2476.670 ;
        RECT 310.930 2297.090 312.110 2298.270 ;
        RECT 310.930 2295.490 312.110 2296.670 ;
        RECT 310.930 2117.090 312.110 2118.270 ;
        RECT 310.930 2115.490 312.110 2116.670 ;
        RECT 310.930 1937.090 312.110 1938.270 ;
        RECT 310.930 1935.490 312.110 1936.670 ;
        RECT 310.930 1757.090 312.110 1758.270 ;
        RECT 310.930 1755.490 312.110 1756.670 ;
        RECT 310.930 1577.090 312.110 1578.270 ;
        RECT 310.930 1575.490 312.110 1576.670 ;
        RECT 310.930 1397.090 312.110 1398.270 ;
        RECT 310.930 1395.490 312.110 1396.670 ;
        RECT 310.930 1217.090 312.110 1218.270 ;
        RECT 310.930 1215.490 312.110 1216.670 ;
        RECT 310.930 1037.090 312.110 1038.270 ;
        RECT 310.930 1035.490 312.110 1036.670 ;
        RECT 310.930 857.090 312.110 858.270 ;
        RECT 310.930 855.490 312.110 856.670 ;
        RECT 310.930 677.090 312.110 678.270 ;
        RECT 310.930 675.490 312.110 676.670 ;
        RECT 310.930 497.090 312.110 498.270 ;
        RECT 310.930 495.490 312.110 496.670 ;
        RECT 310.930 317.090 312.110 318.270 ;
        RECT 310.930 315.490 312.110 316.670 ;
        RECT 310.930 137.090 312.110 138.270 ;
        RECT 310.930 135.490 312.110 136.670 ;
        RECT 310.930 -25.910 312.110 -24.730 ;
        RECT 310.930 -27.510 312.110 -26.330 ;
        RECT 490.930 3546.010 492.110 3547.190 ;
        RECT 490.930 3544.410 492.110 3545.590 ;
        RECT 490.930 3377.090 492.110 3378.270 ;
        RECT 490.930 3375.490 492.110 3376.670 ;
        RECT 490.930 3197.090 492.110 3198.270 ;
        RECT 490.930 3195.490 492.110 3196.670 ;
        RECT 490.930 3017.090 492.110 3018.270 ;
        RECT 490.930 3015.490 492.110 3016.670 ;
        RECT 490.930 2837.090 492.110 2838.270 ;
        RECT 490.930 2835.490 492.110 2836.670 ;
        RECT 490.930 2657.090 492.110 2658.270 ;
        RECT 490.930 2655.490 492.110 2656.670 ;
        RECT 490.930 2477.090 492.110 2478.270 ;
        RECT 490.930 2475.490 492.110 2476.670 ;
        RECT 490.930 2297.090 492.110 2298.270 ;
        RECT 490.930 2295.490 492.110 2296.670 ;
        RECT 490.930 2117.090 492.110 2118.270 ;
        RECT 490.930 2115.490 492.110 2116.670 ;
        RECT 490.930 1937.090 492.110 1938.270 ;
        RECT 490.930 1935.490 492.110 1936.670 ;
        RECT 490.930 1757.090 492.110 1758.270 ;
        RECT 490.930 1755.490 492.110 1756.670 ;
        RECT 490.930 1577.090 492.110 1578.270 ;
        RECT 490.930 1575.490 492.110 1576.670 ;
        RECT 490.930 1397.090 492.110 1398.270 ;
        RECT 490.930 1395.490 492.110 1396.670 ;
        RECT 490.930 1217.090 492.110 1218.270 ;
        RECT 490.930 1215.490 492.110 1216.670 ;
        RECT 490.930 1037.090 492.110 1038.270 ;
        RECT 490.930 1035.490 492.110 1036.670 ;
        RECT 490.930 857.090 492.110 858.270 ;
        RECT 490.930 855.490 492.110 856.670 ;
        RECT 490.930 677.090 492.110 678.270 ;
        RECT 490.930 675.490 492.110 676.670 ;
        RECT 490.930 497.090 492.110 498.270 ;
        RECT 490.930 495.490 492.110 496.670 ;
        RECT 490.930 317.090 492.110 318.270 ;
        RECT 490.930 315.490 492.110 316.670 ;
        RECT 490.930 137.090 492.110 138.270 ;
        RECT 490.930 135.490 492.110 136.670 ;
        RECT 490.930 -25.910 492.110 -24.730 ;
        RECT 490.930 -27.510 492.110 -26.330 ;
        RECT 670.930 3546.010 672.110 3547.190 ;
        RECT 670.930 3544.410 672.110 3545.590 ;
        RECT 670.930 3377.090 672.110 3378.270 ;
        RECT 670.930 3375.490 672.110 3376.670 ;
        RECT 670.930 3197.090 672.110 3198.270 ;
        RECT 670.930 3195.490 672.110 3196.670 ;
        RECT 670.930 3017.090 672.110 3018.270 ;
        RECT 670.930 3015.490 672.110 3016.670 ;
        RECT 670.930 2837.090 672.110 2838.270 ;
        RECT 670.930 2835.490 672.110 2836.670 ;
        RECT 670.930 2657.090 672.110 2658.270 ;
        RECT 670.930 2655.490 672.110 2656.670 ;
        RECT 670.930 2477.090 672.110 2478.270 ;
        RECT 670.930 2475.490 672.110 2476.670 ;
        RECT 670.930 2297.090 672.110 2298.270 ;
        RECT 670.930 2295.490 672.110 2296.670 ;
        RECT 670.930 2117.090 672.110 2118.270 ;
        RECT 670.930 2115.490 672.110 2116.670 ;
        RECT 670.930 1937.090 672.110 1938.270 ;
        RECT 670.930 1935.490 672.110 1936.670 ;
        RECT 670.930 1757.090 672.110 1758.270 ;
        RECT 670.930 1755.490 672.110 1756.670 ;
        RECT 670.930 1577.090 672.110 1578.270 ;
        RECT 670.930 1575.490 672.110 1576.670 ;
        RECT 670.930 1397.090 672.110 1398.270 ;
        RECT 670.930 1395.490 672.110 1396.670 ;
        RECT 670.930 1217.090 672.110 1218.270 ;
        RECT 670.930 1215.490 672.110 1216.670 ;
        RECT 670.930 1037.090 672.110 1038.270 ;
        RECT 670.930 1035.490 672.110 1036.670 ;
        RECT 670.930 857.090 672.110 858.270 ;
        RECT 670.930 855.490 672.110 856.670 ;
        RECT 670.930 677.090 672.110 678.270 ;
        RECT 670.930 675.490 672.110 676.670 ;
        RECT 670.930 497.090 672.110 498.270 ;
        RECT 670.930 495.490 672.110 496.670 ;
        RECT 670.930 317.090 672.110 318.270 ;
        RECT 670.930 315.490 672.110 316.670 ;
        RECT 670.930 137.090 672.110 138.270 ;
        RECT 670.930 135.490 672.110 136.670 ;
        RECT 670.930 -25.910 672.110 -24.730 ;
        RECT 670.930 -27.510 672.110 -26.330 ;
        RECT 850.930 3546.010 852.110 3547.190 ;
        RECT 850.930 3544.410 852.110 3545.590 ;
        RECT 850.930 3377.090 852.110 3378.270 ;
        RECT 850.930 3375.490 852.110 3376.670 ;
        RECT 850.930 3197.090 852.110 3198.270 ;
        RECT 850.930 3195.490 852.110 3196.670 ;
        RECT 850.930 3017.090 852.110 3018.270 ;
        RECT 850.930 3015.490 852.110 3016.670 ;
        RECT 850.930 2837.090 852.110 2838.270 ;
        RECT 850.930 2835.490 852.110 2836.670 ;
        RECT 850.930 2657.090 852.110 2658.270 ;
        RECT 850.930 2655.490 852.110 2656.670 ;
        RECT 850.930 2477.090 852.110 2478.270 ;
        RECT 850.930 2475.490 852.110 2476.670 ;
        RECT 850.930 2297.090 852.110 2298.270 ;
        RECT 850.930 2295.490 852.110 2296.670 ;
        RECT 850.930 2117.090 852.110 2118.270 ;
        RECT 850.930 2115.490 852.110 2116.670 ;
        RECT 850.930 1937.090 852.110 1938.270 ;
        RECT 850.930 1935.490 852.110 1936.670 ;
        RECT 850.930 1757.090 852.110 1758.270 ;
        RECT 850.930 1755.490 852.110 1756.670 ;
        RECT 850.930 1577.090 852.110 1578.270 ;
        RECT 850.930 1575.490 852.110 1576.670 ;
        RECT 850.930 1397.090 852.110 1398.270 ;
        RECT 850.930 1395.490 852.110 1396.670 ;
        RECT 850.930 1217.090 852.110 1218.270 ;
        RECT 850.930 1215.490 852.110 1216.670 ;
        RECT 850.930 1037.090 852.110 1038.270 ;
        RECT 850.930 1035.490 852.110 1036.670 ;
        RECT 850.930 857.090 852.110 858.270 ;
        RECT 850.930 855.490 852.110 856.670 ;
        RECT 850.930 677.090 852.110 678.270 ;
        RECT 850.930 675.490 852.110 676.670 ;
        RECT 850.930 497.090 852.110 498.270 ;
        RECT 850.930 495.490 852.110 496.670 ;
        RECT 850.930 317.090 852.110 318.270 ;
        RECT 850.930 315.490 852.110 316.670 ;
        RECT 850.930 137.090 852.110 138.270 ;
        RECT 850.930 135.490 852.110 136.670 ;
        RECT 850.930 -25.910 852.110 -24.730 ;
        RECT 850.930 -27.510 852.110 -26.330 ;
        RECT 1030.930 3546.010 1032.110 3547.190 ;
        RECT 1030.930 3544.410 1032.110 3545.590 ;
        RECT 1030.930 3377.090 1032.110 3378.270 ;
        RECT 1030.930 3375.490 1032.110 3376.670 ;
        RECT 1030.930 3197.090 1032.110 3198.270 ;
        RECT 1030.930 3195.490 1032.110 3196.670 ;
        RECT 1030.930 3017.090 1032.110 3018.270 ;
        RECT 1030.930 3015.490 1032.110 3016.670 ;
        RECT 1030.930 2837.090 1032.110 2838.270 ;
        RECT 1030.930 2835.490 1032.110 2836.670 ;
        RECT 1030.930 2657.090 1032.110 2658.270 ;
        RECT 1030.930 2655.490 1032.110 2656.670 ;
        RECT 1030.930 2477.090 1032.110 2478.270 ;
        RECT 1030.930 2475.490 1032.110 2476.670 ;
        RECT 1030.930 2297.090 1032.110 2298.270 ;
        RECT 1030.930 2295.490 1032.110 2296.670 ;
        RECT 1030.930 2117.090 1032.110 2118.270 ;
        RECT 1030.930 2115.490 1032.110 2116.670 ;
        RECT 1030.930 1937.090 1032.110 1938.270 ;
        RECT 1030.930 1935.490 1032.110 1936.670 ;
        RECT 1030.930 1757.090 1032.110 1758.270 ;
        RECT 1030.930 1755.490 1032.110 1756.670 ;
        RECT 1030.930 1577.090 1032.110 1578.270 ;
        RECT 1030.930 1575.490 1032.110 1576.670 ;
        RECT 1030.930 1397.090 1032.110 1398.270 ;
        RECT 1030.930 1395.490 1032.110 1396.670 ;
        RECT 1030.930 1217.090 1032.110 1218.270 ;
        RECT 1030.930 1215.490 1032.110 1216.670 ;
        RECT 1030.930 1037.090 1032.110 1038.270 ;
        RECT 1030.930 1035.490 1032.110 1036.670 ;
        RECT 1030.930 857.090 1032.110 858.270 ;
        RECT 1030.930 855.490 1032.110 856.670 ;
        RECT 1030.930 677.090 1032.110 678.270 ;
        RECT 1030.930 675.490 1032.110 676.670 ;
        RECT 1030.930 497.090 1032.110 498.270 ;
        RECT 1030.930 495.490 1032.110 496.670 ;
        RECT 1030.930 317.090 1032.110 318.270 ;
        RECT 1030.930 315.490 1032.110 316.670 ;
        RECT 1030.930 137.090 1032.110 138.270 ;
        RECT 1030.930 135.490 1032.110 136.670 ;
        RECT 1030.930 -25.910 1032.110 -24.730 ;
        RECT 1030.930 -27.510 1032.110 -26.330 ;
        RECT 1210.930 3546.010 1212.110 3547.190 ;
        RECT 1210.930 3544.410 1212.110 3545.590 ;
        RECT 1210.930 3377.090 1212.110 3378.270 ;
        RECT 1210.930 3375.490 1212.110 3376.670 ;
        RECT 1210.930 3197.090 1212.110 3198.270 ;
        RECT 1210.930 3195.490 1212.110 3196.670 ;
        RECT 1210.930 3017.090 1212.110 3018.270 ;
        RECT 1210.930 3015.490 1212.110 3016.670 ;
        RECT 1210.930 2837.090 1212.110 2838.270 ;
        RECT 1210.930 2835.490 1212.110 2836.670 ;
        RECT 1210.930 2657.090 1212.110 2658.270 ;
        RECT 1210.930 2655.490 1212.110 2656.670 ;
        RECT 1210.930 2477.090 1212.110 2478.270 ;
        RECT 1210.930 2475.490 1212.110 2476.670 ;
        RECT 1210.930 2297.090 1212.110 2298.270 ;
        RECT 1210.930 2295.490 1212.110 2296.670 ;
        RECT 1210.930 2117.090 1212.110 2118.270 ;
        RECT 1210.930 2115.490 1212.110 2116.670 ;
        RECT 1210.930 1937.090 1212.110 1938.270 ;
        RECT 1210.930 1935.490 1212.110 1936.670 ;
        RECT 1210.930 1757.090 1212.110 1758.270 ;
        RECT 1210.930 1755.490 1212.110 1756.670 ;
        RECT 1210.930 1577.090 1212.110 1578.270 ;
        RECT 1210.930 1575.490 1212.110 1576.670 ;
        RECT 1210.930 1397.090 1212.110 1398.270 ;
        RECT 1210.930 1395.490 1212.110 1396.670 ;
        RECT 1210.930 1217.090 1212.110 1218.270 ;
        RECT 1210.930 1215.490 1212.110 1216.670 ;
        RECT 1210.930 1037.090 1212.110 1038.270 ;
        RECT 1210.930 1035.490 1212.110 1036.670 ;
        RECT 1210.930 857.090 1212.110 858.270 ;
        RECT 1210.930 855.490 1212.110 856.670 ;
        RECT 1210.930 677.090 1212.110 678.270 ;
        RECT 1210.930 675.490 1212.110 676.670 ;
        RECT 1210.930 497.090 1212.110 498.270 ;
        RECT 1210.930 495.490 1212.110 496.670 ;
        RECT 1210.930 317.090 1212.110 318.270 ;
        RECT 1210.930 315.490 1212.110 316.670 ;
        RECT 1210.930 137.090 1212.110 138.270 ;
        RECT 1210.930 135.490 1212.110 136.670 ;
        RECT 1210.930 -25.910 1212.110 -24.730 ;
        RECT 1210.930 -27.510 1212.110 -26.330 ;
        RECT 1390.930 3546.010 1392.110 3547.190 ;
        RECT 1390.930 3544.410 1392.110 3545.590 ;
        RECT 1390.930 3377.090 1392.110 3378.270 ;
        RECT 1390.930 3375.490 1392.110 3376.670 ;
        RECT 1390.930 3197.090 1392.110 3198.270 ;
        RECT 1390.930 3195.490 1392.110 3196.670 ;
        RECT 1390.930 3017.090 1392.110 3018.270 ;
        RECT 1390.930 3015.490 1392.110 3016.670 ;
        RECT 1390.930 2837.090 1392.110 2838.270 ;
        RECT 1390.930 2835.490 1392.110 2836.670 ;
        RECT 1390.930 2657.090 1392.110 2658.270 ;
        RECT 1390.930 2655.490 1392.110 2656.670 ;
        RECT 1390.930 2477.090 1392.110 2478.270 ;
        RECT 1390.930 2475.490 1392.110 2476.670 ;
        RECT 1390.930 2297.090 1392.110 2298.270 ;
        RECT 1390.930 2295.490 1392.110 2296.670 ;
        RECT 1390.930 2117.090 1392.110 2118.270 ;
        RECT 1390.930 2115.490 1392.110 2116.670 ;
        RECT 1390.930 1937.090 1392.110 1938.270 ;
        RECT 1390.930 1935.490 1392.110 1936.670 ;
        RECT 1390.930 1757.090 1392.110 1758.270 ;
        RECT 1390.930 1755.490 1392.110 1756.670 ;
        RECT 1390.930 1577.090 1392.110 1578.270 ;
        RECT 1390.930 1575.490 1392.110 1576.670 ;
        RECT 1390.930 1397.090 1392.110 1398.270 ;
        RECT 1390.930 1395.490 1392.110 1396.670 ;
        RECT 1390.930 1217.090 1392.110 1218.270 ;
        RECT 1390.930 1215.490 1392.110 1216.670 ;
        RECT 1390.930 1037.090 1392.110 1038.270 ;
        RECT 1390.930 1035.490 1392.110 1036.670 ;
        RECT 1390.930 857.090 1392.110 858.270 ;
        RECT 1390.930 855.490 1392.110 856.670 ;
        RECT 1390.930 677.090 1392.110 678.270 ;
        RECT 1390.930 675.490 1392.110 676.670 ;
        RECT 1390.930 497.090 1392.110 498.270 ;
        RECT 1390.930 495.490 1392.110 496.670 ;
        RECT 1390.930 317.090 1392.110 318.270 ;
        RECT 1390.930 315.490 1392.110 316.670 ;
        RECT 1390.930 137.090 1392.110 138.270 ;
        RECT 1390.930 135.490 1392.110 136.670 ;
        RECT 1390.930 -25.910 1392.110 -24.730 ;
        RECT 1390.930 -27.510 1392.110 -26.330 ;
        RECT 1570.930 3546.010 1572.110 3547.190 ;
        RECT 1570.930 3544.410 1572.110 3545.590 ;
        RECT 1570.930 3377.090 1572.110 3378.270 ;
        RECT 1570.930 3375.490 1572.110 3376.670 ;
        RECT 1570.930 3197.090 1572.110 3198.270 ;
        RECT 1570.930 3195.490 1572.110 3196.670 ;
        RECT 1570.930 3017.090 1572.110 3018.270 ;
        RECT 1570.930 3015.490 1572.110 3016.670 ;
        RECT 1570.930 2837.090 1572.110 2838.270 ;
        RECT 1570.930 2835.490 1572.110 2836.670 ;
        RECT 1570.930 2657.090 1572.110 2658.270 ;
        RECT 1570.930 2655.490 1572.110 2656.670 ;
        RECT 1570.930 2477.090 1572.110 2478.270 ;
        RECT 1570.930 2475.490 1572.110 2476.670 ;
        RECT 1570.930 2297.090 1572.110 2298.270 ;
        RECT 1570.930 2295.490 1572.110 2296.670 ;
        RECT 1570.930 2117.090 1572.110 2118.270 ;
        RECT 1570.930 2115.490 1572.110 2116.670 ;
        RECT 1570.930 1937.090 1572.110 1938.270 ;
        RECT 1570.930 1935.490 1572.110 1936.670 ;
        RECT 1570.930 1757.090 1572.110 1758.270 ;
        RECT 1570.930 1755.490 1572.110 1756.670 ;
        RECT 1570.930 1577.090 1572.110 1578.270 ;
        RECT 1570.930 1575.490 1572.110 1576.670 ;
        RECT 1570.930 1397.090 1572.110 1398.270 ;
        RECT 1570.930 1395.490 1572.110 1396.670 ;
        RECT 1570.930 1217.090 1572.110 1218.270 ;
        RECT 1570.930 1215.490 1572.110 1216.670 ;
        RECT 1570.930 1037.090 1572.110 1038.270 ;
        RECT 1570.930 1035.490 1572.110 1036.670 ;
        RECT 1570.930 857.090 1572.110 858.270 ;
        RECT 1570.930 855.490 1572.110 856.670 ;
        RECT 1570.930 677.090 1572.110 678.270 ;
        RECT 1570.930 675.490 1572.110 676.670 ;
        RECT 1570.930 497.090 1572.110 498.270 ;
        RECT 1570.930 495.490 1572.110 496.670 ;
        RECT 1570.930 317.090 1572.110 318.270 ;
        RECT 1570.930 315.490 1572.110 316.670 ;
        RECT 1570.930 137.090 1572.110 138.270 ;
        RECT 1570.930 135.490 1572.110 136.670 ;
        RECT 1570.930 -25.910 1572.110 -24.730 ;
        RECT 1570.930 -27.510 1572.110 -26.330 ;
        RECT 1750.930 3546.010 1752.110 3547.190 ;
        RECT 1750.930 3544.410 1752.110 3545.590 ;
        RECT 1750.930 3377.090 1752.110 3378.270 ;
        RECT 1750.930 3375.490 1752.110 3376.670 ;
        RECT 1750.930 3197.090 1752.110 3198.270 ;
        RECT 1750.930 3195.490 1752.110 3196.670 ;
        RECT 1750.930 3017.090 1752.110 3018.270 ;
        RECT 1750.930 3015.490 1752.110 3016.670 ;
        RECT 1750.930 2837.090 1752.110 2838.270 ;
        RECT 1750.930 2835.490 1752.110 2836.670 ;
        RECT 1750.930 2657.090 1752.110 2658.270 ;
        RECT 1750.930 2655.490 1752.110 2656.670 ;
        RECT 1750.930 2477.090 1752.110 2478.270 ;
        RECT 1750.930 2475.490 1752.110 2476.670 ;
        RECT 1750.930 2297.090 1752.110 2298.270 ;
        RECT 1750.930 2295.490 1752.110 2296.670 ;
        RECT 1750.930 2117.090 1752.110 2118.270 ;
        RECT 1750.930 2115.490 1752.110 2116.670 ;
        RECT 1750.930 1937.090 1752.110 1938.270 ;
        RECT 1750.930 1935.490 1752.110 1936.670 ;
        RECT 1750.930 1757.090 1752.110 1758.270 ;
        RECT 1750.930 1755.490 1752.110 1756.670 ;
        RECT 1750.930 1577.090 1752.110 1578.270 ;
        RECT 1750.930 1575.490 1752.110 1576.670 ;
        RECT 1750.930 1397.090 1752.110 1398.270 ;
        RECT 1750.930 1395.490 1752.110 1396.670 ;
        RECT 1750.930 1217.090 1752.110 1218.270 ;
        RECT 1750.930 1215.490 1752.110 1216.670 ;
        RECT 1750.930 1037.090 1752.110 1038.270 ;
        RECT 1750.930 1035.490 1752.110 1036.670 ;
        RECT 1750.930 857.090 1752.110 858.270 ;
        RECT 1750.930 855.490 1752.110 856.670 ;
        RECT 1750.930 677.090 1752.110 678.270 ;
        RECT 1750.930 675.490 1752.110 676.670 ;
        RECT 1750.930 497.090 1752.110 498.270 ;
        RECT 1750.930 495.490 1752.110 496.670 ;
        RECT 1750.930 317.090 1752.110 318.270 ;
        RECT 1750.930 315.490 1752.110 316.670 ;
        RECT 1750.930 137.090 1752.110 138.270 ;
        RECT 1750.930 135.490 1752.110 136.670 ;
        RECT 1750.930 -25.910 1752.110 -24.730 ;
        RECT 1750.930 -27.510 1752.110 -26.330 ;
        RECT 1930.930 3546.010 1932.110 3547.190 ;
        RECT 1930.930 3544.410 1932.110 3545.590 ;
        RECT 1930.930 3377.090 1932.110 3378.270 ;
        RECT 1930.930 3375.490 1932.110 3376.670 ;
        RECT 1930.930 3197.090 1932.110 3198.270 ;
        RECT 1930.930 3195.490 1932.110 3196.670 ;
        RECT 1930.930 3017.090 1932.110 3018.270 ;
        RECT 1930.930 3015.490 1932.110 3016.670 ;
        RECT 1930.930 2837.090 1932.110 2838.270 ;
        RECT 1930.930 2835.490 1932.110 2836.670 ;
        RECT 1930.930 2657.090 1932.110 2658.270 ;
        RECT 1930.930 2655.490 1932.110 2656.670 ;
        RECT 1930.930 2477.090 1932.110 2478.270 ;
        RECT 1930.930 2475.490 1932.110 2476.670 ;
        RECT 1930.930 2297.090 1932.110 2298.270 ;
        RECT 1930.930 2295.490 1932.110 2296.670 ;
        RECT 1930.930 2117.090 1932.110 2118.270 ;
        RECT 1930.930 2115.490 1932.110 2116.670 ;
        RECT 1930.930 1937.090 1932.110 1938.270 ;
        RECT 1930.930 1935.490 1932.110 1936.670 ;
        RECT 1930.930 1757.090 1932.110 1758.270 ;
        RECT 1930.930 1755.490 1932.110 1756.670 ;
        RECT 1930.930 1577.090 1932.110 1578.270 ;
        RECT 1930.930 1575.490 1932.110 1576.670 ;
        RECT 1930.930 1397.090 1932.110 1398.270 ;
        RECT 1930.930 1395.490 1932.110 1396.670 ;
        RECT 1930.930 1217.090 1932.110 1218.270 ;
        RECT 1930.930 1215.490 1932.110 1216.670 ;
        RECT 1930.930 1037.090 1932.110 1038.270 ;
        RECT 1930.930 1035.490 1932.110 1036.670 ;
        RECT 1930.930 857.090 1932.110 858.270 ;
        RECT 1930.930 855.490 1932.110 856.670 ;
        RECT 1930.930 677.090 1932.110 678.270 ;
        RECT 1930.930 675.490 1932.110 676.670 ;
        RECT 1930.930 497.090 1932.110 498.270 ;
        RECT 1930.930 495.490 1932.110 496.670 ;
        RECT 1930.930 317.090 1932.110 318.270 ;
        RECT 1930.930 315.490 1932.110 316.670 ;
        RECT 1930.930 137.090 1932.110 138.270 ;
        RECT 1930.930 135.490 1932.110 136.670 ;
        RECT 1930.930 -25.910 1932.110 -24.730 ;
        RECT 1930.930 -27.510 1932.110 -26.330 ;
        RECT 2110.930 3546.010 2112.110 3547.190 ;
        RECT 2110.930 3544.410 2112.110 3545.590 ;
        RECT 2110.930 3377.090 2112.110 3378.270 ;
        RECT 2110.930 3375.490 2112.110 3376.670 ;
        RECT 2110.930 3197.090 2112.110 3198.270 ;
        RECT 2110.930 3195.490 2112.110 3196.670 ;
        RECT 2110.930 3017.090 2112.110 3018.270 ;
        RECT 2110.930 3015.490 2112.110 3016.670 ;
        RECT 2110.930 2837.090 2112.110 2838.270 ;
        RECT 2110.930 2835.490 2112.110 2836.670 ;
        RECT 2110.930 2657.090 2112.110 2658.270 ;
        RECT 2110.930 2655.490 2112.110 2656.670 ;
        RECT 2110.930 2477.090 2112.110 2478.270 ;
        RECT 2110.930 2475.490 2112.110 2476.670 ;
        RECT 2110.930 2297.090 2112.110 2298.270 ;
        RECT 2110.930 2295.490 2112.110 2296.670 ;
        RECT 2110.930 2117.090 2112.110 2118.270 ;
        RECT 2110.930 2115.490 2112.110 2116.670 ;
        RECT 2110.930 1937.090 2112.110 1938.270 ;
        RECT 2110.930 1935.490 2112.110 1936.670 ;
        RECT 2110.930 1757.090 2112.110 1758.270 ;
        RECT 2110.930 1755.490 2112.110 1756.670 ;
        RECT 2110.930 1577.090 2112.110 1578.270 ;
        RECT 2110.930 1575.490 2112.110 1576.670 ;
        RECT 2110.930 1397.090 2112.110 1398.270 ;
        RECT 2110.930 1395.490 2112.110 1396.670 ;
        RECT 2110.930 1217.090 2112.110 1218.270 ;
        RECT 2110.930 1215.490 2112.110 1216.670 ;
        RECT 2110.930 1037.090 2112.110 1038.270 ;
        RECT 2110.930 1035.490 2112.110 1036.670 ;
        RECT 2110.930 857.090 2112.110 858.270 ;
        RECT 2110.930 855.490 2112.110 856.670 ;
        RECT 2110.930 677.090 2112.110 678.270 ;
        RECT 2110.930 675.490 2112.110 676.670 ;
        RECT 2110.930 497.090 2112.110 498.270 ;
        RECT 2110.930 495.490 2112.110 496.670 ;
        RECT 2110.930 317.090 2112.110 318.270 ;
        RECT 2110.930 315.490 2112.110 316.670 ;
        RECT 2110.930 137.090 2112.110 138.270 ;
        RECT 2110.930 135.490 2112.110 136.670 ;
        RECT 2110.930 -25.910 2112.110 -24.730 ;
        RECT 2110.930 -27.510 2112.110 -26.330 ;
        RECT 2290.930 3546.010 2292.110 3547.190 ;
        RECT 2290.930 3544.410 2292.110 3545.590 ;
        RECT 2290.930 3377.090 2292.110 3378.270 ;
        RECT 2290.930 3375.490 2292.110 3376.670 ;
        RECT 2290.930 3197.090 2292.110 3198.270 ;
        RECT 2290.930 3195.490 2292.110 3196.670 ;
        RECT 2290.930 3017.090 2292.110 3018.270 ;
        RECT 2290.930 3015.490 2292.110 3016.670 ;
        RECT 2290.930 2837.090 2292.110 2838.270 ;
        RECT 2290.930 2835.490 2292.110 2836.670 ;
        RECT 2290.930 2657.090 2292.110 2658.270 ;
        RECT 2290.930 2655.490 2292.110 2656.670 ;
        RECT 2290.930 2477.090 2292.110 2478.270 ;
        RECT 2290.930 2475.490 2292.110 2476.670 ;
        RECT 2290.930 2297.090 2292.110 2298.270 ;
        RECT 2290.930 2295.490 2292.110 2296.670 ;
        RECT 2290.930 2117.090 2292.110 2118.270 ;
        RECT 2290.930 2115.490 2292.110 2116.670 ;
        RECT 2290.930 1937.090 2292.110 1938.270 ;
        RECT 2290.930 1935.490 2292.110 1936.670 ;
        RECT 2290.930 1757.090 2292.110 1758.270 ;
        RECT 2290.930 1755.490 2292.110 1756.670 ;
        RECT 2290.930 1577.090 2292.110 1578.270 ;
        RECT 2290.930 1575.490 2292.110 1576.670 ;
        RECT 2290.930 1397.090 2292.110 1398.270 ;
        RECT 2290.930 1395.490 2292.110 1396.670 ;
        RECT 2290.930 1217.090 2292.110 1218.270 ;
        RECT 2290.930 1215.490 2292.110 1216.670 ;
        RECT 2290.930 1037.090 2292.110 1038.270 ;
        RECT 2290.930 1035.490 2292.110 1036.670 ;
        RECT 2290.930 857.090 2292.110 858.270 ;
        RECT 2290.930 855.490 2292.110 856.670 ;
        RECT 2290.930 677.090 2292.110 678.270 ;
        RECT 2290.930 675.490 2292.110 676.670 ;
        RECT 2290.930 497.090 2292.110 498.270 ;
        RECT 2290.930 495.490 2292.110 496.670 ;
        RECT 2290.930 317.090 2292.110 318.270 ;
        RECT 2290.930 315.490 2292.110 316.670 ;
        RECT 2290.930 137.090 2292.110 138.270 ;
        RECT 2290.930 135.490 2292.110 136.670 ;
        RECT 2290.930 -25.910 2292.110 -24.730 ;
        RECT 2290.930 -27.510 2292.110 -26.330 ;
        RECT 2470.930 3546.010 2472.110 3547.190 ;
        RECT 2470.930 3544.410 2472.110 3545.590 ;
        RECT 2470.930 3377.090 2472.110 3378.270 ;
        RECT 2470.930 3375.490 2472.110 3376.670 ;
        RECT 2470.930 3197.090 2472.110 3198.270 ;
        RECT 2470.930 3195.490 2472.110 3196.670 ;
        RECT 2470.930 3017.090 2472.110 3018.270 ;
        RECT 2470.930 3015.490 2472.110 3016.670 ;
        RECT 2470.930 2837.090 2472.110 2838.270 ;
        RECT 2470.930 2835.490 2472.110 2836.670 ;
        RECT 2470.930 2657.090 2472.110 2658.270 ;
        RECT 2470.930 2655.490 2472.110 2656.670 ;
        RECT 2470.930 2477.090 2472.110 2478.270 ;
        RECT 2470.930 2475.490 2472.110 2476.670 ;
        RECT 2470.930 2297.090 2472.110 2298.270 ;
        RECT 2470.930 2295.490 2472.110 2296.670 ;
        RECT 2470.930 2117.090 2472.110 2118.270 ;
        RECT 2470.930 2115.490 2472.110 2116.670 ;
        RECT 2470.930 1937.090 2472.110 1938.270 ;
        RECT 2470.930 1935.490 2472.110 1936.670 ;
        RECT 2470.930 1757.090 2472.110 1758.270 ;
        RECT 2470.930 1755.490 2472.110 1756.670 ;
        RECT 2470.930 1577.090 2472.110 1578.270 ;
        RECT 2470.930 1575.490 2472.110 1576.670 ;
        RECT 2470.930 1397.090 2472.110 1398.270 ;
        RECT 2470.930 1395.490 2472.110 1396.670 ;
        RECT 2470.930 1217.090 2472.110 1218.270 ;
        RECT 2470.930 1215.490 2472.110 1216.670 ;
        RECT 2470.930 1037.090 2472.110 1038.270 ;
        RECT 2470.930 1035.490 2472.110 1036.670 ;
        RECT 2470.930 857.090 2472.110 858.270 ;
        RECT 2470.930 855.490 2472.110 856.670 ;
        RECT 2470.930 677.090 2472.110 678.270 ;
        RECT 2470.930 675.490 2472.110 676.670 ;
        RECT 2470.930 497.090 2472.110 498.270 ;
        RECT 2470.930 495.490 2472.110 496.670 ;
        RECT 2470.930 317.090 2472.110 318.270 ;
        RECT 2470.930 315.490 2472.110 316.670 ;
        RECT 2470.930 137.090 2472.110 138.270 ;
        RECT 2470.930 135.490 2472.110 136.670 ;
        RECT 2470.930 -25.910 2472.110 -24.730 ;
        RECT 2470.930 -27.510 2472.110 -26.330 ;
        RECT 2650.930 3546.010 2652.110 3547.190 ;
        RECT 2650.930 3544.410 2652.110 3545.590 ;
        RECT 2650.930 3377.090 2652.110 3378.270 ;
        RECT 2650.930 3375.490 2652.110 3376.670 ;
        RECT 2650.930 3197.090 2652.110 3198.270 ;
        RECT 2650.930 3195.490 2652.110 3196.670 ;
        RECT 2650.930 3017.090 2652.110 3018.270 ;
        RECT 2650.930 3015.490 2652.110 3016.670 ;
        RECT 2650.930 2837.090 2652.110 2838.270 ;
        RECT 2650.930 2835.490 2652.110 2836.670 ;
        RECT 2650.930 2657.090 2652.110 2658.270 ;
        RECT 2650.930 2655.490 2652.110 2656.670 ;
        RECT 2650.930 2477.090 2652.110 2478.270 ;
        RECT 2650.930 2475.490 2652.110 2476.670 ;
        RECT 2650.930 2297.090 2652.110 2298.270 ;
        RECT 2650.930 2295.490 2652.110 2296.670 ;
        RECT 2650.930 2117.090 2652.110 2118.270 ;
        RECT 2650.930 2115.490 2652.110 2116.670 ;
        RECT 2650.930 1937.090 2652.110 1938.270 ;
        RECT 2650.930 1935.490 2652.110 1936.670 ;
        RECT 2650.930 1757.090 2652.110 1758.270 ;
        RECT 2650.930 1755.490 2652.110 1756.670 ;
        RECT 2650.930 1577.090 2652.110 1578.270 ;
        RECT 2650.930 1575.490 2652.110 1576.670 ;
        RECT 2650.930 1397.090 2652.110 1398.270 ;
        RECT 2650.930 1395.490 2652.110 1396.670 ;
        RECT 2650.930 1217.090 2652.110 1218.270 ;
        RECT 2650.930 1215.490 2652.110 1216.670 ;
        RECT 2650.930 1037.090 2652.110 1038.270 ;
        RECT 2650.930 1035.490 2652.110 1036.670 ;
        RECT 2650.930 857.090 2652.110 858.270 ;
        RECT 2650.930 855.490 2652.110 856.670 ;
        RECT 2650.930 677.090 2652.110 678.270 ;
        RECT 2650.930 675.490 2652.110 676.670 ;
        RECT 2650.930 497.090 2652.110 498.270 ;
        RECT 2650.930 495.490 2652.110 496.670 ;
        RECT 2650.930 317.090 2652.110 318.270 ;
        RECT 2650.930 315.490 2652.110 316.670 ;
        RECT 2650.930 137.090 2652.110 138.270 ;
        RECT 2650.930 135.490 2652.110 136.670 ;
        RECT 2650.930 -25.910 2652.110 -24.730 ;
        RECT 2650.930 -27.510 2652.110 -26.330 ;
        RECT 2830.930 3546.010 2832.110 3547.190 ;
        RECT 2830.930 3544.410 2832.110 3545.590 ;
        RECT 2830.930 3377.090 2832.110 3378.270 ;
        RECT 2830.930 3375.490 2832.110 3376.670 ;
        RECT 2830.930 3197.090 2832.110 3198.270 ;
        RECT 2830.930 3195.490 2832.110 3196.670 ;
        RECT 2830.930 3017.090 2832.110 3018.270 ;
        RECT 2830.930 3015.490 2832.110 3016.670 ;
        RECT 2830.930 2837.090 2832.110 2838.270 ;
        RECT 2830.930 2835.490 2832.110 2836.670 ;
        RECT 2830.930 2657.090 2832.110 2658.270 ;
        RECT 2830.930 2655.490 2832.110 2656.670 ;
        RECT 2830.930 2477.090 2832.110 2478.270 ;
        RECT 2830.930 2475.490 2832.110 2476.670 ;
        RECT 2830.930 2297.090 2832.110 2298.270 ;
        RECT 2830.930 2295.490 2832.110 2296.670 ;
        RECT 2830.930 2117.090 2832.110 2118.270 ;
        RECT 2830.930 2115.490 2832.110 2116.670 ;
        RECT 2830.930 1937.090 2832.110 1938.270 ;
        RECT 2830.930 1935.490 2832.110 1936.670 ;
        RECT 2830.930 1757.090 2832.110 1758.270 ;
        RECT 2830.930 1755.490 2832.110 1756.670 ;
        RECT 2830.930 1577.090 2832.110 1578.270 ;
        RECT 2830.930 1575.490 2832.110 1576.670 ;
        RECT 2830.930 1397.090 2832.110 1398.270 ;
        RECT 2830.930 1395.490 2832.110 1396.670 ;
        RECT 2830.930 1217.090 2832.110 1218.270 ;
        RECT 2830.930 1215.490 2832.110 1216.670 ;
        RECT 2830.930 1037.090 2832.110 1038.270 ;
        RECT 2830.930 1035.490 2832.110 1036.670 ;
        RECT 2830.930 857.090 2832.110 858.270 ;
        RECT 2830.930 855.490 2832.110 856.670 ;
        RECT 2830.930 677.090 2832.110 678.270 ;
        RECT 2830.930 675.490 2832.110 676.670 ;
        RECT 2830.930 497.090 2832.110 498.270 ;
        RECT 2830.930 495.490 2832.110 496.670 ;
        RECT 2830.930 317.090 2832.110 318.270 ;
        RECT 2830.930 315.490 2832.110 316.670 ;
        RECT 2830.930 137.090 2832.110 138.270 ;
        RECT 2830.930 135.490 2832.110 136.670 ;
        RECT 2830.930 -25.910 2832.110 -24.730 ;
        RECT 2830.930 -27.510 2832.110 -26.330 ;
        RECT 2950.510 3546.010 2951.690 3547.190 ;
        RECT 2950.510 3544.410 2951.690 3545.590 ;
        RECT 2950.510 3377.090 2951.690 3378.270 ;
        RECT 2950.510 3375.490 2951.690 3376.670 ;
        RECT 2950.510 3197.090 2951.690 3198.270 ;
        RECT 2950.510 3195.490 2951.690 3196.670 ;
        RECT 2950.510 3017.090 2951.690 3018.270 ;
        RECT 2950.510 3015.490 2951.690 3016.670 ;
        RECT 2950.510 2837.090 2951.690 2838.270 ;
        RECT 2950.510 2835.490 2951.690 2836.670 ;
        RECT 2950.510 2657.090 2951.690 2658.270 ;
        RECT 2950.510 2655.490 2951.690 2656.670 ;
        RECT 2950.510 2477.090 2951.690 2478.270 ;
        RECT 2950.510 2475.490 2951.690 2476.670 ;
        RECT 2950.510 2297.090 2951.690 2298.270 ;
        RECT 2950.510 2295.490 2951.690 2296.670 ;
        RECT 2950.510 2117.090 2951.690 2118.270 ;
        RECT 2950.510 2115.490 2951.690 2116.670 ;
        RECT 2950.510 1937.090 2951.690 1938.270 ;
        RECT 2950.510 1935.490 2951.690 1936.670 ;
        RECT 2950.510 1757.090 2951.690 1758.270 ;
        RECT 2950.510 1755.490 2951.690 1756.670 ;
        RECT 2950.510 1577.090 2951.690 1578.270 ;
        RECT 2950.510 1575.490 2951.690 1576.670 ;
        RECT 2950.510 1397.090 2951.690 1398.270 ;
        RECT 2950.510 1395.490 2951.690 1396.670 ;
        RECT 2950.510 1217.090 2951.690 1218.270 ;
        RECT 2950.510 1215.490 2951.690 1216.670 ;
        RECT 2950.510 1037.090 2951.690 1038.270 ;
        RECT 2950.510 1035.490 2951.690 1036.670 ;
        RECT 2950.510 857.090 2951.690 858.270 ;
        RECT 2950.510 855.490 2951.690 856.670 ;
        RECT 2950.510 677.090 2951.690 678.270 ;
        RECT 2950.510 675.490 2951.690 676.670 ;
        RECT 2950.510 497.090 2951.690 498.270 ;
        RECT 2950.510 495.490 2951.690 496.670 ;
        RECT 2950.510 317.090 2951.690 318.270 ;
        RECT 2950.510 315.490 2951.690 316.670 ;
        RECT 2950.510 137.090 2951.690 138.270 ;
        RECT 2950.510 135.490 2951.690 136.670 ;
        RECT 2950.510 -25.910 2951.690 -24.730 ;
        RECT 2950.510 -27.510 2951.690 -26.330 ;
      LAYER met5 ;
        RECT -32.980 3547.300 -29.980 3547.310 ;
        RECT 130.020 3547.300 133.020 3547.310 ;
        RECT 310.020 3547.300 313.020 3547.310 ;
        RECT 490.020 3547.300 493.020 3547.310 ;
        RECT 670.020 3547.300 673.020 3547.310 ;
        RECT 850.020 3547.300 853.020 3547.310 ;
        RECT 1030.020 3547.300 1033.020 3547.310 ;
        RECT 1210.020 3547.300 1213.020 3547.310 ;
        RECT 1390.020 3547.300 1393.020 3547.310 ;
        RECT 1570.020 3547.300 1573.020 3547.310 ;
        RECT 1750.020 3547.300 1753.020 3547.310 ;
        RECT 1930.020 3547.300 1933.020 3547.310 ;
        RECT 2110.020 3547.300 2113.020 3547.310 ;
        RECT 2290.020 3547.300 2293.020 3547.310 ;
        RECT 2470.020 3547.300 2473.020 3547.310 ;
        RECT 2650.020 3547.300 2653.020 3547.310 ;
        RECT 2830.020 3547.300 2833.020 3547.310 ;
        RECT 2949.600 3547.300 2952.600 3547.310 ;
        RECT -32.980 3544.300 2952.600 3547.300 ;
        RECT -32.980 3544.290 -29.980 3544.300 ;
        RECT 130.020 3544.290 133.020 3544.300 ;
        RECT 310.020 3544.290 313.020 3544.300 ;
        RECT 490.020 3544.290 493.020 3544.300 ;
        RECT 670.020 3544.290 673.020 3544.300 ;
        RECT 850.020 3544.290 853.020 3544.300 ;
        RECT 1030.020 3544.290 1033.020 3544.300 ;
        RECT 1210.020 3544.290 1213.020 3544.300 ;
        RECT 1390.020 3544.290 1393.020 3544.300 ;
        RECT 1570.020 3544.290 1573.020 3544.300 ;
        RECT 1750.020 3544.290 1753.020 3544.300 ;
        RECT 1930.020 3544.290 1933.020 3544.300 ;
        RECT 2110.020 3544.290 2113.020 3544.300 ;
        RECT 2290.020 3544.290 2293.020 3544.300 ;
        RECT 2470.020 3544.290 2473.020 3544.300 ;
        RECT 2650.020 3544.290 2653.020 3544.300 ;
        RECT 2830.020 3544.290 2833.020 3544.300 ;
        RECT 2949.600 3544.290 2952.600 3544.300 ;
        RECT -32.980 3378.380 -29.980 3378.390 ;
        RECT 130.020 3378.380 133.020 3378.390 ;
        RECT 310.020 3378.380 313.020 3378.390 ;
        RECT 490.020 3378.380 493.020 3378.390 ;
        RECT 670.020 3378.380 673.020 3378.390 ;
        RECT 850.020 3378.380 853.020 3378.390 ;
        RECT 1030.020 3378.380 1033.020 3378.390 ;
        RECT 1210.020 3378.380 1213.020 3378.390 ;
        RECT 1390.020 3378.380 1393.020 3378.390 ;
        RECT 1570.020 3378.380 1573.020 3378.390 ;
        RECT 1750.020 3378.380 1753.020 3378.390 ;
        RECT 1930.020 3378.380 1933.020 3378.390 ;
        RECT 2110.020 3378.380 2113.020 3378.390 ;
        RECT 2290.020 3378.380 2293.020 3378.390 ;
        RECT 2470.020 3378.380 2473.020 3378.390 ;
        RECT 2650.020 3378.380 2653.020 3378.390 ;
        RECT 2830.020 3378.380 2833.020 3378.390 ;
        RECT 2949.600 3378.380 2952.600 3378.390 ;
        RECT -32.980 3375.380 2952.600 3378.380 ;
        RECT -32.980 3375.370 -29.980 3375.380 ;
        RECT 130.020 3375.370 133.020 3375.380 ;
        RECT 310.020 3375.370 313.020 3375.380 ;
        RECT 490.020 3375.370 493.020 3375.380 ;
        RECT 670.020 3375.370 673.020 3375.380 ;
        RECT 850.020 3375.370 853.020 3375.380 ;
        RECT 1030.020 3375.370 1033.020 3375.380 ;
        RECT 1210.020 3375.370 1213.020 3375.380 ;
        RECT 1390.020 3375.370 1393.020 3375.380 ;
        RECT 1570.020 3375.370 1573.020 3375.380 ;
        RECT 1750.020 3375.370 1753.020 3375.380 ;
        RECT 1930.020 3375.370 1933.020 3375.380 ;
        RECT 2110.020 3375.370 2113.020 3375.380 ;
        RECT 2290.020 3375.370 2293.020 3375.380 ;
        RECT 2470.020 3375.370 2473.020 3375.380 ;
        RECT 2650.020 3375.370 2653.020 3375.380 ;
        RECT 2830.020 3375.370 2833.020 3375.380 ;
        RECT 2949.600 3375.370 2952.600 3375.380 ;
        RECT -32.980 3198.380 -29.980 3198.390 ;
        RECT 130.020 3198.380 133.020 3198.390 ;
        RECT 310.020 3198.380 313.020 3198.390 ;
        RECT 490.020 3198.380 493.020 3198.390 ;
        RECT 670.020 3198.380 673.020 3198.390 ;
        RECT 850.020 3198.380 853.020 3198.390 ;
        RECT 1030.020 3198.380 1033.020 3198.390 ;
        RECT 1210.020 3198.380 1213.020 3198.390 ;
        RECT 1390.020 3198.380 1393.020 3198.390 ;
        RECT 1570.020 3198.380 1573.020 3198.390 ;
        RECT 1750.020 3198.380 1753.020 3198.390 ;
        RECT 1930.020 3198.380 1933.020 3198.390 ;
        RECT 2110.020 3198.380 2113.020 3198.390 ;
        RECT 2290.020 3198.380 2293.020 3198.390 ;
        RECT 2470.020 3198.380 2473.020 3198.390 ;
        RECT 2650.020 3198.380 2653.020 3198.390 ;
        RECT 2830.020 3198.380 2833.020 3198.390 ;
        RECT 2949.600 3198.380 2952.600 3198.390 ;
        RECT -32.980 3195.380 2952.600 3198.380 ;
        RECT -32.980 3195.370 -29.980 3195.380 ;
        RECT 130.020 3195.370 133.020 3195.380 ;
        RECT 310.020 3195.370 313.020 3195.380 ;
        RECT 490.020 3195.370 493.020 3195.380 ;
        RECT 670.020 3195.370 673.020 3195.380 ;
        RECT 850.020 3195.370 853.020 3195.380 ;
        RECT 1030.020 3195.370 1033.020 3195.380 ;
        RECT 1210.020 3195.370 1213.020 3195.380 ;
        RECT 1390.020 3195.370 1393.020 3195.380 ;
        RECT 1570.020 3195.370 1573.020 3195.380 ;
        RECT 1750.020 3195.370 1753.020 3195.380 ;
        RECT 1930.020 3195.370 1933.020 3195.380 ;
        RECT 2110.020 3195.370 2113.020 3195.380 ;
        RECT 2290.020 3195.370 2293.020 3195.380 ;
        RECT 2470.020 3195.370 2473.020 3195.380 ;
        RECT 2650.020 3195.370 2653.020 3195.380 ;
        RECT 2830.020 3195.370 2833.020 3195.380 ;
        RECT 2949.600 3195.370 2952.600 3195.380 ;
        RECT -32.980 3018.380 -29.980 3018.390 ;
        RECT 130.020 3018.380 133.020 3018.390 ;
        RECT 310.020 3018.380 313.020 3018.390 ;
        RECT 490.020 3018.380 493.020 3018.390 ;
        RECT 670.020 3018.380 673.020 3018.390 ;
        RECT 850.020 3018.380 853.020 3018.390 ;
        RECT 1030.020 3018.380 1033.020 3018.390 ;
        RECT 1210.020 3018.380 1213.020 3018.390 ;
        RECT 1390.020 3018.380 1393.020 3018.390 ;
        RECT 1570.020 3018.380 1573.020 3018.390 ;
        RECT 1750.020 3018.380 1753.020 3018.390 ;
        RECT 1930.020 3018.380 1933.020 3018.390 ;
        RECT 2110.020 3018.380 2113.020 3018.390 ;
        RECT 2290.020 3018.380 2293.020 3018.390 ;
        RECT 2470.020 3018.380 2473.020 3018.390 ;
        RECT 2650.020 3018.380 2653.020 3018.390 ;
        RECT 2830.020 3018.380 2833.020 3018.390 ;
        RECT 2949.600 3018.380 2952.600 3018.390 ;
        RECT -32.980 3015.380 2952.600 3018.380 ;
        RECT -32.980 3015.370 -29.980 3015.380 ;
        RECT 130.020 3015.370 133.020 3015.380 ;
        RECT 310.020 3015.370 313.020 3015.380 ;
        RECT 490.020 3015.370 493.020 3015.380 ;
        RECT 670.020 3015.370 673.020 3015.380 ;
        RECT 850.020 3015.370 853.020 3015.380 ;
        RECT 1030.020 3015.370 1033.020 3015.380 ;
        RECT 1210.020 3015.370 1213.020 3015.380 ;
        RECT 1390.020 3015.370 1393.020 3015.380 ;
        RECT 1570.020 3015.370 1573.020 3015.380 ;
        RECT 1750.020 3015.370 1753.020 3015.380 ;
        RECT 1930.020 3015.370 1933.020 3015.380 ;
        RECT 2110.020 3015.370 2113.020 3015.380 ;
        RECT 2290.020 3015.370 2293.020 3015.380 ;
        RECT 2470.020 3015.370 2473.020 3015.380 ;
        RECT 2650.020 3015.370 2653.020 3015.380 ;
        RECT 2830.020 3015.370 2833.020 3015.380 ;
        RECT 2949.600 3015.370 2952.600 3015.380 ;
        RECT -32.980 2838.380 -29.980 2838.390 ;
        RECT 130.020 2838.380 133.020 2838.390 ;
        RECT 310.020 2838.380 313.020 2838.390 ;
        RECT 490.020 2838.380 493.020 2838.390 ;
        RECT 670.020 2838.380 673.020 2838.390 ;
        RECT 850.020 2838.380 853.020 2838.390 ;
        RECT 1030.020 2838.380 1033.020 2838.390 ;
        RECT 1210.020 2838.380 1213.020 2838.390 ;
        RECT 1390.020 2838.380 1393.020 2838.390 ;
        RECT 1570.020 2838.380 1573.020 2838.390 ;
        RECT 1750.020 2838.380 1753.020 2838.390 ;
        RECT 1930.020 2838.380 1933.020 2838.390 ;
        RECT 2110.020 2838.380 2113.020 2838.390 ;
        RECT 2290.020 2838.380 2293.020 2838.390 ;
        RECT 2470.020 2838.380 2473.020 2838.390 ;
        RECT 2650.020 2838.380 2653.020 2838.390 ;
        RECT 2830.020 2838.380 2833.020 2838.390 ;
        RECT 2949.600 2838.380 2952.600 2838.390 ;
        RECT -32.980 2835.380 2952.600 2838.380 ;
        RECT -32.980 2835.370 -29.980 2835.380 ;
        RECT 130.020 2835.370 133.020 2835.380 ;
        RECT 310.020 2835.370 313.020 2835.380 ;
        RECT 490.020 2835.370 493.020 2835.380 ;
        RECT 670.020 2835.370 673.020 2835.380 ;
        RECT 850.020 2835.370 853.020 2835.380 ;
        RECT 1030.020 2835.370 1033.020 2835.380 ;
        RECT 1210.020 2835.370 1213.020 2835.380 ;
        RECT 1390.020 2835.370 1393.020 2835.380 ;
        RECT 1570.020 2835.370 1573.020 2835.380 ;
        RECT 1750.020 2835.370 1753.020 2835.380 ;
        RECT 1930.020 2835.370 1933.020 2835.380 ;
        RECT 2110.020 2835.370 2113.020 2835.380 ;
        RECT 2290.020 2835.370 2293.020 2835.380 ;
        RECT 2470.020 2835.370 2473.020 2835.380 ;
        RECT 2650.020 2835.370 2653.020 2835.380 ;
        RECT 2830.020 2835.370 2833.020 2835.380 ;
        RECT 2949.600 2835.370 2952.600 2835.380 ;
        RECT -32.980 2658.380 -29.980 2658.390 ;
        RECT 130.020 2658.380 133.020 2658.390 ;
        RECT 310.020 2658.380 313.020 2658.390 ;
        RECT 490.020 2658.380 493.020 2658.390 ;
        RECT 670.020 2658.380 673.020 2658.390 ;
        RECT 850.020 2658.380 853.020 2658.390 ;
        RECT 1030.020 2658.380 1033.020 2658.390 ;
        RECT 1210.020 2658.380 1213.020 2658.390 ;
        RECT 1390.020 2658.380 1393.020 2658.390 ;
        RECT 1570.020 2658.380 1573.020 2658.390 ;
        RECT 1750.020 2658.380 1753.020 2658.390 ;
        RECT 1930.020 2658.380 1933.020 2658.390 ;
        RECT 2110.020 2658.380 2113.020 2658.390 ;
        RECT 2290.020 2658.380 2293.020 2658.390 ;
        RECT 2470.020 2658.380 2473.020 2658.390 ;
        RECT 2650.020 2658.380 2653.020 2658.390 ;
        RECT 2830.020 2658.380 2833.020 2658.390 ;
        RECT 2949.600 2658.380 2952.600 2658.390 ;
        RECT -32.980 2655.380 2952.600 2658.380 ;
        RECT -32.980 2655.370 -29.980 2655.380 ;
        RECT 130.020 2655.370 133.020 2655.380 ;
        RECT 310.020 2655.370 313.020 2655.380 ;
        RECT 490.020 2655.370 493.020 2655.380 ;
        RECT 670.020 2655.370 673.020 2655.380 ;
        RECT 850.020 2655.370 853.020 2655.380 ;
        RECT 1030.020 2655.370 1033.020 2655.380 ;
        RECT 1210.020 2655.370 1213.020 2655.380 ;
        RECT 1390.020 2655.370 1393.020 2655.380 ;
        RECT 1570.020 2655.370 1573.020 2655.380 ;
        RECT 1750.020 2655.370 1753.020 2655.380 ;
        RECT 1930.020 2655.370 1933.020 2655.380 ;
        RECT 2110.020 2655.370 2113.020 2655.380 ;
        RECT 2290.020 2655.370 2293.020 2655.380 ;
        RECT 2470.020 2655.370 2473.020 2655.380 ;
        RECT 2650.020 2655.370 2653.020 2655.380 ;
        RECT 2830.020 2655.370 2833.020 2655.380 ;
        RECT 2949.600 2655.370 2952.600 2655.380 ;
        RECT -32.980 2478.380 -29.980 2478.390 ;
        RECT 130.020 2478.380 133.020 2478.390 ;
        RECT 310.020 2478.380 313.020 2478.390 ;
        RECT 490.020 2478.380 493.020 2478.390 ;
        RECT 670.020 2478.380 673.020 2478.390 ;
        RECT 850.020 2478.380 853.020 2478.390 ;
        RECT 1030.020 2478.380 1033.020 2478.390 ;
        RECT 1210.020 2478.380 1213.020 2478.390 ;
        RECT 1390.020 2478.380 1393.020 2478.390 ;
        RECT 1570.020 2478.380 1573.020 2478.390 ;
        RECT 1750.020 2478.380 1753.020 2478.390 ;
        RECT 1930.020 2478.380 1933.020 2478.390 ;
        RECT 2110.020 2478.380 2113.020 2478.390 ;
        RECT 2290.020 2478.380 2293.020 2478.390 ;
        RECT 2470.020 2478.380 2473.020 2478.390 ;
        RECT 2650.020 2478.380 2653.020 2478.390 ;
        RECT 2830.020 2478.380 2833.020 2478.390 ;
        RECT 2949.600 2478.380 2952.600 2478.390 ;
        RECT -32.980 2475.380 2952.600 2478.380 ;
        RECT -32.980 2475.370 -29.980 2475.380 ;
        RECT 130.020 2475.370 133.020 2475.380 ;
        RECT 310.020 2475.370 313.020 2475.380 ;
        RECT 490.020 2475.370 493.020 2475.380 ;
        RECT 670.020 2475.370 673.020 2475.380 ;
        RECT 850.020 2475.370 853.020 2475.380 ;
        RECT 1030.020 2475.370 1033.020 2475.380 ;
        RECT 1210.020 2475.370 1213.020 2475.380 ;
        RECT 1390.020 2475.370 1393.020 2475.380 ;
        RECT 1570.020 2475.370 1573.020 2475.380 ;
        RECT 1750.020 2475.370 1753.020 2475.380 ;
        RECT 1930.020 2475.370 1933.020 2475.380 ;
        RECT 2110.020 2475.370 2113.020 2475.380 ;
        RECT 2290.020 2475.370 2293.020 2475.380 ;
        RECT 2470.020 2475.370 2473.020 2475.380 ;
        RECT 2650.020 2475.370 2653.020 2475.380 ;
        RECT 2830.020 2475.370 2833.020 2475.380 ;
        RECT 2949.600 2475.370 2952.600 2475.380 ;
        RECT -32.980 2298.380 -29.980 2298.390 ;
        RECT 130.020 2298.380 133.020 2298.390 ;
        RECT 310.020 2298.380 313.020 2298.390 ;
        RECT 490.020 2298.380 493.020 2298.390 ;
        RECT 670.020 2298.380 673.020 2298.390 ;
        RECT 850.020 2298.380 853.020 2298.390 ;
        RECT 1030.020 2298.380 1033.020 2298.390 ;
        RECT 1210.020 2298.380 1213.020 2298.390 ;
        RECT 1390.020 2298.380 1393.020 2298.390 ;
        RECT 1570.020 2298.380 1573.020 2298.390 ;
        RECT 1750.020 2298.380 1753.020 2298.390 ;
        RECT 1930.020 2298.380 1933.020 2298.390 ;
        RECT 2110.020 2298.380 2113.020 2298.390 ;
        RECT 2290.020 2298.380 2293.020 2298.390 ;
        RECT 2470.020 2298.380 2473.020 2298.390 ;
        RECT 2650.020 2298.380 2653.020 2298.390 ;
        RECT 2830.020 2298.380 2833.020 2298.390 ;
        RECT 2949.600 2298.380 2952.600 2298.390 ;
        RECT -32.980 2295.380 2952.600 2298.380 ;
        RECT -32.980 2295.370 -29.980 2295.380 ;
        RECT 130.020 2295.370 133.020 2295.380 ;
        RECT 310.020 2295.370 313.020 2295.380 ;
        RECT 490.020 2295.370 493.020 2295.380 ;
        RECT 670.020 2295.370 673.020 2295.380 ;
        RECT 850.020 2295.370 853.020 2295.380 ;
        RECT 1030.020 2295.370 1033.020 2295.380 ;
        RECT 1210.020 2295.370 1213.020 2295.380 ;
        RECT 1390.020 2295.370 1393.020 2295.380 ;
        RECT 1570.020 2295.370 1573.020 2295.380 ;
        RECT 1750.020 2295.370 1753.020 2295.380 ;
        RECT 1930.020 2295.370 1933.020 2295.380 ;
        RECT 2110.020 2295.370 2113.020 2295.380 ;
        RECT 2290.020 2295.370 2293.020 2295.380 ;
        RECT 2470.020 2295.370 2473.020 2295.380 ;
        RECT 2650.020 2295.370 2653.020 2295.380 ;
        RECT 2830.020 2295.370 2833.020 2295.380 ;
        RECT 2949.600 2295.370 2952.600 2295.380 ;
        RECT -32.980 2118.380 -29.980 2118.390 ;
        RECT 130.020 2118.380 133.020 2118.390 ;
        RECT 310.020 2118.380 313.020 2118.390 ;
        RECT 490.020 2118.380 493.020 2118.390 ;
        RECT 670.020 2118.380 673.020 2118.390 ;
        RECT 850.020 2118.380 853.020 2118.390 ;
        RECT 1030.020 2118.380 1033.020 2118.390 ;
        RECT 1210.020 2118.380 1213.020 2118.390 ;
        RECT 1390.020 2118.380 1393.020 2118.390 ;
        RECT 1570.020 2118.380 1573.020 2118.390 ;
        RECT 1750.020 2118.380 1753.020 2118.390 ;
        RECT 1930.020 2118.380 1933.020 2118.390 ;
        RECT 2110.020 2118.380 2113.020 2118.390 ;
        RECT 2290.020 2118.380 2293.020 2118.390 ;
        RECT 2470.020 2118.380 2473.020 2118.390 ;
        RECT 2650.020 2118.380 2653.020 2118.390 ;
        RECT 2830.020 2118.380 2833.020 2118.390 ;
        RECT 2949.600 2118.380 2952.600 2118.390 ;
        RECT -32.980 2115.380 2952.600 2118.380 ;
        RECT -32.980 2115.370 -29.980 2115.380 ;
        RECT 130.020 2115.370 133.020 2115.380 ;
        RECT 310.020 2115.370 313.020 2115.380 ;
        RECT 490.020 2115.370 493.020 2115.380 ;
        RECT 670.020 2115.370 673.020 2115.380 ;
        RECT 850.020 2115.370 853.020 2115.380 ;
        RECT 1030.020 2115.370 1033.020 2115.380 ;
        RECT 1210.020 2115.370 1213.020 2115.380 ;
        RECT 1390.020 2115.370 1393.020 2115.380 ;
        RECT 1570.020 2115.370 1573.020 2115.380 ;
        RECT 1750.020 2115.370 1753.020 2115.380 ;
        RECT 1930.020 2115.370 1933.020 2115.380 ;
        RECT 2110.020 2115.370 2113.020 2115.380 ;
        RECT 2290.020 2115.370 2293.020 2115.380 ;
        RECT 2470.020 2115.370 2473.020 2115.380 ;
        RECT 2650.020 2115.370 2653.020 2115.380 ;
        RECT 2830.020 2115.370 2833.020 2115.380 ;
        RECT 2949.600 2115.370 2952.600 2115.380 ;
        RECT -32.980 1938.380 -29.980 1938.390 ;
        RECT 130.020 1938.380 133.020 1938.390 ;
        RECT 310.020 1938.380 313.020 1938.390 ;
        RECT 490.020 1938.380 493.020 1938.390 ;
        RECT 670.020 1938.380 673.020 1938.390 ;
        RECT 850.020 1938.380 853.020 1938.390 ;
        RECT 1030.020 1938.380 1033.020 1938.390 ;
        RECT 1210.020 1938.380 1213.020 1938.390 ;
        RECT 1390.020 1938.380 1393.020 1938.390 ;
        RECT 1570.020 1938.380 1573.020 1938.390 ;
        RECT 1750.020 1938.380 1753.020 1938.390 ;
        RECT 1930.020 1938.380 1933.020 1938.390 ;
        RECT 2110.020 1938.380 2113.020 1938.390 ;
        RECT 2290.020 1938.380 2293.020 1938.390 ;
        RECT 2470.020 1938.380 2473.020 1938.390 ;
        RECT 2650.020 1938.380 2653.020 1938.390 ;
        RECT 2830.020 1938.380 2833.020 1938.390 ;
        RECT 2949.600 1938.380 2952.600 1938.390 ;
        RECT -32.980 1935.380 2952.600 1938.380 ;
        RECT -32.980 1935.370 -29.980 1935.380 ;
        RECT 130.020 1935.370 133.020 1935.380 ;
        RECT 310.020 1935.370 313.020 1935.380 ;
        RECT 490.020 1935.370 493.020 1935.380 ;
        RECT 670.020 1935.370 673.020 1935.380 ;
        RECT 850.020 1935.370 853.020 1935.380 ;
        RECT 1030.020 1935.370 1033.020 1935.380 ;
        RECT 1210.020 1935.370 1213.020 1935.380 ;
        RECT 1390.020 1935.370 1393.020 1935.380 ;
        RECT 1570.020 1935.370 1573.020 1935.380 ;
        RECT 1750.020 1935.370 1753.020 1935.380 ;
        RECT 1930.020 1935.370 1933.020 1935.380 ;
        RECT 2110.020 1935.370 2113.020 1935.380 ;
        RECT 2290.020 1935.370 2293.020 1935.380 ;
        RECT 2470.020 1935.370 2473.020 1935.380 ;
        RECT 2650.020 1935.370 2653.020 1935.380 ;
        RECT 2830.020 1935.370 2833.020 1935.380 ;
        RECT 2949.600 1935.370 2952.600 1935.380 ;
        RECT -32.980 1758.380 -29.980 1758.390 ;
        RECT 130.020 1758.380 133.020 1758.390 ;
        RECT 310.020 1758.380 313.020 1758.390 ;
        RECT 490.020 1758.380 493.020 1758.390 ;
        RECT 670.020 1758.380 673.020 1758.390 ;
        RECT 850.020 1758.380 853.020 1758.390 ;
        RECT 1030.020 1758.380 1033.020 1758.390 ;
        RECT 1210.020 1758.380 1213.020 1758.390 ;
        RECT 1390.020 1758.380 1393.020 1758.390 ;
        RECT 1570.020 1758.380 1573.020 1758.390 ;
        RECT 1750.020 1758.380 1753.020 1758.390 ;
        RECT 1930.020 1758.380 1933.020 1758.390 ;
        RECT 2110.020 1758.380 2113.020 1758.390 ;
        RECT 2290.020 1758.380 2293.020 1758.390 ;
        RECT 2470.020 1758.380 2473.020 1758.390 ;
        RECT 2650.020 1758.380 2653.020 1758.390 ;
        RECT 2830.020 1758.380 2833.020 1758.390 ;
        RECT 2949.600 1758.380 2952.600 1758.390 ;
        RECT -32.980 1755.380 2952.600 1758.380 ;
        RECT -32.980 1755.370 -29.980 1755.380 ;
        RECT 130.020 1755.370 133.020 1755.380 ;
        RECT 310.020 1755.370 313.020 1755.380 ;
        RECT 490.020 1755.370 493.020 1755.380 ;
        RECT 670.020 1755.370 673.020 1755.380 ;
        RECT 850.020 1755.370 853.020 1755.380 ;
        RECT 1030.020 1755.370 1033.020 1755.380 ;
        RECT 1210.020 1755.370 1213.020 1755.380 ;
        RECT 1390.020 1755.370 1393.020 1755.380 ;
        RECT 1570.020 1755.370 1573.020 1755.380 ;
        RECT 1750.020 1755.370 1753.020 1755.380 ;
        RECT 1930.020 1755.370 1933.020 1755.380 ;
        RECT 2110.020 1755.370 2113.020 1755.380 ;
        RECT 2290.020 1755.370 2293.020 1755.380 ;
        RECT 2470.020 1755.370 2473.020 1755.380 ;
        RECT 2650.020 1755.370 2653.020 1755.380 ;
        RECT 2830.020 1755.370 2833.020 1755.380 ;
        RECT 2949.600 1755.370 2952.600 1755.380 ;
        RECT -32.980 1578.380 -29.980 1578.390 ;
        RECT 130.020 1578.380 133.020 1578.390 ;
        RECT 310.020 1578.380 313.020 1578.390 ;
        RECT 490.020 1578.380 493.020 1578.390 ;
        RECT 670.020 1578.380 673.020 1578.390 ;
        RECT 850.020 1578.380 853.020 1578.390 ;
        RECT 1030.020 1578.380 1033.020 1578.390 ;
        RECT 1210.020 1578.380 1213.020 1578.390 ;
        RECT 1390.020 1578.380 1393.020 1578.390 ;
        RECT 1570.020 1578.380 1573.020 1578.390 ;
        RECT 1750.020 1578.380 1753.020 1578.390 ;
        RECT 1930.020 1578.380 1933.020 1578.390 ;
        RECT 2110.020 1578.380 2113.020 1578.390 ;
        RECT 2290.020 1578.380 2293.020 1578.390 ;
        RECT 2470.020 1578.380 2473.020 1578.390 ;
        RECT 2650.020 1578.380 2653.020 1578.390 ;
        RECT 2830.020 1578.380 2833.020 1578.390 ;
        RECT 2949.600 1578.380 2952.600 1578.390 ;
        RECT -32.980 1575.380 2952.600 1578.380 ;
        RECT -32.980 1575.370 -29.980 1575.380 ;
        RECT 130.020 1575.370 133.020 1575.380 ;
        RECT 310.020 1575.370 313.020 1575.380 ;
        RECT 490.020 1575.370 493.020 1575.380 ;
        RECT 670.020 1575.370 673.020 1575.380 ;
        RECT 850.020 1575.370 853.020 1575.380 ;
        RECT 1030.020 1575.370 1033.020 1575.380 ;
        RECT 1210.020 1575.370 1213.020 1575.380 ;
        RECT 1390.020 1575.370 1393.020 1575.380 ;
        RECT 1570.020 1575.370 1573.020 1575.380 ;
        RECT 1750.020 1575.370 1753.020 1575.380 ;
        RECT 1930.020 1575.370 1933.020 1575.380 ;
        RECT 2110.020 1575.370 2113.020 1575.380 ;
        RECT 2290.020 1575.370 2293.020 1575.380 ;
        RECT 2470.020 1575.370 2473.020 1575.380 ;
        RECT 2650.020 1575.370 2653.020 1575.380 ;
        RECT 2830.020 1575.370 2833.020 1575.380 ;
        RECT 2949.600 1575.370 2952.600 1575.380 ;
        RECT -32.980 1398.380 -29.980 1398.390 ;
        RECT 130.020 1398.380 133.020 1398.390 ;
        RECT 310.020 1398.380 313.020 1398.390 ;
        RECT 490.020 1398.380 493.020 1398.390 ;
        RECT 670.020 1398.380 673.020 1398.390 ;
        RECT 850.020 1398.380 853.020 1398.390 ;
        RECT 1030.020 1398.380 1033.020 1398.390 ;
        RECT 1210.020 1398.380 1213.020 1398.390 ;
        RECT 1390.020 1398.380 1393.020 1398.390 ;
        RECT 1570.020 1398.380 1573.020 1398.390 ;
        RECT 1750.020 1398.380 1753.020 1398.390 ;
        RECT 1930.020 1398.380 1933.020 1398.390 ;
        RECT 2110.020 1398.380 2113.020 1398.390 ;
        RECT 2290.020 1398.380 2293.020 1398.390 ;
        RECT 2470.020 1398.380 2473.020 1398.390 ;
        RECT 2650.020 1398.380 2653.020 1398.390 ;
        RECT 2830.020 1398.380 2833.020 1398.390 ;
        RECT 2949.600 1398.380 2952.600 1398.390 ;
        RECT -32.980 1395.380 2952.600 1398.380 ;
        RECT -32.980 1395.370 -29.980 1395.380 ;
        RECT 130.020 1395.370 133.020 1395.380 ;
        RECT 310.020 1395.370 313.020 1395.380 ;
        RECT 490.020 1395.370 493.020 1395.380 ;
        RECT 670.020 1395.370 673.020 1395.380 ;
        RECT 850.020 1395.370 853.020 1395.380 ;
        RECT 1030.020 1395.370 1033.020 1395.380 ;
        RECT 1210.020 1395.370 1213.020 1395.380 ;
        RECT 1390.020 1395.370 1393.020 1395.380 ;
        RECT 1570.020 1395.370 1573.020 1395.380 ;
        RECT 1750.020 1395.370 1753.020 1395.380 ;
        RECT 1930.020 1395.370 1933.020 1395.380 ;
        RECT 2110.020 1395.370 2113.020 1395.380 ;
        RECT 2290.020 1395.370 2293.020 1395.380 ;
        RECT 2470.020 1395.370 2473.020 1395.380 ;
        RECT 2650.020 1395.370 2653.020 1395.380 ;
        RECT 2830.020 1395.370 2833.020 1395.380 ;
        RECT 2949.600 1395.370 2952.600 1395.380 ;
        RECT -32.980 1218.380 -29.980 1218.390 ;
        RECT 130.020 1218.380 133.020 1218.390 ;
        RECT 310.020 1218.380 313.020 1218.390 ;
        RECT 490.020 1218.380 493.020 1218.390 ;
        RECT 670.020 1218.380 673.020 1218.390 ;
        RECT 850.020 1218.380 853.020 1218.390 ;
        RECT 1030.020 1218.380 1033.020 1218.390 ;
        RECT 1210.020 1218.380 1213.020 1218.390 ;
        RECT 1390.020 1218.380 1393.020 1218.390 ;
        RECT 1570.020 1218.380 1573.020 1218.390 ;
        RECT 1750.020 1218.380 1753.020 1218.390 ;
        RECT 1930.020 1218.380 1933.020 1218.390 ;
        RECT 2110.020 1218.380 2113.020 1218.390 ;
        RECT 2290.020 1218.380 2293.020 1218.390 ;
        RECT 2470.020 1218.380 2473.020 1218.390 ;
        RECT 2650.020 1218.380 2653.020 1218.390 ;
        RECT 2830.020 1218.380 2833.020 1218.390 ;
        RECT 2949.600 1218.380 2952.600 1218.390 ;
        RECT -32.980 1215.380 2952.600 1218.380 ;
        RECT -32.980 1215.370 -29.980 1215.380 ;
        RECT 130.020 1215.370 133.020 1215.380 ;
        RECT 310.020 1215.370 313.020 1215.380 ;
        RECT 490.020 1215.370 493.020 1215.380 ;
        RECT 670.020 1215.370 673.020 1215.380 ;
        RECT 850.020 1215.370 853.020 1215.380 ;
        RECT 1030.020 1215.370 1033.020 1215.380 ;
        RECT 1210.020 1215.370 1213.020 1215.380 ;
        RECT 1390.020 1215.370 1393.020 1215.380 ;
        RECT 1570.020 1215.370 1573.020 1215.380 ;
        RECT 1750.020 1215.370 1753.020 1215.380 ;
        RECT 1930.020 1215.370 1933.020 1215.380 ;
        RECT 2110.020 1215.370 2113.020 1215.380 ;
        RECT 2290.020 1215.370 2293.020 1215.380 ;
        RECT 2470.020 1215.370 2473.020 1215.380 ;
        RECT 2650.020 1215.370 2653.020 1215.380 ;
        RECT 2830.020 1215.370 2833.020 1215.380 ;
        RECT 2949.600 1215.370 2952.600 1215.380 ;
        RECT -32.980 1038.380 -29.980 1038.390 ;
        RECT 130.020 1038.380 133.020 1038.390 ;
        RECT 310.020 1038.380 313.020 1038.390 ;
        RECT 490.020 1038.380 493.020 1038.390 ;
        RECT 670.020 1038.380 673.020 1038.390 ;
        RECT 850.020 1038.380 853.020 1038.390 ;
        RECT 1030.020 1038.380 1033.020 1038.390 ;
        RECT 1210.020 1038.380 1213.020 1038.390 ;
        RECT 1390.020 1038.380 1393.020 1038.390 ;
        RECT 1570.020 1038.380 1573.020 1038.390 ;
        RECT 1750.020 1038.380 1753.020 1038.390 ;
        RECT 1930.020 1038.380 1933.020 1038.390 ;
        RECT 2110.020 1038.380 2113.020 1038.390 ;
        RECT 2290.020 1038.380 2293.020 1038.390 ;
        RECT 2470.020 1038.380 2473.020 1038.390 ;
        RECT 2650.020 1038.380 2653.020 1038.390 ;
        RECT 2830.020 1038.380 2833.020 1038.390 ;
        RECT 2949.600 1038.380 2952.600 1038.390 ;
        RECT -32.980 1035.380 2952.600 1038.380 ;
        RECT -32.980 1035.370 -29.980 1035.380 ;
        RECT 130.020 1035.370 133.020 1035.380 ;
        RECT 310.020 1035.370 313.020 1035.380 ;
        RECT 490.020 1035.370 493.020 1035.380 ;
        RECT 670.020 1035.370 673.020 1035.380 ;
        RECT 850.020 1035.370 853.020 1035.380 ;
        RECT 1030.020 1035.370 1033.020 1035.380 ;
        RECT 1210.020 1035.370 1213.020 1035.380 ;
        RECT 1390.020 1035.370 1393.020 1035.380 ;
        RECT 1570.020 1035.370 1573.020 1035.380 ;
        RECT 1750.020 1035.370 1753.020 1035.380 ;
        RECT 1930.020 1035.370 1933.020 1035.380 ;
        RECT 2110.020 1035.370 2113.020 1035.380 ;
        RECT 2290.020 1035.370 2293.020 1035.380 ;
        RECT 2470.020 1035.370 2473.020 1035.380 ;
        RECT 2650.020 1035.370 2653.020 1035.380 ;
        RECT 2830.020 1035.370 2833.020 1035.380 ;
        RECT 2949.600 1035.370 2952.600 1035.380 ;
        RECT -32.980 858.380 -29.980 858.390 ;
        RECT 130.020 858.380 133.020 858.390 ;
        RECT 310.020 858.380 313.020 858.390 ;
        RECT 490.020 858.380 493.020 858.390 ;
        RECT 670.020 858.380 673.020 858.390 ;
        RECT 850.020 858.380 853.020 858.390 ;
        RECT 1030.020 858.380 1033.020 858.390 ;
        RECT 1210.020 858.380 1213.020 858.390 ;
        RECT 1390.020 858.380 1393.020 858.390 ;
        RECT 1570.020 858.380 1573.020 858.390 ;
        RECT 1750.020 858.380 1753.020 858.390 ;
        RECT 1930.020 858.380 1933.020 858.390 ;
        RECT 2110.020 858.380 2113.020 858.390 ;
        RECT 2290.020 858.380 2293.020 858.390 ;
        RECT 2470.020 858.380 2473.020 858.390 ;
        RECT 2650.020 858.380 2653.020 858.390 ;
        RECT 2830.020 858.380 2833.020 858.390 ;
        RECT 2949.600 858.380 2952.600 858.390 ;
        RECT -32.980 855.380 2952.600 858.380 ;
        RECT -32.980 855.370 -29.980 855.380 ;
        RECT 130.020 855.370 133.020 855.380 ;
        RECT 310.020 855.370 313.020 855.380 ;
        RECT 490.020 855.370 493.020 855.380 ;
        RECT 670.020 855.370 673.020 855.380 ;
        RECT 850.020 855.370 853.020 855.380 ;
        RECT 1030.020 855.370 1033.020 855.380 ;
        RECT 1210.020 855.370 1213.020 855.380 ;
        RECT 1390.020 855.370 1393.020 855.380 ;
        RECT 1570.020 855.370 1573.020 855.380 ;
        RECT 1750.020 855.370 1753.020 855.380 ;
        RECT 1930.020 855.370 1933.020 855.380 ;
        RECT 2110.020 855.370 2113.020 855.380 ;
        RECT 2290.020 855.370 2293.020 855.380 ;
        RECT 2470.020 855.370 2473.020 855.380 ;
        RECT 2650.020 855.370 2653.020 855.380 ;
        RECT 2830.020 855.370 2833.020 855.380 ;
        RECT 2949.600 855.370 2952.600 855.380 ;
        RECT -32.980 678.380 -29.980 678.390 ;
        RECT 130.020 678.380 133.020 678.390 ;
        RECT 310.020 678.380 313.020 678.390 ;
        RECT 490.020 678.380 493.020 678.390 ;
        RECT 670.020 678.380 673.020 678.390 ;
        RECT 850.020 678.380 853.020 678.390 ;
        RECT 1030.020 678.380 1033.020 678.390 ;
        RECT 1210.020 678.380 1213.020 678.390 ;
        RECT 1390.020 678.380 1393.020 678.390 ;
        RECT 1570.020 678.380 1573.020 678.390 ;
        RECT 1750.020 678.380 1753.020 678.390 ;
        RECT 1930.020 678.380 1933.020 678.390 ;
        RECT 2110.020 678.380 2113.020 678.390 ;
        RECT 2290.020 678.380 2293.020 678.390 ;
        RECT 2470.020 678.380 2473.020 678.390 ;
        RECT 2650.020 678.380 2653.020 678.390 ;
        RECT 2830.020 678.380 2833.020 678.390 ;
        RECT 2949.600 678.380 2952.600 678.390 ;
        RECT -32.980 675.380 2952.600 678.380 ;
        RECT -32.980 675.370 -29.980 675.380 ;
        RECT 130.020 675.370 133.020 675.380 ;
        RECT 310.020 675.370 313.020 675.380 ;
        RECT 490.020 675.370 493.020 675.380 ;
        RECT 670.020 675.370 673.020 675.380 ;
        RECT 850.020 675.370 853.020 675.380 ;
        RECT 1030.020 675.370 1033.020 675.380 ;
        RECT 1210.020 675.370 1213.020 675.380 ;
        RECT 1390.020 675.370 1393.020 675.380 ;
        RECT 1570.020 675.370 1573.020 675.380 ;
        RECT 1750.020 675.370 1753.020 675.380 ;
        RECT 1930.020 675.370 1933.020 675.380 ;
        RECT 2110.020 675.370 2113.020 675.380 ;
        RECT 2290.020 675.370 2293.020 675.380 ;
        RECT 2470.020 675.370 2473.020 675.380 ;
        RECT 2650.020 675.370 2653.020 675.380 ;
        RECT 2830.020 675.370 2833.020 675.380 ;
        RECT 2949.600 675.370 2952.600 675.380 ;
        RECT -32.980 498.380 -29.980 498.390 ;
        RECT 130.020 498.380 133.020 498.390 ;
        RECT 310.020 498.380 313.020 498.390 ;
        RECT 490.020 498.380 493.020 498.390 ;
        RECT 670.020 498.380 673.020 498.390 ;
        RECT 850.020 498.380 853.020 498.390 ;
        RECT 1030.020 498.380 1033.020 498.390 ;
        RECT 1210.020 498.380 1213.020 498.390 ;
        RECT 1390.020 498.380 1393.020 498.390 ;
        RECT 1570.020 498.380 1573.020 498.390 ;
        RECT 1750.020 498.380 1753.020 498.390 ;
        RECT 1930.020 498.380 1933.020 498.390 ;
        RECT 2110.020 498.380 2113.020 498.390 ;
        RECT 2290.020 498.380 2293.020 498.390 ;
        RECT 2470.020 498.380 2473.020 498.390 ;
        RECT 2650.020 498.380 2653.020 498.390 ;
        RECT 2830.020 498.380 2833.020 498.390 ;
        RECT 2949.600 498.380 2952.600 498.390 ;
        RECT -32.980 495.380 2952.600 498.380 ;
        RECT -32.980 495.370 -29.980 495.380 ;
        RECT 130.020 495.370 133.020 495.380 ;
        RECT 310.020 495.370 313.020 495.380 ;
        RECT 490.020 495.370 493.020 495.380 ;
        RECT 670.020 495.370 673.020 495.380 ;
        RECT 850.020 495.370 853.020 495.380 ;
        RECT 1030.020 495.370 1033.020 495.380 ;
        RECT 1210.020 495.370 1213.020 495.380 ;
        RECT 1390.020 495.370 1393.020 495.380 ;
        RECT 1570.020 495.370 1573.020 495.380 ;
        RECT 1750.020 495.370 1753.020 495.380 ;
        RECT 1930.020 495.370 1933.020 495.380 ;
        RECT 2110.020 495.370 2113.020 495.380 ;
        RECT 2290.020 495.370 2293.020 495.380 ;
        RECT 2470.020 495.370 2473.020 495.380 ;
        RECT 2650.020 495.370 2653.020 495.380 ;
        RECT 2830.020 495.370 2833.020 495.380 ;
        RECT 2949.600 495.370 2952.600 495.380 ;
        RECT -32.980 318.380 -29.980 318.390 ;
        RECT 130.020 318.380 133.020 318.390 ;
        RECT 310.020 318.380 313.020 318.390 ;
        RECT 490.020 318.380 493.020 318.390 ;
        RECT 670.020 318.380 673.020 318.390 ;
        RECT 850.020 318.380 853.020 318.390 ;
        RECT 1030.020 318.380 1033.020 318.390 ;
        RECT 1210.020 318.380 1213.020 318.390 ;
        RECT 1390.020 318.380 1393.020 318.390 ;
        RECT 1570.020 318.380 1573.020 318.390 ;
        RECT 1750.020 318.380 1753.020 318.390 ;
        RECT 1930.020 318.380 1933.020 318.390 ;
        RECT 2110.020 318.380 2113.020 318.390 ;
        RECT 2290.020 318.380 2293.020 318.390 ;
        RECT 2470.020 318.380 2473.020 318.390 ;
        RECT 2650.020 318.380 2653.020 318.390 ;
        RECT 2830.020 318.380 2833.020 318.390 ;
        RECT 2949.600 318.380 2952.600 318.390 ;
        RECT -32.980 315.380 2952.600 318.380 ;
        RECT -32.980 315.370 -29.980 315.380 ;
        RECT 130.020 315.370 133.020 315.380 ;
        RECT 310.020 315.370 313.020 315.380 ;
        RECT 490.020 315.370 493.020 315.380 ;
        RECT 670.020 315.370 673.020 315.380 ;
        RECT 850.020 315.370 853.020 315.380 ;
        RECT 1030.020 315.370 1033.020 315.380 ;
        RECT 1210.020 315.370 1213.020 315.380 ;
        RECT 1390.020 315.370 1393.020 315.380 ;
        RECT 1570.020 315.370 1573.020 315.380 ;
        RECT 1750.020 315.370 1753.020 315.380 ;
        RECT 1930.020 315.370 1933.020 315.380 ;
        RECT 2110.020 315.370 2113.020 315.380 ;
        RECT 2290.020 315.370 2293.020 315.380 ;
        RECT 2470.020 315.370 2473.020 315.380 ;
        RECT 2650.020 315.370 2653.020 315.380 ;
        RECT 2830.020 315.370 2833.020 315.380 ;
        RECT 2949.600 315.370 2952.600 315.380 ;
        RECT -32.980 138.380 -29.980 138.390 ;
        RECT 130.020 138.380 133.020 138.390 ;
        RECT 310.020 138.380 313.020 138.390 ;
        RECT 490.020 138.380 493.020 138.390 ;
        RECT 670.020 138.380 673.020 138.390 ;
        RECT 850.020 138.380 853.020 138.390 ;
        RECT 1030.020 138.380 1033.020 138.390 ;
        RECT 1210.020 138.380 1213.020 138.390 ;
        RECT 1390.020 138.380 1393.020 138.390 ;
        RECT 1570.020 138.380 1573.020 138.390 ;
        RECT 1750.020 138.380 1753.020 138.390 ;
        RECT 1930.020 138.380 1933.020 138.390 ;
        RECT 2110.020 138.380 2113.020 138.390 ;
        RECT 2290.020 138.380 2293.020 138.390 ;
        RECT 2470.020 138.380 2473.020 138.390 ;
        RECT 2650.020 138.380 2653.020 138.390 ;
        RECT 2830.020 138.380 2833.020 138.390 ;
        RECT 2949.600 138.380 2952.600 138.390 ;
        RECT -32.980 135.380 2952.600 138.380 ;
        RECT -32.980 135.370 -29.980 135.380 ;
        RECT 130.020 135.370 133.020 135.380 ;
        RECT 310.020 135.370 313.020 135.380 ;
        RECT 490.020 135.370 493.020 135.380 ;
        RECT 670.020 135.370 673.020 135.380 ;
        RECT 850.020 135.370 853.020 135.380 ;
        RECT 1030.020 135.370 1033.020 135.380 ;
        RECT 1210.020 135.370 1213.020 135.380 ;
        RECT 1390.020 135.370 1393.020 135.380 ;
        RECT 1570.020 135.370 1573.020 135.380 ;
        RECT 1750.020 135.370 1753.020 135.380 ;
        RECT 1930.020 135.370 1933.020 135.380 ;
        RECT 2110.020 135.370 2113.020 135.380 ;
        RECT 2290.020 135.370 2293.020 135.380 ;
        RECT 2470.020 135.370 2473.020 135.380 ;
        RECT 2650.020 135.370 2653.020 135.380 ;
        RECT 2830.020 135.370 2833.020 135.380 ;
        RECT 2949.600 135.370 2952.600 135.380 ;
        RECT -32.980 -24.620 -29.980 -24.610 ;
        RECT 130.020 -24.620 133.020 -24.610 ;
        RECT 310.020 -24.620 313.020 -24.610 ;
        RECT 490.020 -24.620 493.020 -24.610 ;
        RECT 670.020 -24.620 673.020 -24.610 ;
        RECT 850.020 -24.620 853.020 -24.610 ;
        RECT 1030.020 -24.620 1033.020 -24.610 ;
        RECT 1210.020 -24.620 1213.020 -24.610 ;
        RECT 1390.020 -24.620 1393.020 -24.610 ;
        RECT 1570.020 -24.620 1573.020 -24.610 ;
        RECT 1750.020 -24.620 1753.020 -24.610 ;
        RECT 1930.020 -24.620 1933.020 -24.610 ;
        RECT 2110.020 -24.620 2113.020 -24.610 ;
        RECT 2290.020 -24.620 2293.020 -24.610 ;
        RECT 2470.020 -24.620 2473.020 -24.610 ;
        RECT 2650.020 -24.620 2653.020 -24.610 ;
        RECT 2830.020 -24.620 2833.020 -24.610 ;
        RECT 2949.600 -24.620 2952.600 -24.610 ;
        RECT -32.980 -27.620 2952.600 -24.620 ;
        RECT -32.980 -27.630 -29.980 -27.620 ;
        RECT 130.020 -27.630 133.020 -27.620 ;
        RECT 310.020 -27.630 313.020 -27.620 ;
        RECT 490.020 -27.630 493.020 -27.620 ;
        RECT 670.020 -27.630 673.020 -27.620 ;
        RECT 850.020 -27.630 853.020 -27.620 ;
        RECT 1030.020 -27.630 1033.020 -27.620 ;
        RECT 1210.020 -27.630 1213.020 -27.620 ;
        RECT 1390.020 -27.630 1393.020 -27.620 ;
        RECT 1570.020 -27.630 1573.020 -27.620 ;
        RECT 1750.020 -27.630 1753.020 -27.620 ;
        RECT 1930.020 -27.630 1933.020 -27.620 ;
        RECT 2110.020 -27.630 2113.020 -27.620 ;
        RECT 2290.020 -27.630 2293.020 -27.620 ;
        RECT 2470.020 -27.630 2473.020 -27.620 ;
        RECT 2650.020 -27.630 2653.020 -27.620 ;
        RECT 2830.020 -27.630 2833.020 -27.620 ;
        RECT 2949.600 -27.630 2952.600 -27.620 ;
    END
  END vssa1
  PIN vdda2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -37.580 -32.220 -34.580 3551.900 ;
        RECT 58.020 -36.820 61.020 3556.500 ;
        RECT 238.020 -36.820 241.020 3556.500 ;
        RECT 418.020 -36.820 421.020 3556.500 ;
        RECT 598.020 -36.820 601.020 3556.500 ;
        RECT 778.020 -36.820 781.020 3556.500 ;
        RECT 958.020 -36.820 961.020 3556.500 ;
        RECT 1138.020 -36.820 1141.020 3556.500 ;
        RECT 1318.020 -36.820 1321.020 3556.500 ;
        RECT 1498.020 -36.820 1501.020 3556.500 ;
        RECT 1678.020 -36.820 1681.020 3556.500 ;
        RECT 1858.020 -36.820 1861.020 3556.500 ;
        RECT 2038.020 -36.820 2041.020 3556.500 ;
        RECT 2218.020 -36.820 2221.020 3556.500 ;
        RECT 2398.020 -36.820 2401.020 3556.500 ;
        RECT 2578.020 -36.820 2581.020 3556.500 ;
        RECT 2758.020 -36.820 2761.020 3556.500 ;
        RECT 2954.200 -32.220 2957.200 3551.900 ;
      LAYER via4 ;
        RECT -36.670 3550.610 -35.490 3551.790 ;
        RECT -36.670 3549.010 -35.490 3550.190 ;
        RECT -36.670 3485.090 -35.490 3486.270 ;
        RECT -36.670 3483.490 -35.490 3484.670 ;
        RECT -36.670 3305.090 -35.490 3306.270 ;
        RECT -36.670 3303.490 -35.490 3304.670 ;
        RECT -36.670 3125.090 -35.490 3126.270 ;
        RECT -36.670 3123.490 -35.490 3124.670 ;
        RECT -36.670 2945.090 -35.490 2946.270 ;
        RECT -36.670 2943.490 -35.490 2944.670 ;
        RECT -36.670 2765.090 -35.490 2766.270 ;
        RECT -36.670 2763.490 -35.490 2764.670 ;
        RECT -36.670 2585.090 -35.490 2586.270 ;
        RECT -36.670 2583.490 -35.490 2584.670 ;
        RECT -36.670 2405.090 -35.490 2406.270 ;
        RECT -36.670 2403.490 -35.490 2404.670 ;
        RECT -36.670 2225.090 -35.490 2226.270 ;
        RECT -36.670 2223.490 -35.490 2224.670 ;
        RECT -36.670 2045.090 -35.490 2046.270 ;
        RECT -36.670 2043.490 -35.490 2044.670 ;
        RECT -36.670 1865.090 -35.490 1866.270 ;
        RECT -36.670 1863.490 -35.490 1864.670 ;
        RECT -36.670 1685.090 -35.490 1686.270 ;
        RECT -36.670 1683.490 -35.490 1684.670 ;
        RECT -36.670 1505.090 -35.490 1506.270 ;
        RECT -36.670 1503.490 -35.490 1504.670 ;
        RECT -36.670 1325.090 -35.490 1326.270 ;
        RECT -36.670 1323.490 -35.490 1324.670 ;
        RECT -36.670 1145.090 -35.490 1146.270 ;
        RECT -36.670 1143.490 -35.490 1144.670 ;
        RECT -36.670 965.090 -35.490 966.270 ;
        RECT -36.670 963.490 -35.490 964.670 ;
        RECT -36.670 785.090 -35.490 786.270 ;
        RECT -36.670 783.490 -35.490 784.670 ;
        RECT -36.670 605.090 -35.490 606.270 ;
        RECT -36.670 603.490 -35.490 604.670 ;
        RECT -36.670 425.090 -35.490 426.270 ;
        RECT -36.670 423.490 -35.490 424.670 ;
        RECT -36.670 245.090 -35.490 246.270 ;
        RECT -36.670 243.490 -35.490 244.670 ;
        RECT -36.670 65.090 -35.490 66.270 ;
        RECT -36.670 63.490 -35.490 64.670 ;
        RECT -36.670 -30.510 -35.490 -29.330 ;
        RECT -36.670 -32.110 -35.490 -30.930 ;
        RECT 58.930 3550.610 60.110 3551.790 ;
        RECT 58.930 3549.010 60.110 3550.190 ;
        RECT 58.930 3485.090 60.110 3486.270 ;
        RECT 58.930 3483.490 60.110 3484.670 ;
        RECT 58.930 3305.090 60.110 3306.270 ;
        RECT 58.930 3303.490 60.110 3304.670 ;
        RECT 58.930 3125.090 60.110 3126.270 ;
        RECT 58.930 3123.490 60.110 3124.670 ;
        RECT 58.930 2945.090 60.110 2946.270 ;
        RECT 58.930 2943.490 60.110 2944.670 ;
        RECT 58.930 2765.090 60.110 2766.270 ;
        RECT 58.930 2763.490 60.110 2764.670 ;
        RECT 58.930 2585.090 60.110 2586.270 ;
        RECT 58.930 2583.490 60.110 2584.670 ;
        RECT 58.930 2405.090 60.110 2406.270 ;
        RECT 58.930 2403.490 60.110 2404.670 ;
        RECT 58.930 2225.090 60.110 2226.270 ;
        RECT 58.930 2223.490 60.110 2224.670 ;
        RECT 58.930 2045.090 60.110 2046.270 ;
        RECT 58.930 2043.490 60.110 2044.670 ;
        RECT 58.930 1865.090 60.110 1866.270 ;
        RECT 58.930 1863.490 60.110 1864.670 ;
        RECT 58.930 1685.090 60.110 1686.270 ;
        RECT 58.930 1683.490 60.110 1684.670 ;
        RECT 58.930 1505.090 60.110 1506.270 ;
        RECT 58.930 1503.490 60.110 1504.670 ;
        RECT 58.930 1325.090 60.110 1326.270 ;
        RECT 58.930 1323.490 60.110 1324.670 ;
        RECT 58.930 1145.090 60.110 1146.270 ;
        RECT 58.930 1143.490 60.110 1144.670 ;
        RECT 58.930 965.090 60.110 966.270 ;
        RECT 58.930 963.490 60.110 964.670 ;
        RECT 58.930 785.090 60.110 786.270 ;
        RECT 58.930 783.490 60.110 784.670 ;
        RECT 58.930 605.090 60.110 606.270 ;
        RECT 58.930 603.490 60.110 604.670 ;
        RECT 58.930 425.090 60.110 426.270 ;
        RECT 58.930 423.490 60.110 424.670 ;
        RECT 58.930 245.090 60.110 246.270 ;
        RECT 58.930 243.490 60.110 244.670 ;
        RECT 58.930 65.090 60.110 66.270 ;
        RECT 58.930 63.490 60.110 64.670 ;
        RECT 58.930 -30.510 60.110 -29.330 ;
        RECT 58.930 -32.110 60.110 -30.930 ;
        RECT 238.930 3550.610 240.110 3551.790 ;
        RECT 238.930 3549.010 240.110 3550.190 ;
        RECT 238.930 3485.090 240.110 3486.270 ;
        RECT 238.930 3483.490 240.110 3484.670 ;
        RECT 238.930 3305.090 240.110 3306.270 ;
        RECT 238.930 3303.490 240.110 3304.670 ;
        RECT 238.930 3125.090 240.110 3126.270 ;
        RECT 238.930 3123.490 240.110 3124.670 ;
        RECT 238.930 2945.090 240.110 2946.270 ;
        RECT 238.930 2943.490 240.110 2944.670 ;
        RECT 238.930 2765.090 240.110 2766.270 ;
        RECT 238.930 2763.490 240.110 2764.670 ;
        RECT 238.930 2585.090 240.110 2586.270 ;
        RECT 238.930 2583.490 240.110 2584.670 ;
        RECT 238.930 2405.090 240.110 2406.270 ;
        RECT 238.930 2403.490 240.110 2404.670 ;
        RECT 238.930 2225.090 240.110 2226.270 ;
        RECT 238.930 2223.490 240.110 2224.670 ;
        RECT 238.930 2045.090 240.110 2046.270 ;
        RECT 238.930 2043.490 240.110 2044.670 ;
        RECT 238.930 1865.090 240.110 1866.270 ;
        RECT 238.930 1863.490 240.110 1864.670 ;
        RECT 238.930 1685.090 240.110 1686.270 ;
        RECT 238.930 1683.490 240.110 1684.670 ;
        RECT 238.930 1505.090 240.110 1506.270 ;
        RECT 238.930 1503.490 240.110 1504.670 ;
        RECT 238.930 1325.090 240.110 1326.270 ;
        RECT 238.930 1323.490 240.110 1324.670 ;
        RECT 238.930 1145.090 240.110 1146.270 ;
        RECT 238.930 1143.490 240.110 1144.670 ;
        RECT 238.930 965.090 240.110 966.270 ;
        RECT 238.930 963.490 240.110 964.670 ;
        RECT 238.930 785.090 240.110 786.270 ;
        RECT 238.930 783.490 240.110 784.670 ;
        RECT 238.930 605.090 240.110 606.270 ;
        RECT 238.930 603.490 240.110 604.670 ;
        RECT 238.930 425.090 240.110 426.270 ;
        RECT 238.930 423.490 240.110 424.670 ;
        RECT 238.930 245.090 240.110 246.270 ;
        RECT 238.930 243.490 240.110 244.670 ;
        RECT 238.930 65.090 240.110 66.270 ;
        RECT 238.930 63.490 240.110 64.670 ;
        RECT 238.930 -30.510 240.110 -29.330 ;
        RECT 238.930 -32.110 240.110 -30.930 ;
        RECT 418.930 3550.610 420.110 3551.790 ;
        RECT 418.930 3549.010 420.110 3550.190 ;
        RECT 418.930 3485.090 420.110 3486.270 ;
        RECT 418.930 3483.490 420.110 3484.670 ;
        RECT 418.930 3305.090 420.110 3306.270 ;
        RECT 418.930 3303.490 420.110 3304.670 ;
        RECT 418.930 3125.090 420.110 3126.270 ;
        RECT 418.930 3123.490 420.110 3124.670 ;
        RECT 418.930 2945.090 420.110 2946.270 ;
        RECT 418.930 2943.490 420.110 2944.670 ;
        RECT 418.930 2765.090 420.110 2766.270 ;
        RECT 418.930 2763.490 420.110 2764.670 ;
        RECT 418.930 2585.090 420.110 2586.270 ;
        RECT 418.930 2583.490 420.110 2584.670 ;
        RECT 418.930 2405.090 420.110 2406.270 ;
        RECT 418.930 2403.490 420.110 2404.670 ;
        RECT 418.930 2225.090 420.110 2226.270 ;
        RECT 418.930 2223.490 420.110 2224.670 ;
        RECT 418.930 2045.090 420.110 2046.270 ;
        RECT 418.930 2043.490 420.110 2044.670 ;
        RECT 418.930 1865.090 420.110 1866.270 ;
        RECT 418.930 1863.490 420.110 1864.670 ;
        RECT 418.930 1685.090 420.110 1686.270 ;
        RECT 418.930 1683.490 420.110 1684.670 ;
        RECT 418.930 1505.090 420.110 1506.270 ;
        RECT 418.930 1503.490 420.110 1504.670 ;
        RECT 418.930 1325.090 420.110 1326.270 ;
        RECT 418.930 1323.490 420.110 1324.670 ;
        RECT 418.930 1145.090 420.110 1146.270 ;
        RECT 418.930 1143.490 420.110 1144.670 ;
        RECT 418.930 965.090 420.110 966.270 ;
        RECT 418.930 963.490 420.110 964.670 ;
        RECT 418.930 785.090 420.110 786.270 ;
        RECT 418.930 783.490 420.110 784.670 ;
        RECT 418.930 605.090 420.110 606.270 ;
        RECT 418.930 603.490 420.110 604.670 ;
        RECT 418.930 425.090 420.110 426.270 ;
        RECT 418.930 423.490 420.110 424.670 ;
        RECT 418.930 245.090 420.110 246.270 ;
        RECT 418.930 243.490 420.110 244.670 ;
        RECT 418.930 65.090 420.110 66.270 ;
        RECT 418.930 63.490 420.110 64.670 ;
        RECT 418.930 -30.510 420.110 -29.330 ;
        RECT 418.930 -32.110 420.110 -30.930 ;
        RECT 598.930 3550.610 600.110 3551.790 ;
        RECT 598.930 3549.010 600.110 3550.190 ;
        RECT 598.930 3485.090 600.110 3486.270 ;
        RECT 598.930 3483.490 600.110 3484.670 ;
        RECT 598.930 3305.090 600.110 3306.270 ;
        RECT 598.930 3303.490 600.110 3304.670 ;
        RECT 598.930 3125.090 600.110 3126.270 ;
        RECT 598.930 3123.490 600.110 3124.670 ;
        RECT 598.930 2945.090 600.110 2946.270 ;
        RECT 598.930 2943.490 600.110 2944.670 ;
        RECT 598.930 2765.090 600.110 2766.270 ;
        RECT 598.930 2763.490 600.110 2764.670 ;
        RECT 598.930 2585.090 600.110 2586.270 ;
        RECT 598.930 2583.490 600.110 2584.670 ;
        RECT 598.930 2405.090 600.110 2406.270 ;
        RECT 598.930 2403.490 600.110 2404.670 ;
        RECT 598.930 2225.090 600.110 2226.270 ;
        RECT 598.930 2223.490 600.110 2224.670 ;
        RECT 598.930 2045.090 600.110 2046.270 ;
        RECT 598.930 2043.490 600.110 2044.670 ;
        RECT 598.930 1865.090 600.110 1866.270 ;
        RECT 598.930 1863.490 600.110 1864.670 ;
        RECT 598.930 1685.090 600.110 1686.270 ;
        RECT 598.930 1683.490 600.110 1684.670 ;
        RECT 598.930 1505.090 600.110 1506.270 ;
        RECT 598.930 1503.490 600.110 1504.670 ;
        RECT 598.930 1325.090 600.110 1326.270 ;
        RECT 598.930 1323.490 600.110 1324.670 ;
        RECT 598.930 1145.090 600.110 1146.270 ;
        RECT 598.930 1143.490 600.110 1144.670 ;
        RECT 598.930 965.090 600.110 966.270 ;
        RECT 598.930 963.490 600.110 964.670 ;
        RECT 598.930 785.090 600.110 786.270 ;
        RECT 598.930 783.490 600.110 784.670 ;
        RECT 598.930 605.090 600.110 606.270 ;
        RECT 598.930 603.490 600.110 604.670 ;
        RECT 598.930 425.090 600.110 426.270 ;
        RECT 598.930 423.490 600.110 424.670 ;
        RECT 598.930 245.090 600.110 246.270 ;
        RECT 598.930 243.490 600.110 244.670 ;
        RECT 598.930 65.090 600.110 66.270 ;
        RECT 598.930 63.490 600.110 64.670 ;
        RECT 598.930 -30.510 600.110 -29.330 ;
        RECT 598.930 -32.110 600.110 -30.930 ;
        RECT 778.930 3550.610 780.110 3551.790 ;
        RECT 778.930 3549.010 780.110 3550.190 ;
        RECT 778.930 3485.090 780.110 3486.270 ;
        RECT 778.930 3483.490 780.110 3484.670 ;
        RECT 778.930 3305.090 780.110 3306.270 ;
        RECT 778.930 3303.490 780.110 3304.670 ;
        RECT 778.930 3125.090 780.110 3126.270 ;
        RECT 778.930 3123.490 780.110 3124.670 ;
        RECT 778.930 2945.090 780.110 2946.270 ;
        RECT 778.930 2943.490 780.110 2944.670 ;
        RECT 778.930 2765.090 780.110 2766.270 ;
        RECT 778.930 2763.490 780.110 2764.670 ;
        RECT 778.930 2585.090 780.110 2586.270 ;
        RECT 778.930 2583.490 780.110 2584.670 ;
        RECT 778.930 2405.090 780.110 2406.270 ;
        RECT 778.930 2403.490 780.110 2404.670 ;
        RECT 778.930 2225.090 780.110 2226.270 ;
        RECT 778.930 2223.490 780.110 2224.670 ;
        RECT 778.930 2045.090 780.110 2046.270 ;
        RECT 778.930 2043.490 780.110 2044.670 ;
        RECT 778.930 1865.090 780.110 1866.270 ;
        RECT 778.930 1863.490 780.110 1864.670 ;
        RECT 778.930 1685.090 780.110 1686.270 ;
        RECT 778.930 1683.490 780.110 1684.670 ;
        RECT 778.930 1505.090 780.110 1506.270 ;
        RECT 778.930 1503.490 780.110 1504.670 ;
        RECT 778.930 1325.090 780.110 1326.270 ;
        RECT 778.930 1323.490 780.110 1324.670 ;
        RECT 778.930 1145.090 780.110 1146.270 ;
        RECT 778.930 1143.490 780.110 1144.670 ;
        RECT 778.930 965.090 780.110 966.270 ;
        RECT 778.930 963.490 780.110 964.670 ;
        RECT 778.930 785.090 780.110 786.270 ;
        RECT 778.930 783.490 780.110 784.670 ;
        RECT 778.930 605.090 780.110 606.270 ;
        RECT 778.930 603.490 780.110 604.670 ;
        RECT 778.930 425.090 780.110 426.270 ;
        RECT 778.930 423.490 780.110 424.670 ;
        RECT 778.930 245.090 780.110 246.270 ;
        RECT 778.930 243.490 780.110 244.670 ;
        RECT 778.930 65.090 780.110 66.270 ;
        RECT 778.930 63.490 780.110 64.670 ;
        RECT 778.930 -30.510 780.110 -29.330 ;
        RECT 778.930 -32.110 780.110 -30.930 ;
        RECT 958.930 3550.610 960.110 3551.790 ;
        RECT 958.930 3549.010 960.110 3550.190 ;
        RECT 958.930 3485.090 960.110 3486.270 ;
        RECT 958.930 3483.490 960.110 3484.670 ;
        RECT 958.930 3305.090 960.110 3306.270 ;
        RECT 958.930 3303.490 960.110 3304.670 ;
        RECT 958.930 3125.090 960.110 3126.270 ;
        RECT 958.930 3123.490 960.110 3124.670 ;
        RECT 958.930 2945.090 960.110 2946.270 ;
        RECT 958.930 2943.490 960.110 2944.670 ;
        RECT 958.930 2765.090 960.110 2766.270 ;
        RECT 958.930 2763.490 960.110 2764.670 ;
        RECT 958.930 2585.090 960.110 2586.270 ;
        RECT 958.930 2583.490 960.110 2584.670 ;
        RECT 958.930 2405.090 960.110 2406.270 ;
        RECT 958.930 2403.490 960.110 2404.670 ;
        RECT 958.930 2225.090 960.110 2226.270 ;
        RECT 958.930 2223.490 960.110 2224.670 ;
        RECT 958.930 2045.090 960.110 2046.270 ;
        RECT 958.930 2043.490 960.110 2044.670 ;
        RECT 958.930 1865.090 960.110 1866.270 ;
        RECT 958.930 1863.490 960.110 1864.670 ;
        RECT 958.930 1685.090 960.110 1686.270 ;
        RECT 958.930 1683.490 960.110 1684.670 ;
        RECT 958.930 1505.090 960.110 1506.270 ;
        RECT 958.930 1503.490 960.110 1504.670 ;
        RECT 958.930 1325.090 960.110 1326.270 ;
        RECT 958.930 1323.490 960.110 1324.670 ;
        RECT 958.930 1145.090 960.110 1146.270 ;
        RECT 958.930 1143.490 960.110 1144.670 ;
        RECT 958.930 965.090 960.110 966.270 ;
        RECT 958.930 963.490 960.110 964.670 ;
        RECT 958.930 785.090 960.110 786.270 ;
        RECT 958.930 783.490 960.110 784.670 ;
        RECT 958.930 605.090 960.110 606.270 ;
        RECT 958.930 603.490 960.110 604.670 ;
        RECT 958.930 425.090 960.110 426.270 ;
        RECT 958.930 423.490 960.110 424.670 ;
        RECT 958.930 245.090 960.110 246.270 ;
        RECT 958.930 243.490 960.110 244.670 ;
        RECT 958.930 65.090 960.110 66.270 ;
        RECT 958.930 63.490 960.110 64.670 ;
        RECT 958.930 -30.510 960.110 -29.330 ;
        RECT 958.930 -32.110 960.110 -30.930 ;
        RECT 1138.930 3550.610 1140.110 3551.790 ;
        RECT 1138.930 3549.010 1140.110 3550.190 ;
        RECT 1138.930 3485.090 1140.110 3486.270 ;
        RECT 1138.930 3483.490 1140.110 3484.670 ;
        RECT 1138.930 3305.090 1140.110 3306.270 ;
        RECT 1138.930 3303.490 1140.110 3304.670 ;
        RECT 1138.930 3125.090 1140.110 3126.270 ;
        RECT 1138.930 3123.490 1140.110 3124.670 ;
        RECT 1138.930 2945.090 1140.110 2946.270 ;
        RECT 1138.930 2943.490 1140.110 2944.670 ;
        RECT 1138.930 2765.090 1140.110 2766.270 ;
        RECT 1138.930 2763.490 1140.110 2764.670 ;
        RECT 1138.930 2585.090 1140.110 2586.270 ;
        RECT 1138.930 2583.490 1140.110 2584.670 ;
        RECT 1138.930 2405.090 1140.110 2406.270 ;
        RECT 1138.930 2403.490 1140.110 2404.670 ;
        RECT 1138.930 2225.090 1140.110 2226.270 ;
        RECT 1138.930 2223.490 1140.110 2224.670 ;
        RECT 1138.930 2045.090 1140.110 2046.270 ;
        RECT 1138.930 2043.490 1140.110 2044.670 ;
        RECT 1138.930 1865.090 1140.110 1866.270 ;
        RECT 1138.930 1863.490 1140.110 1864.670 ;
        RECT 1138.930 1685.090 1140.110 1686.270 ;
        RECT 1138.930 1683.490 1140.110 1684.670 ;
        RECT 1138.930 1505.090 1140.110 1506.270 ;
        RECT 1138.930 1503.490 1140.110 1504.670 ;
        RECT 1138.930 1325.090 1140.110 1326.270 ;
        RECT 1138.930 1323.490 1140.110 1324.670 ;
        RECT 1138.930 1145.090 1140.110 1146.270 ;
        RECT 1138.930 1143.490 1140.110 1144.670 ;
        RECT 1138.930 965.090 1140.110 966.270 ;
        RECT 1138.930 963.490 1140.110 964.670 ;
        RECT 1138.930 785.090 1140.110 786.270 ;
        RECT 1138.930 783.490 1140.110 784.670 ;
        RECT 1138.930 605.090 1140.110 606.270 ;
        RECT 1138.930 603.490 1140.110 604.670 ;
        RECT 1138.930 425.090 1140.110 426.270 ;
        RECT 1138.930 423.490 1140.110 424.670 ;
        RECT 1138.930 245.090 1140.110 246.270 ;
        RECT 1138.930 243.490 1140.110 244.670 ;
        RECT 1138.930 65.090 1140.110 66.270 ;
        RECT 1138.930 63.490 1140.110 64.670 ;
        RECT 1138.930 -30.510 1140.110 -29.330 ;
        RECT 1138.930 -32.110 1140.110 -30.930 ;
        RECT 1318.930 3550.610 1320.110 3551.790 ;
        RECT 1318.930 3549.010 1320.110 3550.190 ;
        RECT 1318.930 3485.090 1320.110 3486.270 ;
        RECT 1318.930 3483.490 1320.110 3484.670 ;
        RECT 1318.930 3305.090 1320.110 3306.270 ;
        RECT 1318.930 3303.490 1320.110 3304.670 ;
        RECT 1318.930 3125.090 1320.110 3126.270 ;
        RECT 1318.930 3123.490 1320.110 3124.670 ;
        RECT 1318.930 2945.090 1320.110 2946.270 ;
        RECT 1318.930 2943.490 1320.110 2944.670 ;
        RECT 1318.930 2765.090 1320.110 2766.270 ;
        RECT 1318.930 2763.490 1320.110 2764.670 ;
        RECT 1318.930 2585.090 1320.110 2586.270 ;
        RECT 1318.930 2583.490 1320.110 2584.670 ;
        RECT 1318.930 2405.090 1320.110 2406.270 ;
        RECT 1318.930 2403.490 1320.110 2404.670 ;
        RECT 1318.930 2225.090 1320.110 2226.270 ;
        RECT 1318.930 2223.490 1320.110 2224.670 ;
        RECT 1318.930 2045.090 1320.110 2046.270 ;
        RECT 1318.930 2043.490 1320.110 2044.670 ;
        RECT 1318.930 1865.090 1320.110 1866.270 ;
        RECT 1318.930 1863.490 1320.110 1864.670 ;
        RECT 1318.930 1685.090 1320.110 1686.270 ;
        RECT 1318.930 1683.490 1320.110 1684.670 ;
        RECT 1318.930 1505.090 1320.110 1506.270 ;
        RECT 1318.930 1503.490 1320.110 1504.670 ;
        RECT 1318.930 1325.090 1320.110 1326.270 ;
        RECT 1318.930 1323.490 1320.110 1324.670 ;
        RECT 1318.930 1145.090 1320.110 1146.270 ;
        RECT 1318.930 1143.490 1320.110 1144.670 ;
        RECT 1318.930 965.090 1320.110 966.270 ;
        RECT 1318.930 963.490 1320.110 964.670 ;
        RECT 1318.930 785.090 1320.110 786.270 ;
        RECT 1318.930 783.490 1320.110 784.670 ;
        RECT 1318.930 605.090 1320.110 606.270 ;
        RECT 1318.930 603.490 1320.110 604.670 ;
        RECT 1318.930 425.090 1320.110 426.270 ;
        RECT 1318.930 423.490 1320.110 424.670 ;
        RECT 1318.930 245.090 1320.110 246.270 ;
        RECT 1318.930 243.490 1320.110 244.670 ;
        RECT 1318.930 65.090 1320.110 66.270 ;
        RECT 1318.930 63.490 1320.110 64.670 ;
        RECT 1318.930 -30.510 1320.110 -29.330 ;
        RECT 1318.930 -32.110 1320.110 -30.930 ;
        RECT 1498.930 3550.610 1500.110 3551.790 ;
        RECT 1498.930 3549.010 1500.110 3550.190 ;
        RECT 1498.930 3485.090 1500.110 3486.270 ;
        RECT 1498.930 3483.490 1500.110 3484.670 ;
        RECT 1498.930 3305.090 1500.110 3306.270 ;
        RECT 1498.930 3303.490 1500.110 3304.670 ;
        RECT 1498.930 3125.090 1500.110 3126.270 ;
        RECT 1498.930 3123.490 1500.110 3124.670 ;
        RECT 1498.930 2945.090 1500.110 2946.270 ;
        RECT 1498.930 2943.490 1500.110 2944.670 ;
        RECT 1498.930 2765.090 1500.110 2766.270 ;
        RECT 1498.930 2763.490 1500.110 2764.670 ;
        RECT 1498.930 2585.090 1500.110 2586.270 ;
        RECT 1498.930 2583.490 1500.110 2584.670 ;
        RECT 1498.930 2405.090 1500.110 2406.270 ;
        RECT 1498.930 2403.490 1500.110 2404.670 ;
        RECT 1498.930 2225.090 1500.110 2226.270 ;
        RECT 1498.930 2223.490 1500.110 2224.670 ;
        RECT 1498.930 2045.090 1500.110 2046.270 ;
        RECT 1498.930 2043.490 1500.110 2044.670 ;
        RECT 1498.930 1865.090 1500.110 1866.270 ;
        RECT 1498.930 1863.490 1500.110 1864.670 ;
        RECT 1498.930 1685.090 1500.110 1686.270 ;
        RECT 1498.930 1683.490 1500.110 1684.670 ;
        RECT 1498.930 1505.090 1500.110 1506.270 ;
        RECT 1498.930 1503.490 1500.110 1504.670 ;
        RECT 1498.930 1325.090 1500.110 1326.270 ;
        RECT 1498.930 1323.490 1500.110 1324.670 ;
        RECT 1498.930 1145.090 1500.110 1146.270 ;
        RECT 1498.930 1143.490 1500.110 1144.670 ;
        RECT 1498.930 965.090 1500.110 966.270 ;
        RECT 1498.930 963.490 1500.110 964.670 ;
        RECT 1498.930 785.090 1500.110 786.270 ;
        RECT 1498.930 783.490 1500.110 784.670 ;
        RECT 1498.930 605.090 1500.110 606.270 ;
        RECT 1498.930 603.490 1500.110 604.670 ;
        RECT 1498.930 425.090 1500.110 426.270 ;
        RECT 1498.930 423.490 1500.110 424.670 ;
        RECT 1498.930 245.090 1500.110 246.270 ;
        RECT 1498.930 243.490 1500.110 244.670 ;
        RECT 1498.930 65.090 1500.110 66.270 ;
        RECT 1498.930 63.490 1500.110 64.670 ;
        RECT 1498.930 -30.510 1500.110 -29.330 ;
        RECT 1498.930 -32.110 1500.110 -30.930 ;
        RECT 1678.930 3550.610 1680.110 3551.790 ;
        RECT 1678.930 3549.010 1680.110 3550.190 ;
        RECT 1678.930 3485.090 1680.110 3486.270 ;
        RECT 1678.930 3483.490 1680.110 3484.670 ;
        RECT 1678.930 3305.090 1680.110 3306.270 ;
        RECT 1678.930 3303.490 1680.110 3304.670 ;
        RECT 1678.930 3125.090 1680.110 3126.270 ;
        RECT 1678.930 3123.490 1680.110 3124.670 ;
        RECT 1678.930 2945.090 1680.110 2946.270 ;
        RECT 1678.930 2943.490 1680.110 2944.670 ;
        RECT 1678.930 2765.090 1680.110 2766.270 ;
        RECT 1678.930 2763.490 1680.110 2764.670 ;
        RECT 1678.930 2585.090 1680.110 2586.270 ;
        RECT 1678.930 2583.490 1680.110 2584.670 ;
        RECT 1678.930 2405.090 1680.110 2406.270 ;
        RECT 1678.930 2403.490 1680.110 2404.670 ;
        RECT 1678.930 2225.090 1680.110 2226.270 ;
        RECT 1678.930 2223.490 1680.110 2224.670 ;
        RECT 1678.930 2045.090 1680.110 2046.270 ;
        RECT 1678.930 2043.490 1680.110 2044.670 ;
        RECT 1678.930 1865.090 1680.110 1866.270 ;
        RECT 1678.930 1863.490 1680.110 1864.670 ;
        RECT 1678.930 1685.090 1680.110 1686.270 ;
        RECT 1678.930 1683.490 1680.110 1684.670 ;
        RECT 1678.930 1505.090 1680.110 1506.270 ;
        RECT 1678.930 1503.490 1680.110 1504.670 ;
        RECT 1678.930 1325.090 1680.110 1326.270 ;
        RECT 1678.930 1323.490 1680.110 1324.670 ;
        RECT 1678.930 1145.090 1680.110 1146.270 ;
        RECT 1678.930 1143.490 1680.110 1144.670 ;
        RECT 1678.930 965.090 1680.110 966.270 ;
        RECT 1678.930 963.490 1680.110 964.670 ;
        RECT 1678.930 785.090 1680.110 786.270 ;
        RECT 1678.930 783.490 1680.110 784.670 ;
        RECT 1678.930 605.090 1680.110 606.270 ;
        RECT 1678.930 603.490 1680.110 604.670 ;
        RECT 1678.930 425.090 1680.110 426.270 ;
        RECT 1678.930 423.490 1680.110 424.670 ;
        RECT 1678.930 245.090 1680.110 246.270 ;
        RECT 1678.930 243.490 1680.110 244.670 ;
        RECT 1678.930 65.090 1680.110 66.270 ;
        RECT 1678.930 63.490 1680.110 64.670 ;
        RECT 1678.930 -30.510 1680.110 -29.330 ;
        RECT 1678.930 -32.110 1680.110 -30.930 ;
        RECT 1858.930 3550.610 1860.110 3551.790 ;
        RECT 1858.930 3549.010 1860.110 3550.190 ;
        RECT 1858.930 3485.090 1860.110 3486.270 ;
        RECT 1858.930 3483.490 1860.110 3484.670 ;
        RECT 1858.930 3305.090 1860.110 3306.270 ;
        RECT 1858.930 3303.490 1860.110 3304.670 ;
        RECT 1858.930 3125.090 1860.110 3126.270 ;
        RECT 1858.930 3123.490 1860.110 3124.670 ;
        RECT 1858.930 2945.090 1860.110 2946.270 ;
        RECT 1858.930 2943.490 1860.110 2944.670 ;
        RECT 1858.930 2765.090 1860.110 2766.270 ;
        RECT 1858.930 2763.490 1860.110 2764.670 ;
        RECT 1858.930 2585.090 1860.110 2586.270 ;
        RECT 1858.930 2583.490 1860.110 2584.670 ;
        RECT 1858.930 2405.090 1860.110 2406.270 ;
        RECT 1858.930 2403.490 1860.110 2404.670 ;
        RECT 1858.930 2225.090 1860.110 2226.270 ;
        RECT 1858.930 2223.490 1860.110 2224.670 ;
        RECT 1858.930 2045.090 1860.110 2046.270 ;
        RECT 1858.930 2043.490 1860.110 2044.670 ;
        RECT 1858.930 1865.090 1860.110 1866.270 ;
        RECT 1858.930 1863.490 1860.110 1864.670 ;
        RECT 1858.930 1685.090 1860.110 1686.270 ;
        RECT 1858.930 1683.490 1860.110 1684.670 ;
        RECT 1858.930 1505.090 1860.110 1506.270 ;
        RECT 1858.930 1503.490 1860.110 1504.670 ;
        RECT 1858.930 1325.090 1860.110 1326.270 ;
        RECT 1858.930 1323.490 1860.110 1324.670 ;
        RECT 1858.930 1145.090 1860.110 1146.270 ;
        RECT 1858.930 1143.490 1860.110 1144.670 ;
        RECT 1858.930 965.090 1860.110 966.270 ;
        RECT 1858.930 963.490 1860.110 964.670 ;
        RECT 1858.930 785.090 1860.110 786.270 ;
        RECT 1858.930 783.490 1860.110 784.670 ;
        RECT 1858.930 605.090 1860.110 606.270 ;
        RECT 1858.930 603.490 1860.110 604.670 ;
        RECT 1858.930 425.090 1860.110 426.270 ;
        RECT 1858.930 423.490 1860.110 424.670 ;
        RECT 1858.930 245.090 1860.110 246.270 ;
        RECT 1858.930 243.490 1860.110 244.670 ;
        RECT 1858.930 65.090 1860.110 66.270 ;
        RECT 1858.930 63.490 1860.110 64.670 ;
        RECT 1858.930 -30.510 1860.110 -29.330 ;
        RECT 1858.930 -32.110 1860.110 -30.930 ;
        RECT 2038.930 3550.610 2040.110 3551.790 ;
        RECT 2038.930 3549.010 2040.110 3550.190 ;
        RECT 2038.930 3485.090 2040.110 3486.270 ;
        RECT 2038.930 3483.490 2040.110 3484.670 ;
        RECT 2038.930 3305.090 2040.110 3306.270 ;
        RECT 2038.930 3303.490 2040.110 3304.670 ;
        RECT 2038.930 3125.090 2040.110 3126.270 ;
        RECT 2038.930 3123.490 2040.110 3124.670 ;
        RECT 2038.930 2945.090 2040.110 2946.270 ;
        RECT 2038.930 2943.490 2040.110 2944.670 ;
        RECT 2038.930 2765.090 2040.110 2766.270 ;
        RECT 2038.930 2763.490 2040.110 2764.670 ;
        RECT 2038.930 2585.090 2040.110 2586.270 ;
        RECT 2038.930 2583.490 2040.110 2584.670 ;
        RECT 2038.930 2405.090 2040.110 2406.270 ;
        RECT 2038.930 2403.490 2040.110 2404.670 ;
        RECT 2038.930 2225.090 2040.110 2226.270 ;
        RECT 2038.930 2223.490 2040.110 2224.670 ;
        RECT 2038.930 2045.090 2040.110 2046.270 ;
        RECT 2038.930 2043.490 2040.110 2044.670 ;
        RECT 2038.930 1865.090 2040.110 1866.270 ;
        RECT 2038.930 1863.490 2040.110 1864.670 ;
        RECT 2038.930 1685.090 2040.110 1686.270 ;
        RECT 2038.930 1683.490 2040.110 1684.670 ;
        RECT 2038.930 1505.090 2040.110 1506.270 ;
        RECT 2038.930 1503.490 2040.110 1504.670 ;
        RECT 2038.930 1325.090 2040.110 1326.270 ;
        RECT 2038.930 1323.490 2040.110 1324.670 ;
        RECT 2038.930 1145.090 2040.110 1146.270 ;
        RECT 2038.930 1143.490 2040.110 1144.670 ;
        RECT 2038.930 965.090 2040.110 966.270 ;
        RECT 2038.930 963.490 2040.110 964.670 ;
        RECT 2038.930 785.090 2040.110 786.270 ;
        RECT 2038.930 783.490 2040.110 784.670 ;
        RECT 2038.930 605.090 2040.110 606.270 ;
        RECT 2038.930 603.490 2040.110 604.670 ;
        RECT 2038.930 425.090 2040.110 426.270 ;
        RECT 2038.930 423.490 2040.110 424.670 ;
        RECT 2038.930 245.090 2040.110 246.270 ;
        RECT 2038.930 243.490 2040.110 244.670 ;
        RECT 2038.930 65.090 2040.110 66.270 ;
        RECT 2038.930 63.490 2040.110 64.670 ;
        RECT 2038.930 -30.510 2040.110 -29.330 ;
        RECT 2038.930 -32.110 2040.110 -30.930 ;
        RECT 2218.930 3550.610 2220.110 3551.790 ;
        RECT 2218.930 3549.010 2220.110 3550.190 ;
        RECT 2218.930 3485.090 2220.110 3486.270 ;
        RECT 2218.930 3483.490 2220.110 3484.670 ;
        RECT 2218.930 3305.090 2220.110 3306.270 ;
        RECT 2218.930 3303.490 2220.110 3304.670 ;
        RECT 2218.930 3125.090 2220.110 3126.270 ;
        RECT 2218.930 3123.490 2220.110 3124.670 ;
        RECT 2218.930 2945.090 2220.110 2946.270 ;
        RECT 2218.930 2943.490 2220.110 2944.670 ;
        RECT 2218.930 2765.090 2220.110 2766.270 ;
        RECT 2218.930 2763.490 2220.110 2764.670 ;
        RECT 2218.930 2585.090 2220.110 2586.270 ;
        RECT 2218.930 2583.490 2220.110 2584.670 ;
        RECT 2218.930 2405.090 2220.110 2406.270 ;
        RECT 2218.930 2403.490 2220.110 2404.670 ;
        RECT 2218.930 2225.090 2220.110 2226.270 ;
        RECT 2218.930 2223.490 2220.110 2224.670 ;
        RECT 2218.930 2045.090 2220.110 2046.270 ;
        RECT 2218.930 2043.490 2220.110 2044.670 ;
        RECT 2218.930 1865.090 2220.110 1866.270 ;
        RECT 2218.930 1863.490 2220.110 1864.670 ;
        RECT 2218.930 1685.090 2220.110 1686.270 ;
        RECT 2218.930 1683.490 2220.110 1684.670 ;
        RECT 2218.930 1505.090 2220.110 1506.270 ;
        RECT 2218.930 1503.490 2220.110 1504.670 ;
        RECT 2218.930 1325.090 2220.110 1326.270 ;
        RECT 2218.930 1323.490 2220.110 1324.670 ;
        RECT 2218.930 1145.090 2220.110 1146.270 ;
        RECT 2218.930 1143.490 2220.110 1144.670 ;
        RECT 2218.930 965.090 2220.110 966.270 ;
        RECT 2218.930 963.490 2220.110 964.670 ;
        RECT 2218.930 785.090 2220.110 786.270 ;
        RECT 2218.930 783.490 2220.110 784.670 ;
        RECT 2218.930 605.090 2220.110 606.270 ;
        RECT 2218.930 603.490 2220.110 604.670 ;
        RECT 2218.930 425.090 2220.110 426.270 ;
        RECT 2218.930 423.490 2220.110 424.670 ;
        RECT 2218.930 245.090 2220.110 246.270 ;
        RECT 2218.930 243.490 2220.110 244.670 ;
        RECT 2218.930 65.090 2220.110 66.270 ;
        RECT 2218.930 63.490 2220.110 64.670 ;
        RECT 2218.930 -30.510 2220.110 -29.330 ;
        RECT 2218.930 -32.110 2220.110 -30.930 ;
        RECT 2398.930 3550.610 2400.110 3551.790 ;
        RECT 2398.930 3549.010 2400.110 3550.190 ;
        RECT 2398.930 3485.090 2400.110 3486.270 ;
        RECT 2398.930 3483.490 2400.110 3484.670 ;
        RECT 2398.930 3305.090 2400.110 3306.270 ;
        RECT 2398.930 3303.490 2400.110 3304.670 ;
        RECT 2398.930 3125.090 2400.110 3126.270 ;
        RECT 2398.930 3123.490 2400.110 3124.670 ;
        RECT 2398.930 2945.090 2400.110 2946.270 ;
        RECT 2398.930 2943.490 2400.110 2944.670 ;
        RECT 2398.930 2765.090 2400.110 2766.270 ;
        RECT 2398.930 2763.490 2400.110 2764.670 ;
        RECT 2398.930 2585.090 2400.110 2586.270 ;
        RECT 2398.930 2583.490 2400.110 2584.670 ;
        RECT 2398.930 2405.090 2400.110 2406.270 ;
        RECT 2398.930 2403.490 2400.110 2404.670 ;
        RECT 2398.930 2225.090 2400.110 2226.270 ;
        RECT 2398.930 2223.490 2400.110 2224.670 ;
        RECT 2398.930 2045.090 2400.110 2046.270 ;
        RECT 2398.930 2043.490 2400.110 2044.670 ;
        RECT 2398.930 1865.090 2400.110 1866.270 ;
        RECT 2398.930 1863.490 2400.110 1864.670 ;
        RECT 2398.930 1685.090 2400.110 1686.270 ;
        RECT 2398.930 1683.490 2400.110 1684.670 ;
        RECT 2398.930 1505.090 2400.110 1506.270 ;
        RECT 2398.930 1503.490 2400.110 1504.670 ;
        RECT 2398.930 1325.090 2400.110 1326.270 ;
        RECT 2398.930 1323.490 2400.110 1324.670 ;
        RECT 2398.930 1145.090 2400.110 1146.270 ;
        RECT 2398.930 1143.490 2400.110 1144.670 ;
        RECT 2398.930 965.090 2400.110 966.270 ;
        RECT 2398.930 963.490 2400.110 964.670 ;
        RECT 2398.930 785.090 2400.110 786.270 ;
        RECT 2398.930 783.490 2400.110 784.670 ;
        RECT 2398.930 605.090 2400.110 606.270 ;
        RECT 2398.930 603.490 2400.110 604.670 ;
        RECT 2398.930 425.090 2400.110 426.270 ;
        RECT 2398.930 423.490 2400.110 424.670 ;
        RECT 2398.930 245.090 2400.110 246.270 ;
        RECT 2398.930 243.490 2400.110 244.670 ;
        RECT 2398.930 65.090 2400.110 66.270 ;
        RECT 2398.930 63.490 2400.110 64.670 ;
        RECT 2398.930 -30.510 2400.110 -29.330 ;
        RECT 2398.930 -32.110 2400.110 -30.930 ;
        RECT 2578.930 3550.610 2580.110 3551.790 ;
        RECT 2578.930 3549.010 2580.110 3550.190 ;
        RECT 2578.930 3485.090 2580.110 3486.270 ;
        RECT 2578.930 3483.490 2580.110 3484.670 ;
        RECT 2578.930 3305.090 2580.110 3306.270 ;
        RECT 2578.930 3303.490 2580.110 3304.670 ;
        RECT 2578.930 3125.090 2580.110 3126.270 ;
        RECT 2578.930 3123.490 2580.110 3124.670 ;
        RECT 2578.930 2945.090 2580.110 2946.270 ;
        RECT 2578.930 2943.490 2580.110 2944.670 ;
        RECT 2578.930 2765.090 2580.110 2766.270 ;
        RECT 2578.930 2763.490 2580.110 2764.670 ;
        RECT 2578.930 2585.090 2580.110 2586.270 ;
        RECT 2578.930 2583.490 2580.110 2584.670 ;
        RECT 2578.930 2405.090 2580.110 2406.270 ;
        RECT 2578.930 2403.490 2580.110 2404.670 ;
        RECT 2578.930 2225.090 2580.110 2226.270 ;
        RECT 2578.930 2223.490 2580.110 2224.670 ;
        RECT 2578.930 2045.090 2580.110 2046.270 ;
        RECT 2578.930 2043.490 2580.110 2044.670 ;
        RECT 2578.930 1865.090 2580.110 1866.270 ;
        RECT 2578.930 1863.490 2580.110 1864.670 ;
        RECT 2578.930 1685.090 2580.110 1686.270 ;
        RECT 2578.930 1683.490 2580.110 1684.670 ;
        RECT 2578.930 1505.090 2580.110 1506.270 ;
        RECT 2578.930 1503.490 2580.110 1504.670 ;
        RECT 2578.930 1325.090 2580.110 1326.270 ;
        RECT 2578.930 1323.490 2580.110 1324.670 ;
        RECT 2578.930 1145.090 2580.110 1146.270 ;
        RECT 2578.930 1143.490 2580.110 1144.670 ;
        RECT 2578.930 965.090 2580.110 966.270 ;
        RECT 2578.930 963.490 2580.110 964.670 ;
        RECT 2578.930 785.090 2580.110 786.270 ;
        RECT 2578.930 783.490 2580.110 784.670 ;
        RECT 2578.930 605.090 2580.110 606.270 ;
        RECT 2578.930 603.490 2580.110 604.670 ;
        RECT 2578.930 425.090 2580.110 426.270 ;
        RECT 2578.930 423.490 2580.110 424.670 ;
        RECT 2578.930 245.090 2580.110 246.270 ;
        RECT 2578.930 243.490 2580.110 244.670 ;
        RECT 2578.930 65.090 2580.110 66.270 ;
        RECT 2578.930 63.490 2580.110 64.670 ;
        RECT 2578.930 -30.510 2580.110 -29.330 ;
        RECT 2578.930 -32.110 2580.110 -30.930 ;
        RECT 2758.930 3550.610 2760.110 3551.790 ;
        RECT 2758.930 3549.010 2760.110 3550.190 ;
        RECT 2758.930 3485.090 2760.110 3486.270 ;
        RECT 2758.930 3483.490 2760.110 3484.670 ;
        RECT 2758.930 3305.090 2760.110 3306.270 ;
        RECT 2758.930 3303.490 2760.110 3304.670 ;
        RECT 2758.930 3125.090 2760.110 3126.270 ;
        RECT 2758.930 3123.490 2760.110 3124.670 ;
        RECT 2758.930 2945.090 2760.110 2946.270 ;
        RECT 2758.930 2943.490 2760.110 2944.670 ;
        RECT 2758.930 2765.090 2760.110 2766.270 ;
        RECT 2758.930 2763.490 2760.110 2764.670 ;
        RECT 2758.930 2585.090 2760.110 2586.270 ;
        RECT 2758.930 2583.490 2760.110 2584.670 ;
        RECT 2758.930 2405.090 2760.110 2406.270 ;
        RECT 2758.930 2403.490 2760.110 2404.670 ;
        RECT 2758.930 2225.090 2760.110 2226.270 ;
        RECT 2758.930 2223.490 2760.110 2224.670 ;
        RECT 2758.930 2045.090 2760.110 2046.270 ;
        RECT 2758.930 2043.490 2760.110 2044.670 ;
        RECT 2758.930 1865.090 2760.110 1866.270 ;
        RECT 2758.930 1863.490 2760.110 1864.670 ;
        RECT 2758.930 1685.090 2760.110 1686.270 ;
        RECT 2758.930 1683.490 2760.110 1684.670 ;
        RECT 2758.930 1505.090 2760.110 1506.270 ;
        RECT 2758.930 1503.490 2760.110 1504.670 ;
        RECT 2758.930 1325.090 2760.110 1326.270 ;
        RECT 2758.930 1323.490 2760.110 1324.670 ;
        RECT 2758.930 1145.090 2760.110 1146.270 ;
        RECT 2758.930 1143.490 2760.110 1144.670 ;
        RECT 2758.930 965.090 2760.110 966.270 ;
        RECT 2758.930 963.490 2760.110 964.670 ;
        RECT 2758.930 785.090 2760.110 786.270 ;
        RECT 2758.930 783.490 2760.110 784.670 ;
        RECT 2758.930 605.090 2760.110 606.270 ;
        RECT 2758.930 603.490 2760.110 604.670 ;
        RECT 2758.930 425.090 2760.110 426.270 ;
        RECT 2758.930 423.490 2760.110 424.670 ;
        RECT 2758.930 245.090 2760.110 246.270 ;
        RECT 2758.930 243.490 2760.110 244.670 ;
        RECT 2758.930 65.090 2760.110 66.270 ;
        RECT 2758.930 63.490 2760.110 64.670 ;
        RECT 2758.930 -30.510 2760.110 -29.330 ;
        RECT 2758.930 -32.110 2760.110 -30.930 ;
        RECT 2955.110 3550.610 2956.290 3551.790 ;
        RECT 2955.110 3549.010 2956.290 3550.190 ;
        RECT 2955.110 3485.090 2956.290 3486.270 ;
        RECT 2955.110 3483.490 2956.290 3484.670 ;
        RECT 2955.110 3305.090 2956.290 3306.270 ;
        RECT 2955.110 3303.490 2956.290 3304.670 ;
        RECT 2955.110 3125.090 2956.290 3126.270 ;
        RECT 2955.110 3123.490 2956.290 3124.670 ;
        RECT 2955.110 2945.090 2956.290 2946.270 ;
        RECT 2955.110 2943.490 2956.290 2944.670 ;
        RECT 2955.110 2765.090 2956.290 2766.270 ;
        RECT 2955.110 2763.490 2956.290 2764.670 ;
        RECT 2955.110 2585.090 2956.290 2586.270 ;
        RECT 2955.110 2583.490 2956.290 2584.670 ;
        RECT 2955.110 2405.090 2956.290 2406.270 ;
        RECT 2955.110 2403.490 2956.290 2404.670 ;
        RECT 2955.110 2225.090 2956.290 2226.270 ;
        RECT 2955.110 2223.490 2956.290 2224.670 ;
        RECT 2955.110 2045.090 2956.290 2046.270 ;
        RECT 2955.110 2043.490 2956.290 2044.670 ;
        RECT 2955.110 1865.090 2956.290 1866.270 ;
        RECT 2955.110 1863.490 2956.290 1864.670 ;
        RECT 2955.110 1685.090 2956.290 1686.270 ;
        RECT 2955.110 1683.490 2956.290 1684.670 ;
        RECT 2955.110 1505.090 2956.290 1506.270 ;
        RECT 2955.110 1503.490 2956.290 1504.670 ;
        RECT 2955.110 1325.090 2956.290 1326.270 ;
        RECT 2955.110 1323.490 2956.290 1324.670 ;
        RECT 2955.110 1145.090 2956.290 1146.270 ;
        RECT 2955.110 1143.490 2956.290 1144.670 ;
        RECT 2955.110 965.090 2956.290 966.270 ;
        RECT 2955.110 963.490 2956.290 964.670 ;
        RECT 2955.110 785.090 2956.290 786.270 ;
        RECT 2955.110 783.490 2956.290 784.670 ;
        RECT 2955.110 605.090 2956.290 606.270 ;
        RECT 2955.110 603.490 2956.290 604.670 ;
        RECT 2955.110 425.090 2956.290 426.270 ;
        RECT 2955.110 423.490 2956.290 424.670 ;
        RECT 2955.110 245.090 2956.290 246.270 ;
        RECT 2955.110 243.490 2956.290 244.670 ;
        RECT 2955.110 65.090 2956.290 66.270 ;
        RECT 2955.110 63.490 2956.290 64.670 ;
        RECT 2955.110 -30.510 2956.290 -29.330 ;
        RECT 2955.110 -32.110 2956.290 -30.930 ;
      LAYER met5 ;
        RECT -37.580 3551.900 -34.580 3551.910 ;
        RECT 58.020 3551.900 61.020 3551.910 ;
        RECT 238.020 3551.900 241.020 3551.910 ;
        RECT 418.020 3551.900 421.020 3551.910 ;
        RECT 598.020 3551.900 601.020 3551.910 ;
        RECT 778.020 3551.900 781.020 3551.910 ;
        RECT 958.020 3551.900 961.020 3551.910 ;
        RECT 1138.020 3551.900 1141.020 3551.910 ;
        RECT 1318.020 3551.900 1321.020 3551.910 ;
        RECT 1498.020 3551.900 1501.020 3551.910 ;
        RECT 1678.020 3551.900 1681.020 3551.910 ;
        RECT 1858.020 3551.900 1861.020 3551.910 ;
        RECT 2038.020 3551.900 2041.020 3551.910 ;
        RECT 2218.020 3551.900 2221.020 3551.910 ;
        RECT 2398.020 3551.900 2401.020 3551.910 ;
        RECT 2578.020 3551.900 2581.020 3551.910 ;
        RECT 2758.020 3551.900 2761.020 3551.910 ;
        RECT 2954.200 3551.900 2957.200 3551.910 ;
        RECT -37.580 3548.900 2957.200 3551.900 ;
        RECT -37.580 3548.890 -34.580 3548.900 ;
        RECT 58.020 3548.890 61.020 3548.900 ;
        RECT 238.020 3548.890 241.020 3548.900 ;
        RECT 418.020 3548.890 421.020 3548.900 ;
        RECT 598.020 3548.890 601.020 3548.900 ;
        RECT 778.020 3548.890 781.020 3548.900 ;
        RECT 958.020 3548.890 961.020 3548.900 ;
        RECT 1138.020 3548.890 1141.020 3548.900 ;
        RECT 1318.020 3548.890 1321.020 3548.900 ;
        RECT 1498.020 3548.890 1501.020 3548.900 ;
        RECT 1678.020 3548.890 1681.020 3548.900 ;
        RECT 1858.020 3548.890 1861.020 3548.900 ;
        RECT 2038.020 3548.890 2041.020 3548.900 ;
        RECT 2218.020 3548.890 2221.020 3548.900 ;
        RECT 2398.020 3548.890 2401.020 3548.900 ;
        RECT 2578.020 3548.890 2581.020 3548.900 ;
        RECT 2758.020 3548.890 2761.020 3548.900 ;
        RECT 2954.200 3548.890 2957.200 3548.900 ;
        RECT -37.580 3486.380 -34.580 3486.390 ;
        RECT 58.020 3486.380 61.020 3486.390 ;
        RECT 238.020 3486.380 241.020 3486.390 ;
        RECT 418.020 3486.380 421.020 3486.390 ;
        RECT 598.020 3486.380 601.020 3486.390 ;
        RECT 778.020 3486.380 781.020 3486.390 ;
        RECT 958.020 3486.380 961.020 3486.390 ;
        RECT 1138.020 3486.380 1141.020 3486.390 ;
        RECT 1318.020 3486.380 1321.020 3486.390 ;
        RECT 1498.020 3486.380 1501.020 3486.390 ;
        RECT 1678.020 3486.380 1681.020 3486.390 ;
        RECT 1858.020 3486.380 1861.020 3486.390 ;
        RECT 2038.020 3486.380 2041.020 3486.390 ;
        RECT 2218.020 3486.380 2221.020 3486.390 ;
        RECT 2398.020 3486.380 2401.020 3486.390 ;
        RECT 2578.020 3486.380 2581.020 3486.390 ;
        RECT 2758.020 3486.380 2761.020 3486.390 ;
        RECT 2954.200 3486.380 2957.200 3486.390 ;
        RECT -42.180 3483.380 2961.800 3486.380 ;
        RECT -37.580 3483.370 -34.580 3483.380 ;
        RECT 58.020 3483.370 61.020 3483.380 ;
        RECT 238.020 3483.370 241.020 3483.380 ;
        RECT 418.020 3483.370 421.020 3483.380 ;
        RECT 598.020 3483.370 601.020 3483.380 ;
        RECT 778.020 3483.370 781.020 3483.380 ;
        RECT 958.020 3483.370 961.020 3483.380 ;
        RECT 1138.020 3483.370 1141.020 3483.380 ;
        RECT 1318.020 3483.370 1321.020 3483.380 ;
        RECT 1498.020 3483.370 1501.020 3483.380 ;
        RECT 1678.020 3483.370 1681.020 3483.380 ;
        RECT 1858.020 3483.370 1861.020 3483.380 ;
        RECT 2038.020 3483.370 2041.020 3483.380 ;
        RECT 2218.020 3483.370 2221.020 3483.380 ;
        RECT 2398.020 3483.370 2401.020 3483.380 ;
        RECT 2578.020 3483.370 2581.020 3483.380 ;
        RECT 2758.020 3483.370 2761.020 3483.380 ;
        RECT 2954.200 3483.370 2957.200 3483.380 ;
        RECT -37.580 3306.380 -34.580 3306.390 ;
        RECT 58.020 3306.380 61.020 3306.390 ;
        RECT 238.020 3306.380 241.020 3306.390 ;
        RECT 418.020 3306.380 421.020 3306.390 ;
        RECT 598.020 3306.380 601.020 3306.390 ;
        RECT 778.020 3306.380 781.020 3306.390 ;
        RECT 958.020 3306.380 961.020 3306.390 ;
        RECT 1138.020 3306.380 1141.020 3306.390 ;
        RECT 1318.020 3306.380 1321.020 3306.390 ;
        RECT 1498.020 3306.380 1501.020 3306.390 ;
        RECT 1678.020 3306.380 1681.020 3306.390 ;
        RECT 1858.020 3306.380 1861.020 3306.390 ;
        RECT 2038.020 3306.380 2041.020 3306.390 ;
        RECT 2218.020 3306.380 2221.020 3306.390 ;
        RECT 2398.020 3306.380 2401.020 3306.390 ;
        RECT 2578.020 3306.380 2581.020 3306.390 ;
        RECT 2758.020 3306.380 2761.020 3306.390 ;
        RECT 2954.200 3306.380 2957.200 3306.390 ;
        RECT -42.180 3303.380 2961.800 3306.380 ;
        RECT -37.580 3303.370 -34.580 3303.380 ;
        RECT 58.020 3303.370 61.020 3303.380 ;
        RECT 238.020 3303.370 241.020 3303.380 ;
        RECT 418.020 3303.370 421.020 3303.380 ;
        RECT 598.020 3303.370 601.020 3303.380 ;
        RECT 778.020 3303.370 781.020 3303.380 ;
        RECT 958.020 3303.370 961.020 3303.380 ;
        RECT 1138.020 3303.370 1141.020 3303.380 ;
        RECT 1318.020 3303.370 1321.020 3303.380 ;
        RECT 1498.020 3303.370 1501.020 3303.380 ;
        RECT 1678.020 3303.370 1681.020 3303.380 ;
        RECT 1858.020 3303.370 1861.020 3303.380 ;
        RECT 2038.020 3303.370 2041.020 3303.380 ;
        RECT 2218.020 3303.370 2221.020 3303.380 ;
        RECT 2398.020 3303.370 2401.020 3303.380 ;
        RECT 2578.020 3303.370 2581.020 3303.380 ;
        RECT 2758.020 3303.370 2761.020 3303.380 ;
        RECT 2954.200 3303.370 2957.200 3303.380 ;
        RECT -37.580 3126.380 -34.580 3126.390 ;
        RECT 58.020 3126.380 61.020 3126.390 ;
        RECT 238.020 3126.380 241.020 3126.390 ;
        RECT 418.020 3126.380 421.020 3126.390 ;
        RECT 598.020 3126.380 601.020 3126.390 ;
        RECT 778.020 3126.380 781.020 3126.390 ;
        RECT 958.020 3126.380 961.020 3126.390 ;
        RECT 1138.020 3126.380 1141.020 3126.390 ;
        RECT 1318.020 3126.380 1321.020 3126.390 ;
        RECT 1498.020 3126.380 1501.020 3126.390 ;
        RECT 1678.020 3126.380 1681.020 3126.390 ;
        RECT 1858.020 3126.380 1861.020 3126.390 ;
        RECT 2038.020 3126.380 2041.020 3126.390 ;
        RECT 2218.020 3126.380 2221.020 3126.390 ;
        RECT 2398.020 3126.380 2401.020 3126.390 ;
        RECT 2578.020 3126.380 2581.020 3126.390 ;
        RECT 2758.020 3126.380 2761.020 3126.390 ;
        RECT 2954.200 3126.380 2957.200 3126.390 ;
        RECT -42.180 3123.380 2961.800 3126.380 ;
        RECT -37.580 3123.370 -34.580 3123.380 ;
        RECT 58.020 3123.370 61.020 3123.380 ;
        RECT 238.020 3123.370 241.020 3123.380 ;
        RECT 418.020 3123.370 421.020 3123.380 ;
        RECT 598.020 3123.370 601.020 3123.380 ;
        RECT 778.020 3123.370 781.020 3123.380 ;
        RECT 958.020 3123.370 961.020 3123.380 ;
        RECT 1138.020 3123.370 1141.020 3123.380 ;
        RECT 1318.020 3123.370 1321.020 3123.380 ;
        RECT 1498.020 3123.370 1501.020 3123.380 ;
        RECT 1678.020 3123.370 1681.020 3123.380 ;
        RECT 1858.020 3123.370 1861.020 3123.380 ;
        RECT 2038.020 3123.370 2041.020 3123.380 ;
        RECT 2218.020 3123.370 2221.020 3123.380 ;
        RECT 2398.020 3123.370 2401.020 3123.380 ;
        RECT 2578.020 3123.370 2581.020 3123.380 ;
        RECT 2758.020 3123.370 2761.020 3123.380 ;
        RECT 2954.200 3123.370 2957.200 3123.380 ;
        RECT -37.580 2946.380 -34.580 2946.390 ;
        RECT 58.020 2946.380 61.020 2946.390 ;
        RECT 238.020 2946.380 241.020 2946.390 ;
        RECT 418.020 2946.380 421.020 2946.390 ;
        RECT 598.020 2946.380 601.020 2946.390 ;
        RECT 778.020 2946.380 781.020 2946.390 ;
        RECT 958.020 2946.380 961.020 2946.390 ;
        RECT 1138.020 2946.380 1141.020 2946.390 ;
        RECT 1318.020 2946.380 1321.020 2946.390 ;
        RECT 1498.020 2946.380 1501.020 2946.390 ;
        RECT 1678.020 2946.380 1681.020 2946.390 ;
        RECT 1858.020 2946.380 1861.020 2946.390 ;
        RECT 2038.020 2946.380 2041.020 2946.390 ;
        RECT 2218.020 2946.380 2221.020 2946.390 ;
        RECT 2398.020 2946.380 2401.020 2946.390 ;
        RECT 2578.020 2946.380 2581.020 2946.390 ;
        RECT 2758.020 2946.380 2761.020 2946.390 ;
        RECT 2954.200 2946.380 2957.200 2946.390 ;
        RECT -42.180 2943.380 2961.800 2946.380 ;
        RECT -37.580 2943.370 -34.580 2943.380 ;
        RECT 58.020 2943.370 61.020 2943.380 ;
        RECT 238.020 2943.370 241.020 2943.380 ;
        RECT 418.020 2943.370 421.020 2943.380 ;
        RECT 598.020 2943.370 601.020 2943.380 ;
        RECT 778.020 2943.370 781.020 2943.380 ;
        RECT 958.020 2943.370 961.020 2943.380 ;
        RECT 1138.020 2943.370 1141.020 2943.380 ;
        RECT 1318.020 2943.370 1321.020 2943.380 ;
        RECT 1498.020 2943.370 1501.020 2943.380 ;
        RECT 1678.020 2943.370 1681.020 2943.380 ;
        RECT 1858.020 2943.370 1861.020 2943.380 ;
        RECT 2038.020 2943.370 2041.020 2943.380 ;
        RECT 2218.020 2943.370 2221.020 2943.380 ;
        RECT 2398.020 2943.370 2401.020 2943.380 ;
        RECT 2578.020 2943.370 2581.020 2943.380 ;
        RECT 2758.020 2943.370 2761.020 2943.380 ;
        RECT 2954.200 2943.370 2957.200 2943.380 ;
        RECT -37.580 2766.380 -34.580 2766.390 ;
        RECT 58.020 2766.380 61.020 2766.390 ;
        RECT 238.020 2766.380 241.020 2766.390 ;
        RECT 418.020 2766.380 421.020 2766.390 ;
        RECT 598.020 2766.380 601.020 2766.390 ;
        RECT 778.020 2766.380 781.020 2766.390 ;
        RECT 958.020 2766.380 961.020 2766.390 ;
        RECT 1138.020 2766.380 1141.020 2766.390 ;
        RECT 1318.020 2766.380 1321.020 2766.390 ;
        RECT 1498.020 2766.380 1501.020 2766.390 ;
        RECT 1678.020 2766.380 1681.020 2766.390 ;
        RECT 1858.020 2766.380 1861.020 2766.390 ;
        RECT 2038.020 2766.380 2041.020 2766.390 ;
        RECT 2218.020 2766.380 2221.020 2766.390 ;
        RECT 2398.020 2766.380 2401.020 2766.390 ;
        RECT 2578.020 2766.380 2581.020 2766.390 ;
        RECT 2758.020 2766.380 2761.020 2766.390 ;
        RECT 2954.200 2766.380 2957.200 2766.390 ;
        RECT -42.180 2763.380 2961.800 2766.380 ;
        RECT -37.580 2763.370 -34.580 2763.380 ;
        RECT 58.020 2763.370 61.020 2763.380 ;
        RECT 238.020 2763.370 241.020 2763.380 ;
        RECT 418.020 2763.370 421.020 2763.380 ;
        RECT 598.020 2763.370 601.020 2763.380 ;
        RECT 778.020 2763.370 781.020 2763.380 ;
        RECT 958.020 2763.370 961.020 2763.380 ;
        RECT 1138.020 2763.370 1141.020 2763.380 ;
        RECT 1318.020 2763.370 1321.020 2763.380 ;
        RECT 1498.020 2763.370 1501.020 2763.380 ;
        RECT 1678.020 2763.370 1681.020 2763.380 ;
        RECT 1858.020 2763.370 1861.020 2763.380 ;
        RECT 2038.020 2763.370 2041.020 2763.380 ;
        RECT 2218.020 2763.370 2221.020 2763.380 ;
        RECT 2398.020 2763.370 2401.020 2763.380 ;
        RECT 2578.020 2763.370 2581.020 2763.380 ;
        RECT 2758.020 2763.370 2761.020 2763.380 ;
        RECT 2954.200 2763.370 2957.200 2763.380 ;
        RECT -37.580 2586.380 -34.580 2586.390 ;
        RECT 58.020 2586.380 61.020 2586.390 ;
        RECT 238.020 2586.380 241.020 2586.390 ;
        RECT 418.020 2586.380 421.020 2586.390 ;
        RECT 598.020 2586.380 601.020 2586.390 ;
        RECT 778.020 2586.380 781.020 2586.390 ;
        RECT 958.020 2586.380 961.020 2586.390 ;
        RECT 1138.020 2586.380 1141.020 2586.390 ;
        RECT 1318.020 2586.380 1321.020 2586.390 ;
        RECT 1498.020 2586.380 1501.020 2586.390 ;
        RECT 1678.020 2586.380 1681.020 2586.390 ;
        RECT 1858.020 2586.380 1861.020 2586.390 ;
        RECT 2038.020 2586.380 2041.020 2586.390 ;
        RECT 2218.020 2586.380 2221.020 2586.390 ;
        RECT 2398.020 2586.380 2401.020 2586.390 ;
        RECT 2578.020 2586.380 2581.020 2586.390 ;
        RECT 2758.020 2586.380 2761.020 2586.390 ;
        RECT 2954.200 2586.380 2957.200 2586.390 ;
        RECT -42.180 2583.380 2961.800 2586.380 ;
        RECT -37.580 2583.370 -34.580 2583.380 ;
        RECT 58.020 2583.370 61.020 2583.380 ;
        RECT 238.020 2583.370 241.020 2583.380 ;
        RECT 418.020 2583.370 421.020 2583.380 ;
        RECT 598.020 2583.370 601.020 2583.380 ;
        RECT 778.020 2583.370 781.020 2583.380 ;
        RECT 958.020 2583.370 961.020 2583.380 ;
        RECT 1138.020 2583.370 1141.020 2583.380 ;
        RECT 1318.020 2583.370 1321.020 2583.380 ;
        RECT 1498.020 2583.370 1501.020 2583.380 ;
        RECT 1678.020 2583.370 1681.020 2583.380 ;
        RECT 1858.020 2583.370 1861.020 2583.380 ;
        RECT 2038.020 2583.370 2041.020 2583.380 ;
        RECT 2218.020 2583.370 2221.020 2583.380 ;
        RECT 2398.020 2583.370 2401.020 2583.380 ;
        RECT 2578.020 2583.370 2581.020 2583.380 ;
        RECT 2758.020 2583.370 2761.020 2583.380 ;
        RECT 2954.200 2583.370 2957.200 2583.380 ;
        RECT -37.580 2406.380 -34.580 2406.390 ;
        RECT 58.020 2406.380 61.020 2406.390 ;
        RECT 238.020 2406.380 241.020 2406.390 ;
        RECT 418.020 2406.380 421.020 2406.390 ;
        RECT 598.020 2406.380 601.020 2406.390 ;
        RECT 778.020 2406.380 781.020 2406.390 ;
        RECT 958.020 2406.380 961.020 2406.390 ;
        RECT 1138.020 2406.380 1141.020 2406.390 ;
        RECT 1318.020 2406.380 1321.020 2406.390 ;
        RECT 1498.020 2406.380 1501.020 2406.390 ;
        RECT 1678.020 2406.380 1681.020 2406.390 ;
        RECT 1858.020 2406.380 1861.020 2406.390 ;
        RECT 2038.020 2406.380 2041.020 2406.390 ;
        RECT 2218.020 2406.380 2221.020 2406.390 ;
        RECT 2398.020 2406.380 2401.020 2406.390 ;
        RECT 2578.020 2406.380 2581.020 2406.390 ;
        RECT 2758.020 2406.380 2761.020 2406.390 ;
        RECT 2954.200 2406.380 2957.200 2406.390 ;
        RECT -42.180 2403.380 2961.800 2406.380 ;
        RECT -37.580 2403.370 -34.580 2403.380 ;
        RECT 58.020 2403.370 61.020 2403.380 ;
        RECT 238.020 2403.370 241.020 2403.380 ;
        RECT 418.020 2403.370 421.020 2403.380 ;
        RECT 598.020 2403.370 601.020 2403.380 ;
        RECT 778.020 2403.370 781.020 2403.380 ;
        RECT 958.020 2403.370 961.020 2403.380 ;
        RECT 1138.020 2403.370 1141.020 2403.380 ;
        RECT 1318.020 2403.370 1321.020 2403.380 ;
        RECT 1498.020 2403.370 1501.020 2403.380 ;
        RECT 1678.020 2403.370 1681.020 2403.380 ;
        RECT 1858.020 2403.370 1861.020 2403.380 ;
        RECT 2038.020 2403.370 2041.020 2403.380 ;
        RECT 2218.020 2403.370 2221.020 2403.380 ;
        RECT 2398.020 2403.370 2401.020 2403.380 ;
        RECT 2578.020 2403.370 2581.020 2403.380 ;
        RECT 2758.020 2403.370 2761.020 2403.380 ;
        RECT 2954.200 2403.370 2957.200 2403.380 ;
        RECT -37.580 2226.380 -34.580 2226.390 ;
        RECT 58.020 2226.380 61.020 2226.390 ;
        RECT 238.020 2226.380 241.020 2226.390 ;
        RECT 418.020 2226.380 421.020 2226.390 ;
        RECT 598.020 2226.380 601.020 2226.390 ;
        RECT 778.020 2226.380 781.020 2226.390 ;
        RECT 958.020 2226.380 961.020 2226.390 ;
        RECT 1138.020 2226.380 1141.020 2226.390 ;
        RECT 1318.020 2226.380 1321.020 2226.390 ;
        RECT 1498.020 2226.380 1501.020 2226.390 ;
        RECT 1678.020 2226.380 1681.020 2226.390 ;
        RECT 1858.020 2226.380 1861.020 2226.390 ;
        RECT 2038.020 2226.380 2041.020 2226.390 ;
        RECT 2218.020 2226.380 2221.020 2226.390 ;
        RECT 2398.020 2226.380 2401.020 2226.390 ;
        RECT 2578.020 2226.380 2581.020 2226.390 ;
        RECT 2758.020 2226.380 2761.020 2226.390 ;
        RECT 2954.200 2226.380 2957.200 2226.390 ;
        RECT -42.180 2223.380 2961.800 2226.380 ;
        RECT -37.580 2223.370 -34.580 2223.380 ;
        RECT 58.020 2223.370 61.020 2223.380 ;
        RECT 238.020 2223.370 241.020 2223.380 ;
        RECT 418.020 2223.370 421.020 2223.380 ;
        RECT 598.020 2223.370 601.020 2223.380 ;
        RECT 778.020 2223.370 781.020 2223.380 ;
        RECT 958.020 2223.370 961.020 2223.380 ;
        RECT 1138.020 2223.370 1141.020 2223.380 ;
        RECT 1318.020 2223.370 1321.020 2223.380 ;
        RECT 1498.020 2223.370 1501.020 2223.380 ;
        RECT 1678.020 2223.370 1681.020 2223.380 ;
        RECT 1858.020 2223.370 1861.020 2223.380 ;
        RECT 2038.020 2223.370 2041.020 2223.380 ;
        RECT 2218.020 2223.370 2221.020 2223.380 ;
        RECT 2398.020 2223.370 2401.020 2223.380 ;
        RECT 2578.020 2223.370 2581.020 2223.380 ;
        RECT 2758.020 2223.370 2761.020 2223.380 ;
        RECT 2954.200 2223.370 2957.200 2223.380 ;
        RECT -37.580 2046.380 -34.580 2046.390 ;
        RECT 58.020 2046.380 61.020 2046.390 ;
        RECT 238.020 2046.380 241.020 2046.390 ;
        RECT 418.020 2046.380 421.020 2046.390 ;
        RECT 598.020 2046.380 601.020 2046.390 ;
        RECT 778.020 2046.380 781.020 2046.390 ;
        RECT 958.020 2046.380 961.020 2046.390 ;
        RECT 1138.020 2046.380 1141.020 2046.390 ;
        RECT 1318.020 2046.380 1321.020 2046.390 ;
        RECT 1498.020 2046.380 1501.020 2046.390 ;
        RECT 1678.020 2046.380 1681.020 2046.390 ;
        RECT 1858.020 2046.380 1861.020 2046.390 ;
        RECT 2038.020 2046.380 2041.020 2046.390 ;
        RECT 2218.020 2046.380 2221.020 2046.390 ;
        RECT 2398.020 2046.380 2401.020 2046.390 ;
        RECT 2578.020 2046.380 2581.020 2046.390 ;
        RECT 2758.020 2046.380 2761.020 2046.390 ;
        RECT 2954.200 2046.380 2957.200 2046.390 ;
        RECT -42.180 2043.380 2961.800 2046.380 ;
        RECT -37.580 2043.370 -34.580 2043.380 ;
        RECT 58.020 2043.370 61.020 2043.380 ;
        RECT 238.020 2043.370 241.020 2043.380 ;
        RECT 418.020 2043.370 421.020 2043.380 ;
        RECT 598.020 2043.370 601.020 2043.380 ;
        RECT 778.020 2043.370 781.020 2043.380 ;
        RECT 958.020 2043.370 961.020 2043.380 ;
        RECT 1138.020 2043.370 1141.020 2043.380 ;
        RECT 1318.020 2043.370 1321.020 2043.380 ;
        RECT 1498.020 2043.370 1501.020 2043.380 ;
        RECT 1678.020 2043.370 1681.020 2043.380 ;
        RECT 1858.020 2043.370 1861.020 2043.380 ;
        RECT 2038.020 2043.370 2041.020 2043.380 ;
        RECT 2218.020 2043.370 2221.020 2043.380 ;
        RECT 2398.020 2043.370 2401.020 2043.380 ;
        RECT 2578.020 2043.370 2581.020 2043.380 ;
        RECT 2758.020 2043.370 2761.020 2043.380 ;
        RECT 2954.200 2043.370 2957.200 2043.380 ;
        RECT -37.580 1866.380 -34.580 1866.390 ;
        RECT 58.020 1866.380 61.020 1866.390 ;
        RECT 238.020 1866.380 241.020 1866.390 ;
        RECT 418.020 1866.380 421.020 1866.390 ;
        RECT 598.020 1866.380 601.020 1866.390 ;
        RECT 778.020 1866.380 781.020 1866.390 ;
        RECT 958.020 1866.380 961.020 1866.390 ;
        RECT 1138.020 1866.380 1141.020 1866.390 ;
        RECT 1318.020 1866.380 1321.020 1866.390 ;
        RECT 1498.020 1866.380 1501.020 1866.390 ;
        RECT 1678.020 1866.380 1681.020 1866.390 ;
        RECT 1858.020 1866.380 1861.020 1866.390 ;
        RECT 2038.020 1866.380 2041.020 1866.390 ;
        RECT 2218.020 1866.380 2221.020 1866.390 ;
        RECT 2398.020 1866.380 2401.020 1866.390 ;
        RECT 2578.020 1866.380 2581.020 1866.390 ;
        RECT 2758.020 1866.380 2761.020 1866.390 ;
        RECT 2954.200 1866.380 2957.200 1866.390 ;
        RECT -42.180 1863.380 2961.800 1866.380 ;
        RECT -37.580 1863.370 -34.580 1863.380 ;
        RECT 58.020 1863.370 61.020 1863.380 ;
        RECT 238.020 1863.370 241.020 1863.380 ;
        RECT 418.020 1863.370 421.020 1863.380 ;
        RECT 598.020 1863.370 601.020 1863.380 ;
        RECT 778.020 1863.370 781.020 1863.380 ;
        RECT 958.020 1863.370 961.020 1863.380 ;
        RECT 1138.020 1863.370 1141.020 1863.380 ;
        RECT 1318.020 1863.370 1321.020 1863.380 ;
        RECT 1498.020 1863.370 1501.020 1863.380 ;
        RECT 1678.020 1863.370 1681.020 1863.380 ;
        RECT 1858.020 1863.370 1861.020 1863.380 ;
        RECT 2038.020 1863.370 2041.020 1863.380 ;
        RECT 2218.020 1863.370 2221.020 1863.380 ;
        RECT 2398.020 1863.370 2401.020 1863.380 ;
        RECT 2578.020 1863.370 2581.020 1863.380 ;
        RECT 2758.020 1863.370 2761.020 1863.380 ;
        RECT 2954.200 1863.370 2957.200 1863.380 ;
        RECT -37.580 1686.380 -34.580 1686.390 ;
        RECT 58.020 1686.380 61.020 1686.390 ;
        RECT 238.020 1686.380 241.020 1686.390 ;
        RECT 418.020 1686.380 421.020 1686.390 ;
        RECT 598.020 1686.380 601.020 1686.390 ;
        RECT 778.020 1686.380 781.020 1686.390 ;
        RECT 958.020 1686.380 961.020 1686.390 ;
        RECT 1138.020 1686.380 1141.020 1686.390 ;
        RECT 1318.020 1686.380 1321.020 1686.390 ;
        RECT 1498.020 1686.380 1501.020 1686.390 ;
        RECT 1678.020 1686.380 1681.020 1686.390 ;
        RECT 1858.020 1686.380 1861.020 1686.390 ;
        RECT 2038.020 1686.380 2041.020 1686.390 ;
        RECT 2218.020 1686.380 2221.020 1686.390 ;
        RECT 2398.020 1686.380 2401.020 1686.390 ;
        RECT 2578.020 1686.380 2581.020 1686.390 ;
        RECT 2758.020 1686.380 2761.020 1686.390 ;
        RECT 2954.200 1686.380 2957.200 1686.390 ;
        RECT -42.180 1683.380 2961.800 1686.380 ;
        RECT -37.580 1683.370 -34.580 1683.380 ;
        RECT 58.020 1683.370 61.020 1683.380 ;
        RECT 238.020 1683.370 241.020 1683.380 ;
        RECT 418.020 1683.370 421.020 1683.380 ;
        RECT 598.020 1683.370 601.020 1683.380 ;
        RECT 778.020 1683.370 781.020 1683.380 ;
        RECT 958.020 1683.370 961.020 1683.380 ;
        RECT 1138.020 1683.370 1141.020 1683.380 ;
        RECT 1318.020 1683.370 1321.020 1683.380 ;
        RECT 1498.020 1683.370 1501.020 1683.380 ;
        RECT 1678.020 1683.370 1681.020 1683.380 ;
        RECT 1858.020 1683.370 1861.020 1683.380 ;
        RECT 2038.020 1683.370 2041.020 1683.380 ;
        RECT 2218.020 1683.370 2221.020 1683.380 ;
        RECT 2398.020 1683.370 2401.020 1683.380 ;
        RECT 2578.020 1683.370 2581.020 1683.380 ;
        RECT 2758.020 1683.370 2761.020 1683.380 ;
        RECT 2954.200 1683.370 2957.200 1683.380 ;
        RECT -37.580 1506.380 -34.580 1506.390 ;
        RECT 58.020 1506.380 61.020 1506.390 ;
        RECT 238.020 1506.380 241.020 1506.390 ;
        RECT 418.020 1506.380 421.020 1506.390 ;
        RECT 598.020 1506.380 601.020 1506.390 ;
        RECT 778.020 1506.380 781.020 1506.390 ;
        RECT 958.020 1506.380 961.020 1506.390 ;
        RECT 1138.020 1506.380 1141.020 1506.390 ;
        RECT 1318.020 1506.380 1321.020 1506.390 ;
        RECT 1498.020 1506.380 1501.020 1506.390 ;
        RECT 1678.020 1506.380 1681.020 1506.390 ;
        RECT 1858.020 1506.380 1861.020 1506.390 ;
        RECT 2038.020 1506.380 2041.020 1506.390 ;
        RECT 2218.020 1506.380 2221.020 1506.390 ;
        RECT 2398.020 1506.380 2401.020 1506.390 ;
        RECT 2578.020 1506.380 2581.020 1506.390 ;
        RECT 2758.020 1506.380 2761.020 1506.390 ;
        RECT 2954.200 1506.380 2957.200 1506.390 ;
        RECT -42.180 1503.380 2961.800 1506.380 ;
        RECT -37.580 1503.370 -34.580 1503.380 ;
        RECT 58.020 1503.370 61.020 1503.380 ;
        RECT 238.020 1503.370 241.020 1503.380 ;
        RECT 418.020 1503.370 421.020 1503.380 ;
        RECT 598.020 1503.370 601.020 1503.380 ;
        RECT 778.020 1503.370 781.020 1503.380 ;
        RECT 958.020 1503.370 961.020 1503.380 ;
        RECT 1138.020 1503.370 1141.020 1503.380 ;
        RECT 1318.020 1503.370 1321.020 1503.380 ;
        RECT 1498.020 1503.370 1501.020 1503.380 ;
        RECT 1678.020 1503.370 1681.020 1503.380 ;
        RECT 1858.020 1503.370 1861.020 1503.380 ;
        RECT 2038.020 1503.370 2041.020 1503.380 ;
        RECT 2218.020 1503.370 2221.020 1503.380 ;
        RECT 2398.020 1503.370 2401.020 1503.380 ;
        RECT 2578.020 1503.370 2581.020 1503.380 ;
        RECT 2758.020 1503.370 2761.020 1503.380 ;
        RECT 2954.200 1503.370 2957.200 1503.380 ;
        RECT -37.580 1326.380 -34.580 1326.390 ;
        RECT 58.020 1326.380 61.020 1326.390 ;
        RECT 238.020 1326.380 241.020 1326.390 ;
        RECT 418.020 1326.380 421.020 1326.390 ;
        RECT 598.020 1326.380 601.020 1326.390 ;
        RECT 778.020 1326.380 781.020 1326.390 ;
        RECT 958.020 1326.380 961.020 1326.390 ;
        RECT 1138.020 1326.380 1141.020 1326.390 ;
        RECT 1318.020 1326.380 1321.020 1326.390 ;
        RECT 1498.020 1326.380 1501.020 1326.390 ;
        RECT 1678.020 1326.380 1681.020 1326.390 ;
        RECT 1858.020 1326.380 1861.020 1326.390 ;
        RECT 2038.020 1326.380 2041.020 1326.390 ;
        RECT 2218.020 1326.380 2221.020 1326.390 ;
        RECT 2398.020 1326.380 2401.020 1326.390 ;
        RECT 2578.020 1326.380 2581.020 1326.390 ;
        RECT 2758.020 1326.380 2761.020 1326.390 ;
        RECT 2954.200 1326.380 2957.200 1326.390 ;
        RECT -42.180 1323.380 2961.800 1326.380 ;
        RECT -37.580 1323.370 -34.580 1323.380 ;
        RECT 58.020 1323.370 61.020 1323.380 ;
        RECT 238.020 1323.370 241.020 1323.380 ;
        RECT 418.020 1323.370 421.020 1323.380 ;
        RECT 598.020 1323.370 601.020 1323.380 ;
        RECT 778.020 1323.370 781.020 1323.380 ;
        RECT 958.020 1323.370 961.020 1323.380 ;
        RECT 1138.020 1323.370 1141.020 1323.380 ;
        RECT 1318.020 1323.370 1321.020 1323.380 ;
        RECT 1498.020 1323.370 1501.020 1323.380 ;
        RECT 1678.020 1323.370 1681.020 1323.380 ;
        RECT 1858.020 1323.370 1861.020 1323.380 ;
        RECT 2038.020 1323.370 2041.020 1323.380 ;
        RECT 2218.020 1323.370 2221.020 1323.380 ;
        RECT 2398.020 1323.370 2401.020 1323.380 ;
        RECT 2578.020 1323.370 2581.020 1323.380 ;
        RECT 2758.020 1323.370 2761.020 1323.380 ;
        RECT 2954.200 1323.370 2957.200 1323.380 ;
        RECT -37.580 1146.380 -34.580 1146.390 ;
        RECT 58.020 1146.380 61.020 1146.390 ;
        RECT 238.020 1146.380 241.020 1146.390 ;
        RECT 418.020 1146.380 421.020 1146.390 ;
        RECT 598.020 1146.380 601.020 1146.390 ;
        RECT 778.020 1146.380 781.020 1146.390 ;
        RECT 958.020 1146.380 961.020 1146.390 ;
        RECT 1138.020 1146.380 1141.020 1146.390 ;
        RECT 1318.020 1146.380 1321.020 1146.390 ;
        RECT 1498.020 1146.380 1501.020 1146.390 ;
        RECT 1678.020 1146.380 1681.020 1146.390 ;
        RECT 1858.020 1146.380 1861.020 1146.390 ;
        RECT 2038.020 1146.380 2041.020 1146.390 ;
        RECT 2218.020 1146.380 2221.020 1146.390 ;
        RECT 2398.020 1146.380 2401.020 1146.390 ;
        RECT 2578.020 1146.380 2581.020 1146.390 ;
        RECT 2758.020 1146.380 2761.020 1146.390 ;
        RECT 2954.200 1146.380 2957.200 1146.390 ;
        RECT -42.180 1143.380 2961.800 1146.380 ;
        RECT -37.580 1143.370 -34.580 1143.380 ;
        RECT 58.020 1143.370 61.020 1143.380 ;
        RECT 238.020 1143.370 241.020 1143.380 ;
        RECT 418.020 1143.370 421.020 1143.380 ;
        RECT 598.020 1143.370 601.020 1143.380 ;
        RECT 778.020 1143.370 781.020 1143.380 ;
        RECT 958.020 1143.370 961.020 1143.380 ;
        RECT 1138.020 1143.370 1141.020 1143.380 ;
        RECT 1318.020 1143.370 1321.020 1143.380 ;
        RECT 1498.020 1143.370 1501.020 1143.380 ;
        RECT 1678.020 1143.370 1681.020 1143.380 ;
        RECT 1858.020 1143.370 1861.020 1143.380 ;
        RECT 2038.020 1143.370 2041.020 1143.380 ;
        RECT 2218.020 1143.370 2221.020 1143.380 ;
        RECT 2398.020 1143.370 2401.020 1143.380 ;
        RECT 2578.020 1143.370 2581.020 1143.380 ;
        RECT 2758.020 1143.370 2761.020 1143.380 ;
        RECT 2954.200 1143.370 2957.200 1143.380 ;
        RECT -37.580 966.380 -34.580 966.390 ;
        RECT 58.020 966.380 61.020 966.390 ;
        RECT 238.020 966.380 241.020 966.390 ;
        RECT 418.020 966.380 421.020 966.390 ;
        RECT 598.020 966.380 601.020 966.390 ;
        RECT 778.020 966.380 781.020 966.390 ;
        RECT 958.020 966.380 961.020 966.390 ;
        RECT 1138.020 966.380 1141.020 966.390 ;
        RECT 1318.020 966.380 1321.020 966.390 ;
        RECT 1498.020 966.380 1501.020 966.390 ;
        RECT 1678.020 966.380 1681.020 966.390 ;
        RECT 1858.020 966.380 1861.020 966.390 ;
        RECT 2038.020 966.380 2041.020 966.390 ;
        RECT 2218.020 966.380 2221.020 966.390 ;
        RECT 2398.020 966.380 2401.020 966.390 ;
        RECT 2578.020 966.380 2581.020 966.390 ;
        RECT 2758.020 966.380 2761.020 966.390 ;
        RECT 2954.200 966.380 2957.200 966.390 ;
        RECT -42.180 963.380 2961.800 966.380 ;
        RECT -37.580 963.370 -34.580 963.380 ;
        RECT 58.020 963.370 61.020 963.380 ;
        RECT 238.020 963.370 241.020 963.380 ;
        RECT 418.020 963.370 421.020 963.380 ;
        RECT 598.020 963.370 601.020 963.380 ;
        RECT 778.020 963.370 781.020 963.380 ;
        RECT 958.020 963.370 961.020 963.380 ;
        RECT 1138.020 963.370 1141.020 963.380 ;
        RECT 1318.020 963.370 1321.020 963.380 ;
        RECT 1498.020 963.370 1501.020 963.380 ;
        RECT 1678.020 963.370 1681.020 963.380 ;
        RECT 1858.020 963.370 1861.020 963.380 ;
        RECT 2038.020 963.370 2041.020 963.380 ;
        RECT 2218.020 963.370 2221.020 963.380 ;
        RECT 2398.020 963.370 2401.020 963.380 ;
        RECT 2578.020 963.370 2581.020 963.380 ;
        RECT 2758.020 963.370 2761.020 963.380 ;
        RECT 2954.200 963.370 2957.200 963.380 ;
        RECT -37.580 786.380 -34.580 786.390 ;
        RECT 58.020 786.380 61.020 786.390 ;
        RECT 238.020 786.380 241.020 786.390 ;
        RECT 418.020 786.380 421.020 786.390 ;
        RECT 598.020 786.380 601.020 786.390 ;
        RECT 778.020 786.380 781.020 786.390 ;
        RECT 958.020 786.380 961.020 786.390 ;
        RECT 1138.020 786.380 1141.020 786.390 ;
        RECT 1318.020 786.380 1321.020 786.390 ;
        RECT 1498.020 786.380 1501.020 786.390 ;
        RECT 1678.020 786.380 1681.020 786.390 ;
        RECT 1858.020 786.380 1861.020 786.390 ;
        RECT 2038.020 786.380 2041.020 786.390 ;
        RECT 2218.020 786.380 2221.020 786.390 ;
        RECT 2398.020 786.380 2401.020 786.390 ;
        RECT 2578.020 786.380 2581.020 786.390 ;
        RECT 2758.020 786.380 2761.020 786.390 ;
        RECT 2954.200 786.380 2957.200 786.390 ;
        RECT -42.180 783.380 2961.800 786.380 ;
        RECT -37.580 783.370 -34.580 783.380 ;
        RECT 58.020 783.370 61.020 783.380 ;
        RECT 238.020 783.370 241.020 783.380 ;
        RECT 418.020 783.370 421.020 783.380 ;
        RECT 598.020 783.370 601.020 783.380 ;
        RECT 778.020 783.370 781.020 783.380 ;
        RECT 958.020 783.370 961.020 783.380 ;
        RECT 1138.020 783.370 1141.020 783.380 ;
        RECT 1318.020 783.370 1321.020 783.380 ;
        RECT 1498.020 783.370 1501.020 783.380 ;
        RECT 1678.020 783.370 1681.020 783.380 ;
        RECT 1858.020 783.370 1861.020 783.380 ;
        RECT 2038.020 783.370 2041.020 783.380 ;
        RECT 2218.020 783.370 2221.020 783.380 ;
        RECT 2398.020 783.370 2401.020 783.380 ;
        RECT 2578.020 783.370 2581.020 783.380 ;
        RECT 2758.020 783.370 2761.020 783.380 ;
        RECT 2954.200 783.370 2957.200 783.380 ;
        RECT -37.580 606.380 -34.580 606.390 ;
        RECT 58.020 606.380 61.020 606.390 ;
        RECT 238.020 606.380 241.020 606.390 ;
        RECT 418.020 606.380 421.020 606.390 ;
        RECT 598.020 606.380 601.020 606.390 ;
        RECT 778.020 606.380 781.020 606.390 ;
        RECT 958.020 606.380 961.020 606.390 ;
        RECT 1138.020 606.380 1141.020 606.390 ;
        RECT 1318.020 606.380 1321.020 606.390 ;
        RECT 1498.020 606.380 1501.020 606.390 ;
        RECT 1678.020 606.380 1681.020 606.390 ;
        RECT 1858.020 606.380 1861.020 606.390 ;
        RECT 2038.020 606.380 2041.020 606.390 ;
        RECT 2218.020 606.380 2221.020 606.390 ;
        RECT 2398.020 606.380 2401.020 606.390 ;
        RECT 2578.020 606.380 2581.020 606.390 ;
        RECT 2758.020 606.380 2761.020 606.390 ;
        RECT 2954.200 606.380 2957.200 606.390 ;
        RECT -42.180 603.380 2961.800 606.380 ;
        RECT -37.580 603.370 -34.580 603.380 ;
        RECT 58.020 603.370 61.020 603.380 ;
        RECT 238.020 603.370 241.020 603.380 ;
        RECT 418.020 603.370 421.020 603.380 ;
        RECT 598.020 603.370 601.020 603.380 ;
        RECT 778.020 603.370 781.020 603.380 ;
        RECT 958.020 603.370 961.020 603.380 ;
        RECT 1138.020 603.370 1141.020 603.380 ;
        RECT 1318.020 603.370 1321.020 603.380 ;
        RECT 1498.020 603.370 1501.020 603.380 ;
        RECT 1678.020 603.370 1681.020 603.380 ;
        RECT 1858.020 603.370 1861.020 603.380 ;
        RECT 2038.020 603.370 2041.020 603.380 ;
        RECT 2218.020 603.370 2221.020 603.380 ;
        RECT 2398.020 603.370 2401.020 603.380 ;
        RECT 2578.020 603.370 2581.020 603.380 ;
        RECT 2758.020 603.370 2761.020 603.380 ;
        RECT 2954.200 603.370 2957.200 603.380 ;
        RECT -37.580 426.380 -34.580 426.390 ;
        RECT 58.020 426.380 61.020 426.390 ;
        RECT 238.020 426.380 241.020 426.390 ;
        RECT 418.020 426.380 421.020 426.390 ;
        RECT 598.020 426.380 601.020 426.390 ;
        RECT 778.020 426.380 781.020 426.390 ;
        RECT 958.020 426.380 961.020 426.390 ;
        RECT 1138.020 426.380 1141.020 426.390 ;
        RECT 1318.020 426.380 1321.020 426.390 ;
        RECT 1498.020 426.380 1501.020 426.390 ;
        RECT 1678.020 426.380 1681.020 426.390 ;
        RECT 1858.020 426.380 1861.020 426.390 ;
        RECT 2038.020 426.380 2041.020 426.390 ;
        RECT 2218.020 426.380 2221.020 426.390 ;
        RECT 2398.020 426.380 2401.020 426.390 ;
        RECT 2578.020 426.380 2581.020 426.390 ;
        RECT 2758.020 426.380 2761.020 426.390 ;
        RECT 2954.200 426.380 2957.200 426.390 ;
        RECT -42.180 423.380 2961.800 426.380 ;
        RECT -37.580 423.370 -34.580 423.380 ;
        RECT 58.020 423.370 61.020 423.380 ;
        RECT 238.020 423.370 241.020 423.380 ;
        RECT 418.020 423.370 421.020 423.380 ;
        RECT 598.020 423.370 601.020 423.380 ;
        RECT 778.020 423.370 781.020 423.380 ;
        RECT 958.020 423.370 961.020 423.380 ;
        RECT 1138.020 423.370 1141.020 423.380 ;
        RECT 1318.020 423.370 1321.020 423.380 ;
        RECT 1498.020 423.370 1501.020 423.380 ;
        RECT 1678.020 423.370 1681.020 423.380 ;
        RECT 1858.020 423.370 1861.020 423.380 ;
        RECT 2038.020 423.370 2041.020 423.380 ;
        RECT 2218.020 423.370 2221.020 423.380 ;
        RECT 2398.020 423.370 2401.020 423.380 ;
        RECT 2578.020 423.370 2581.020 423.380 ;
        RECT 2758.020 423.370 2761.020 423.380 ;
        RECT 2954.200 423.370 2957.200 423.380 ;
        RECT -37.580 246.380 -34.580 246.390 ;
        RECT 58.020 246.380 61.020 246.390 ;
        RECT 238.020 246.380 241.020 246.390 ;
        RECT 418.020 246.380 421.020 246.390 ;
        RECT 598.020 246.380 601.020 246.390 ;
        RECT 778.020 246.380 781.020 246.390 ;
        RECT 958.020 246.380 961.020 246.390 ;
        RECT 1138.020 246.380 1141.020 246.390 ;
        RECT 1318.020 246.380 1321.020 246.390 ;
        RECT 1498.020 246.380 1501.020 246.390 ;
        RECT 1678.020 246.380 1681.020 246.390 ;
        RECT 1858.020 246.380 1861.020 246.390 ;
        RECT 2038.020 246.380 2041.020 246.390 ;
        RECT 2218.020 246.380 2221.020 246.390 ;
        RECT 2398.020 246.380 2401.020 246.390 ;
        RECT 2578.020 246.380 2581.020 246.390 ;
        RECT 2758.020 246.380 2761.020 246.390 ;
        RECT 2954.200 246.380 2957.200 246.390 ;
        RECT -42.180 243.380 2961.800 246.380 ;
        RECT -37.580 243.370 -34.580 243.380 ;
        RECT 58.020 243.370 61.020 243.380 ;
        RECT 238.020 243.370 241.020 243.380 ;
        RECT 418.020 243.370 421.020 243.380 ;
        RECT 598.020 243.370 601.020 243.380 ;
        RECT 778.020 243.370 781.020 243.380 ;
        RECT 958.020 243.370 961.020 243.380 ;
        RECT 1138.020 243.370 1141.020 243.380 ;
        RECT 1318.020 243.370 1321.020 243.380 ;
        RECT 1498.020 243.370 1501.020 243.380 ;
        RECT 1678.020 243.370 1681.020 243.380 ;
        RECT 1858.020 243.370 1861.020 243.380 ;
        RECT 2038.020 243.370 2041.020 243.380 ;
        RECT 2218.020 243.370 2221.020 243.380 ;
        RECT 2398.020 243.370 2401.020 243.380 ;
        RECT 2578.020 243.370 2581.020 243.380 ;
        RECT 2758.020 243.370 2761.020 243.380 ;
        RECT 2954.200 243.370 2957.200 243.380 ;
        RECT -37.580 66.380 -34.580 66.390 ;
        RECT 58.020 66.380 61.020 66.390 ;
        RECT 238.020 66.380 241.020 66.390 ;
        RECT 418.020 66.380 421.020 66.390 ;
        RECT 598.020 66.380 601.020 66.390 ;
        RECT 778.020 66.380 781.020 66.390 ;
        RECT 958.020 66.380 961.020 66.390 ;
        RECT 1138.020 66.380 1141.020 66.390 ;
        RECT 1318.020 66.380 1321.020 66.390 ;
        RECT 1498.020 66.380 1501.020 66.390 ;
        RECT 1678.020 66.380 1681.020 66.390 ;
        RECT 1858.020 66.380 1861.020 66.390 ;
        RECT 2038.020 66.380 2041.020 66.390 ;
        RECT 2218.020 66.380 2221.020 66.390 ;
        RECT 2398.020 66.380 2401.020 66.390 ;
        RECT 2578.020 66.380 2581.020 66.390 ;
        RECT 2758.020 66.380 2761.020 66.390 ;
        RECT 2954.200 66.380 2957.200 66.390 ;
        RECT -42.180 63.380 2961.800 66.380 ;
        RECT -37.580 63.370 -34.580 63.380 ;
        RECT 58.020 63.370 61.020 63.380 ;
        RECT 238.020 63.370 241.020 63.380 ;
        RECT 418.020 63.370 421.020 63.380 ;
        RECT 598.020 63.370 601.020 63.380 ;
        RECT 778.020 63.370 781.020 63.380 ;
        RECT 958.020 63.370 961.020 63.380 ;
        RECT 1138.020 63.370 1141.020 63.380 ;
        RECT 1318.020 63.370 1321.020 63.380 ;
        RECT 1498.020 63.370 1501.020 63.380 ;
        RECT 1678.020 63.370 1681.020 63.380 ;
        RECT 1858.020 63.370 1861.020 63.380 ;
        RECT 2038.020 63.370 2041.020 63.380 ;
        RECT 2218.020 63.370 2221.020 63.380 ;
        RECT 2398.020 63.370 2401.020 63.380 ;
        RECT 2578.020 63.370 2581.020 63.380 ;
        RECT 2758.020 63.370 2761.020 63.380 ;
        RECT 2954.200 63.370 2957.200 63.380 ;
        RECT -37.580 -29.220 -34.580 -29.210 ;
        RECT 58.020 -29.220 61.020 -29.210 ;
        RECT 238.020 -29.220 241.020 -29.210 ;
        RECT 418.020 -29.220 421.020 -29.210 ;
        RECT 598.020 -29.220 601.020 -29.210 ;
        RECT 778.020 -29.220 781.020 -29.210 ;
        RECT 958.020 -29.220 961.020 -29.210 ;
        RECT 1138.020 -29.220 1141.020 -29.210 ;
        RECT 1318.020 -29.220 1321.020 -29.210 ;
        RECT 1498.020 -29.220 1501.020 -29.210 ;
        RECT 1678.020 -29.220 1681.020 -29.210 ;
        RECT 1858.020 -29.220 1861.020 -29.210 ;
        RECT 2038.020 -29.220 2041.020 -29.210 ;
        RECT 2218.020 -29.220 2221.020 -29.210 ;
        RECT 2398.020 -29.220 2401.020 -29.210 ;
        RECT 2578.020 -29.220 2581.020 -29.210 ;
        RECT 2758.020 -29.220 2761.020 -29.210 ;
        RECT 2954.200 -29.220 2957.200 -29.210 ;
        RECT -37.580 -32.220 2957.200 -29.220 ;
        RECT -37.580 -32.230 -34.580 -32.220 ;
        RECT 58.020 -32.230 61.020 -32.220 ;
        RECT 238.020 -32.230 241.020 -32.220 ;
        RECT 418.020 -32.230 421.020 -32.220 ;
        RECT 598.020 -32.230 601.020 -32.220 ;
        RECT 778.020 -32.230 781.020 -32.220 ;
        RECT 958.020 -32.230 961.020 -32.220 ;
        RECT 1138.020 -32.230 1141.020 -32.220 ;
        RECT 1318.020 -32.230 1321.020 -32.220 ;
        RECT 1498.020 -32.230 1501.020 -32.220 ;
        RECT 1678.020 -32.230 1681.020 -32.220 ;
        RECT 1858.020 -32.230 1861.020 -32.220 ;
        RECT 2038.020 -32.230 2041.020 -32.220 ;
        RECT 2218.020 -32.230 2221.020 -32.220 ;
        RECT 2398.020 -32.230 2401.020 -32.220 ;
        RECT 2578.020 -32.230 2581.020 -32.220 ;
        RECT 2758.020 -32.230 2761.020 -32.220 ;
        RECT 2954.200 -32.230 2957.200 -32.220 ;
    END
  END vdda2
  PIN vssa2
    DIRECTION INPUT ;
    PORT
      LAYER met4 ;
        RECT -42.180 -36.820 -39.180 3556.500 ;
        RECT 148.020 -36.820 151.020 3556.500 ;
        RECT 328.020 -36.820 331.020 3556.500 ;
        RECT 508.020 -36.820 511.020 3556.500 ;
        RECT 688.020 -36.820 691.020 3556.500 ;
        RECT 868.020 -36.820 871.020 3556.500 ;
        RECT 1048.020 -36.820 1051.020 3556.500 ;
        RECT 1228.020 -36.820 1231.020 3556.500 ;
        RECT 1408.020 -36.820 1411.020 3556.500 ;
        RECT 1588.020 -36.820 1591.020 3556.500 ;
        RECT 1768.020 -36.820 1771.020 3556.500 ;
        RECT 1948.020 -36.820 1951.020 3556.500 ;
        RECT 2128.020 -36.820 2131.020 3556.500 ;
        RECT 2308.020 -36.820 2311.020 3556.500 ;
        RECT 2488.020 -36.820 2491.020 3556.500 ;
        RECT 2668.020 -36.820 2671.020 3556.500 ;
        RECT 2848.020 -36.820 2851.020 3556.500 ;
        RECT 2958.800 -36.820 2961.800 3556.500 ;
      LAYER via4 ;
        RECT -41.270 3555.210 -40.090 3556.390 ;
        RECT -41.270 3553.610 -40.090 3554.790 ;
        RECT -41.270 3395.090 -40.090 3396.270 ;
        RECT -41.270 3393.490 -40.090 3394.670 ;
        RECT -41.270 3215.090 -40.090 3216.270 ;
        RECT -41.270 3213.490 -40.090 3214.670 ;
        RECT -41.270 3035.090 -40.090 3036.270 ;
        RECT -41.270 3033.490 -40.090 3034.670 ;
        RECT -41.270 2855.090 -40.090 2856.270 ;
        RECT -41.270 2853.490 -40.090 2854.670 ;
        RECT -41.270 2675.090 -40.090 2676.270 ;
        RECT -41.270 2673.490 -40.090 2674.670 ;
        RECT -41.270 2495.090 -40.090 2496.270 ;
        RECT -41.270 2493.490 -40.090 2494.670 ;
        RECT -41.270 2315.090 -40.090 2316.270 ;
        RECT -41.270 2313.490 -40.090 2314.670 ;
        RECT -41.270 2135.090 -40.090 2136.270 ;
        RECT -41.270 2133.490 -40.090 2134.670 ;
        RECT -41.270 1955.090 -40.090 1956.270 ;
        RECT -41.270 1953.490 -40.090 1954.670 ;
        RECT -41.270 1775.090 -40.090 1776.270 ;
        RECT -41.270 1773.490 -40.090 1774.670 ;
        RECT -41.270 1595.090 -40.090 1596.270 ;
        RECT -41.270 1593.490 -40.090 1594.670 ;
        RECT -41.270 1415.090 -40.090 1416.270 ;
        RECT -41.270 1413.490 -40.090 1414.670 ;
        RECT -41.270 1235.090 -40.090 1236.270 ;
        RECT -41.270 1233.490 -40.090 1234.670 ;
        RECT -41.270 1055.090 -40.090 1056.270 ;
        RECT -41.270 1053.490 -40.090 1054.670 ;
        RECT -41.270 875.090 -40.090 876.270 ;
        RECT -41.270 873.490 -40.090 874.670 ;
        RECT -41.270 695.090 -40.090 696.270 ;
        RECT -41.270 693.490 -40.090 694.670 ;
        RECT -41.270 515.090 -40.090 516.270 ;
        RECT -41.270 513.490 -40.090 514.670 ;
        RECT -41.270 335.090 -40.090 336.270 ;
        RECT -41.270 333.490 -40.090 334.670 ;
        RECT -41.270 155.090 -40.090 156.270 ;
        RECT -41.270 153.490 -40.090 154.670 ;
        RECT -41.270 -35.110 -40.090 -33.930 ;
        RECT -41.270 -36.710 -40.090 -35.530 ;
        RECT 148.930 3555.210 150.110 3556.390 ;
        RECT 148.930 3553.610 150.110 3554.790 ;
        RECT 148.930 3395.090 150.110 3396.270 ;
        RECT 148.930 3393.490 150.110 3394.670 ;
        RECT 148.930 3215.090 150.110 3216.270 ;
        RECT 148.930 3213.490 150.110 3214.670 ;
        RECT 148.930 3035.090 150.110 3036.270 ;
        RECT 148.930 3033.490 150.110 3034.670 ;
        RECT 148.930 2855.090 150.110 2856.270 ;
        RECT 148.930 2853.490 150.110 2854.670 ;
        RECT 148.930 2675.090 150.110 2676.270 ;
        RECT 148.930 2673.490 150.110 2674.670 ;
        RECT 148.930 2495.090 150.110 2496.270 ;
        RECT 148.930 2493.490 150.110 2494.670 ;
        RECT 148.930 2315.090 150.110 2316.270 ;
        RECT 148.930 2313.490 150.110 2314.670 ;
        RECT 148.930 2135.090 150.110 2136.270 ;
        RECT 148.930 2133.490 150.110 2134.670 ;
        RECT 148.930 1955.090 150.110 1956.270 ;
        RECT 148.930 1953.490 150.110 1954.670 ;
        RECT 148.930 1775.090 150.110 1776.270 ;
        RECT 148.930 1773.490 150.110 1774.670 ;
        RECT 148.930 1595.090 150.110 1596.270 ;
        RECT 148.930 1593.490 150.110 1594.670 ;
        RECT 148.930 1415.090 150.110 1416.270 ;
        RECT 148.930 1413.490 150.110 1414.670 ;
        RECT 148.930 1235.090 150.110 1236.270 ;
        RECT 148.930 1233.490 150.110 1234.670 ;
        RECT 148.930 1055.090 150.110 1056.270 ;
        RECT 148.930 1053.490 150.110 1054.670 ;
        RECT 148.930 875.090 150.110 876.270 ;
        RECT 148.930 873.490 150.110 874.670 ;
        RECT 148.930 695.090 150.110 696.270 ;
        RECT 148.930 693.490 150.110 694.670 ;
        RECT 148.930 515.090 150.110 516.270 ;
        RECT 148.930 513.490 150.110 514.670 ;
        RECT 148.930 335.090 150.110 336.270 ;
        RECT 148.930 333.490 150.110 334.670 ;
        RECT 148.930 155.090 150.110 156.270 ;
        RECT 148.930 153.490 150.110 154.670 ;
        RECT 148.930 -35.110 150.110 -33.930 ;
        RECT 148.930 -36.710 150.110 -35.530 ;
        RECT 328.930 3555.210 330.110 3556.390 ;
        RECT 328.930 3553.610 330.110 3554.790 ;
        RECT 328.930 3395.090 330.110 3396.270 ;
        RECT 328.930 3393.490 330.110 3394.670 ;
        RECT 328.930 3215.090 330.110 3216.270 ;
        RECT 328.930 3213.490 330.110 3214.670 ;
        RECT 328.930 3035.090 330.110 3036.270 ;
        RECT 328.930 3033.490 330.110 3034.670 ;
        RECT 328.930 2855.090 330.110 2856.270 ;
        RECT 328.930 2853.490 330.110 2854.670 ;
        RECT 328.930 2675.090 330.110 2676.270 ;
        RECT 328.930 2673.490 330.110 2674.670 ;
        RECT 328.930 2495.090 330.110 2496.270 ;
        RECT 328.930 2493.490 330.110 2494.670 ;
        RECT 328.930 2315.090 330.110 2316.270 ;
        RECT 328.930 2313.490 330.110 2314.670 ;
        RECT 328.930 2135.090 330.110 2136.270 ;
        RECT 328.930 2133.490 330.110 2134.670 ;
        RECT 328.930 1955.090 330.110 1956.270 ;
        RECT 328.930 1953.490 330.110 1954.670 ;
        RECT 328.930 1775.090 330.110 1776.270 ;
        RECT 328.930 1773.490 330.110 1774.670 ;
        RECT 328.930 1595.090 330.110 1596.270 ;
        RECT 328.930 1593.490 330.110 1594.670 ;
        RECT 328.930 1415.090 330.110 1416.270 ;
        RECT 328.930 1413.490 330.110 1414.670 ;
        RECT 328.930 1235.090 330.110 1236.270 ;
        RECT 328.930 1233.490 330.110 1234.670 ;
        RECT 328.930 1055.090 330.110 1056.270 ;
        RECT 328.930 1053.490 330.110 1054.670 ;
        RECT 328.930 875.090 330.110 876.270 ;
        RECT 328.930 873.490 330.110 874.670 ;
        RECT 328.930 695.090 330.110 696.270 ;
        RECT 328.930 693.490 330.110 694.670 ;
        RECT 328.930 515.090 330.110 516.270 ;
        RECT 328.930 513.490 330.110 514.670 ;
        RECT 328.930 335.090 330.110 336.270 ;
        RECT 328.930 333.490 330.110 334.670 ;
        RECT 328.930 155.090 330.110 156.270 ;
        RECT 328.930 153.490 330.110 154.670 ;
        RECT 328.930 -35.110 330.110 -33.930 ;
        RECT 328.930 -36.710 330.110 -35.530 ;
        RECT 508.930 3555.210 510.110 3556.390 ;
        RECT 508.930 3553.610 510.110 3554.790 ;
        RECT 508.930 3395.090 510.110 3396.270 ;
        RECT 508.930 3393.490 510.110 3394.670 ;
        RECT 508.930 3215.090 510.110 3216.270 ;
        RECT 508.930 3213.490 510.110 3214.670 ;
        RECT 508.930 3035.090 510.110 3036.270 ;
        RECT 508.930 3033.490 510.110 3034.670 ;
        RECT 508.930 2855.090 510.110 2856.270 ;
        RECT 508.930 2853.490 510.110 2854.670 ;
        RECT 508.930 2675.090 510.110 2676.270 ;
        RECT 508.930 2673.490 510.110 2674.670 ;
        RECT 508.930 2495.090 510.110 2496.270 ;
        RECT 508.930 2493.490 510.110 2494.670 ;
        RECT 508.930 2315.090 510.110 2316.270 ;
        RECT 508.930 2313.490 510.110 2314.670 ;
        RECT 508.930 2135.090 510.110 2136.270 ;
        RECT 508.930 2133.490 510.110 2134.670 ;
        RECT 508.930 1955.090 510.110 1956.270 ;
        RECT 508.930 1953.490 510.110 1954.670 ;
        RECT 508.930 1775.090 510.110 1776.270 ;
        RECT 508.930 1773.490 510.110 1774.670 ;
        RECT 508.930 1595.090 510.110 1596.270 ;
        RECT 508.930 1593.490 510.110 1594.670 ;
        RECT 508.930 1415.090 510.110 1416.270 ;
        RECT 508.930 1413.490 510.110 1414.670 ;
        RECT 508.930 1235.090 510.110 1236.270 ;
        RECT 508.930 1233.490 510.110 1234.670 ;
        RECT 508.930 1055.090 510.110 1056.270 ;
        RECT 508.930 1053.490 510.110 1054.670 ;
        RECT 508.930 875.090 510.110 876.270 ;
        RECT 508.930 873.490 510.110 874.670 ;
        RECT 508.930 695.090 510.110 696.270 ;
        RECT 508.930 693.490 510.110 694.670 ;
        RECT 508.930 515.090 510.110 516.270 ;
        RECT 508.930 513.490 510.110 514.670 ;
        RECT 508.930 335.090 510.110 336.270 ;
        RECT 508.930 333.490 510.110 334.670 ;
        RECT 508.930 155.090 510.110 156.270 ;
        RECT 508.930 153.490 510.110 154.670 ;
        RECT 508.930 -35.110 510.110 -33.930 ;
        RECT 508.930 -36.710 510.110 -35.530 ;
        RECT 688.930 3555.210 690.110 3556.390 ;
        RECT 688.930 3553.610 690.110 3554.790 ;
        RECT 688.930 3395.090 690.110 3396.270 ;
        RECT 688.930 3393.490 690.110 3394.670 ;
        RECT 688.930 3215.090 690.110 3216.270 ;
        RECT 688.930 3213.490 690.110 3214.670 ;
        RECT 688.930 3035.090 690.110 3036.270 ;
        RECT 688.930 3033.490 690.110 3034.670 ;
        RECT 688.930 2855.090 690.110 2856.270 ;
        RECT 688.930 2853.490 690.110 2854.670 ;
        RECT 688.930 2675.090 690.110 2676.270 ;
        RECT 688.930 2673.490 690.110 2674.670 ;
        RECT 688.930 2495.090 690.110 2496.270 ;
        RECT 688.930 2493.490 690.110 2494.670 ;
        RECT 688.930 2315.090 690.110 2316.270 ;
        RECT 688.930 2313.490 690.110 2314.670 ;
        RECT 688.930 2135.090 690.110 2136.270 ;
        RECT 688.930 2133.490 690.110 2134.670 ;
        RECT 688.930 1955.090 690.110 1956.270 ;
        RECT 688.930 1953.490 690.110 1954.670 ;
        RECT 688.930 1775.090 690.110 1776.270 ;
        RECT 688.930 1773.490 690.110 1774.670 ;
        RECT 688.930 1595.090 690.110 1596.270 ;
        RECT 688.930 1593.490 690.110 1594.670 ;
        RECT 688.930 1415.090 690.110 1416.270 ;
        RECT 688.930 1413.490 690.110 1414.670 ;
        RECT 688.930 1235.090 690.110 1236.270 ;
        RECT 688.930 1233.490 690.110 1234.670 ;
        RECT 688.930 1055.090 690.110 1056.270 ;
        RECT 688.930 1053.490 690.110 1054.670 ;
        RECT 688.930 875.090 690.110 876.270 ;
        RECT 688.930 873.490 690.110 874.670 ;
        RECT 688.930 695.090 690.110 696.270 ;
        RECT 688.930 693.490 690.110 694.670 ;
        RECT 688.930 515.090 690.110 516.270 ;
        RECT 688.930 513.490 690.110 514.670 ;
        RECT 688.930 335.090 690.110 336.270 ;
        RECT 688.930 333.490 690.110 334.670 ;
        RECT 688.930 155.090 690.110 156.270 ;
        RECT 688.930 153.490 690.110 154.670 ;
        RECT 688.930 -35.110 690.110 -33.930 ;
        RECT 688.930 -36.710 690.110 -35.530 ;
        RECT 868.930 3555.210 870.110 3556.390 ;
        RECT 868.930 3553.610 870.110 3554.790 ;
        RECT 868.930 3395.090 870.110 3396.270 ;
        RECT 868.930 3393.490 870.110 3394.670 ;
        RECT 868.930 3215.090 870.110 3216.270 ;
        RECT 868.930 3213.490 870.110 3214.670 ;
        RECT 868.930 3035.090 870.110 3036.270 ;
        RECT 868.930 3033.490 870.110 3034.670 ;
        RECT 868.930 2855.090 870.110 2856.270 ;
        RECT 868.930 2853.490 870.110 2854.670 ;
        RECT 868.930 2675.090 870.110 2676.270 ;
        RECT 868.930 2673.490 870.110 2674.670 ;
        RECT 868.930 2495.090 870.110 2496.270 ;
        RECT 868.930 2493.490 870.110 2494.670 ;
        RECT 868.930 2315.090 870.110 2316.270 ;
        RECT 868.930 2313.490 870.110 2314.670 ;
        RECT 868.930 2135.090 870.110 2136.270 ;
        RECT 868.930 2133.490 870.110 2134.670 ;
        RECT 868.930 1955.090 870.110 1956.270 ;
        RECT 868.930 1953.490 870.110 1954.670 ;
        RECT 868.930 1775.090 870.110 1776.270 ;
        RECT 868.930 1773.490 870.110 1774.670 ;
        RECT 868.930 1595.090 870.110 1596.270 ;
        RECT 868.930 1593.490 870.110 1594.670 ;
        RECT 868.930 1415.090 870.110 1416.270 ;
        RECT 868.930 1413.490 870.110 1414.670 ;
        RECT 868.930 1235.090 870.110 1236.270 ;
        RECT 868.930 1233.490 870.110 1234.670 ;
        RECT 868.930 1055.090 870.110 1056.270 ;
        RECT 868.930 1053.490 870.110 1054.670 ;
        RECT 868.930 875.090 870.110 876.270 ;
        RECT 868.930 873.490 870.110 874.670 ;
        RECT 868.930 695.090 870.110 696.270 ;
        RECT 868.930 693.490 870.110 694.670 ;
        RECT 868.930 515.090 870.110 516.270 ;
        RECT 868.930 513.490 870.110 514.670 ;
        RECT 868.930 335.090 870.110 336.270 ;
        RECT 868.930 333.490 870.110 334.670 ;
        RECT 868.930 155.090 870.110 156.270 ;
        RECT 868.930 153.490 870.110 154.670 ;
        RECT 868.930 -35.110 870.110 -33.930 ;
        RECT 868.930 -36.710 870.110 -35.530 ;
        RECT 1048.930 3555.210 1050.110 3556.390 ;
        RECT 1048.930 3553.610 1050.110 3554.790 ;
        RECT 1048.930 3395.090 1050.110 3396.270 ;
        RECT 1048.930 3393.490 1050.110 3394.670 ;
        RECT 1048.930 3215.090 1050.110 3216.270 ;
        RECT 1048.930 3213.490 1050.110 3214.670 ;
        RECT 1048.930 3035.090 1050.110 3036.270 ;
        RECT 1048.930 3033.490 1050.110 3034.670 ;
        RECT 1048.930 2855.090 1050.110 2856.270 ;
        RECT 1048.930 2853.490 1050.110 2854.670 ;
        RECT 1048.930 2675.090 1050.110 2676.270 ;
        RECT 1048.930 2673.490 1050.110 2674.670 ;
        RECT 1048.930 2495.090 1050.110 2496.270 ;
        RECT 1048.930 2493.490 1050.110 2494.670 ;
        RECT 1048.930 2315.090 1050.110 2316.270 ;
        RECT 1048.930 2313.490 1050.110 2314.670 ;
        RECT 1048.930 2135.090 1050.110 2136.270 ;
        RECT 1048.930 2133.490 1050.110 2134.670 ;
        RECT 1048.930 1955.090 1050.110 1956.270 ;
        RECT 1048.930 1953.490 1050.110 1954.670 ;
        RECT 1048.930 1775.090 1050.110 1776.270 ;
        RECT 1048.930 1773.490 1050.110 1774.670 ;
        RECT 1048.930 1595.090 1050.110 1596.270 ;
        RECT 1048.930 1593.490 1050.110 1594.670 ;
        RECT 1048.930 1415.090 1050.110 1416.270 ;
        RECT 1048.930 1413.490 1050.110 1414.670 ;
        RECT 1048.930 1235.090 1050.110 1236.270 ;
        RECT 1048.930 1233.490 1050.110 1234.670 ;
        RECT 1048.930 1055.090 1050.110 1056.270 ;
        RECT 1048.930 1053.490 1050.110 1054.670 ;
        RECT 1048.930 875.090 1050.110 876.270 ;
        RECT 1048.930 873.490 1050.110 874.670 ;
        RECT 1048.930 695.090 1050.110 696.270 ;
        RECT 1048.930 693.490 1050.110 694.670 ;
        RECT 1048.930 515.090 1050.110 516.270 ;
        RECT 1048.930 513.490 1050.110 514.670 ;
        RECT 1048.930 335.090 1050.110 336.270 ;
        RECT 1048.930 333.490 1050.110 334.670 ;
        RECT 1048.930 155.090 1050.110 156.270 ;
        RECT 1048.930 153.490 1050.110 154.670 ;
        RECT 1048.930 -35.110 1050.110 -33.930 ;
        RECT 1048.930 -36.710 1050.110 -35.530 ;
        RECT 1228.930 3555.210 1230.110 3556.390 ;
        RECT 1228.930 3553.610 1230.110 3554.790 ;
        RECT 1228.930 3395.090 1230.110 3396.270 ;
        RECT 1228.930 3393.490 1230.110 3394.670 ;
        RECT 1228.930 3215.090 1230.110 3216.270 ;
        RECT 1228.930 3213.490 1230.110 3214.670 ;
        RECT 1228.930 3035.090 1230.110 3036.270 ;
        RECT 1228.930 3033.490 1230.110 3034.670 ;
        RECT 1228.930 2855.090 1230.110 2856.270 ;
        RECT 1228.930 2853.490 1230.110 2854.670 ;
        RECT 1228.930 2675.090 1230.110 2676.270 ;
        RECT 1228.930 2673.490 1230.110 2674.670 ;
        RECT 1228.930 2495.090 1230.110 2496.270 ;
        RECT 1228.930 2493.490 1230.110 2494.670 ;
        RECT 1228.930 2315.090 1230.110 2316.270 ;
        RECT 1228.930 2313.490 1230.110 2314.670 ;
        RECT 1228.930 2135.090 1230.110 2136.270 ;
        RECT 1228.930 2133.490 1230.110 2134.670 ;
        RECT 1228.930 1955.090 1230.110 1956.270 ;
        RECT 1228.930 1953.490 1230.110 1954.670 ;
        RECT 1228.930 1775.090 1230.110 1776.270 ;
        RECT 1228.930 1773.490 1230.110 1774.670 ;
        RECT 1228.930 1595.090 1230.110 1596.270 ;
        RECT 1228.930 1593.490 1230.110 1594.670 ;
        RECT 1228.930 1415.090 1230.110 1416.270 ;
        RECT 1228.930 1413.490 1230.110 1414.670 ;
        RECT 1228.930 1235.090 1230.110 1236.270 ;
        RECT 1228.930 1233.490 1230.110 1234.670 ;
        RECT 1228.930 1055.090 1230.110 1056.270 ;
        RECT 1228.930 1053.490 1230.110 1054.670 ;
        RECT 1228.930 875.090 1230.110 876.270 ;
        RECT 1228.930 873.490 1230.110 874.670 ;
        RECT 1228.930 695.090 1230.110 696.270 ;
        RECT 1228.930 693.490 1230.110 694.670 ;
        RECT 1228.930 515.090 1230.110 516.270 ;
        RECT 1228.930 513.490 1230.110 514.670 ;
        RECT 1228.930 335.090 1230.110 336.270 ;
        RECT 1228.930 333.490 1230.110 334.670 ;
        RECT 1228.930 155.090 1230.110 156.270 ;
        RECT 1228.930 153.490 1230.110 154.670 ;
        RECT 1228.930 -35.110 1230.110 -33.930 ;
        RECT 1228.930 -36.710 1230.110 -35.530 ;
        RECT 1408.930 3555.210 1410.110 3556.390 ;
        RECT 1408.930 3553.610 1410.110 3554.790 ;
        RECT 1408.930 3395.090 1410.110 3396.270 ;
        RECT 1408.930 3393.490 1410.110 3394.670 ;
        RECT 1408.930 3215.090 1410.110 3216.270 ;
        RECT 1408.930 3213.490 1410.110 3214.670 ;
        RECT 1408.930 3035.090 1410.110 3036.270 ;
        RECT 1408.930 3033.490 1410.110 3034.670 ;
        RECT 1408.930 2855.090 1410.110 2856.270 ;
        RECT 1408.930 2853.490 1410.110 2854.670 ;
        RECT 1408.930 2675.090 1410.110 2676.270 ;
        RECT 1408.930 2673.490 1410.110 2674.670 ;
        RECT 1408.930 2495.090 1410.110 2496.270 ;
        RECT 1408.930 2493.490 1410.110 2494.670 ;
        RECT 1408.930 2315.090 1410.110 2316.270 ;
        RECT 1408.930 2313.490 1410.110 2314.670 ;
        RECT 1408.930 2135.090 1410.110 2136.270 ;
        RECT 1408.930 2133.490 1410.110 2134.670 ;
        RECT 1408.930 1955.090 1410.110 1956.270 ;
        RECT 1408.930 1953.490 1410.110 1954.670 ;
        RECT 1408.930 1775.090 1410.110 1776.270 ;
        RECT 1408.930 1773.490 1410.110 1774.670 ;
        RECT 1408.930 1595.090 1410.110 1596.270 ;
        RECT 1408.930 1593.490 1410.110 1594.670 ;
        RECT 1408.930 1415.090 1410.110 1416.270 ;
        RECT 1408.930 1413.490 1410.110 1414.670 ;
        RECT 1408.930 1235.090 1410.110 1236.270 ;
        RECT 1408.930 1233.490 1410.110 1234.670 ;
        RECT 1408.930 1055.090 1410.110 1056.270 ;
        RECT 1408.930 1053.490 1410.110 1054.670 ;
        RECT 1408.930 875.090 1410.110 876.270 ;
        RECT 1408.930 873.490 1410.110 874.670 ;
        RECT 1408.930 695.090 1410.110 696.270 ;
        RECT 1408.930 693.490 1410.110 694.670 ;
        RECT 1408.930 515.090 1410.110 516.270 ;
        RECT 1408.930 513.490 1410.110 514.670 ;
        RECT 1408.930 335.090 1410.110 336.270 ;
        RECT 1408.930 333.490 1410.110 334.670 ;
        RECT 1408.930 155.090 1410.110 156.270 ;
        RECT 1408.930 153.490 1410.110 154.670 ;
        RECT 1408.930 -35.110 1410.110 -33.930 ;
        RECT 1408.930 -36.710 1410.110 -35.530 ;
        RECT 1588.930 3555.210 1590.110 3556.390 ;
        RECT 1588.930 3553.610 1590.110 3554.790 ;
        RECT 1588.930 3395.090 1590.110 3396.270 ;
        RECT 1588.930 3393.490 1590.110 3394.670 ;
        RECT 1588.930 3215.090 1590.110 3216.270 ;
        RECT 1588.930 3213.490 1590.110 3214.670 ;
        RECT 1588.930 3035.090 1590.110 3036.270 ;
        RECT 1588.930 3033.490 1590.110 3034.670 ;
        RECT 1588.930 2855.090 1590.110 2856.270 ;
        RECT 1588.930 2853.490 1590.110 2854.670 ;
        RECT 1588.930 2675.090 1590.110 2676.270 ;
        RECT 1588.930 2673.490 1590.110 2674.670 ;
        RECT 1588.930 2495.090 1590.110 2496.270 ;
        RECT 1588.930 2493.490 1590.110 2494.670 ;
        RECT 1588.930 2315.090 1590.110 2316.270 ;
        RECT 1588.930 2313.490 1590.110 2314.670 ;
        RECT 1588.930 2135.090 1590.110 2136.270 ;
        RECT 1588.930 2133.490 1590.110 2134.670 ;
        RECT 1588.930 1955.090 1590.110 1956.270 ;
        RECT 1588.930 1953.490 1590.110 1954.670 ;
        RECT 1588.930 1775.090 1590.110 1776.270 ;
        RECT 1588.930 1773.490 1590.110 1774.670 ;
        RECT 1588.930 1595.090 1590.110 1596.270 ;
        RECT 1588.930 1593.490 1590.110 1594.670 ;
        RECT 1588.930 1415.090 1590.110 1416.270 ;
        RECT 1588.930 1413.490 1590.110 1414.670 ;
        RECT 1588.930 1235.090 1590.110 1236.270 ;
        RECT 1588.930 1233.490 1590.110 1234.670 ;
        RECT 1588.930 1055.090 1590.110 1056.270 ;
        RECT 1588.930 1053.490 1590.110 1054.670 ;
        RECT 1588.930 875.090 1590.110 876.270 ;
        RECT 1588.930 873.490 1590.110 874.670 ;
        RECT 1588.930 695.090 1590.110 696.270 ;
        RECT 1588.930 693.490 1590.110 694.670 ;
        RECT 1588.930 515.090 1590.110 516.270 ;
        RECT 1588.930 513.490 1590.110 514.670 ;
        RECT 1588.930 335.090 1590.110 336.270 ;
        RECT 1588.930 333.490 1590.110 334.670 ;
        RECT 1588.930 155.090 1590.110 156.270 ;
        RECT 1588.930 153.490 1590.110 154.670 ;
        RECT 1588.930 -35.110 1590.110 -33.930 ;
        RECT 1588.930 -36.710 1590.110 -35.530 ;
        RECT 1768.930 3555.210 1770.110 3556.390 ;
        RECT 1768.930 3553.610 1770.110 3554.790 ;
        RECT 1768.930 3395.090 1770.110 3396.270 ;
        RECT 1768.930 3393.490 1770.110 3394.670 ;
        RECT 1768.930 3215.090 1770.110 3216.270 ;
        RECT 1768.930 3213.490 1770.110 3214.670 ;
        RECT 1768.930 3035.090 1770.110 3036.270 ;
        RECT 1768.930 3033.490 1770.110 3034.670 ;
        RECT 1768.930 2855.090 1770.110 2856.270 ;
        RECT 1768.930 2853.490 1770.110 2854.670 ;
        RECT 1768.930 2675.090 1770.110 2676.270 ;
        RECT 1768.930 2673.490 1770.110 2674.670 ;
        RECT 1768.930 2495.090 1770.110 2496.270 ;
        RECT 1768.930 2493.490 1770.110 2494.670 ;
        RECT 1768.930 2315.090 1770.110 2316.270 ;
        RECT 1768.930 2313.490 1770.110 2314.670 ;
        RECT 1768.930 2135.090 1770.110 2136.270 ;
        RECT 1768.930 2133.490 1770.110 2134.670 ;
        RECT 1768.930 1955.090 1770.110 1956.270 ;
        RECT 1768.930 1953.490 1770.110 1954.670 ;
        RECT 1768.930 1775.090 1770.110 1776.270 ;
        RECT 1768.930 1773.490 1770.110 1774.670 ;
        RECT 1768.930 1595.090 1770.110 1596.270 ;
        RECT 1768.930 1593.490 1770.110 1594.670 ;
        RECT 1768.930 1415.090 1770.110 1416.270 ;
        RECT 1768.930 1413.490 1770.110 1414.670 ;
        RECT 1768.930 1235.090 1770.110 1236.270 ;
        RECT 1768.930 1233.490 1770.110 1234.670 ;
        RECT 1768.930 1055.090 1770.110 1056.270 ;
        RECT 1768.930 1053.490 1770.110 1054.670 ;
        RECT 1768.930 875.090 1770.110 876.270 ;
        RECT 1768.930 873.490 1770.110 874.670 ;
        RECT 1768.930 695.090 1770.110 696.270 ;
        RECT 1768.930 693.490 1770.110 694.670 ;
        RECT 1768.930 515.090 1770.110 516.270 ;
        RECT 1768.930 513.490 1770.110 514.670 ;
        RECT 1768.930 335.090 1770.110 336.270 ;
        RECT 1768.930 333.490 1770.110 334.670 ;
        RECT 1768.930 155.090 1770.110 156.270 ;
        RECT 1768.930 153.490 1770.110 154.670 ;
        RECT 1768.930 -35.110 1770.110 -33.930 ;
        RECT 1768.930 -36.710 1770.110 -35.530 ;
        RECT 1948.930 3555.210 1950.110 3556.390 ;
        RECT 1948.930 3553.610 1950.110 3554.790 ;
        RECT 1948.930 3395.090 1950.110 3396.270 ;
        RECT 1948.930 3393.490 1950.110 3394.670 ;
        RECT 1948.930 3215.090 1950.110 3216.270 ;
        RECT 1948.930 3213.490 1950.110 3214.670 ;
        RECT 1948.930 3035.090 1950.110 3036.270 ;
        RECT 1948.930 3033.490 1950.110 3034.670 ;
        RECT 1948.930 2855.090 1950.110 2856.270 ;
        RECT 1948.930 2853.490 1950.110 2854.670 ;
        RECT 1948.930 2675.090 1950.110 2676.270 ;
        RECT 1948.930 2673.490 1950.110 2674.670 ;
        RECT 1948.930 2495.090 1950.110 2496.270 ;
        RECT 1948.930 2493.490 1950.110 2494.670 ;
        RECT 1948.930 2315.090 1950.110 2316.270 ;
        RECT 1948.930 2313.490 1950.110 2314.670 ;
        RECT 1948.930 2135.090 1950.110 2136.270 ;
        RECT 1948.930 2133.490 1950.110 2134.670 ;
        RECT 1948.930 1955.090 1950.110 1956.270 ;
        RECT 1948.930 1953.490 1950.110 1954.670 ;
        RECT 1948.930 1775.090 1950.110 1776.270 ;
        RECT 1948.930 1773.490 1950.110 1774.670 ;
        RECT 1948.930 1595.090 1950.110 1596.270 ;
        RECT 1948.930 1593.490 1950.110 1594.670 ;
        RECT 1948.930 1415.090 1950.110 1416.270 ;
        RECT 1948.930 1413.490 1950.110 1414.670 ;
        RECT 1948.930 1235.090 1950.110 1236.270 ;
        RECT 1948.930 1233.490 1950.110 1234.670 ;
        RECT 1948.930 1055.090 1950.110 1056.270 ;
        RECT 1948.930 1053.490 1950.110 1054.670 ;
        RECT 1948.930 875.090 1950.110 876.270 ;
        RECT 1948.930 873.490 1950.110 874.670 ;
        RECT 1948.930 695.090 1950.110 696.270 ;
        RECT 1948.930 693.490 1950.110 694.670 ;
        RECT 1948.930 515.090 1950.110 516.270 ;
        RECT 1948.930 513.490 1950.110 514.670 ;
        RECT 1948.930 335.090 1950.110 336.270 ;
        RECT 1948.930 333.490 1950.110 334.670 ;
        RECT 1948.930 155.090 1950.110 156.270 ;
        RECT 1948.930 153.490 1950.110 154.670 ;
        RECT 1948.930 -35.110 1950.110 -33.930 ;
        RECT 1948.930 -36.710 1950.110 -35.530 ;
        RECT 2128.930 3555.210 2130.110 3556.390 ;
        RECT 2128.930 3553.610 2130.110 3554.790 ;
        RECT 2128.930 3395.090 2130.110 3396.270 ;
        RECT 2128.930 3393.490 2130.110 3394.670 ;
        RECT 2128.930 3215.090 2130.110 3216.270 ;
        RECT 2128.930 3213.490 2130.110 3214.670 ;
        RECT 2128.930 3035.090 2130.110 3036.270 ;
        RECT 2128.930 3033.490 2130.110 3034.670 ;
        RECT 2128.930 2855.090 2130.110 2856.270 ;
        RECT 2128.930 2853.490 2130.110 2854.670 ;
        RECT 2128.930 2675.090 2130.110 2676.270 ;
        RECT 2128.930 2673.490 2130.110 2674.670 ;
        RECT 2128.930 2495.090 2130.110 2496.270 ;
        RECT 2128.930 2493.490 2130.110 2494.670 ;
        RECT 2128.930 2315.090 2130.110 2316.270 ;
        RECT 2128.930 2313.490 2130.110 2314.670 ;
        RECT 2128.930 2135.090 2130.110 2136.270 ;
        RECT 2128.930 2133.490 2130.110 2134.670 ;
        RECT 2128.930 1955.090 2130.110 1956.270 ;
        RECT 2128.930 1953.490 2130.110 1954.670 ;
        RECT 2128.930 1775.090 2130.110 1776.270 ;
        RECT 2128.930 1773.490 2130.110 1774.670 ;
        RECT 2128.930 1595.090 2130.110 1596.270 ;
        RECT 2128.930 1593.490 2130.110 1594.670 ;
        RECT 2128.930 1415.090 2130.110 1416.270 ;
        RECT 2128.930 1413.490 2130.110 1414.670 ;
        RECT 2128.930 1235.090 2130.110 1236.270 ;
        RECT 2128.930 1233.490 2130.110 1234.670 ;
        RECT 2128.930 1055.090 2130.110 1056.270 ;
        RECT 2128.930 1053.490 2130.110 1054.670 ;
        RECT 2128.930 875.090 2130.110 876.270 ;
        RECT 2128.930 873.490 2130.110 874.670 ;
        RECT 2128.930 695.090 2130.110 696.270 ;
        RECT 2128.930 693.490 2130.110 694.670 ;
        RECT 2128.930 515.090 2130.110 516.270 ;
        RECT 2128.930 513.490 2130.110 514.670 ;
        RECT 2128.930 335.090 2130.110 336.270 ;
        RECT 2128.930 333.490 2130.110 334.670 ;
        RECT 2128.930 155.090 2130.110 156.270 ;
        RECT 2128.930 153.490 2130.110 154.670 ;
        RECT 2128.930 -35.110 2130.110 -33.930 ;
        RECT 2128.930 -36.710 2130.110 -35.530 ;
        RECT 2308.930 3555.210 2310.110 3556.390 ;
        RECT 2308.930 3553.610 2310.110 3554.790 ;
        RECT 2308.930 3395.090 2310.110 3396.270 ;
        RECT 2308.930 3393.490 2310.110 3394.670 ;
        RECT 2308.930 3215.090 2310.110 3216.270 ;
        RECT 2308.930 3213.490 2310.110 3214.670 ;
        RECT 2308.930 3035.090 2310.110 3036.270 ;
        RECT 2308.930 3033.490 2310.110 3034.670 ;
        RECT 2308.930 2855.090 2310.110 2856.270 ;
        RECT 2308.930 2853.490 2310.110 2854.670 ;
        RECT 2308.930 2675.090 2310.110 2676.270 ;
        RECT 2308.930 2673.490 2310.110 2674.670 ;
        RECT 2308.930 2495.090 2310.110 2496.270 ;
        RECT 2308.930 2493.490 2310.110 2494.670 ;
        RECT 2308.930 2315.090 2310.110 2316.270 ;
        RECT 2308.930 2313.490 2310.110 2314.670 ;
        RECT 2308.930 2135.090 2310.110 2136.270 ;
        RECT 2308.930 2133.490 2310.110 2134.670 ;
        RECT 2308.930 1955.090 2310.110 1956.270 ;
        RECT 2308.930 1953.490 2310.110 1954.670 ;
        RECT 2308.930 1775.090 2310.110 1776.270 ;
        RECT 2308.930 1773.490 2310.110 1774.670 ;
        RECT 2308.930 1595.090 2310.110 1596.270 ;
        RECT 2308.930 1593.490 2310.110 1594.670 ;
        RECT 2308.930 1415.090 2310.110 1416.270 ;
        RECT 2308.930 1413.490 2310.110 1414.670 ;
        RECT 2308.930 1235.090 2310.110 1236.270 ;
        RECT 2308.930 1233.490 2310.110 1234.670 ;
        RECT 2308.930 1055.090 2310.110 1056.270 ;
        RECT 2308.930 1053.490 2310.110 1054.670 ;
        RECT 2308.930 875.090 2310.110 876.270 ;
        RECT 2308.930 873.490 2310.110 874.670 ;
        RECT 2308.930 695.090 2310.110 696.270 ;
        RECT 2308.930 693.490 2310.110 694.670 ;
        RECT 2308.930 515.090 2310.110 516.270 ;
        RECT 2308.930 513.490 2310.110 514.670 ;
        RECT 2308.930 335.090 2310.110 336.270 ;
        RECT 2308.930 333.490 2310.110 334.670 ;
        RECT 2308.930 155.090 2310.110 156.270 ;
        RECT 2308.930 153.490 2310.110 154.670 ;
        RECT 2308.930 -35.110 2310.110 -33.930 ;
        RECT 2308.930 -36.710 2310.110 -35.530 ;
        RECT 2488.930 3555.210 2490.110 3556.390 ;
        RECT 2488.930 3553.610 2490.110 3554.790 ;
        RECT 2488.930 3395.090 2490.110 3396.270 ;
        RECT 2488.930 3393.490 2490.110 3394.670 ;
        RECT 2488.930 3215.090 2490.110 3216.270 ;
        RECT 2488.930 3213.490 2490.110 3214.670 ;
        RECT 2488.930 3035.090 2490.110 3036.270 ;
        RECT 2488.930 3033.490 2490.110 3034.670 ;
        RECT 2488.930 2855.090 2490.110 2856.270 ;
        RECT 2488.930 2853.490 2490.110 2854.670 ;
        RECT 2488.930 2675.090 2490.110 2676.270 ;
        RECT 2488.930 2673.490 2490.110 2674.670 ;
        RECT 2488.930 2495.090 2490.110 2496.270 ;
        RECT 2488.930 2493.490 2490.110 2494.670 ;
        RECT 2488.930 2315.090 2490.110 2316.270 ;
        RECT 2488.930 2313.490 2490.110 2314.670 ;
        RECT 2488.930 2135.090 2490.110 2136.270 ;
        RECT 2488.930 2133.490 2490.110 2134.670 ;
        RECT 2488.930 1955.090 2490.110 1956.270 ;
        RECT 2488.930 1953.490 2490.110 1954.670 ;
        RECT 2488.930 1775.090 2490.110 1776.270 ;
        RECT 2488.930 1773.490 2490.110 1774.670 ;
        RECT 2488.930 1595.090 2490.110 1596.270 ;
        RECT 2488.930 1593.490 2490.110 1594.670 ;
        RECT 2488.930 1415.090 2490.110 1416.270 ;
        RECT 2488.930 1413.490 2490.110 1414.670 ;
        RECT 2488.930 1235.090 2490.110 1236.270 ;
        RECT 2488.930 1233.490 2490.110 1234.670 ;
        RECT 2488.930 1055.090 2490.110 1056.270 ;
        RECT 2488.930 1053.490 2490.110 1054.670 ;
        RECT 2488.930 875.090 2490.110 876.270 ;
        RECT 2488.930 873.490 2490.110 874.670 ;
        RECT 2488.930 695.090 2490.110 696.270 ;
        RECT 2488.930 693.490 2490.110 694.670 ;
        RECT 2488.930 515.090 2490.110 516.270 ;
        RECT 2488.930 513.490 2490.110 514.670 ;
        RECT 2488.930 335.090 2490.110 336.270 ;
        RECT 2488.930 333.490 2490.110 334.670 ;
        RECT 2488.930 155.090 2490.110 156.270 ;
        RECT 2488.930 153.490 2490.110 154.670 ;
        RECT 2488.930 -35.110 2490.110 -33.930 ;
        RECT 2488.930 -36.710 2490.110 -35.530 ;
        RECT 2668.930 3555.210 2670.110 3556.390 ;
        RECT 2668.930 3553.610 2670.110 3554.790 ;
        RECT 2668.930 3395.090 2670.110 3396.270 ;
        RECT 2668.930 3393.490 2670.110 3394.670 ;
        RECT 2668.930 3215.090 2670.110 3216.270 ;
        RECT 2668.930 3213.490 2670.110 3214.670 ;
        RECT 2668.930 3035.090 2670.110 3036.270 ;
        RECT 2668.930 3033.490 2670.110 3034.670 ;
        RECT 2668.930 2855.090 2670.110 2856.270 ;
        RECT 2668.930 2853.490 2670.110 2854.670 ;
        RECT 2668.930 2675.090 2670.110 2676.270 ;
        RECT 2668.930 2673.490 2670.110 2674.670 ;
        RECT 2668.930 2495.090 2670.110 2496.270 ;
        RECT 2668.930 2493.490 2670.110 2494.670 ;
        RECT 2668.930 2315.090 2670.110 2316.270 ;
        RECT 2668.930 2313.490 2670.110 2314.670 ;
        RECT 2668.930 2135.090 2670.110 2136.270 ;
        RECT 2668.930 2133.490 2670.110 2134.670 ;
        RECT 2668.930 1955.090 2670.110 1956.270 ;
        RECT 2668.930 1953.490 2670.110 1954.670 ;
        RECT 2668.930 1775.090 2670.110 1776.270 ;
        RECT 2668.930 1773.490 2670.110 1774.670 ;
        RECT 2668.930 1595.090 2670.110 1596.270 ;
        RECT 2668.930 1593.490 2670.110 1594.670 ;
        RECT 2668.930 1415.090 2670.110 1416.270 ;
        RECT 2668.930 1413.490 2670.110 1414.670 ;
        RECT 2668.930 1235.090 2670.110 1236.270 ;
        RECT 2668.930 1233.490 2670.110 1234.670 ;
        RECT 2668.930 1055.090 2670.110 1056.270 ;
        RECT 2668.930 1053.490 2670.110 1054.670 ;
        RECT 2668.930 875.090 2670.110 876.270 ;
        RECT 2668.930 873.490 2670.110 874.670 ;
        RECT 2668.930 695.090 2670.110 696.270 ;
        RECT 2668.930 693.490 2670.110 694.670 ;
        RECT 2668.930 515.090 2670.110 516.270 ;
        RECT 2668.930 513.490 2670.110 514.670 ;
        RECT 2668.930 335.090 2670.110 336.270 ;
        RECT 2668.930 333.490 2670.110 334.670 ;
        RECT 2668.930 155.090 2670.110 156.270 ;
        RECT 2668.930 153.490 2670.110 154.670 ;
        RECT 2668.930 -35.110 2670.110 -33.930 ;
        RECT 2668.930 -36.710 2670.110 -35.530 ;
        RECT 2848.930 3555.210 2850.110 3556.390 ;
        RECT 2848.930 3553.610 2850.110 3554.790 ;
        RECT 2848.930 3395.090 2850.110 3396.270 ;
        RECT 2848.930 3393.490 2850.110 3394.670 ;
        RECT 2848.930 3215.090 2850.110 3216.270 ;
        RECT 2848.930 3213.490 2850.110 3214.670 ;
        RECT 2848.930 3035.090 2850.110 3036.270 ;
        RECT 2848.930 3033.490 2850.110 3034.670 ;
        RECT 2848.930 2855.090 2850.110 2856.270 ;
        RECT 2848.930 2853.490 2850.110 2854.670 ;
        RECT 2848.930 2675.090 2850.110 2676.270 ;
        RECT 2848.930 2673.490 2850.110 2674.670 ;
        RECT 2848.930 2495.090 2850.110 2496.270 ;
        RECT 2848.930 2493.490 2850.110 2494.670 ;
        RECT 2848.930 2315.090 2850.110 2316.270 ;
        RECT 2848.930 2313.490 2850.110 2314.670 ;
        RECT 2848.930 2135.090 2850.110 2136.270 ;
        RECT 2848.930 2133.490 2850.110 2134.670 ;
        RECT 2848.930 1955.090 2850.110 1956.270 ;
        RECT 2848.930 1953.490 2850.110 1954.670 ;
        RECT 2848.930 1775.090 2850.110 1776.270 ;
        RECT 2848.930 1773.490 2850.110 1774.670 ;
        RECT 2848.930 1595.090 2850.110 1596.270 ;
        RECT 2848.930 1593.490 2850.110 1594.670 ;
        RECT 2848.930 1415.090 2850.110 1416.270 ;
        RECT 2848.930 1413.490 2850.110 1414.670 ;
        RECT 2848.930 1235.090 2850.110 1236.270 ;
        RECT 2848.930 1233.490 2850.110 1234.670 ;
        RECT 2848.930 1055.090 2850.110 1056.270 ;
        RECT 2848.930 1053.490 2850.110 1054.670 ;
        RECT 2848.930 875.090 2850.110 876.270 ;
        RECT 2848.930 873.490 2850.110 874.670 ;
        RECT 2848.930 695.090 2850.110 696.270 ;
        RECT 2848.930 693.490 2850.110 694.670 ;
        RECT 2848.930 515.090 2850.110 516.270 ;
        RECT 2848.930 513.490 2850.110 514.670 ;
        RECT 2848.930 335.090 2850.110 336.270 ;
        RECT 2848.930 333.490 2850.110 334.670 ;
        RECT 2848.930 155.090 2850.110 156.270 ;
        RECT 2848.930 153.490 2850.110 154.670 ;
        RECT 2848.930 -35.110 2850.110 -33.930 ;
        RECT 2848.930 -36.710 2850.110 -35.530 ;
        RECT 2959.710 3555.210 2960.890 3556.390 ;
        RECT 2959.710 3553.610 2960.890 3554.790 ;
        RECT 2959.710 3395.090 2960.890 3396.270 ;
        RECT 2959.710 3393.490 2960.890 3394.670 ;
        RECT 2959.710 3215.090 2960.890 3216.270 ;
        RECT 2959.710 3213.490 2960.890 3214.670 ;
        RECT 2959.710 3035.090 2960.890 3036.270 ;
        RECT 2959.710 3033.490 2960.890 3034.670 ;
        RECT 2959.710 2855.090 2960.890 2856.270 ;
        RECT 2959.710 2853.490 2960.890 2854.670 ;
        RECT 2959.710 2675.090 2960.890 2676.270 ;
        RECT 2959.710 2673.490 2960.890 2674.670 ;
        RECT 2959.710 2495.090 2960.890 2496.270 ;
        RECT 2959.710 2493.490 2960.890 2494.670 ;
        RECT 2959.710 2315.090 2960.890 2316.270 ;
        RECT 2959.710 2313.490 2960.890 2314.670 ;
        RECT 2959.710 2135.090 2960.890 2136.270 ;
        RECT 2959.710 2133.490 2960.890 2134.670 ;
        RECT 2959.710 1955.090 2960.890 1956.270 ;
        RECT 2959.710 1953.490 2960.890 1954.670 ;
        RECT 2959.710 1775.090 2960.890 1776.270 ;
        RECT 2959.710 1773.490 2960.890 1774.670 ;
        RECT 2959.710 1595.090 2960.890 1596.270 ;
        RECT 2959.710 1593.490 2960.890 1594.670 ;
        RECT 2959.710 1415.090 2960.890 1416.270 ;
        RECT 2959.710 1413.490 2960.890 1414.670 ;
        RECT 2959.710 1235.090 2960.890 1236.270 ;
        RECT 2959.710 1233.490 2960.890 1234.670 ;
        RECT 2959.710 1055.090 2960.890 1056.270 ;
        RECT 2959.710 1053.490 2960.890 1054.670 ;
        RECT 2959.710 875.090 2960.890 876.270 ;
        RECT 2959.710 873.490 2960.890 874.670 ;
        RECT 2959.710 695.090 2960.890 696.270 ;
        RECT 2959.710 693.490 2960.890 694.670 ;
        RECT 2959.710 515.090 2960.890 516.270 ;
        RECT 2959.710 513.490 2960.890 514.670 ;
        RECT 2959.710 335.090 2960.890 336.270 ;
        RECT 2959.710 333.490 2960.890 334.670 ;
        RECT 2959.710 155.090 2960.890 156.270 ;
        RECT 2959.710 153.490 2960.890 154.670 ;
        RECT 2959.710 -35.110 2960.890 -33.930 ;
        RECT 2959.710 -36.710 2960.890 -35.530 ;
      LAYER met5 ;
        RECT -42.180 3556.500 -39.180 3556.510 ;
        RECT 148.020 3556.500 151.020 3556.510 ;
        RECT 328.020 3556.500 331.020 3556.510 ;
        RECT 508.020 3556.500 511.020 3556.510 ;
        RECT 688.020 3556.500 691.020 3556.510 ;
        RECT 868.020 3556.500 871.020 3556.510 ;
        RECT 1048.020 3556.500 1051.020 3556.510 ;
        RECT 1228.020 3556.500 1231.020 3556.510 ;
        RECT 1408.020 3556.500 1411.020 3556.510 ;
        RECT 1588.020 3556.500 1591.020 3556.510 ;
        RECT 1768.020 3556.500 1771.020 3556.510 ;
        RECT 1948.020 3556.500 1951.020 3556.510 ;
        RECT 2128.020 3556.500 2131.020 3556.510 ;
        RECT 2308.020 3556.500 2311.020 3556.510 ;
        RECT 2488.020 3556.500 2491.020 3556.510 ;
        RECT 2668.020 3556.500 2671.020 3556.510 ;
        RECT 2848.020 3556.500 2851.020 3556.510 ;
        RECT 2958.800 3556.500 2961.800 3556.510 ;
        RECT -42.180 3553.500 2961.800 3556.500 ;
        RECT -42.180 3553.490 -39.180 3553.500 ;
        RECT 148.020 3553.490 151.020 3553.500 ;
        RECT 328.020 3553.490 331.020 3553.500 ;
        RECT 508.020 3553.490 511.020 3553.500 ;
        RECT 688.020 3553.490 691.020 3553.500 ;
        RECT 868.020 3553.490 871.020 3553.500 ;
        RECT 1048.020 3553.490 1051.020 3553.500 ;
        RECT 1228.020 3553.490 1231.020 3553.500 ;
        RECT 1408.020 3553.490 1411.020 3553.500 ;
        RECT 1588.020 3553.490 1591.020 3553.500 ;
        RECT 1768.020 3553.490 1771.020 3553.500 ;
        RECT 1948.020 3553.490 1951.020 3553.500 ;
        RECT 2128.020 3553.490 2131.020 3553.500 ;
        RECT 2308.020 3553.490 2311.020 3553.500 ;
        RECT 2488.020 3553.490 2491.020 3553.500 ;
        RECT 2668.020 3553.490 2671.020 3553.500 ;
        RECT 2848.020 3553.490 2851.020 3553.500 ;
        RECT 2958.800 3553.490 2961.800 3553.500 ;
        RECT -42.180 3396.380 -39.180 3396.390 ;
        RECT 148.020 3396.380 151.020 3396.390 ;
        RECT 328.020 3396.380 331.020 3396.390 ;
        RECT 508.020 3396.380 511.020 3396.390 ;
        RECT 688.020 3396.380 691.020 3396.390 ;
        RECT 868.020 3396.380 871.020 3396.390 ;
        RECT 1048.020 3396.380 1051.020 3396.390 ;
        RECT 1228.020 3396.380 1231.020 3396.390 ;
        RECT 1408.020 3396.380 1411.020 3396.390 ;
        RECT 1588.020 3396.380 1591.020 3396.390 ;
        RECT 1768.020 3396.380 1771.020 3396.390 ;
        RECT 1948.020 3396.380 1951.020 3396.390 ;
        RECT 2128.020 3396.380 2131.020 3396.390 ;
        RECT 2308.020 3396.380 2311.020 3396.390 ;
        RECT 2488.020 3396.380 2491.020 3396.390 ;
        RECT 2668.020 3396.380 2671.020 3396.390 ;
        RECT 2848.020 3396.380 2851.020 3396.390 ;
        RECT 2958.800 3396.380 2961.800 3396.390 ;
        RECT -42.180 3393.380 2961.800 3396.380 ;
        RECT -42.180 3393.370 -39.180 3393.380 ;
        RECT 148.020 3393.370 151.020 3393.380 ;
        RECT 328.020 3393.370 331.020 3393.380 ;
        RECT 508.020 3393.370 511.020 3393.380 ;
        RECT 688.020 3393.370 691.020 3393.380 ;
        RECT 868.020 3393.370 871.020 3393.380 ;
        RECT 1048.020 3393.370 1051.020 3393.380 ;
        RECT 1228.020 3393.370 1231.020 3393.380 ;
        RECT 1408.020 3393.370 1411.020 3393.380 ;
        RECT 1588.020 3393.370 1591.020 3393.380 ;
        RECT 1768.020 3393.370 1771.020 3393.380 ;
        RECT 1948.020 3393.370 1951.020 3393.380 ;
        RECT 2128.020 3393.370 2131.020 3393.380 ;
        RECT 2308.020 3393.370 2311.020 3393.380 ;
        RECT 2488.020 3393.370 2491.020 3393.380 ;
        RECT 2668.020 3393.370 2671.020 3393.380 ;
        RECT 2848.020 3393.370 2851.020 3393.380 ;
        RECT 2958.800 3393.370 2961.800 3393.380 ;
        RECT -42.180 3216.380 -39.180 3216.390 ;
        RECT 148.020 3216.380 151.020 3216.390 ;
        RECT 328.020 3216.380 331.020 3216.390 ;
        RECT 508.020 3216.380 511.020 3216.390 ;
        RECT 688.020 3216.380 691.020 3216.390 ;
        RECT 868.020 3216.380 871.020 3216.390 ;
        RECT 1048.020 3216.380 1051.020 3216.390 ;
        RECT 1228.020 3216.380 1231.020 3216.390 ;
        RECT 1408.020 3216.380 1411.020 3216.390 ;
        RECT 1588.020 3216.380 1591.020 3216.390 ;
        RECT 1768.020 3216.380 1771.020 3216.390 ;
        RECT 1948.020 3216.380 1951.020 3216.390 ;
        RECT 2128.020 3216.380 2131.020 3216.390 ;
        RECT 2308.020 3216.380 2311.020 3216.390 ;
        RECT 2488.020 3216.380 2491.020 3216.390 ;
        RECT 2668.020 3216.380 2671.020 3216.390 ;
        RECT 2848.020 3216.380 2851.020 3216.390 ;
        RECT 2958.800 3216.380 2961.800 3216.390 ;
        RECT -42.180 3213.380 2961.800 3216.380 ;
        RECT -42.180 3213.370 -39.180 3213.380 ;
        RECT 148.020 3213.370 151.020 3213.380 ;
        RECT 328.020 3213.370 331.020 3213.380 ;
        RECT 508.020 3213.370 511.020 3213.380 ;
        RECT 688.020 3213.370 691.020 3213.380 ;
        RECT 868.020 3213.370 871.020 3213.380 ;
        RECT 1048.020 3213.370 1051.020 3213.380 ;
        RECT 1228.020 3213.370 1231.020 3213.380 ;
        RECT 1408.020 3213.370 1411.020 3213.380 ;
        RECT 1588.020 3213.370 1591.020 3213.380 ;
        RECT 1768.020 3213.370 1771.020 3213.380 ;
        RECT 1948.020 3213.370 1951.020 3213.380 ;
        RECT 2128.020 3213.370 2131.020 3213.380 ;
        RECT 2308.020 3213.370 2311.020 3213.380 ;
        RECT 2488.020 3213.370 2491.020 3213.380 ;
        RECT 2668.020 3213.370 2671.020 3213.380 ;
        RECT 2848.020 3213.370 2851.020 3213.380 ;
        RECT 2958.800 3213.370 2961.800 3213.380 ;
        RECT -42.180 3036.380 -39.180 3036.390 ;
        RECT 148.020 3036.380 151.020 3036.390 ;
        RECT 328.020 3036.380 331.020 3036.390 ;
        RECT 508.020 3036.380 511.020 3036.390 ;
        RECT 688.020 3036.380 691.020 3036.390 ;
        RECT 868.020 3036.380 871.020 3036.390 ;
        RECT 1048.020 3036.380 1051.020 3036.390 ;
        RECT 1228.020 3036.380 1231.020 3036.390 ;
        RECT 1408.020 3036.380 1411.020 3036.390 ;
        RECT 1588.020 3036.380 1591.020 3036.390 ;
        RECT 1768.020 3036.380 1771.020 3036.390 ;
        RECT 1948.020 3036.380 1951.020 3036.390 ;
        RECT 2128.020 3036.380 2131.020 3036.390 ;
        RECT 2308.020 3036.380 2311.020 3036.390 ;
        RECT 2488.020 3036.380 2491.020 3036.390 ;
        RECT 2668.020 3036.380 2671.020 3036.390 ;
        RECT 2848.020 3036.380 2851.020 3036.390 ;
        RECT 2958.800 3036.380 2961.800 3036.390 ;
        RECT -42.180 3033.380 2961.800 3036.380 ;
        RECT -42.180 3033.370 -39.180 3033.380 ;
        RECT 148.020 3033.370 151.020 3033.380 ;
        RECT 328.020 3033.370 331.020 3033.380 ;
        RECT 508.020 3033.370 511.020 3033.380 ;
        RECT 688.020 3033.370 691.020 3033.380 ;
        RECT 868.020 3033.370 871.020 3033.380 ;
        RECT 1048.020 3033.370 1051.020 3033.380 ;
        RECT 1228.020 3033.370 1231.020 3033.380 ;
        RECT 1408.020 3033.370 1411.020 3033.380 ;
        RECT 1588.020 3033.370 1591.020 3033.380 ;
        RECT 1768.020 3033.370 1771.020 3033.380 ;
        RECT 1948.020 3033.370 1951.020 3033.380 ;
        RECT 2128.020 3033.370 2131.020 3033.380 ;
        RECT 2308.020 3033.370 2311.020 3033.380 ;
        RECT 2488.020 3033.370 2491.020 3033.380 ;
        RECT 2668.020 3033.370 2671.020 3033.380 ;
        RECT 2848.020 3033.370 2851.020 3033.380 ;
        RECT 2958.800 3033.370 2961.800 3033.380 ;
        RECT -42.180 2856.380 -39.180 2856.390 ;
        RECT 148.020 2856.380 151.020 2856.390 ;
        RECT 328.020 2856.380 331.020 2856.390 ;
        RECT 508.020 2856.380 511.020 2856.390 ;
        RECT 688.020 2856.380 691.020 2856.390 ;
        RECT 868.020 2856.380 871.020 2856.390 ;
        RECT 1048.020 2856.380 1051.020 2856.390 ;
        RECT 1228.020 2856.380 1231.020 2856.390 ;
        RECT 1408.020 2856.380 1411.020 2856.390 ;
        RECT 1588.020 2856.380 1591.020 2856.390 ;
        RECT 1768.020 2856.380 1771.020 2856.390 ;
        RECT 1948.020 2856.380 1951.020 2856.390 ;
        RECT 2128.020 2856.380 2131.020 2856.390 ;
        RECT 2308.020 2856.380 2311.020 2856.390 ;
        RECT 2488.020 2856.380 2491.020 2856.390 ;
        RECT 2668.020 2856.380 2671.020 2856.390 ;
        RECT 2848.020 2856.380 2851.020 2856.390 ;
        RECT 2958.800 2856.380 2961.800 2856.390 ;
        RECT -42.180 2853.380 2961.800 2856.380 ;
        RECT -42.180 2853.370 -39.180 2853.380 ;
        RECT 148.020 2853.370 151.020 2853.380 ;
        RECT 328.020 2853.370 331.020 2853.380 ;
        RECT 508.020 2853.370 511.020 2853.380 ;
        RECT 688.020 2853.370 691.020 2853.380 ;
        RECT 868.020 2853.370 871.020 2853.380 ;
        RECT 1048.020 2853.370 1051.020 2853.380 ;
        RECT 1228.020 2853.370 1231.020 2853.380 ;
        RECT 1408.020 2853.370 1411.020 2853.380 ;
        RECT 1588.020 2853.370 1591.020 2853.380 ;
        RECT 1768.020 2853.370 1771.020 2853.380 ;
        RECT 1948.020 2853.370 1951.020 2853.380 ;
        RECT 2128.020 2853.370 2131.020 2853.380 ;
        RECT 2308.020 2853.370 2311.020 2853.380 ;
        RECT 2488.020 2853.370 2491.020 2853.380 ;
        RECT 2668.020 2853.370 2671.020 2853.380 ;
        RECT 2848.020 2853.370 2851.020 2853.380 ;
        RECT 2958.800 2853.370 2961.800 2853.380 ;
        RECT -42.180 2676.380 -39.180 2676.390 ;
        RECT 148.020 2676.380 151.020 2676.390 ;
        RECT 328.020 2676.380 331.020 2676.390 ;
        RECT 508.020 2676.380 511.020 2676.390 ;
        RECT 688.020 2676.380 691.020 2676.390 ;
        RECT 868.020 2676.380 871.020 2676.390 ;
        RECT 1048.020 2676.380 1051.020 2676.390 ;
        RECT 1228.020 2676.380 1231.020 2676.390 ;
        RECT 1408.020 2676.380 1411.020 2676.390 ;
        RECT 1588.020 2676.380 1591.020 2676.390 ;
        RECT 1768.020 2676.380 1771.020 2676.390 ;
        RECT 1948.020 2676.380 1951.020 2676.390 ;
        RECT 2128.020 2676.380 2131.020 2676.390 ;
        RECT 2308.020 2676.380 2311.020 2676.390 ;
        RECT 2488.020 2676.380 2491.020 2676.390 ;
        RECT 2668.020 2676.380 2671.020 2676.390 ;
        RECT 2848.020 2676.380 2851.020 2676.390 ;
        RECT 2958.800 2676.380 2961.800 2676.390 ;
        RECT -42.180 2673.380 2961.800 2676.380 ;
        RECT -42.180 2673.370 -39.180 2673.380 ;
        RECT 148.020 2673.370 151.020 2673.380 ;
        RECT 328.020 2673.370 331.020 2673.380 ;
        RECT 508.020 2673.370 511.020 2673.380 ;
        RECT 688.020 2673.370 691.020 2673.380 ;
        RECT 868.020 2673.370 871.020 2673.380 ;
        RECT 1048.020 2673.370 1051.020 2673.380 ;
        RECT 1228.020 2673.370 1231.020 2673.380 ;
        RECT 1408.020 2673.370 1411.020 2673.380 ;
        RECT 1588.020 2673.370 1591.020 2673.380 ;
        RECT 1768.020 2673.370 1771.020 2673.380 ;
        RECT 1948.020 2673.370 1951.020 2673.380 ;
        RECT 2128.020 2673.370 2131.020 2673.380 ;
        RECT 2308.020 2673.370 2311.020 2673.380 ;
        RECT 2488.020 2673.370 2491.020 2673.380 ;
        RECT 2668.020 2673.370 2671.020 2673.380 ;
        RECT 2848.020 2673.370 2851.020 2673.380 ;
        RECT 2958.800 2673.370 2961.800 2673.380 ;
        RECT -42.180 2496.380 -39.180 2496.390 ;
        RECT 148.020 2496.380 151.020 2496.390 ;
        RECT 328.020 2496.380 331.020 2496.390 ;
        RECT 508.020 2496.380 511.020 2496.390 ;
        RECT 688.020 2496.380 691.020 2496.390 ;
        RECT 868.020 2496.380 871.020 2496.390 ;
        RECT 1048.020 2496.380 1051.020 2496.390 ;
        RECT 1228.020 2496.380 1231.020 2496.390 ;
        RECT 1408.020 2496.380 1411.020 2496.390 ;
        RECT 1588.020 2496.380 1591.020 2496.390 ;
        RECT 1768.020 2496.380 1771.020 2496.390 ;
        RECT 1948.020 2496.380 1951.020 2496.390 ;
        RECT 2128.020 2496.380 2131.020 2496.390 ;
        RECT 2308.020 2496.380 2311.020 2496.390 ;
        RECT 2488.020 2496.380 2491.020 2496.390 ;
        RECT 2668.020 2496.380 2671.020 2496.390 ;
        RECT 2848.020 2496.380 2851.020 2496.390 ;
        RECT 2958.800 2496.380 2961.800 2496.390 ;
        RECT -42.180 2493.380 2961.800 2496.380 ;
        RECT -42.180 2493.370 -39.180 2493.380 ;
        RECT 148.020 2493.370 151.020 2493.380 ;
        RECT 328.020 2493.370 331.020 2493.380 ;
        RECT 508.020 2493.370 511.020 2493.380 ;
        RECT 688.020 2493.370 691.020 2493.380 ;
        RECT 868.020 2493.370 871.020 2493.380 ;
        RECT 1048.020 2493.370 1051.020 2493.380 ;
        RECT 1228.020 2493.370 1231.020 2493.380 ;
        RECT 1408.020 2493.370 1411.020 2493.380 ;
        RECT 1588.020 2493.370 1591.020 2493.380 ;
        RECT 1768.020 2493.370 1771.020 2493.380 ;
        RECT 1948.020 2493.370 1951.020 2493.380 ;
        RECT 2128.020 2493.370 2131.020 2493.380 ;
        RECT 2308.020 2493.370 2311.020 2493.380 ;
        RECT 2488.020 2493.370 2491.020 2493.380 ;
        RECT 2668.020 2493.370 2671.020 2493.380 ;
        RECT 2848.020 2493.370 2851.020 2493.380 ;
        RECT 2958.800 2493.370 2961.800 2493.380 ;
        RECT -42.180 2316.380 -39.180 2316.390 ;
        RECT 148.020 2316.380 151.020 2316.390 ;
        RECT 328.020 2316.380 331.020 2316.390 ;
        RECT 508.020 2316.380 511.020 2316.390 ;
        RECT 688.020 2316.380 691.020 2316.390 ;
        RECT 868.020 2316.380 871.020 2316.390 ;
        RECT 1048.020 2316.380 1051.020 2316.390 ;
        RECT 1228.020 2316.380 1231.020 2316.390 ;
        RECT 1408.020 2316.380 1411.020 2316.390 ;
        RECT 1588.020 2316.380 1591.020 2316.390 ;
        RECT 1768.020 2316.380 1771.020 2316.390 ;
        RECT 1948.020 2316.380 1951.020 2316.390 ;
        RECT 2128.020 2316.380 2131.020 2316.390 ;
        RECT 2308.020 2316.380 2311.020 2316.390 ;
        RECT 2488.020 2316.380 2491.020 2316.390 ;
        RECT 2668.020 2316.380 2671.020 2316.390 ;
        RECT 2848.020 2316.380 2851.020 2316.390 ;
        RECT 2958.800 2316.380 2961.800 2316.390 ;
        RECT -42.180 2313.380 2961.800 2316.380 ;
        RECT -42.180 2313.370 -39.180 2313.380 ;
        RECT 148.020 2313.370 151.020 2313.380 ;
        RECT 328.020 2313.370 331.020 2313.380 ;
        RECT 508.020 2313.370 511.020 2313.380 ;
        RECT 688.020 2313.370 691.020 2313.380 ;
        RECT 868.020 2313.370 871.020 2313.380 ;
        RECT 1048.020 2313.370 1051.020 2313.380 ;
        RECT 1228.020 2313.370 1231.020 2313.380 ;
        RECT 1408.020 2313.370 1411.020 2313.380 ;
        RECT 1588.020 2313.370 1591.020 2313.380 ;
        RECT 1768.020 2313.370 1771.020 2313.380 ;
        RECT 1948.020 2313.370 1951.020 2313.380 ;
        RECT 2128.020 2313.370 2131.020 2313.380 ;
        RECT 2308.020 2313.370 2311.020 2313.380 ;
        RECT 2488.020 2313.370 2491.020 2313.380 ;
        RECT 2668.020 2313.370 2671.020 2313.380 ;
        RECT 2848.020 2313.370 2851.020 2313.380 ;
        RECT 2958.800 2313.370 2961.800 2313.380 ;
        RECT -42.180 2136.380 -39.180 2136.390 ;
        RECT 148.020 2136.380 151.020 2136.390 ;
        RECT 328.020 2136.380 331.020 2136.390 ;
        RECT 508.020 2136.380 511.020 2136.390 ;
        RECT 688.020 2136.380 691.020 2136.390 ;
        RECT 868.020 2136.380 871.020 2136.390 ;
        RECT 1048.020 2136.380 1051.020 2136.390 ;
        RECT 1228.020 2136.380 1231.020 2136.390 ;
        RECT 1408.020 2136.380 1411.020 2136.390 ;
        RECT 1588.020 2136.380 1591.020 2136.390 ;
        RECT 1768.020 2136.380 1771.020 2136.390 ;
        RECT 1948.020 2136.380 1951.020 2136.390 ;
        RECT 2128.020 2136.380 2131.020 2136.390 ;
        RECT 2308.020 2136.380 2311.020 2136.390 ;
        RECT 2488.020 2136.380 2491.020 2136.390 ;
        RECT 2668.020 2136.380 2671.020 2136.390 ;
        RECT 2848.020 2136.380 2851.020 2136.390 ;
        RECT 2958.800 2136.380 2961.800 2136.390 ;
        RECT -42.180 2133.380 2961.800 2136.380 ;
        RECT -42.180 2133.370 -39.180 2133.380 ;
        RECT 148.020 2133.370 151.020 2133.380 ;
        RECT 328.020 2133.370 331.020 2133.380 ;
        RECT 508.020 2133.370 511.020 2133.380 ;
        RECT 688.020 2133.370 691.020 2133.380 ;
        RECT 868.020 2133.370 871.020 2133.380 ;
        RECT 1048.020 2133.370 1051.020 2133.380 ;
        RECT 1228.020 2133.370 1231.020 2133.380 ;
        RECT 1408.020 2133.370 1411.020 2133.380 ;
        RECT 1588.020 2133.370 1591.020 2133.380 ;
        RECT 1768.020 2133.370 1771.020 2133.380 ;
        RECT 1948.020 2133.370 1951.020 2133.380 ;
        RECT 2128.020 2133.370 2131.020 2133.380 ;
        RECT 2308.020 2133.370 2311.020 2133.380 ;
        RECT 2488.020 2133.370 2491.020 2133.380 ;
        RECT 2668.020 2133.370 2671.020 2133.380 ;
        RECT 2848.020 2133.370 2851.020 2133.380 ;
        RECT 2958.800 2133.370 2961.800 2133.380 ;
        RECT -42.180 1956.380 -39.180 1956.390 ;
        RECT 148.020 1956.380 151.020 1956.390 ;
        RECT 328.020 1956.380 331.020 1956.390 ;
        RECT 508.020 1956.380 511.020 1956.390 ;
        RECT 688.020 1956.380 691.020 1956.390 ;
        RECT 868.020 1956.380 871.020 1956.390 ;
        RECT 1048.020 1956.380 1051.020 1956.390 ;
        RECT 1228.020 1956.380 1231.020 1956.390 ;
        RECT 1408.020 1956.380 1411.020 1956.390 ;
        RECT 1588.020 1956.380 1591.020 1956.390 ;
        RECT 1768.020 1956.380 1771.020 1956.390 ;
        RECT 1948.020 1956.380 1951.020 1956.390 ;
        RECT 2128.020 1956.380 2131.020 1956.390 ;
        RECT 2308.020 1956.380 2311.020 1956.390 ;
        RECT 2488.020 1956.380 2491.020 1956.390 ;
        RECT 2668.020 1956.380 2671.020 1956.390 ;
        RECT 2848.020 1956.380 2851.020 1956.390 ;
        RECT 2958.800 1956.380 2961.800 1956.390 ;
        RECT -42.180 1953.380 2961.800 1956.380 ;
        RECT -42.180 1953.370 -39.180 1953.380 ;
        RECT 148.020 1953.370 151.020 1953.380 ;
        RECT 328.020 1953.370 331.020 1953.380 ;
        RECT 508.020 1953.370 511.020 1953.380 ;
        RECT 688.020 1953.370 691.020 1953.380 ;
        RECT 868.020 1953.370 871.020 1953.380 ;
        RECT 1048.020 1953.370 1051.020 1953.380 ;
        RECT 1228.020 1953.370 1231.020 1953.380 ;
        RECT 1408.020 1953.370 1411.020 1953.380 ;
        RECT 1588.020 1953.370 1591.020 1953.380 ;
        RECT 1768.020 1953.370 1771.020 1953.380 ;
        RECT 1948.020 1953.370 1951.020 1953.380 ;
        RECT 2128.020 1953.370 2131.020 1953.380 ;
        RECT 2308.020 1953.370 2311.020 1953.380 ;
        RECT 2488.020 1953.370 2491.020 1953.380 ;
        RECT 2668.020 1953.370 2671.020 1953.380 ;
        RECT 2848.020 1953.370 2851.020 1953.380 ;
        RECT 2958.800 1953.370 2961.800 1953.380 ;
        RECT -42.180 1776.380 -39.180 1776.390 ;
        RECT 148.020 1776.380 151.020 1776.390 ;
        RECT 328.020 1776.380 331.020 1776.390 ;
        RECT 508.020 1776.380 511.020 1776.390 ;
        RECT 688.020 1776.380 691.020 1776.390 ;
        RECT 868.020 1776.380 871.020 1776.390 ;
        RECT 1048.020 1776.380 1051.020 1776.390 ;
        RECT 1228.020 1776.380 1231.020 1776.390 ;
        RECT 1408.020 1776.380 1411.020 1776.390 ;
        RECT 1588.020 1776.380 1591.020 1776.390 ;
        RECT 1768.020 1776.380 1771.020 1776.390 ;
        RECT 1948.020 1776.380 1951.020 1776.390 ;
        RECT 2128.020 1776.380 2131.020 1776.390 ;
        RECT 2308.020 1776.380 2311.020 1776.390 ;
        RECT 2488.020 1776.380 2491.020 1776.390 ;
        RECT 2668.020 1776.380 2671.020 1776.390 ;
        RECT 2848.020 1776.380 2851.020 1776.390 ;
        RECT 2958.800 1776.380 2961.800 1776.390 ;
        RECT -42.180 1773.380 2961.800 1776.380 ;
        RECT -42.180 1773.370 -39.180 1773.380 ;
        RECT 148.020 1773.370 151.020 1773.380 ;
        RECT 328.020 1773.370 331.020 1773.380 ;
        RECT 508.020 1773.370 511.020 1773.380 ;
        RECT 688.020 1773.370 691.020 1773.380 ;
        RECT 868.020 1773.370 871.020 1773.380 ;
        RECT 1048.020 1773.370 1051.020 1773.380 ;
        RECT 1228.020 1773.370 1231.020 1773.380 ;
        RECT 1408.020 1773.370 1411.020 1773.380 ;
        RECT 1588.020 1773.370 1591.020 1773.380 ;
        RECT 1768.020 1773.370 1771.020 1773.380 ;
        RECT 1948.020 1773.370 1951.020 1773.380 ;
        RECT 2128.020 1773.370 2131.020 1773.380 ;
        RECT 2308.020 1773.370 2311.020 1773.380 ;
        RECT 2488.020 1773.370 2491.020 1773.380 ;
        RECT 2668.020 1773.370 2671.020 1773.380 ;
        RECT 2848.020 1773.370 2851.020 1773.380 ;
        RECT 2958.800 1773.370 2961.800 1773.380 ;
        RECT -42.180 1596.380 -39.180 1596.390 ;
        RECT 148.020 1596.380 151.020 1596.390 ;
        RECT 328.020 1596.380 331.020 1596.390 ;
        RECT 508.020 1596.380 511.020 1596.390 ;
        RECT 688.020 1596.380 691.020 1596.390 ;
        RECT 868.020 1596.380 871.020 1596.390 ;
        RECT 1048.020 1596.380 1051.020 1596.390 ;
        RECT 1228.020 1596.380 1231.020 1596.390 ;
        RECT 1408.020 1596.380 1411.020 1596.390 ;
        RECT 1588.020 1596.380 1591.020 1596.390 ;
        RECT 1768.020 1596.380 1771.020 1596.390 ;
        RECT 1948.020 1596.380 1951.020 1596.390 ;
        RECT 2128.020 1596.380 2131.020 1596.390 ;
        RECT 2308.020 1596.380 2311.020 1596.390 ;
        RECT 2488.020 1596.380 2491.020 1596.390 ;
        RECT 2668.020 1596.380 2671.020 1596.390 ;
        RECT 2848.020 1596.380 2851.020 1596.390 ;
        RECT 2958.800 1596.380 2961.800 1596.390 ;
        RECT -42.180 1593.380 2961.800 1596.380 ;
        RECT -42.180 1593.370 -39.180 1593.380 ;
        RECT 148.020 1593.370 151.020 1593.380 ;
        RECT 328.020 1593.370 331.020 1593.380 ;
        RECT 508.020 1593.370 511.020 1593.380 ;
        RECT 688.020 1593.370 691.020 1593.380 ;
        RECT 868.020 1593.370 871.020 1593.380 ;
        RECT 1048.020 1593.370 1051.020 1593.380 ;
        RECT 1228.020 1593.370 1231.020 1593.380 ;
        RECT 1408.020 1593.370 1411.020 1593.380 ;
        RECT 1588.020 1593.370 1591.020 1593.380 ;
        RECT 1768.020 1593.370 1771.020 1593.380 ;
        RECT 1948.020 1593.370 1951.020 1593.380 ;
        RECT 2128.020 1593.370 2131.020 1593.380 ;
        RECT 2308.020 1593.370 2311.020 1593.380 ;
        RECT 2488.020 1593.370 2491.020 1593.380 ;
        RECT 2668.020 1593.370 2671.020 1593.380 ;
        RECT 2848.020 1593.370 2851.020 1593.380 ;
        RECT 2958.800 1593.370 2961.800 1593.380 ;
        RECT -42.180 1416.380 -39.180 1416.390 ;
        RECT 148.020 1416.380 151.020 1416.390 ;
        RECT 328.020 1416.380 331.020 1416.390 ;
        RECT 508.020 1416.380 511.020 1416.390 ;
        RECT 688.020 1416.380 691.020 1416.390 ;
        RECT 868.020 1416.380 871.020 1416.390 ;
        RECT 1048.020 1416.380 1051.020 1416.390 ;
        RECT 1228.020 1416.380 1231.020 1416.390 ;
        RECT 1408.020 1416.380 1411.020 1416.390 ;
        RECT 1588.020 1416.380 1591.020 1416.390 ;
        RECT 1768.020 1416.380 1771.020 1416.390 ;
        RECT 1948.020 1416.380 1951.020 1416.390 ;
        RECT 2128.020 1416.380 2131.020 1416.390 ;
        RECT 2308.020 1416.380 2311.020 1416.390 ;
        RECT 2488.020 1416.380 2491.020 1416.390 ;
        RECT 2668.020 1416.380 2671.020 1416.390 ;
        RECT 2848.020 1416.380 2851.020 1416.390 ;
        RECT 2958.800 1416.380 2961.800 1416.390 ;
        RECT -42.180 1413.380 2961.800 1416.380 ;
        RECT -42.180 1413.370 -39.180 1413.380 ;
        RECT 148.020 1413.370 151.020 1413.380 ;
        RECT 328.020 1413.370 331.020 1413.380 ;
        RECT 508.020 1413.370 511.020 1413.380 ;
        RECT 688.020 1413.370 691.020 1413.380 ;
        RECT 868.020 1413.370 871.020 1413.380 ;
        RECT 1048.020 1413.370 1051.020 1413.380 ;
        RECT 1228.020 1413.370 1231.020 1413.380 ;
        RECT 1408.020 1413.370 1411.020 1413.380 ;
        RECT 1588.020 1413.370 1591.020 1413.380 ;
        RECT 1768.020 1413.370 1771.020 1413.380 ;
        RECT 1948.020 1413.370 1951.020 1413.380 ;
        RECT 2128.020 1413.370 2131.020 1413.380 ;
        RECT 2308.020 1413.370 2311.020 1413.380 ;
        RECT 2488.020 1413.370 2491.020 1413.380 ;
        RECT 2668.020 1413.370 2671.020 1413.380 ;
        RECT 2848.020 1413.370 2851.020 1413.380 ;
        RECT 2958.800 1413.370 2961.800 1413.380 ;
        RECT -42.180 1236.380 -39.180 1236.390 ;
        RECT 148.020 1236.380 151.020 1236.390 ;
        RECT 328.020 1236.380 331.020 1236.390 ;
        RECT 508.020 1236.380 511.020 1236.390 ;
        RECT 688.020 1236.380 691.020 1236.390 ;
        RECT 868.020 1236.380 871.020 1236.390 ;
        RECT 1048.020 1236.380 1051.020 1236.390 ;
        RECT 1228.020 1236.380 1231.020 1236.390 ;
        RECT 1408.020 1236.380 1411.020 1236.390 ;
        RECT 1588.020 1236.380 1591.020 1236.390 ;
        RECT 1768.020 1236.380 1771.020 1236.390 ;
        RECT 1948.020 1236.380 1951.020 1236.390 ;
        RECT 2128.020 1236.380 2131.020 1236.390 ;
        RECT 2308.020 1236.380 2311.020 1236.390 ;
        RECT 2488.020 1236.380 2491.020 1236.390 ;
        RECT 2668.020 1236.380 2671.020 1236.390 ;
        RECT 2848.020 1236.380 2851.020 1236.390 ;
        RECT 2958.800 1236.380 2961.800 1236.390 ;
        RECT -42.180 1233.380 2961.800 1236.380 ;
        RECT -42.180 1233.370 -39.180 1233.380 ;
        RECT 148.020 1233.370 151.020 1233.380 ;
        RECT 328.020 1233.370 331.020 1233.380 ;
        RECT 508.020 1233.370 511.020 1233.380 ;
        RECT 688.020 1233.370 691.020 1233.380 ;
        RECT 868.020 1233.370 871.020 1233.380 ;
        RECT 1048.020 1233.370 1051.020 1233.380 ;
        RECT 1228.020 1233.370 1231.020 1233.380 ;
        RECT 1408.020 1233.370 1411.020 1233.380 ;
        RECT 1588.020 1233.370 1591.020 1233.380 ;
        RECT 1768.020 1233.370 1771.020 1233.380 ;
        RECT 1948.020 1233.370 1951.020 1233.380 ;
        RECT 2128.020 1233.370 2131.020 1233.380 ;
        RECT 2308.020 1233.370 2311.020 1233.380 ;
        RECT 2488.020 1233.370 2491.020 1233.380 ;
        RECT 2668.020 1233.370 2671.020 1233.380 ;
        RECT 2848.020 1233.370 2851.020 1233.380 ;
        RECT 2958.800 1233.370 2961.800 1233.380 ;
        RECT -42.180 1056.380 -39.180 1056.390 ;
        RECT 148.020 1056.380 151.020 1056.390 ;
        RECT 328.020 1056.380 331.020 1056.390 ;
        RECT 508.020 1056.380 511.020 1056.390 ;
        RECT 688.020 1056.380 691.020 1056.390 ;
        RECT 868.020 1056.380 871.020 1056.390 ;
        RECT 1048.020 1056.380 1051.020 1056.390 ;
        RECT 1228.020 1056.380 1231.020 1056.390 ;
        RECT 1408.020 1056.380 1411.020 1056.390 ;
        RECT 1588.020 1056.380 1591.020 1056.390 ;
        RECT 1768.020 1056.380 1771.020 1056.390 ;
        RECT 1948.020 1056.380 1951.020 1056.390 ;
        RECT 2128.020 1056.380 2131.020 1056.390 ;
        RECT 2308.020 1056.380 2311.020 1056.390 ;
        RECT 2488.020 1056.380 2491.020 1056.390 ;
        RECT 2668.020 1056.380 2671.020 1056.390 ;
        RECT 2848.020 1056.380 2851.020 1056.390 ;
        RECT 2958.800 1056.380 2961.800 1056.390 ;
        RECT -42.180 1053.380 2961.800 1056.380 ;
        RECT -42.180 1053.370 -39.180 1053.380 ;
        RECT 148.020 1053.370 151.020 1053.380 ;
        RECT 328.020 1053.370 331.020 1053.380 ;
        RECT 508.020 1053.370 511.020 1053.380 ;
        RECT 688.020 1053.370 691.020 1053.380 ;
        RECT 868.020 1053.370 871.020 1053.380 ;
        RECT 1048.020 1053.370 1051.020 1053.380 ;
        RECT 1228.020 1053.370 1231.020 1053.380 ;
        RECT 1408.020 1053.370 1411.020 1053.380 ;
        RECT 1588.020 1053.370 1591.020 1053.380 ;
        RECT 1768.020 1053.370 1771.020 1053.380 ;
        RECT 1948.020 1053.370 1951.020 1053.380 ;
        RECT 2128.020 1053.370 2131.020 1053.380 ;
        RECT 2308.020 1053.370 2311.020 1053.380 ;
        RECT 2488.020 1053.370 2491.020 1053.380 ;
        RECT 2668.020 1053.370 2671.020 1053.380 ;
        RECT 2848.020 1053.370 2851.020 1053.380 ;
        RECT 2958.800 1053.370 2961.800 1053.380 ;
        RECT -42.180 876.380 -39.180 876.390 ;
        RECT 148.020 876.380 151.020 876.390 ;
        RECT 328.020 876.380 331.020 876.390 ;
        RECT 508.020 876.380 511.020 876.390 ;
        RECT 688.020 876.380 691.020 876.390 ;
        RECT 868.020 876.380 871.020 876.390 ;
        RECT 1048.020 876.380 1051.020 876.390 ;
        RECT 1228.020 876.380 1231.020 876.390 ;
        RECT 1408.020 876.380 1411.020 876.390 ;
        RECT 1588.020 876.380 1591.020 876.390 ;
        RECT 1768.020 876.380 1771.020 876.390 ;
        RECT 1948.020 876.380 1951.020 876.390 ;
        RECT 2128.020 876.380 2131.020 876.390 ;
        RECT 2308.020 876.380 2311.020 876.390 ;
        RECT 2488.020 876.380 2491.020 876.390 ;
        RECT 2668.020 876.380 2671.020 876.390 ;
        RECT 2848.020 876.380 2851.020 876.390 ;
        RECT 2958.800 876.380 2961.800 876.390 ;
        RECT -42.180 873.380 2961.800 876.380 ;
        RECT -42.180 873.370 -39.180 873.380 ;
        RECT 148.020 873.370 151.020 873.380 ;
        RECT 328.020 873.370 331.020 873.380 ;
        RECT 508.020 873.370 511.020 873.380 ;
        RECT 688.020 873.370 691.020 873.380 ;
        RECT 868.020 873.370 871.020 873.380 ;
        RECT 1048.020 873.370 1051.020 873.380 ;
        RECT 1228.020 873.370 1231.020 873.380 ;
        RECT 1408.020 873.370 1411.020 873.380 ;
        RECT 1588.020 873.370 1591.020 873.380 ;
        RECT 1768.020 873.370 1771.020 873.380 ;
        RECT 1948.020 873.370 1951.020 873.380 ;
        RECT 2128.020 873.370 2131.020 873.380 ;
        RECT 2308.020 873.370 2311.020 873.380 ;
        RECT 2488.020 873.370 2491.020 873.380 ;
        RECT 2668.020 873.370 2671.020 873.380 ;
        RECT 2848.020 873.370 2851.020 873.380 ;
        RECT 2958.800 873.370 2961.800 873.380 ;
        RECT -42.180 696.380 -39.180 696.390 ;
        RECT 148.020 696.380 151.020 696.390 ;
        RECT 328.020 696.380 331.020 696.390 ;
        RECT 508.020 696.380 511.020 696.390 ;
        RECT 688.020 696.380 691.020 696.390 ;
        RECT 868.020 696.380 871.020 696.390 ;
        RECT 1048.020 696.380 1051.020 696.390 ;
        RECT 1228.020 696.380 1231.020 696.390 ;
        RECT 1408.020 696.380 1411.020 696.390 ;
        RECT 1588.020 696.380 1591.020 696.390 ;
        RECT 1768.020 696.380 1771.020 696.390 ;
        RECT 1948.020 696.380 1951.020 696.390 ;
        RECT 2128.020 696.380 2131.020 696.390 ;
        RECT 2308.020 696.380 2311.020 696.390 ;
        RECT 2488.020 696.380 2491.020 696.390 ;
        RECT 2668.020 696.380 2671.020 696.390 ;
        RECT 2848.020 696.380 2851.020 696.390 ;
        RECT 2958.800 696.380 2961.800 696.390 ;
        RECT -42.180 693.380 2961.800 696.380 ;
        RECT -42.180 693.370 -39.180 693.380 ;
        RECT 148.020 693.370 151.020 693.380 ;
        RECT 328.020 693.370 331.020 693.380 ;
        RECT 508.020 693.370 511.020 693.380 ;
        RECT 688.020 693.370 691.020 693.380 ;
        RECT 868.020 693.370 871.020 693.380 ;
        RECT 1048.020 693.370 1051.020 693.380 ;
        RECT 1228.020 693.370 1231.020 693.380 ;
        RECT 1408.020 693.370 1411.020 693.380 ;
        RECT 1588.020 693.370 1591.020 693.380 ;
        RECT 1768.020 693.370 1771.020 693.380 ;
        RECT 1948.020 693.370 1951.020 693.380 ;
        RECT 2128.020 693.370 2131.020 693.380 ;
        RECT 2308.020 693.370 2311.020 693.380 ;
        RECT 2488.020 693.370 2491.020 693.380 ;
        RECT 2668.020 693.370 2671.020 693.380 ;
        RECT 2848.020 693.370 2851.020 693.380 ;
        RECT 2958.800 693.370 2961.800 693.380 ;
        RECT -42.180 516.380 -39.180 516.390 ;
        RECT 148.020 516.380 151.020 516.390 ;
        RECT 328.020 516.380 331.020 516.390 ;
        RECT 508.020 516.380 511.020 516.390 ;
        RECT 688.020 516.380 691.020 516.390 ;
        RECT 868.020 516.380 871.020 516.390 ;
        RECT 1048.020 516.380 1051.020 516.390 ;
        RECT 1228.020 516.380 1231.020 516.390 ;
        RECT 1408.020 516.380 1411.020 516.390 ;
        RECT 1588.020 516.380 1591.020 516.390 ;
        RECT 1768.020 516.380 1771.020 516.390 ;
        RECT 1948.020 516.380 1951.020 516.390 ;
        RECT 2128.020 516.380 2131.020 516.390 ;
        RECT 2308.020 516.380 2311.020 516.390 ;
        RECT 2488.020 516.380 2491.020 516.390 ;
        RECT 2668.020 516.380 2671.020 516.390 ;
        RECT 2848.020 516.380 2851.020 516.390 ;
        RECT 2958.800 516.380 2961.800 516.390 ;
        RECT -42.180 513.380 2961.800 516.380 ;
        RECT -42.180 513.370 -39.180 513.380 ;
        RECT 148.020 513.370 151.020 513.380 ;
        RECT 328.020 513.370 331.020 513.380 ;
        RECT 508.020 513.370 511.020 513.380 ;
        RECT 688.020 513.370 691.020 513.380 ;
        RECT 868.020 513.370 871.020 513.380 ;
        RECT 1048.020 513.370 1051.020 513.380 ;
        RECT 1228.020 513.370 1231.020 513.380 ;
        RECT 1408.020 513.370 1411.020 513.380 ;
        RECT 1588.020 513.370 1591.020 513.380 ;
        RECT 1768.020 513.370 1771.020 513.380 ;
        RECT 1948.020 513.370 1951.020 513.380 ;
        RECT 2128.020 513.370 2131.020 513.380 ;
        RECT 2308.020 513.370 2311.020 513.380 ;
        RECT 2488.020 513.370 2491.020 513.380 ;
        RECT 2668.020 513.370 2671.020 513.380 ;
        RECT 2848.020 513.370 2851.020 513.380 ;
        RECT 2958.800 513.370 2961.800 513.380 ;
        RECT -42.180 336.380 -39.180 336.390 ;
        RECT 148.020 336.380 151.020 336.390 ;
        RECT 328.020 336.380 331.020 336.390 ;
        RECT 508.020 336.380 511.020 336.390 ;
        RECT 688.020 336.380 691.020 336.390 ;
        RECT 868.020 336.380 871.020 336.390 ;
        RECT 1048.020 336.380 1051.020 336.390 ;
        RECT 1228.020 336.380 1231.020 336.390 ;
        RECT 1408.020 336.380 1411.020 336.390 ;
        RECT 1588.020 336.380 1591.020 336.390 ;
        RECT 1768.020 336.380 1771.020 336.390 ;
        RECT 1948.020 336.380 1951.020 336.390 ;
        RECT 2128.020 336.380 2131.020 336.390 ;
        RECT 2308.020 336.380 2311.020 336.390 ;
        RECT 2488.020 336.380 2491.020 336.390 ;
        RECT 2668.020 336.380 2671.020 336.390 ;
        RECT 2848.020 336.380 2851.020 336.390 ;
        RECT 2958.800 336.380 2961.800 336.390 ;
        RECT -42.180 333.380 2961.800 336.380 ;
        RECT -42.180 333.370 -39.180 333.380 ;
        RECT 148.020 333.370 151.020 333.380 ;
        RECT 328.020 333.370 331.020 333.380 ;
        RECT 508.020 333.370 511.020 333.380 ;
        RECT 688.020 333.370 691.020 333.380 ;
        RECT 868.020 333.370 871.020 333.380 ;
        RECT 1048.020 333.370 1051.020 333.380 ;
        RECT 1228.020 333.370 1231.020 333.380 ;
        RECT 1408.020 333.370 1411.020 333.380 ;
        RECT 1588.020 333.370 1591.020 333.380 ;
        RECT 1768.020 333.370 1771.020 333.380 ;
        RECT 1948.020 333.370 1951.020 333.380 ;
        RECT 2128.020 333.370 2131.020 333.380 ;
        RECT 2308.020 333.370 2311.020 333.380 ;
        RECT 2488.020 333.370 2491.020 333.380 ;
        RECT 2668.020 333.370 2671.020 333.380 ;
        RECT 2848.020 333.370 2851.020 333.380 ;
        RECT 2958.800 333.370 2961.800 333.380 ;
        RECT -42.180 156.380 -39.180 156.390 ;
        RECT 148.020 156.380 151.020 156.390 ;
        RECT 328.020 156.380 331.020 156.390 ;
        RECT 508.020 156.380 511.020 156.390 ;
        RECT 688.020 156.380 691.020 156.390 ;
        RECT 868.020 156.380 871.020 156.390 ;
        RECT 1048.020 156.380 1051.020 156.390 ;
        RECT 1228.020 156.380 1231.020 156.390 ;
        RECT 1408.020 156.380 1411.020 156.390 ;
        RECT 1588.020 156.380 1591.020 156.390 ;
        RECT 1768.020 156.380 1771.020 156.390 ;
        RECT 1948.020 156.380 1951.020 156.390 ;
        RECT 2128.020 156.380 2131.020 156.390 ;
        RECT 2308.020 156.380 2311.020 156.390 ;
        RECT 2488.020 156.380 2491.020 156.390 ;
        RECT 2668.020 156.380 2671.020 156.390 ;
        RECT 2848.020 156.380 2851.020 156.390 ;
        RECT 2958.800 156.380 2961.800 156.390 ;
        RECT -42.180 153.380 2961.800 156.380 ;
        RECT -42.180 153.370 -39.180 153.380 ;
        RECT 148.020 153.370 151.020 153.380 ;
        RECT 328.020 153.370 331.020 153.380 ;
        RECT 508.020 153.370 511.020 153.380 ;
        RECT 688.020 153.370 691.020 153.380 ;
        RECT 868.020 153.370 871.020 153.380 ;
        RECT 1048.020 153.370 1051.020 153.380 ;
        RECT 1228.020 153.370 1231.020 153.380 ;
        RECT 1408.020 153.370 1411.020 153.380 ;
        RECT 1588.020 153.370 1591.020 153.380 ;
        RECT 1768.020 153.370 1771.020 153.380 ;
        RECT 1948.020 153.370 1951.020 153.380 ;
        RECT 2128.020 153.370 2131.020 153.380 ;
        RECT 2308.020 153.370 2311.020 153.380 ;
        RECT 2488.020 153.370 2491.020 153.380 ;
        RECT 2668.020 153.370 2671.020 153.380 ;
        RECT 2848.020 153.370 2851.020 153.380 ;
        RECT 2958.800 153.370 2961.800 153.380 ;
        RECT -42.180 -33.820 -39.180 -33.810 ;
        RECT 148.020 -33.820 151.020 -33.810 ;
        RECT 328.020 -33.820 331.020 -33.810 ;
        RECT 508.020 -33.820 511.020 -33.810 ;
        RECT 688.020 -33.820 691.020 -33.810 ;
        RECT 868.020 -33.820 871.020 -33.810 ;
        RECT 1048.020 -33.820 1051.020 -33.810 ;
        RECT 1228.020 -33.820 1231.020 -33.810 ;
        RECT 1408.020 -33.820 1411.020 -33.810 ;
        RECT 1588.020 -33.820 1591.020 -33.810 ;
        RECT 1768.020 -33.820 1771.020 -33.810 ;
        RECT 1948.020 -33.820 1951.020 -33.810 ;
        RECT 2128.020 -33.820 2131.020 -33.810 ;
        RECT 2308.020 -33.820 2311.020 -33.810 ;
        RECT 2488.020 -33.820 2491.020 -33.810 ;
        RECT 2668.020 -33.820 2671.020 -33.810 ;
        RECT 2848.020 -33.820 2851.020 -33.810 ;
        RECT 2958.800 -33.820 2961.800 -33.810 ;
        RECT -42.180 -36.820 2961.800 -33.820 ;
        RECT -42.180 -36.830 -39.180 -36.820 ;
        RECT 148.020 -36.830 151.020 -36.820 ;
        RECT 328.020 -36.830 331.020 -36.820 ;
        RECT 508.020 -36.830 511.020 -36.820 ;
        RECT 688.020 -36.830 691.020 -36.820 ;
        RECT 868.020 -36.830 871.020 -36.820 ;
        RECT 1048.020 -36.830 1051.020 -36.820 ;
        RECT 1228.020 -36.830 1231.020 -36.820 ;
        RECT 1408.020 -36.830 1411.020 -36.820 ;
        RECT 1588.020 -36.830 1591.020 -36.820 ;
        RECT 1768.020 -36.830 1771.020 -36.820 ;
        RECT 1948.020 -36.830 1951.020 -36.820 ;
        RECT 2128.020 -36.830 2131.020 -36.820 ;
        RECT 2308.020 -36.830 2311.020 -36.820 ;
        RECT 2488.020 -36.830 2491.020 -36.820 ;
        RECT 2668.020 -36.830 2671.020 -36.820 ;
        RECT 2848.020 -36.830 2851.020 -36.820 ;
        RECT 2958.800 -36.830 2961.800 -36.820 ;
    END
  END vssa2
  OBS
      LAYER li1 ;
        RECT 1155.430 1710.795 1444.310 1995.715 ;
      LAYER met1 ;
        RECT 1150.900 1705.480 1448.840 1995.760 ;
      LAYER met2 ;
        RECT 1151.480 1995.720 1152.940 1996.000 ;
        RECT 1153.780 1995.720 1155.700 1996.000 ;
        RECT 1156.540 1995.720 1158.460 1996.000 ;
        RECT 1159.300 1995.720 1160.760 1996.000 ;
        RECT 1161.600 1995.720 1163.520 1996.000 ;
        RECT 1164.360 1995.720 1166.280 1996.000 ;
        RECT 1167.120 1995.720 1169.040 1996.000 ;
        RECT 1169.880 1995.720 1171.340 1996.000 ;
        RECT 1172.180 1995.720 1174.100 1996.000 ;
        RECT 1174.940 1995.720 1176.860 1996.000 ;
        RECT 1177.700 1995.720 1179.160 1996.000 ;
        RECT 1180.000 1995.720 1181.920 1996.000 ;
        RECT 1182.760 1995.720 1184.680 1996.000 ;
        RECT 1185.520 1995.720 1187.440 1996.000 ;
        RECT 1188.280 1995.720 1189.740 1996.000 ;
        RECT 1190.580 1995.720 1192.500 1996.000 ;
        RECT 1193.340 1995.720 1195.260 1996.000 ;
        RECT 1196.100 1995.720 1197.560 1996.000 ;
        RECT 1198.400 1995.720 1200.320 1996.000 ;
        RECT 1201.160 1995.720 1203.080 1996.000 ;
        RECT 1203.920 1995.720 1205.840 1996.000 ;
        RECT 1206.680 1995.720 1208.140 1996.000 ;
        RECT 1208.980 1995.720 1210.900 1996.000 ;
        RECT 1211.740 1995.720 1213.660 1996.000 ;
        RECT 1214.500 1995.720 1215.960 1996.000 ;
        RECT 1216.800 1995.720 1218.720 1996.000 ;
        RECT 1219.560 1995.720 1221.480 1996.000 ;
        RECT 1222.320 1995.720 1224.240 1996.000 ;
        RECT 1225.080 1995.720 1226.540 1996.000 ;
        RECT 1227.380 1995.720 1229.300 1996.000 ;
        RECT 1230.140 1995.720 1232.060 1996.000 ;
        RECT 1232.900 1995.720 1234.820 1996.000 ;
        RECT 1235.660 1995.720 1237.120 1996.000 ;
        RECT 1237.960 1995.720 1239.880 1996.000 ;
        RECT 1240.720 1995.720 1242.640 1996.000 ;
        RECT 1243.480 1995.720 1244.940 1996.000 ;
        RECT 1245.780 1995.720 1247.700 1996.000 ;
        RECT 1248.540 1995.720 1250.460 1996.000 ;
        RECT 1251.300 1995.720 1253.220 1996.000 ;
        RECT 1254.060 1995.720 1255.520 1996.000 ;
        RECT 1256.360 1995.720 1258.280 1996.000 ;
        RECT 1259.120 1995.720 1261.040 1996.000 ;
        RECT 1261.880 1995.720 1263.340 1996.000 ;
        RECT 1264.180 1995.720 1266.100 1996.000 ;
        RECT 1266.940 1995.720 1268.860 1996.000 ;
        RECT 1269.700 1995.720 1271.620 1996.000 ;
        RECT 1272.460 1995.720 1273.920 1996.000 ;
        RECT 1274.760 1995.720 1276.680 1996.000 ;
        RECT 1277.520 1995.720 1279.440 1996.000 ;
        RECT 1280.280 1995.720 1281.740 1996.000 ;
        RECT 1282.580 1995.720 1284.500 1996.000 ;
        RECT 1285.340 1995.720 1287.260 1996.000 ;
        RECT 1288.100 1995.720 1290.020 1996.000 ;
        RECT 1290.860 1995.720 1292.320 1996.000 ;
        RECT 1293.160 1995.720 1295.080 1996.000 ;
        RECT 1295.920 1995.720 1297.840 1996.000 ;
        RECT 1298.680 1995.720 1300.600 1996.000 ;
        RECT 1301.440 1995.720 1302.900 1996.000 ;
        RECT 1303.740 1995.720 1305.660 1996.000 ;
        RECT 1306.500 1995.720 1308.420 1996.000 ;
        RECT 1309.260 1995.720 1310.720 1996.000 ;
        RECT 1311.560 1995.720 1313.480 1996.000 ;
        RECT 1314.320 1995.720 1316.240 1996.000 ;
        RECT 1317.080 1995.720 1319.000 1996.000 ;
        RECT 1319.840 1995.720 1321.300 1996.000 ;
        RECT 1322.140 1995.720 1324.060 1996.000 ;
        RECT 1324.900 1995.720 1326.820 1996.000 ;
        RECT 1327.660 1995.720 1329.120 1996.000 ;
        RECT 1329.960 1995.720 1331.880 1996.000 ;
        RECT 1332.720 1995.720 1334.640 1996.000 ;
        RECT 1335.480 1995.720 1337.400 1996.000 ;
        RECT 1338.240 1995.720 1339.700 1996.000 ;
        RECT 1340.540 1995.720 1342.460 1996.000 ;
        RECT 1343.300 1995.720 1345.220 1996.000 ;
        RECT 1346.060 1995.720 1347.520 1996.000 ;
        RECT 1348.360 1995.720 1350.280 1996.000 ;
        RECT 1351.120 1995.720 1353.040 1996.000 ;
        RECT 1353.880 1995.720 1355.800 1996.000 ;
        RECT 1356.640 1995.720 1358.100 1996.000 ;
        RECT 1358.940 1995.720 1360.860 1996.000 ;
        RECT 1361.700 1995.720 1363.620 1996.000 ;
        RECT 1364.460 1995.720 1365.920 1996.000 ;
        RECT 1366.760 1995.720 1368.680 1996.000 ;
        RECT 1369.520 1995.720 1371.440 1996.000 ;
        RECT 1372.280 1995.720 1374.200 1996.000 ;
        RECT 1375.040 1995.720 1376.500 1996.000 ;
        RECT 1377.340 1995.720 1379.260 1996.000 ;
        RECT 1380.100 1995.720 1382.020 1996.000 ;
        RECT 1382.860 1995.720 1384.780 1996.000 ;
        RECT 1385.620 1995.720 1387.080 1996.000 ;
        RECT 1387.920 1995.720 1389.840 1996.000 ;
        RECT 1390.680 1995.720 1392.600 1996.000 ;
        RECT 1393.440 1995.720 1394.900 1996.000 ;
        RECT 1395.740 1995.720 1397.660 1996.000 ;
        RECT 1398.500 1995.720 1400.420 1996.000 ;
        RECT 1401.260 1995.720 1403.180 1996.000 ;
        RECT 1404.020 1995.720 1405.480 1996.000 ;
        RECT 1406.320 1995.720 1408.240 1996.000 ;
        RECT 1409.080 1995.720 1411.000 1996.000 ;
        RECT 1411.840 1995.720 1413.300 1996.000 ;
        RECT 1414.140 1995.720 1416.060 1996.000 ;
        RECT 1416.900 1995.720 1418.820 1996.000 ;
        RECT 1419.660 1995.720 1421.580 1996.000 ;
        RECT 1422.420 1995.720 1423.880 1996.000 ;
        RECT 1424.720 1995.720 1426.640 1996.000 ;
        RECT 1427.480 1995.720 1429.400 1996.000 ;
        RECT 1430.240 1995.720 1431.700 1996.000 ;
        RECT 1432.540 1995.720 1434.460 1996.000 ;
        RECT 1435.300 1995.720 1437.220 1996.000 ;
        RECT 1438.060 1995.720 1439.980 1996.000 ;
        RECT 1440.820 1995.720 1442.280 1996.000 ;
        RECT 1443.120 1995.720 1445.040 1996.000 ;
        RECT 1445.880 1995.720 1447.800 1996.000 ;
        RECT 1448.640 1995.720 1448.810 1996.000 ;
        RECT 1150.930 1704.280 1448.810 1995.720 ;
        RECT 1151.940 1704.000 1152.020 1704.280 ;
        RECT 1153.780 1704.000 1153.860 1704.280 ;
        RECT 1155.620 1704.000 1155.700 1704.280 ;
        RECT 1157.460 1704.000 1157.540 1704.280 ;
        RECT 1159.300 1704.000 1159.380 1704.280 ;
        RECT 1161.140 1704.000 1161.220 1704.280 ;
        RECT 1162.980 1704.000 1163.060 1704.280 ;
        RECT 1164.820 1704.000 1164.900 1704.280 ;
        RECT 1166.660 1704.000 1166.740 1704.280 ;
        RECT 1168.500 1704.000 1168.580 1704.280 ;
        RECT 1170.340 1704.000 1170.420 1704.280 ;
        RECT 1172.180 1704.000 1172.260 1704.280 ;
        RECT 1174.020 1704.000 1174.100 1704.280 ;
        RECT 1175.860 1704.000 1175.940 1704.280 ;
        RECT 1177.700 1704.000 1177.780 1704.280 ;
        RECT 1179.540 1704.000 1179.620 1704.280 ;
        RECT 1181.380 1704.000 1181.460 1704.280 ;
        RECT 1183.220 1704.000 1183.300 1704.280 ;
        RECT 1185.060 1704.000 1185.140 1704.280 ;
        RECT 1186.900 1704.000 1186.980 1704.280 ;
        RECT 1188.740 1704.000 1188.820 1704.280 ;
        RECT 1190.580 1704.000 1190.660 1704.280 ;
        RECT 1192.420 1704.000 1192.500 1704.280 ;
        RECT 1194.260 1704.000 1194.340 1704.280 ;
        RECT 1196.100 1704.000 1196.180 1704.280 ;
        RECT 1197.940 1704.000 1198.020 1704.280 ;
        RECT 1199.780 1704.000 1199.860 1704.280 ;
        RECT 1201.620 1704.000 1201.700 1704.280 ;
        RECT 1203.460 1704.000 1203.540 1704.280 ;
        RECT 1205.300 1704.000 1205.380 1704.280 ;
        RECT 1207.140 1704.000 1207.220 1704.280 ;
        RECT 1208.980 1704.000 1209.060 1704.280 ;
        RECT 1210.820 1704.000 1210.900 1704.280 ;
        RECT 1212.660 1704.000 1212.740 1704.280 ;
        RECT 1214.500 1704.000 1214.580 1704.280 ;
        RECT 1216.340 1704.000 1216.420 1704.280 ;
        RECT 1218.180 1704.000 1218.260 1704.280 ;
        RECT 1220.020 1704.000 1220.100 1704.280 ;
        RECT 1221.860 1704.000 1221.940 1704.280 ;
        RECT 1223.700 1704.000 1223.780 1704.280 ;
        RECT 1226.000 1704.000 1226.080 1704.280 ;
        RECT 1227.840 1704.000 1227.920 1704.280 ;
        RECT 1229.680 1704.000 1229.760 1704.280 ;
        RECT 1231.520 1704.000 1231.600 1704.280 ;
        RECT 1233.360 1704.000 1233.440 1704.280 ;
        RECT 1235.200 1704.000 1235.280 1704.280 ;
        RECT 1237.040 1704.000 1237.120 1704.280 ;
        RECT 1238.880 1704.000 1238.960 1704.280 ;
        RECT 1240.720 1704.000 1240.800 1704.280 ;
        RECT 1242.560 1704.000 1242.640 1704.280 ;
        RECT 1244.400 1704.000 1244.480 1704.280 ;
        RECT 1246.240 1704.000 1246.320 1704.280 ;
        RECT 1248.080 1704.000 1248.160 1704.280 ;
        RECT 1249.920 1704.000 1250.000 1704.280 ;
        RECT 1251.760 1704.000 1251.840 1704.280 ;
        RECT 1253.600 1704.000 1253.680 1704.280 ;
        RECT 1255.440 1704.000 1255.520 1704.280 ;
        RECT 1257.280 1704.000 1257.360 1704.280 ;
        RECT 1259.120 1704.000 1259.200 1704.280 ;
        RECT 1260.960 1704.000 1261.040 1704.280 ;
        RECT 1262.800 1704.000 1262.880 1704.280 ;
        RECT 1264.640 1704.000 1264.720 1704.280 ;
        RECT 1266.480 1704.000 1266.560 1704.280 ;
        RECT 1268.320 1704.000 1268.400 1704.280 ;
        RECT 1270.160 1704.000 1270.240 1704.280 ;
        RECT 1272.000 1704.000 1272.080 1704.280 ;
        RECT 1273.840 1704.000 1273.920 1704.280 ;
        RECT 1275.680 1704.000 1275.760 1704.280 ;
        RECT 1277.520 1704.000 1277.600 1704.280 ;
        RECT 1279.360 1704.000 1279.440 1704.280 ;
        RECT 1281.200 1704.000 1281.280 1704.280 ;
        RECT 1283.040 1704.000 1283.120 1704.280 ;
        RECT 1284.880 1704.000 1284.960 1704.280 ;
        RECT 1286.720 1704.000 1286.800 1704.280 ;
        RECT 1288.560 1704.000 1288.640 1704.280 ;
        RECT 1290.400 1704.000 1290.480 1704.280 ;
        RECT 1292.240 1704.000 1292.320 1704.280 ;
        RECT 1294.080 1704.000 1294.160 1704.280 ;
        RECT 1295.920 1704.000 1296.000 1704.280 ;
        RECT 1297.760 1704.000 1297.840 1704.280 ;
        RECT 1299.600 1704.000 1299.680 1704.280 ;
        RECT 1301.900 1704.000 1301.980 1704.280 ;
        RECT 1303.740 1704.000 1303.820 1704.280 ;
        RECT 1305.580 1704.000 1305.660 1704.280 ;
        RECT 1307.420 1704.000 1307.500 1704.280 ;
        RECT 1309.260 1704.000 1309.340 1704.280 ;
        RECT 1311.100 1704.000 1311.180 1704.280 ;
        RECT 1312.940 1704.000 1313.020 1704.280 ;
        RECT 1314.780 1704.000 1314.860 1704.280 ;
        RECT 1316.620 1704.000 1316.700 1704.280 ;
        RECT 1318.460 1704.000 1318.540 1704.280 ;
        RECT 1320.300 1704.000 1320.380 1704.280 ;
        RECT 1322.140 1704.000 1322.220 1704.280 ;
        RECT 1323.980 1704.000 1324.060 1704.280 ;
        RECT 1325.820 1704.000 1325.900 1704.280 ;
        RECT 1327.660 1704.000 1327.740 1704.280 ;
        RECT 1329.500 1704.000 1329.580 1704.280 ;
        RECT 1331.340 1704.000 1331.420 1704.280 ;
        RECT 1333.180 1704.000 1333.260 1704.280 ;
        RECT 1335.020 1704.000 1335.100 1704.280 ;
        RECT 1336.860 1704.000 1336.940 1704.280 ;
        RECT 1338.700 1704.000 1338.780 1704.280 ;
        RECT 1340.540 1704.000 1340.620 1704.280 ;
        RECT 1342.380 1704.000 1342.460 1704.280 ;
        RECT 1344.220 1704.000 1344.300 1704.280 ;
        RECT 1346.060 1704.000 1346.140 1704.280 ;
        RECT 1347.900 1704.000 1347.980 1704.280 ;
        RECT 1349.740 1704.000 1349.820 1704.280 ;
        RECT 1351.580 1704.000 1351.660 1704.280 ;
        RECT 1353.420 1704.000 1353.500 1704.280 ;
        RECT 1355.260 1704.000 1355.340 1704.280 ;
        RECT 1357.100 1704.000 1357.180 1704.280 ;
        RECT 1358.940 1704.000 1359.020 1704.280 ;
        RECT 1360.780 1704.000 1360.860 1704.280 ;
        RECT 1362.620 1704.000 1362.700 1704.280 ;
        RECT 1364.460 1704.000 1364.540 1704.280 ;
        RECT 1366.300 1704.000 1366.380 1704.280 ;
        RECT 1368.140 1704.000 1368.220 1704.280 ;
        RECT 1369.980 1704.000 1370.060 1704.280 ;
        RECT 1371.820 1704.000 1371.900 1704.280 ;
        RECT 1373.660 1704.000 1373.740 1704.280 ;
        RECT 1375.960 1704.000 1376.040 1704.280 ;
        RECT 1377.800 1704.000 1377.880 1704.280 ;
        RECT 1379.640 1704.000 1379.720 1704.280 ;
        RECT 1381.480 1704.000 1381.560 1704.280 ;
        RECT 1383.320 1704.000 1383.400 1704.280 ;
        RECT 1385.160 1704.000 1385.240 1704.280 ;
        RECT 1387.000 1704.000 1387.080 1704.280 ;
        RECT 1388.840 1704.000 1388.920 1704.280 ;
        RECT 1390.680 1704.000 1390.760 1704.280 ;
        RECT 1392.520 1704.000 1392.600 1704.280 ;
        RECT 1394.360 1704.000 1394.440 1704.280 ;
        RECT 1396.200 1704.000 1396.280 1704.280 ;
        RECT 1398.040 1704.000 1398.120 1704.280 ;
        RECT 1399.880 1704.000 1399.960 1704.280 ;
        RECT 1401.720 1704.000 1401.800 1704.280 ;
        RECT 1403.560 1704.000 1403.640 1704.280 ;
        RECT 1405.400 1704.000 1405.480 1704.280 ;
        RECT 1407.240 1704.000 1407.320 1704.280 ;
        RECT 1409.080 1704.000 1409.160 1704.280 ;
        RECT 1410.920 1704.000 1411.000 1704.280 ;
        RECT 1412.760 1704.000 1412.840 1704.280 ;
        RECT 1414.600 1704.000 1414.680 1704.280 ;
        RECT 1416.440 1704.000 1416.520 1704.280 ;
        RECT 1418.280 1704.000 1418.360 1704.280 ;
        RECT 1420.120 1704.000 1420.200 1704.280 ;
        RECT 1421.960 1704.000 1422.040 1704.280 ;
        RECT 1423.800 1704.000 1423.880 1704.280 ;
        RECT 1425.640 1704.000 1425.720 1704.280 ;
        RECT 1427.480 1704.000 1427.560 1704.280 ;
        RECT 1429.320 1704.000 1429.400 1704.280 ;
        RECT 1431.160 1704.000 1431.240 1704.280 ;
        RECT 1433.000 1704.000 1433.080 1704.280 ;
        RECT 1434.840 1704.000 1434.920 1704.280 ;
        RECT 1436.680 1704.000 1436.760 1704.280 ;
        RECT 1438.520 1704.000 1438.600 1704.280 ;
        RECT 1440.360 1704.000 1440.440 1704.280 ;
        RECT 1442.200 1704.000 1442.280 1704.280 ;
        RECT 1444.040 1704.000 1444.120 1704.280 ;
        RECT 1445.880 1704.000 1445.960 1704.280 ;
        RECT 1447.720 1704.000 1447.800 1704.280 ;
      LAYER met3 ;
        RECT 1160.555 1704.255 1411.585 1988.485 ;
      LAYER met4 ;
        RECT 1170.950 1710.640 1172.550 1988.560 ;
        RECT 1247.750 1710.640 1249.350 1988.560 ;
      LAYER met4 ;
        RECT 1324.550 1710.640 1354.020 1988.560 ;
        RECT 1357.020 1710.640 1372.020 1988.560 ;
        RECT 1375.020 1710.640 1390.020 1988.560 ;
        RECT 1393.020 1710.640 1402.950 1988.560 ;
  END
END user_project_wrapper
END LIBRARY

