magic
tech sky130A
magscale 1 2
timestamp 1607945491
<< obsli1 >>
rect 1086 2159 58862 57681
<< obsm1 >>
rect 180 892 59768 59152
<< metal2 >>
rect 184 59200 240 60000
rect 644 59200 700 60000
rect 1196 59200 1252 60000
rect 1748 59200 1804 60000
rect 2208 59200 2264 60000
rect 2760 59200 2816 60000
rect 3312 59200 3368 60000
rect 3864 59200 3920 60000
rect 4324 59200 4380 60000
rect 4876 59200 4932 60000
rect 5428 59200 5484 60000
rect 5888 59200 5944 60000
rect 6440 59200 6496 60000
rect 6992 59200 7048 60000
rect 7544 59200 7600 60000
rect 8004 59200 8060 60000
rect 8556 59200 8612 60000
rect 9108 59200 9164 60000
rect 9568 59200 9624 60000
rect 10120 59200 10176 60000
rect 10672 59200 10728 60000
rect 11224 59200 11280 60000
rect 11684 59200 11740 60000
rect 12236 59200 12292 60000
rect 12788 59200 12844 60000
rect 13248 59200 13304 60000
rect 13800 59200 13856 60000
rect 14352 59200 14408 60000
rect 14904 59200 14960 60000
rect 15364 59200 15420 60000
rect 15916 59200 15972 60000
rect 16468 59200 16524 60000
rect 17020 59200 17076 60000
rect 17480 59200 17536 60000
rect 18032 59200 18088 60000
rect 18584 59200 18640 60000
rect 19044 59200 19100 60000
rect 19596 59200 19652 60000
rect 20148 59200 20204 60000
rect 20700 59200 20756 60000
rect 21160 59200 21216 60000
rect 21712 59200 21768 60000
rect 22264 59200 22320 60000
rect 22724 59200 22780 60000
rect 23276 59200 23332 60000
rect 23828 59200 23884 60000
rect 24380 59200 24436 60000
rect 24840 59200 24896 60000
rect 25392 59200 25448 60000
rect 25944 59200 26000 60000
rect 26404 59200 26460 60000
rect 26956 59200 27012 60000
rect 27508 59200 27564 60000
rect 28060 59200 28116 60000
rect 28520 59200 28576 60000
rect 29072 59200 29128 60000
rect 29624 59200 29680 60000
rect 30176 59200 30232 60000
rect 30636 59200 30692 60000
rect 31188 59200 31244 60000
rect 31740 59200 31796 60000
rect 32200 59200 32256 60000
rect 32752 59200 32808 60000
rect 33304 59200 33360 60000
rect 33856 59200 33912 60000
rect 34316 59200 34372 60000
rect 34868 59200 34924 60000
rect 35420 59200 35476 60000
rect 35880 59200 35936 60000
rect 36432 59200 36488 60000
rect 36984 59200 37040 60000
rect 37536 59200 37592 60000
rect 37996 59200 38052 60000
rect 38548 59200 38604 60000
rect 39100 59200 39156 60000
rect 39560 59200 39616 60000
rect 40112 59200 40168 60000
rect 40664 59200 40720 60000
rect 41216 59200 41272 60000
rect 41676 59200 41732 60000
rect 42228 59200 42284 60000
rect 42780 59200 42836 60000
rect 43240 59200 43296 60000
rect 43792 59200 43848 60000
rect 44344 59200 44400 60000
rect 44896 59200 44952 60000
rect 45356 59200 45412 60000
rect 45908 59200 45964 60000
rect 46460 59200 46516 60000
rect 47012 59200 47068 60000
rect 47472 59200 47528 60000
rect 48024 59200 48080 60000
rect 48576 59200 48632 60000
rect 49036 59200 49092 60000
rect 49588 59200 49644 60000
rect 50140 59200 50196 60000
rect 50692 59200 50748 60000
rect 51152 59200 51208 60000
rect 51704 59200 51760 60000
rect 52256 59200 52312 60000
rect 52716 59200 52772 60000
rect 53268 59200 53324 60000
rect 53820 59200 53876 60000
rect 54372 59200 54428 60000
rect 54832 59200 54888 60000
rect 55384 59200 55440 60000
rect 55936 59200 55992 60000
rect 56396 59200 56452 60000
rect 56948 59200 57004 60000
rect 57500 59200 57556 60000
rect 58052 59200 58108 60000
rect 58512 59200 58568 60000
rect 59064 59200 59120 60000
rect 59616 59200 59672 60000
rect 0 0 56 800
rect 92 0 148 800
rect 184 0 240 800
rect 276 0 332 800
rect 460 0 516 800
rect 552 0 608 800
rect 644 0 700 800
rect 828 0 884 800
rect 920 0 976 800
rect 1012 0 1068 800
rect 1196 0 1252 800
rect 1288 0 1344 800
rect 1380 0 1436 800
rect 1564 0 1620 800
rect 1656 0 1712 800
rect 1748 0 1804 800
rect 1932 0 1988 800
rect 2024 0 2080 800
rect 2116 0 2172 800
rect 2300 0 2356 800
rect 2392 0 2448 800
rect 2484 0 2540 800
rect 2668 0 2724 800
rect 2760 0 2816 800
rect 2852 0 2908 800
rect 3036 0 3092 800
rect 3128 0 3184 800
rect 3220 0 3276 800
rect 3404 0 3460 800
rect 3496 0 3552 800
rect 3588 0 3644 800
rect 3772 0 3828 800
rect 3864 0 3920 800
rect 3956 0 4012 800
rect 4140 0 4196 800
rect 4232 0 4288 800
rect 4324 0 4380 800
rect 4508 0 4564 800
rect 4600 0 4656 800
rect 4692 0 4748 800
rect 4876 0 4932 800
rect 4968 0 5024 800
rect 5060 0 5116 800
rect 5244 0 5300 800
rect 5336 0 5392 800
rect 5428 0 5484 800
rect 5612 0 5668 800
rect 5704 0 5760 800
rect 5796 0 5852 800
rect 5980 0 6036 800
rect 6072 0 6128 800
rect 6164 0 6220 800
rect 6348 0 6404 800
rect 6440 0 6496 800
rect 6532 0 6588 800
rect 6716 0 6772 800
rect 6808 0 6864 800
rect 6900 0 6956 800
rect 7084 0 7140 800
rect 7176 0 7232 800
rect 7268 0 7324 800
rect 7452 0 7508 800
rect 7544 0 7600 800
rect 7636 0 7692 800
rect 7820 0 7876 800
rect 7912 0 7968 800
rect 8004 0 8060 800
rect 8188 0 8244 800
rect 8280 0 8336 800
rect 8372 0 8428 800
rect 8556 0 8612 800
rect 8648 0 8704 800
rect 8740 0 8796 800
rect 8924 0 8980 800
rect 9016 0 9072 800
rect 9108 0 9164 800
rect 9292 0 9348 800
rect 9384 0 9440 800
rect 9476 0 9532 800
rect 9660 0 9716 800
rect 9752 0 9808 800
rect 9844 0 9900 800
rect 10028 0 10084 800
rect 10120 0 10176 800
rect 10212 0 10268 800
rect 10396 0 10452 800
rect 10488 0 10544 800
rect 10580 0 10636 800
rect 10764 0 10820 800
rect 10856 0 10912 800
rect 10948 0 11004 800
rect 11132 0 11188 800
rect 11224 0 11280 800
rect 11316 0 11372 800
rect 11500 0 11556 800
rect 11592 0 11648 800
rect 11684 0 11740 800
rect 11868 0 11924 800
rect 11960 0 12016 800
rect 12052 0 12108 800
rect 12236 0 12292 800
rect 12328 0 12384 800
rect 12420 0 12476 800
rect 12604 0 12660 800
rect 12696 0 12752 800
rect 12788 0 12844 800
rect 12972 0 13028 800
rect 13064 0 13120 800
rect 13156 0 13212 800
rect 13340 0 13396 800
rect 13432 0 13488 800
rect 13524 0 13580 800
rect 13708 0 13764 800
rect 13800 0 13856 800
rect 13892 0 13948 800
rect 14076 0 14132 800
rect 14168 0 14224 800
rect 14260 0 14316 800
rect 14444 0 14500 800
rect 14536 0 14592 800
rect 14628 0 14684 800
rect 14812 0 14868 800
rect 14904 0 14960 800
rect 14996 0 15052 800
rect 15088 0 15144 800
rect 15272 0 15328 800
rect 15364 0 15420 800
rect 15456 0 15512 800
rect 15640 0 15696 800
rect 15732 0 15788 800
rect 15824 0 15880 800
rect 16008 0 16064 800
rect 16100 0 16156 800
rect 16192 0 16248 800
rect 16376 0 16432 800
rect 16468 0 16524 800
rect 16560 0 16616 800
rect 16744 0 16800 800
rect 16836 0 16892 800
rect 16928 0 16984 800
rect 17112 0 17168 800
rect 17204 0 17260 800
rect 17296 0 17352 800
rect 17480 0 17536 800
rect 17572 0 17628 800
rect 17664 0 17720 800
rect 17848 0 17904 800
rect 17940 0 17996 800
rect 18032 0 18088 800
rect 18216 0 18272 800
rect 18308 0 18364 800
rect 18400 0 18456 800
rect 18584 0 18640 800
rect 18676 0 18732 800
rect 18768 0 18824 800
rect 18952 0 19008 800
rect 19044 0 19100 800
rect 19136 0 19192 800
rect 19320 0 19376 800
rect 19412 0 19468 800
rect 19504 0 19560 800
rect 19688 0 19744 800
rect 19780 0 19836 800
rect 19872 0 19928 800
rect 20056 0 20112 800
rect 20148 0 20204 800
rect 20240 0 20296 800
rect 20424 0 20480 800
rect 20516 0 20572 800
rect 20608 0 20664 800
rect 20792 0 20848 800
rect 20884 0 20940 800
rect 20976 0 21032 800
rect 21160 0 21216 800
rect 21252 0 21308 800
rect 21344 0 21400 800
rect 21528 0 21584 800
rect 21620 0 21676 800
rect 21712 0 21768 800
rect 21896 0 21952 800
rect 21988 0 22044 800
rect 22080 0 22136 800
rect 22264 0 22320 800
rect 22356 0 22412 800
rect 22448 0 22504 800
rect 22632 0 22688 800
rect 22724 0 22780 800
rect 22816 0 22872 800
rect 23000 0 23056 800
rect 23092 0 23148 800
rect 23184 0 23240 800
rect 23368 0 23424 800
rect 23460 0 23516 800
rect 23552 0 23608 800
rect 23736 0 23792 800
rect 23828 0 23884 800
rect 23920 0 23976 800
rect 24104 0 24160 800
rect 24196 0 24252 800
rect 24288 0 24344 800
rect 24472 0 24528 800
rect 24564 0 24620 800
rect 24656 0 24712 800
rect 24840 0 24896 800
rect 24932 0 24988 800
rect 25024 0 25080 800
rect 25208 0 25264 800
rect 25300 0 25356 800
rect 25392 0 25448 800
rect 25576 0 25632 800
rect 25668 0 25724 800
rect 25760 0 25816 800
rect 25944 0 26000 800
rect 26036 0 26092 800
rect 26128 0 26184 800
rect 26312 0 26368 800
rect 26404 0 26460 800
rect 26496 0 26552 800
rect 26680 0 26736 800
rect 26772 0 26828 800
rect 26864 0 26920 800
rect 27048 0 27104 800
rect 27140 0 27196 800
rect 27232 0 27288 800
rect 27416 0 27472 800
rect 27508 0 27564 800
rect 27600 0 27656 800
rect 27784 0 27840 800
rect 27876 0 27932 800
rect 27968 0 28024 800
rect 28152 0 28208 800
rect 28244 0 28300 800
rect 28336 0 28392 800
rect 28520 0 28576 800
rect 28612 0 28668 800
rect 28704 0 28760 800
rect 28888 0 28944 800
rect 28980 0 29036 800
rect 29072 0 29128 800
rect 29256 0 29312 800
rect 29348 0 29404 800
rect 29440 0 29496 800
rect 29624 0 29680 800
rect 29716 0 29772 800
rect 29808 0 29864 800
rect 29992 0 30048 800
rect 30084 0 30140 800
rect 30176 0 30232 800
rect 30268 0 30324 800
rect 30452 0 30508 800
rect 30544 0 30600 800
rect 30636 0 30692 800
rect 30820 0 30876 800
rect 30912 0 30968 800
rect 31004 0 31060 800
rect 31188 0 31244 800
rect 31280 0 31336 800
rect 31372 0 31428 800
rect 31556 0 31612 800
rect 31648 0 31704 800
rect 31740 0 31796 800
rect 31924 0 31980 800
rect 32016 0 32072 800
rect 32108 0 32164 800
rect 32292 0 32348 800
rect 32384 0 32440 800
rect 32476 0 32532 800
rect 32660 0 32716 800
rect 32752 0 32808 800
rect 32844 0 32900 800
rect 33028 0 33084 800
rect 33120 0 33176 800
rect 33212 0 33268 800
rect 33396 0 33452 800
rect 33488 0 33544 800
rect 33580 0 33636 800
rect 33764 0 33820 800
rect 33856 0 33912 800
rect 33948 0 34004 800
rect 34132 0 34188 800
rect 34224 0 34280 800
rect 34316 0 34372 800
rect 34500 0 34556 800
rect 34592 0 34648 800
rect 34684 0 34740 800
rect 34868 0 34924 800
rect 34960 0 35016 800
rect 35052 0 35108 800
rect 35236 0 35292 800
rect 35328 0 35384 800
rect 35420 0 35476 800
rect 35604 0 35660 800
rect 35696 0 35752 800
rect 35788 0 35844 800
rect 35972 0 36028 800
rect 36064 0 36120 800
rect 36156 0 36212 800
rect 36340 0 36396 800
rect 36432 0 36488 800
rect 36524 0 36580 800
rect 36708 0 36764 800
rect 36800 0 36856 800
rect 36892 0 36948 800
rect 37076 0 37132 800
rect 37168 0 37224 800
rect 37260 0 37316 800
rect 37444 0 37500 800
rect 37536 0 37592 800
rect 37628 0 37684 800
rect 37812 0 37868 800
rect 37904 0 37960 800
rect 37996 0 38052 800
rect 38180 0 38236 800
rect 38272 0 38328 800
rect 38364 0 38420 800
rect 38548 0 38604 800
rect 38640 0 38696 800
rect 38732 0 38788 800
rect 38916 0 38972 800
rect 39008 0 39064 800
rect 39100 0 39156 800
rect 39284 0 39340 800
rect 39376 0 39432 800
rect 39468 0 39524 800
rect 39652 0 39708 800
rect 39744 0 39800 800
rect 39836 0 39892 800
rect 40020 0 40076 800
rect 40112 0 40168 800
rect 40204 0 40260 800
rect 40388 0 40444 800
rect 40480 0 40536 800
rect 40572 0 40628 800
rect 40756 0 40812 800
rect 40848 0 40904 800
rect 40940 0 40996 800
rect 41124 0 41180 800
rect 41216 0 41272 800
rect 41308 0 41364 800
rect 41492 0 41548 800
rect 41584 0 41640 800
rect 41676 0 41732 800
rect 41860 0 41916 800
rect 41952 0 42008 800
rect 42044 0 42100 800
rect 42228 0 42284 800
rect 42320 0 42376 800
rect 42412 0 42468 800
rect 42596 0 42652 800
rect 42688 0 42744 800
rect 42780 0 42836 800
rect 42964 0 43020 800
rect 43056 0 43112 800
rect 43148 0 43204 800
rect 43332 0 43388 800
rect 43424 0 43480 800
rect 43516 0 43572 800
rect 43700 0 43756 800
rect 43792 0 43848 800
rect 43884 0 43940 800
rect 44068 0 44124 800
rect 44160 0 44216 800
rect 44252 0 44308 800
rect 44436 0 44492 800
rect 44528 0 44584 800
rect 44620 0 44676 800
rect 44804 0 44860 800
rect 44896 0 44952 800
rect 44988 0 45044 800
rect 45080 0 45136 800
rect 45264 0 45320 800
rect 45356 0 45412 800
rect 45448 0 45504 800
rect 45632 0 45688 800
rect 45724 0 45780 800
rect 45816 0 45872 800
rect 46000 0 46056 800
rect 46092 0 46148 800
rect 46184 0 46240 800
rect 46368 0 46424 800
rect 46460 0 46516 800
rect 46552 0 46608 800
rect 46736 0 46792 800
rect 46828 0 46884 800
rect 46920 0 46976 800
rect 47104 0 47160 800
rect 47196 0 47252 800
rect 47288 0 47344 800
rect 47472 0 47528 800
rect 47564 0 47620 800
rect 47656 0 47712 800
rect 47840 0 47896 800
rect 47932 0 47988 800
rect 48024 0 48080 800
rect 48208 0 48264 800
rect 48300 0 48356 800
rect 48392 0 48448 800
rect 48576 0 48632 800
rect 48668 0 48724 800
rect 48760 0 48816 800
rect 48944 0 49000 800
rect 49036 0 49092 800
rect 49128 0 49184 800
rect 49312 0 49368 800
rect 49404 0 49460 800
rect 49496 0 49552 800
rect 49680 0 49736 800
rect 49772 0 49828 800
rect 49864 0 49920 800
rect 50048 0 50104 800
rect 50140 0 50196 800
rect 50232 0 50288 800
rect 50416 0 50472 800
rect 50508 0 50564 800
rect 50600 0 50656 800
rect 50784 0 50840 800
rect 50876 0 50932 800
rect 50968 0 51024 800
rect 51152 0 51208 800
rect 51244 0 51300 800
rect 51336 0 51392 800
rect 51520 0 51576 800
rect 51612 0 51668 800
rect 51704 0 51760 800
rect 51888 0 51944 800
rect 51980 0 52036 800
rect 52072 0 52128 800
rect 52256 0 52312 800
rect 52348 0 52404 800
rect 52440 0 52496 800
rect 52624 0 52680 800
rect 52716 0 52772 800
rect 52808 0 52864 800
rect 52992 0 53048 800
rect 53084 0 53140 800
rect 53176 0 53232 800
rect 53360 0 53416 800
rect 53452 0 53508 800
rect 53544 0 53600 800
rect 53728 0 53784 800
rect 53820 0 53876 800
rect 53912 0 53968 800
rect 54096 0 54152 800
rect 54188 0 54244 800
rect 54280 0 54336 800
rect 54464 0 54520 800
rect 54556 0 54612 800
rect 54648 0 54704 800
rect 54832 0 54888 800
rect 54924 0 54980 800
rect 55016 0 55072 800
rect 55200 0 55256 800
rect 55292 0 55348 800
rect 55384 0 55440 800
rect 55568 0 55624 800
rect 55660 0 55716 800
rect 55752 0 55808 800
rect 55936 0 55992 800
rect 56028 0 56084 800
rect 56120 0 56176 800
rect 56304 0 56360 800
rect 56396 0 56452 800
rect 56488 0 56544 800
rect 56672 0 56728 800
rect 56764 0 56820 800
rect 56856 0 56912 800
rect 57040 0 57096 800
rect 57132 0 57188 800
rect 57224 0 57280 800
rect 57408 0 57464 800
rect 57500 0 57556 800
rect 57592 0 57648 800
rect 57776 0 57832 800
rect 57868 0 57924 800
rect 57960 0 58016 800
rect 58144 0 58200 800
rect 58236 0 58292 800
rect 58328 0 58384 800
rect 58512 0 58568 800
rect 58604 0 58660 800
rect 58696 0 58752 800
rect 58880 0 58936 800
rect 58972 0 59028 800
rect 59064 0 59120 800
rect 59248 0 59304 800
rect 59340 0 59396 800
rect 59432 0 59488 800
rect 59616 0 59672 800
rect 59708 0 59764 800
rect 59800 0 59856 800
<< obsm2 >>
rect 296 59144 588 59200
rect 756 59144 1140 59200
rect 1308 59144 1692 59200
rect 1860 59144 2152 59200
rect 2320 59144 2704 59200
rect 2872 59144 3256 59200
rect 3424 59144 3808 59200
rect 3976 59144 4268 59200
rect 4436 59144 4820 59200
rect 4988 59144 5372 59200
rect 5540 59144 5832 59200
rect 6000 59144 6384 59200
rect 6552 59144 6936 59200
rect 7104 59144 7488 59200
rect 7656 59144 7948 59200
rect 8116 59144 8500 59200
rect 8668 59144 9052 59200
rect 9220 59144 9512 59200
rect 9680 59144 10064 59200
rect 10232 59144 10616 59200
rect 10784 59144 11168 59200
rect 11336 59144 11628 59200
rect 11796 59144 12180 59200
rect 12348 59144 12732 59200
rect 12900 59144 13192 59200
rect 13360 59144 13744 59200
rect 13912 59144 14296 59200
rect 14464 59144 14848 59200
rect 15016 59144 15308 59200
rect 15476 59144 15860 59200
rect 16028 59144 16412 59200
rect 16580 59144 16964 59200
rect 17132 59144 17424 59200
rect 17592 59144 17976 59200
rect 18144 59144 18528 59200
rect 18696 59144 18988 59200
rect 19156 59144 19540 59200
rect 19708 59144 20092 59200
rect 20260 59144 20644 59200
rect 20812 59144 21104 59200
rect 21272 59144 21656 59200
rect 21824 59144 22208 59200
rect 22376 59144 22668 59200
rect 22836 59144 23220 59200
rect 23388 59144 23772 59200
rect 23940 59144 24324 59200
rect 24492 59144 24784 59200
rect 24952 59144 25336 59200
rect 25504 59144 25888 59200
rect 26056 59144 26348 59200
rect 26516 59144 26900 59200
rect 27068 59144 27452 59200
rect 27620 59144 28004 59200
rect 28172 59144 28464 59200
rect 28632 59144 29016 59200
rect 29184 59144 29568 59200
rect 29736 59144 30120 59200
rect 30288 59144 30580 59200
rect 30748 59144 31132 59200
rect 31300 59144 31684 59200
rect 31852 59144 32144 59200
rect 32312 59144 32696 59200
rect 32864 59144 33248 59200
rect 33416 59144 33800 59200
rect 33968 59144 34260 59200
rect 34428 59144 34812 59200
rect 34980 59144 35364 59200
rect 35532 59144 35824 59200
rect 35992 59144 36376 59200
rect 36544 59144 36928 59200
rect 37096 59144 37480 59200
rect 37648 59144 37940 59200
rect 38108 59144 38492 59200
rect 38660 59144 39044 59200
rect 39212 59144 39504 59200
rect 39672 59144 40056 59200
rect 40224 59144 40608 59200
rect 40776 59144 41160 59200
rect 41328 59144 41620 59200
rect 41788 59144 42172 59200
rect 42340 59144 42724 59200
rect 42892 59144 43184 59200
rect 43352 59144 43736 59200
rect 43904 59144 44288 59200
rect 44456 59144 44840 59200
rect 45008 59144 45300 59200
rect 45468 59144 45852 59200
rect 46020 59144 46404 59200
rect 46572 59144 46956 59200
rect 47124 59144 47416 59200
rect 47584 59144 47968 59200
rect 48136 59144 48520 59200
rect 48688 59144 48980 59200
rect 49148 59144 49532 59200
rect 49700 59144 50084 59200
rect 50252 59144 50636 59200
rect 50804 59144 51096 59200
rect 51264 59144 51648 59200
rect 51816 59144 52200 59200
rect 52368 59144 52660 59200
rect 52828 59144 53212 59200
rect 53380 59144 53764 59200
rect 53932 59144 54316 59200
rect 54484 59144 54776 59200
rect 54944 59144 55328 59200
rect 55496 59144 55880 59200
rect 56048 59144 56340 59200
rect 56508 59144 56892 59200
rect 57060 59144 57444 59200
rect 57612 59144 57996 59200
rect 58164 59144 58456 59200
rect 58624 59144 59008 59200
rect 59176 59144 59560 59200
rect 59728 59144 59762 59200
rect 186 856 59762 59144
rect 388 800 404 856
rect 756 800 772 856
rect 1124 800 1140 856
rect 1492 800 1508 856
rect 1860 800 1876 856
rect 2228 800 2244 856
rect 2596 800 2612 856
rect 2964 800 2980 856
rect 3332 800 3348 856
rect 3700 800 3716 856
rect 4068 800 4084 856
rect 4436 800 4452 856
rect 4804 800 4820 856
rect 5172 800 5188 856
rect 5540 800 5556 856
rect 5908 800 5924 856
rect 6276 800 6292 856
rect 6644 800 6660 856
rect 7012 800 7028 856
rect 7380 800 7396 856
rect 7748 800 7764 856
rect 8116 800 8132 856
rect 8484 800 8500 856
rect 8852 800 8868 856
rect 9220 800 9236 856
rect 9588 800 9604 856
rect 9956 800 9972 856
rect 10324 800 10340 856
rect 10692 800 10708 856
rect 11060 800 11076 856
rect 11428 800 11444 856
rect 11796 800 11812 856
rect 12164 800 12180 856
rect 12532 800 12548 856
rect 12900 800 12916 856
rect 13268 800 13284 856
rect 13636 800 13652 856
rect 14004 800 14020 856
rect 14372 800 14388 856
rect 14740 800 14756 856
rect 15200 800 15216 856
rect 15568 800 15584 856
rect 15936 800 15952 856
rect 16304 800 16320 856
rect 16672 800 16688 856
rect 17040 800 17056 856
rect 17408 800 17424 856
rect 17776 800 17792 856
rect 18144 800 18160 856
rect 18512 800 18528 856
rect 18880 800 18896 856
rect 19248 800 19264 856
rect 19616 800 19632 856
rect 19984 800 20000 856
rect 20352 800 20368 856
rect 20720 800 20736 856
rect 21088 800 21104 856
rect 21456 800 21472 856
rect 21824 800 21840 856
rect 22192 800 22208 856
rect 22560 800 22576 856
rect 22928 800 22944 856
rect 23296 800 23312 856
rect 23664 800 23680 856
rect 24032 800 24048 856
rect 24400 800 24416 856
rect 24768 800 24784 856
rect 25136 800 25152 856
rect 25504 800 25520 856
rect 25872 800 25888 856
rect 26240 800 26256 856
rect 26608 800 26624 856
rect 26976 800 26992 856
rect 27344 800 27360 856
rect 27712 800 27728 856
rect 28080 800 28096 856
rect 28448 800 28464 856
rect 28816 800 28832 856
rect 29184 800 29200 856
rect 29552 800 29568 856
rect 29920 800 29936 856
rect 30380 800 30396 856
rect 30748 800 30764 856
rect 31116 800 31132 856
rect 31484 800 31500 856
rect 31852 800 31868 856
rect 32220 800 32236 856
rect 32588 800 32604 856
rect 32956 800 32972 856
rect 33324 800 33340 856
rect 33692 800 33708 856
rect 34060 800 34076 856
rect 34428 800 34444 856
rect 34796 800 34812 856
rect 35164 800 35180 856
rect 35532 800 35548 856
rect 35900 800 35916 856
rect 36268 800 36284 856
rect 36636 800 36652 856
rect 37004 800 37020 856
rect 37372 800 37388 856
rect 37740 800 37756 856
rect 38108 800 38124 856
rect 38476 800 38492 856
rect 38844 800 38860 856
rect 39212 800 39228 856
rect 39580 800 39596 856
rect 39948 800 39964 856
rect 40316 800 40332 856
rect 40684 800 40700 856
rect 41052 800 41068 856
rect 41420 800 41436 856
rect 41788 800 41804 856
rect 42156 800 42172 856
rect 42524 800 42540 856
rect 42892 800 42908 856
rect 43260 800 43276 856
rect 43628 800 43644 856
rect 43996 800 44012 856
rect 44364 800 44380 856
rect 44732 800 44748 856
rect 45192 800 45208 856
rect 45560 800 45576 856
rect 45928 800 45944 856
rect 46296 800 46312 856
rect 46664 800 46680 856
rect 47032 800 47048 856
rect 47400 800 47416 856
rect 47768 800 47784 856
rect 48136 800 48152 856
rect 48504 800 48520 856
rect 48872 800 48888 856
rect 49240 800 49256 856
rect 49608 800 49624 856
rect 49976 800 49992 856
rect 50344 800 50360 856
rect 50712 800 50728 856
rect 51080 800 51096 856
rect 51448 800 51464 856
rect 51816 800 51832 856
rect 52184 800 52200 856
rect 52552 800 52568 856
rect 52920 800 52936 856
rect 53288 800 53304 856
rect 53656 800 53672 856
rect 54024 800 54040 856
rect 54392 800 54408 856
rect 54760 800 54776 856
rect 55128 800 55144 856
rect 55496 800 55512 856
rect 55864 800 55880 856
rect 56232 800 56248 856
rect 56600 800 56616 856
rect 56968 800 56984 856
rect 57336 800 57352 856
rect 57704 800 57720 856
rect 58072 800 58088 856
rect 58440 800 58456 856
rect 58808 800 58824 856
rect 59176 800 59192 856
rect 59544 800 59560 856
<< obsm3 >>
rect 3767 851 55169 57697
<< metal4 >>
rect 4190 2128 4510 57712
rect 19550 2128 19870 57712
<< obsm4 >>
rect 16417 2128 19470 57712
rect 19950 2128 50590 57712
<< labels >>
rlabel metal2 s 184 59200 240 60000 6 io_in[0]
port 1 nsew default input
rlabel metal2 s 15916 59200 15972 60000 6 io_in[10]
port 2 nsew default input
rlabel metal2 s 17480 59200 17536 60000 6 io_in[11]
port 3 nsew default input
rlabel metal2 s 19044 59200 19100 60000 6 io_in[12]
port 4 nsew default input
rlabel metal2 s 20700 59200 20756 60000 6 io_in[13]
port 5 nsew default input
rlabel metal2 s 22264 59200 22320 60000 6 io_in[14]
port 6 nsew default input
rlabel metal2 s 23828 59200 23884 60000 6 io_in[15]
port 7 nsew default input
rlabel metal2 s 25392 59200 25448 60000 6 io_in[16]
port 8 nsew default input
rlabel metal2 s 26956 59200 27012 60000 6 io_in[17]
port 9 nsew default input
rlabel metal2 s 28520 59200 28576 60000 6 io_in[18]
port 10 nsew default input
rlabel metal2 s 30176 59200 30232 60000 6 io_in[19]
port 11 nsew default input
rlabel metal2 s 1748 59200 1804 60000 6 io_in[1]
port 12 nsew default input
rlabel metal2 s 31740 59200 31796 60000 6 io_in[20]
port 13 nsew default input
rlabel metal2 s 33304 59200 33360 60000 6 io_in[21]
port 14 nsew default input
rlabel metal2 s 34868 59200 34924 60000 6 io_in[22]
port 15 nsew default input
rlabel metal2 s 36432 59200 36488 60000 6 io_in[23]
port 16 nsew default input
rlabel metal2 s 37996 59200 38052 60000 6 io_in[24]
port 17 nsew default input
rlabel metal2 s 39560 59200 39616 60000 6 io_in[25]
port 18 nsew default input
rlabel metal2 s 41216 59200 41272 60000 6 io_in[26]
port 19 nsew default input
rlabel metal2 s 42780 59200 42836 60000 6 io_in[27]
port 20 nsew default input
rlabel metal2 s 44344 59200 44400 60000 6 io_in[28]
port 21 nsew default input
rlabel metal2 s 45908 59200 45964 60000 6 io_in[29]
port 22 nsew default input
rlabel metal2 s 3312 59200 3368 60000 6 io_in[2]
port 23 nsew default input
rlabel metal2 s 47472 59200 47528 60000 6 io_in[30]
port 24 nsew default input
rlabel metal2 s 49036 59200 49092 60000 6 io_in[31]
port 25 nsew default input
rlabel metal2 s 50692 59200 50748 60000 6 io_in[32]
port 26 nsew default input
rlabel metal2 s 52256 59200 52312 60000 6 io_in[33]
port 27 nsew default input
rlabel metal2 s 53820 59200 53876 60000 6 io_in[34]
port 28 nsew default input
rlabel metal2 s 55384 59200 55440 60000 6 io_in[35]
port 29 nsew default input
rlabel metal2 s 56948 59200 57004 60000 6 io_in[36]
port 30 nsew default input
rlabel metal2 s 58512 59200 58568 60000 6 io_in[37]
port 31 nsew default input
rlabel metal2 s 4876 59200 4932 60000 6 io_in[3]
port 32 nsew default input
rlabel metal2 s 6440 59200 6496 60000 6 io_in[4]
port 33 nsew default input
rlabel metal2 s 8004 59200 8060 60000 6 io_in[5]
port 34 nsew default input
rlabel metal2 s 9568 59200 9624 60000 6 io_in[6]
port 35 nsew default input
rlabel metal2 s 11224 59200 11280 60000 6 io_in[7]
port 36 nsew default input
rlabel metal2 s 12788 59200 12844 60000 6 io_in[8]
port 37 nsew default input
rlabel metal2 s 14352 59200 14408 60000 6 io_in[9]
port 38 nsew default input
rlabel metal2 s 644 59200 700 60000 6 io_oeb[0]
port 39 nsew default output
rlabel metal2 s 16468 59200 16524 60000 6 io_oeb[10]
port 40 nsew default output
rlabel metal2 s 18032 59200 18088 60000 6 io_oeb[11]
port 41 nsew default output
rlabel metal2 s 19596 59200 19652 60000 6 io_oeb[12]
port 42 nsew default output
rlabel metal2 s 21160 59200 21216 60000 6 io_oeb[13]
port 43 nsew default output
rlabel metal2 s 22724 59200 22780 60000 6 io_oeb[14]
port 44 nsew default output
rlabel metal2 s 24380 59200 24436 60000 6 io_oeb[15]
port 45 nsew default output
rlabel metal2 s 25944 59200 26000 60000 6 io_oeb[16]
port 46 nsew default output
rlabel metal2 s 27508 59200 27564 60000 6 io_oeb[17]
port 47 nsew default output
rlabel metal2 s 29072 59200 29128 60000 6 io_oeb[18]
port 48 nsew default output
rlabel metal2 s 30636 59200 30692 60000 6 io_oeb[19]
port 49 nsew default output
rlabel metal2 s 2208 59200 2264 60000 6 io_oeb[1]
port 50 nsew default output
rlabel metal2 s 32200 59200 32256 60000 6 io_oeb[20]
port 51 nsew default output
rlabel metal2 s 33856 59200 33912 60000 6 io_oeb[21]
port 52 nsew default output
rlabel metal2 s 35420 59200 35476 60000 6 io_oeb[22]
port 53 nsew default output
rlabel metal2 s 36984 59200 37040 60000 6 io_oeb[23]
port 54 nsew default output
rlabel metal2 s 38548 59200 38604 60000 6 io_oeb[24]
port 55 nsew default output
rlabel metal2 s 40112 59200 40168 60000 6 io_oeb[25]
port 56 nsew default output
rlabel metal2 s 41676 59200 41732 60000 6 io_oeb[26]
port 57 nsew default output
rlabel metal2 s 43240 59200 43296 60000 6 io_oeb[27]
port 58 nsew default output
rlabel metal2 s 44896 59200 44952 60000 6 io_oeb[28]
port 59 nsew default output
rlabel metal2 s 46460 59200 46516 60000 6 io_oeb[29]
port 60 nsew default output
rlabel metal2 s 3864 59200 3920 60000 6 io_oeb[2]
port 61 nsew default output
rlabel metal2 s 48024 59200 48080 60000 6 io_oeb[30]
port 62 nsew default output
rlabel metal2 s 49588 59200 49644 60000 6 io_oeb[31]
port 63 nsew default output
rlabel metal2 s 51152 59200 51208 60000 6 io_oeb[32]
port 64 nsew default output
rlabel metal2 s 52716 59200 52772 60000 6 io_oeb[33]
port 65 nsew default output
rlabel metal2 s 54372 59200 54428 60000 6 io_oeb[34]
port 66 nsew default output
rlabel metal2 s 55936 59200 55992 60000 6 io_oeb[35]
port 67 nsew default output
rlabel metal2 s 57500 59200 57556 60000 6 io_oeb[36]
port 68 nsew default output
rlabel metal2 s 59064 59200 59120 60000 6 io_oeb[37]
port 69 nsew default output
rlabel metal2 s 5428 59200 5484 60000 6 io_oeb[3]
port 70 nsew default output
rlabel metal2 s 6992 59200 7048 60000 6 io_oeb[4]
port 71 nsew default output
rlabel metal2 s 8556 59200 8612 60000 6 io_oeb[5]
port 72 nsew default output
rlabel metal2 s 10120 59200 10176 60000 6 io_oeb[6]
port 73 nsew default output
rlabel metal2 s 11684 59200 11740 60000 6 io_oeb[7]
port 74 nsew default output
rlabel metal2 s 13248 59200 13304 60000 6 io_oeb[8]
port 75 nsew default output
rlabel metal2 s 14904 59200 14960 60000 6 io_oeb[9]
port 76 nsew default output
rlabel metal2 s 1196 59200 1252 60000 6 io_out[0]
port 77 nsew default output
rlabel metal2 s 17020 59200 17076 60000 6 io_out[10]
port 78 nsew default output
rlabel metal2 s 18584 59200 18640 60000 6 io_out[11]
port 79 nsew default output
rlabel metal2 s 20148 59200 20204 60000 6 io_out[12]
port 80 nsew default output
rlabel metal2 s 21712 59200 21768 60000 6 io_out[13]
port 81 nsew default output
rlabel metal2 s 23276 59200 23332 60000 6 io_out[14]
port 82 nsew default output
rlabel metal2 s 24840 59200 24896 60000 6 io_out[15]
port 83 nsew default output
rlabel metal2 s 26404 59200 26460 60000 6 io_out[16]
port 84 nsew default output
rlabel metal2 s 28060 59200 28116 60000 6 io_out[17]
port 85 nsew default output
rlabel metal2 s 29624 59200 29680 60000 6 io_out[18]
port 86 nsew default output
rlabel metal2 s 31188 59200 31244 60000 6 io_out[19]
port 87 nsew default output
rlabel metal2 s 2760 59200 2816 60000 6 io_out[1]
port 88 nsew default output
rlabel metal2 s 32752 59200 32808 60000 6 io_out[20]
port 89 nsew default output
rlabel metal2 s 34316 59200 34372 60000 6 io_out[21]
port 90 nsew default output
rlabel metal2 s 35880 59200 35936 60000 6 io_out[22]
port 91 nsew default output
rlabel metal2 s 37536 59200 37592 60000 6 io_out[23]
port 92 nsew default output
rlabel metal2 s 39100 59200 39156 60000 6 io_out[24]
port 93 nsew default output
rlabel metal2 s 40664 59200 40720 60000 6 io_out[25]
port 94 nsew default output
rlabel metal2 s 42228 59200 42284 60000 6 io_out[26]
port 95 nsew default output
rlabel metal2 s 43792 59200 43848 60000 6 io_out[27]
port 96 nsew default output
rlabel metal2 s 45356 59200 45412 60000 6 io_out[28]
port 97 nsew default output
rlabel metal2 s 47012 59200 47068 60000 6 io_out[29]
port 98 nsew default output
rlabel metal2 s 4324 59200 4380 60000 6 io_out[2]
port 99 nsew default output
rlabel metal2 s 48576 59200 48632 60000 6 io_out[30]
port 100 nsew default output
rlabel metal2 s 50140 59200 50196 60000 6 io_out[31]
port 101 nsew default output
rlabel metal2 s 51704 59200 51760 60000 6 io_out[32]
port 102 nsew default output
rlabel metal2 s 53268 59200 53324 60000 6 io_out[33]
port 103 nsew default output
rlabel metal2 s 54832 59200 54888 60000 6 io_out[34]
port 104 nsew default output
rlabel metal2 s 56396 59200 56452 60000 6 io_out[35]
port 105 nsew default output
rlabel metal2 s 58052 59200 58108 60000 6 io_out[36]
port 106 nsew default output
rlabel metal2 s 59616 59200 59672 60000 6 io_out[37]
port 107 nsew default output
rlabel metal2 s 5888 59200 5944 60000 6 io_out[3]
port 108 nsew default output
rlabel metal2 s 7544 59200 7600 60000 6 io_out[4]
port 109 nsew default output
rlabel metal2 s 9108 59200 9164 60000 6 io_out[5]
port 110 nsew default output
rlabel metal2 s 10672 59200 10728 60000 6 io_out[6]
port 111 nsew default output
rlabel metal2 s 12236 59200 12292 60000 6 io_out[7]
port 112 nsew default output
rlabel metal2 s 13800 59200 13856 60000 6 io_out[8]
port 113 nsew default output
rlabel metal2 s 15364 59200 15420 60000 6 io_out[9]
port 114 nsew default output
rlabel metal2 s 12972 0 13028 800 6 la_data_in[0]
port 115 nsew default input
rlabel metal2 s 49680 0 49736 800 6 la_data_in[100]
port 116 nsew default input
rlabel metal2 s 50048 0 50104 800 6 la_data_in[101]
port 117 nsew default input
rlabel metal2 s 50416 0 50472 800 6 la_data_in[102]
port 118 nsew default input
rlabel metal2 s 50784 0 50840 800 6 la_data_in[103]
port 119 nsew default input
rlabel metal2 s 51152 0 51208 800 6 la_data_in[104]
port 120 nsew default input
rlabel metal2 s 51520 0 51576 800 6 la_data_in[105]
port 121 nsew default input
rlabel metal2 s 51888 0 51944 800 6 la_data_in[106]
port 122 nsew default input
rlabel metal2 s 52256 0 52312 800 6 la_data_in[107]
port 123 nsew default input
rlabel metal2 s 52624 0 52680 800 6 la_data_in[108]
port 124 nsew default input
rlabel metal2 s 52992 0 53048 800 6 la_data_in[109]
port 125 nsew default input
rlabel metal2 s 16560 0 16616 800 6 la_data_in[10]
port 126 nsew default input
rlabel metal2 s 53360 0 53416 800 6 la_data_in[110]
port 127 nsew default input
rlabel metal2 s 53728 0 53784 800 6 la_data_in[111]
port 128 nsew default input
rlabel metal2 s 54096 0 54152 800 6 la_data_in[112]
port 129 nsew default input
rlabel metal2 s 54464 0 54520 800 6 la_data_in[113]
port 130 nsew default input
rlabel metal2 s 54832 0 54888 800 6 la_data_in[114]
port 131 nsew default input
rlabel metal2 s 55200 0 55256 800 6 la_data_in[115]
port 132 nsew default input
rlabel metal2 s 55568 0 55624 800 6 la_data_in[116]
port 133 nsew default input
rlabel metal2 s 55936 0 55992 800 6 la_data_in[117]
port 134 nsew default input
rlabel metal2 s 56304 0 56360 800 6 la_data_in[118]
port 135 nsew default input
rlabel metal2 s 56672 0 56728 800 6 la_data_in[119]
port 136 nsew default input
rlabel metal2 s 16928 0 16984 800 6 la_data_in[11]
port 137 nsew default input
rlabel metal2 s 57040 0 57096 800 6 la_data_in[120]
port 138 nsew default input
rlabel metal2 s 57408 0 57464 800 6 la_data_in[121]
port 139 nsew default input
rlabel metal2 s 57776 0 57832 800 6 la_data_in[122]
port 140 nsew default input
rlabel metal2 s 58144 0 58200 800 6 la_data_in[123]
port 141 nsew default input
rlabel metal2 s 58512 0 58568 800 6 la_data_in[124]
port 142 nsew default input
rlabel metal2 s 58880 0 58936 800 6 la_data_in[125]
port 143 nsew default input
rlabel metal2 s 59248 0 59304 800 6 la_data_in[126]
port 144 nsew default input
rlabel metal2 s 59616 0 59672 800 6 la_data_in[127]
port 145 nsew default input
rlabel metal2 s 17296 0 17352 800 6 la_data_in[12]
port 146 nsew default input
rlabel metal2 s 17664 0 17720 800 6 la_data_in[13]
port 147 nsew default input
rlabel metal2 s 18032 0 18088 800 6 la_data_in[14]
port 148 nsew default input
rlabel metal2 s 18400 0 18456 800 6 la_data_in[15]
port 149 nsew default input
rlabel metal2 s 18768 0 18824 800 6 la_data_in[16]
port 150 nsew default input
rlabel metal2 s 19136 0 19192 800 6 la_data_in[17]
port 151 nsew default input
rlabel metal2 s 19504 0 19560 800 6 la_data_in[18]
port 152 nsew default input
rlabel metal2 s 19872 0 19928 800 6 la_data_in[19]
port 153 nsew default input
rlabel metal2 s 13340 0 13396 800 6 la_data_in[1]
port 154 nsew default input
rlabel metal2 s 20240 0 20296 800 6 la_data_in[20]
port 155 nsew default input
rlabel metal2 s 20608 0 20664 800 6 la_data_in[21]
port 156 nsew default input
rlabel metal2 s 20976 0 21032 800 6 la_data_in[22]
port 157 nsew default input
rlabel metal2 s 21344 0 21400 800 6 la_data_in[23]
port 158 nsew default input
rlabel metal2 s 21712 0 21768 800 6 la_data_in[24]
port 159 nsew default input
rlabel metal2 s 22080 0 22136 800 6 la_data_in[25]
port 160 nsew default input
rlabel metal2 s 22448 0 22504 800 6 la_data_in[26]
port 161 nsew default input
rlabel metal2 s 22816 0 22872 800 6 la_data_in[27]
port 162 nsew default input
rlabel metal2 s 23184 0 23240 800 6 la_data_in[28]
port 163 nsew default input
rlabel metal2 s 23552 0 23608 800 6 la_data_in[29]
port 164 nsew default input
rlabel metal2 s 13708 0 13764 800 6 la_data_in[2]
port 165 nsew default input
rlabel metal2 s 23920 0 23976 800 6 la_data_in[30]
port 166 nsew default input
rlabel metal2 s 24288 0 24344 800 6 la_data_in[31]
port 167 nsew default input
rlabel metal2 s 24656 0 24712 800 6 la_data_in[32]
port 168 nsew default input
rlabel metal2 s 25024 0 25080 800 6 la_data_in[33]
port 169 nsew default input
rlabel metal2 s 25392 0 25448 800 6 la_data_in[34]
port 170 nsew default input
rlabel metal2 s 25760 0 25816 800 6 la_data_in[35]
port 171 nsew default input
rlabel metal2 s 26128 0 26184 800 6 la_data_in[36]
port 172 nsew default input
rlabel metal2 s 26496 0 26552 800 6 la_data_in[37]
port 173 nsew default input
rlabel metal2 s 26864 0 26920 800 6 la_data_in[38]
port 174 nsew default input
rlabel metal2 s 27232 0 27288 800 6 la_data_in[39]
port 175 nsew default input
rlabel metal2 s 14076 0 14132 800 6 la_data_in[3]
port 176 nsew default input
rlabel metal2 s 27600 0 27656 800 6 la_data_in[40]
port 177 nsew default input
rlabel metal2 s 27968 0 28024 800 6 la_data_in[41]
port 178 nsew default input
rlabel metal2 s 28336 0 28392 800 6 la_data_in[42]
port 179 nsew default input
rlabel metal2 s 28704 0 28760 800 6 la_data_in[43]
port 180 nsew default input
rlabel metal2 s 29072 0 29128 800 6 la_data_in[44]
port 181 nsew default input
rlabel metal2 s 29440 0 29496 800 6 la_data_in[45]
port 182 nsew default input
rlabel metal2 s 29808 0 29864 800 6 la_data_in[46]
port 183 nsew default input
rlabel metal2 s 30176 0 30232 800 6 la_data_in[47]
port 184 nsew default input
rlabel metal2 s 30544 0 30600 800 6 la_data_in[48]
port 185 nsew default input
rlabel metal2 s 30912 0 30968 800 6 la_data_in[49]
port 186 nsew default input
rlabel metal2 s 14444 0 14500 800 6 la_data_in[4]
port 187 nsew default input
rlabel metal2 s 31280 0 31336 800 6 la_data_in[50]
port 188 nsew default input
rlabel metal2 s 31648 0 31704 800 6 la_data_in[51]
port 189 nsew default input
rlabel metal2 s 32016 0 32072 800 6 la_data_in[52]
port 190 nsew default input
rlabel metal2 s 32384 0 32440 800 6 la_data_in[53]
port 191 nsew default input
rlabel metal2 s 32752 0 32808 800 6 la_data_in[54]
port 192 nsew default input
rlabel metal2 s 33120 0 33176 800 6 la_data_in[55]
port 193 nsew default input
rlabel metal2 s 33488 0 33544 800 6 la_data_in[56]
port 194 nsew default input
rlabel metal2 s 33856 0 33912 800 6 la_data_in[57]
port 195 nsew default input
rlabel metal2 s 34224 0 34280 800 6 la_data_in[58]
port 196 nsew default input
rlabel metal2 s 34592 0 34648 800 6 la_data_in[59]
port 197 nsew default input
rlabel metal2 s 14812 0 14868 800 6 la_data_in[5]
port 198 nsew default input
rlabel metal2 s 34960 0 35016 800 6 la_data_in[60]
port 199 nsew default input
rlabel metal2 s 35328 0 35384 800 6 la_data_in[61]
port 200 nsew default input
rlabel metal2 s 35696 0 35752 800 6 la_data_in[62]
port 201 nsew default input
rlabel metal2 s 36064 0 36120 800 6 la_data_in[63]
port 202 nsew default input
rlabel metal2 s 36432 0 36488 800 6 la_data_in[64]
port 203 nsew default input
rlabel metal2 s 36800 0 36856 800 6 la_data_in[65]
port 204 nsew default input
rlabel metal2 s 37168 0 37224 800 6 la_data_in[66]
port 205 nsew default input
rlabel metal2 s 37536 0 37592 800 6 la_data_in[67]
port 206 nsew default input
rlabel metal2 s 37904 0 37960 800 6 la_data_in[68]
port 207 nsew default input
rlabel metal2 s 38272 0 38328 800 6 la_data_in[69]
port 208 nsew default input
rlabel metal2 s 15088 0 15144 800 6 la_data_in[6]
port 209 nsew default input
rlabel metal2 s 38640 0 38696 800 6 la_data_in[70]
port 210 nsew default input
rlabel metal2 s 39008 0 39064 800 6 la_data_in[71]
port 211 nsew default input
rlabel metal2 s 39376 0 39432 800 6 la_data_in[72]
port 212 nsew default input
rlabel metal2 s 39744 0 39800 800 6 la_data_in[73]
port 213 nsew default input
rlabel metal2 s 40112 0 40168 800 6 la_data_in[74]
port 214 nsew default input
rlabel metal2 s 40480 0 40536 800 6 la_data_in[75]
port 215 nsew default input
rlabel metal2 s 40848 0 40904 800 6 la_data_in[76]
port 216 nsew default input
rlabel metal2 s 41216 0 41272 800 6 la_data_in[77]
port 217 nsew default input
rlabel metal2 s 41584 0 41640 800 6 la_data_in[78]
port 218 nsew default input
rlabel metal2 s 41952 0 42008 800 6 la_data_in[79]
port 219 nsew default input
rlabel metal2 s 15456 0 15512 800 6 la_data_in[7]
port 220 nsew default input
rlabel metal2 s 42320 0 42376 800 6 la_data_in[80]
port 221 nsew default input
rlabel metal2 s 42688 0 42744 800 6 la_data_in[81]
port 222 nsew default input
rlabel metal2 s 43056 0 43112 800 6 la_data_in[82]
port 223 nsew default input
rlabel metal2 s 43424 0 43480 800 6 la_data_in[83]
port 224 nsew default input
rlabel metal2 s 43792 0 43848 800 6 la_data_in[84]
port 225 nsew default input
rlabel metal2 s 44160 0 44216 800 6 la_data_in[85]
port 226 nsew default input
rlabel metal2 s 44528 0 44584 800 6 la_data_in[86]
port 227 nsew default input
rlabel metal2 s 44896 0 44952 800 6 la_data_in[87]
port 228 nsew default input
rlabel metal2 s 45264 0 45320 800 6 la_data_in[88]
port 229 nsew default input
rlabel metal2 s 45632 0 45688 800 6 la_data_in[89]
port 230 nsew default input
rlabel metal2 s 15824 0 15880 800 6 la_data_in[8]
port 231 nsew default input
rlabel metal2 s 46000 0 46056 800 6 la_data_in[90]
port 232 nsew default input
rlabel metal2 s 46368 0 46424 800 6 la_data_in[91]
port 233 nsew default input
rlabel metal2 s 46736 0 46792 800 6 la_data_in[92]
port 234 nsew default input
rlabel metal2 s 47104 0 47160 800 6 la_data_in[93]
port 235 nsew default input
rlabel metal2 s 47472 0 47528 800 6 la_data_in[94]
port 236 nsew default input
rlabel metal2 s 47840 0 47896 800 6 la_data_in[95]
port 237 nsew default input
rlabel metal2 s 48208 0 48264 800 6 la_data_in[96]
port 238 nsew default input
rlabel metal2 s 48576 0 48632 800 6 la_data_in[97]
port 239 nsew default input
rlabel metal2 s 48944 0 49000 800 6 la_data_in[98]
port 240 nsew default input
rlabel metal2 s 49312 0 49368 800 6 la_data_in[99]
port 241 nsew default input
rlabel metal2 s 16192 0 16248 800 6 la_data_in[9]
port 242 nsew default input
rlabel metal2 s 13064 0 13120 800 6 la_data_out[0]
port 243 nsew default output
rlabel metal2 s 49772 0 49828 800 6 la_data_out[100]
port 244 nsew default output
rlabel metal2 s 50140 0 50196 800 6 la_data_out[101]
port 245 nsew default output
rlabel metal2 s 50508 0 50564 800 6 la_data_out[102]
port 246 nsew default output
rlabel metal2 s 50876 0 50932 800 6 la_data_out[103]
port 247 nsew default output
rlabel metal2 s 51244 0 51300 800 6 la_data_out[104]
port 248 nsew default output
rlabel metal2 s 51612 0 51668 800 6 la_data_out[105]
port 249 nsew default output
rlabel metal2 s 51980 0 52036 800 6 la_data_out[106]
port 250 nsew default output
rlabel metal2 s 52348 0 52404 800 6 la_data_out[107]
port 251 nsew default output
rlabel metal2 s 52716 0 52772 800 6 la_data_out[108]
port 252 nsew default output
rlabel metal2 s 53084 0 53140 800 6 la_data_out[109]
port 253 nsew default output
rlabel metal2 s 16744 0 16800 800 6 la_data_out[10]
port 254 nsew default output
rlabel metal2 s 53452 0 53508 800 6 la_data_out[110]
port 255 nsew default output
rlabel metal2 s 53820 0 53876 800 6 la_data_out[111]
port 256 nsew default output
rlabel metal2 s 54188 0 54244 800 6 la_data_out[112]
port 257 nsew default output
rlabel metal2 s 54556 0 54612 800 6 la_data_out[113]
port 258 nsew default output
rlabel metal2 s 54924 0 54980 800 6 la_data_out[114]
port 259 nsew default output
rlabel metal2 s 55292 0 55348 800 6 la_data_out[115]
port 260 nsew default output
rlabel metal2 s 55660 0 55716 800 6 la_data_out[116]
port 261 nsew default output
rlabel metal2 s 56028 0 56084 800 6 la_data_out[117]
port 262 nsew default output
rlabel metal2 s 56396 0 56452 800 6 la_data_out[118]
port 263 nsew default output
rlabel metal2 s 56764 0 56820 800 6 la_data_out[119]
port 264 nsew default output
rlabel metal2 s 17112 0 17168 800 6 la_data_out[11]
port 265 nsew default output
rlabel metal2 s 57132 0 57188 800 6 la_data_out[120]
port 266 nsew default output
rlabel metal2 s 57500 0 57556 800 6 la_data_out[121]
port 267 nsew default output
rlabel metal2 s 57868 0 57924 800 6 la_data_out[122]
port 268 nsew default output
rlabel metal2 s 58236 0 58292 800 6 la_data_out[123]
port 269 nsew default output
rlabel metal2 s 58604 0 58660 800 6 la_data_out[124]
port 270 nsew default output
rlabel metal2 s 58972 0 59028 800 6 la_data_out[125]
port 271 nsew default output
rlabel metal2 s 59340 0 59396 800 6 la_data_out[126]
port 272 nsew default output
rlabel metal2 s 59708 0 59764 800 6 la_data_out[127]
port 273 nsew default output
rlabel metal2 s 17480 0 17536 800 6 la_data_out[12]
port 274 nsew default output
rlabel metal2 s 17848 0 17904 800 6 la_data_out[13]
port 275 nsew default output
rlabel metal2 s 18216 0 18272 800 6 la_data_out[14]
port 276 nsew default output
rlabel metal2 s 18584 0 18640 800 6 la_data_out[15]
port 277 nsew default output
rlabel metal2 s 18952 0 19008 800 6 la_data_out[16]
port 278 nsew default output
rlabel metal2 s 19320 0 19376 800 6 la_data_out[17]
port 279 nsew default output
rlabel metal2 s 19688 0 19744 800 6 la_data_out[18]
port 280 nsew default output
rlabel metal2 s 20056 0 20112 800 6 la_data_out[19]
port 281 nsew default output
rlabel metal2 s 13432 0 13488 800 6 la_data_out[1]
port 282 nsew default output
rlabel metal2 s 20424 0 20480 800 6 la_data_out[20]
port 283 nsew default output
rlabel metal2 s 20792 0 20848 800 6 la_data_out[21]
port 284 nsew default output
rlabel metal2 s 21160 0 21216 800 6 la_data_out[22]
port 285 nsew default output
rlabel metal2 s 21528 0 21584 800 6 la_data_out[23]
port 286 nsew default output
rlabel metal2 s 21896 0 21952 800 6 la_data_out[24]
port 287 nsew default output
rlabel metal2 s 22264 0 22320 800 6 la_data_out[25]
port 288 nsew default output
rlabel metal2 s 22632 0 22688 800 6 la_data_out[26]
port 289 nsew default output
rlabel metal2 s 23000 0 23056 800 6 la_data_out[27]
port 290 nsew default output
rlabel metal2 s 23368 0 23424 800 6 la_data_out[28]
port 291 nsew default output
rlabel metal2 s 23736 0 23792 800 6 la_data_out[29]
port 292 nsew default output
rlabel metal2 s 13800 0 13856 800 6 la_data_out[2]
port 293 nsew default output
rlabel metal2 s 24104 0 24160 800 6 la_data_out[30]
port 294 nsew default output
rlabel metal2 s 24472 0 24528 800 6 la_data_out[31]
port 295 nsew default output
rlabel metal2 s 24840 0 24896 800 6 la_data_out[32]
port 296 nsew default output
rlabel metal2 s 25208 0 25264 800 6 la_data_out[33]
port 297 nsew default output
rlabel metal2 s 25576 0 25632 800 6 la_data_out[34]
port 298 nsew default output
rlabel metal2 s 25944 0 26000 800 6 la_data_out[35]
port 299 nsew default output
rlabel metal2 s 26312 0 26368 800 6 la_data_out[36]
port 300 nsew default output
rlabel metal2 s 26680 0 26736 800 6 la_data_out[37]
port 301 nsew default output
rlabel metal2 s 27048 0 27104 800 6 la_data_out[38]
port 302 nsew default output
rlabel metal2 s 27416 0 27472 800 6 la_data_out[39]
port 303 nsew default output
rlabel metal2 s 14168 0 14224 800 6 la_data_out[3]
port 304 nsew default output
rlabel metal2 s 27784 0 27840 800 6 la_data_out[40]
port 305 nsew default output
rlabel metal2 s 28152 0 28208 800 6 la_data_out[41]
port 306 nsew default output
rlabel metal2 s 28520 0 28576 800 6 la_data_out[42]
port 307 nsew default output
rlabel metal2 s 28888 0 28944 800 6 la_data_out[43]
port 308 nsew default output
rlabel metal2 s 29256 0 29312 800 6 la_data_out[44]
port 309 nsew default output
rlabel metal2 s 29624 0 29680 800 6 la_data_out[45]
port 310 nsew default output
rlabel metal2 s 29992 0 30048 800 6 la_data_out[46]
port 311 nsew default output
rlabel metal2 s 30268 0 30324 800 6 la_data_out[47]
port 312 nsew default output
rlabel metal2 s 30636 0 30692 800 6 la_data_out[48]
port 313 nsew default output
rlabel metal2 s 31004 0 31060 800 6 la_data_out[49]
port 314 nsew default output
rlabel metal2 s 14536 0 14592 800 6 la_data_out[4]
port 315 nsew default output
rlabel metal2 s 31372 0 31428 800 6 la_data_out[50]
port 316 nsew default output
rlabel metal2 s 31740 0 31796 800 6 la_data_out[51]
port 317 nsew default output
rlabel metal2 s 32108 0 32164 800 6 la_data_out[52]
port 318 nsew default output
rlabel metal2 s 32476 0 32532 800 6 la_data_out[53]
port 319 nsew default output
rlabel metal2 s 32844 0 32900 800 6 la_data_out[54]
port 320 nsew default output
rlabel metal2 s 33212 0 33268 800 6 la_data_out[55]
port 321 nsew default output
rlabel metal2 s 33580 0 33636 800 6 la_data_out[56]
port 322 nsew default output
rlabel metal2 s 33948 0 34004 800 6 la_data_out[57]
port 323 nsew default output
rlabel metal2 s 34316 0 34372 800 6 la_data_out[58]
port 324 nsew default output
rlabel metal2 s 34684 0 34740 800 6 la_data_out[59]
port 325 nsew default output
rlabel metal2 s 14904 0 14960 800 6 la_data_out[5]
port 326 nsew default output
rlabel metal2 s 35052 0 35108 800 6 la_data_out[60]
port 327 nsew default output
rlabel metal2 s 35420 0 35476 800 6 la_data_out[61]
port 328 nsew default output
rlabel metal2 s 35788 0 35844 800 6 la_data_out[62]
port 329 nsew default output
rlabel metal2 s 36156 0 36212 800 6 la_data_out[63]
port 330 nsew default output
rlabel metal2 s 36524 0 36580 800 6 la_data_out[64]
port 331 nsew default output
rlabel metal2 s 36892 0 36948 800 6 la_data_out[65]
port 332 nsew default output
rlabel metal2 s 37260 0 37316 800 6 la_data_out[66]
port 333 nsew default output
rlabel metal2 s 37628 0 37684 800 6 la_data_out[67]
port 334 nsew default output
rlabel metal2 s 37996 0 38052 800 6 la_data_out[68]
port 335 nsew default output
rlabel metal2 s 38364 0 38420 800 6 la_data_out[69]
port 336 nsew default output
rlabel metal2 s 15272 0 15328 800 6 la_data_out[6]
port 337 nsew default output
rlabel metal2 s 38732 0 38788 800 6 la_data_out[70]
port 338 nsew default output
rlabel metal2 s 39100 0 39156 800 6 la_data_out[71]
port 339 nsew default output
rlabel metal2 s 39468 0 39524 800 6 la_data_out[72]
port 340 nsew default output
rlabel metal2 s 39836 0 39892 800 6 la_data_out[73]
port 341 nsew default output
rlabel metal2 s 40204 0 40260 800 6 la_data_out[74]
port 342 nsew default output
rlabel metal2 s 40572 0 40628 800 6 la_data_out[75]
port 343 nsew default output
rlabel metal2 s 40940 0 40996 800 6 la_data_out[76]
port 344 nsew default output
rlabel metal2 s 41308 0 41364 800 6 la_data_out[77]
port 345 nsew default output
rlabel metal2 s 41676 0 41732 800 6 la_data_out[78]
port 346 nsew default output
rlabel metal2 s 42044 0 42100 800 6 la_data_out[79]
port 347 nsew default output
rlabel metal2 s 15640 0 15696 800 6 la_data_out[7]
port 348 nsew default output
rlabel metal2 s 42412 0 42468 800 6 la_data_out[80]
port 349 nsew default output
rlabel metal2 s 42780 0 42836 800 6 la_data_out[81]
port 350 nsew default output
rlabel metal2 s 43148 0 43204 800 6 la_data_out[82]
port 351 nsew default output
rlabel metal2 s 43516 0 43572 800 6 la_data_out[83]
port 352 nsew default output
rlabel metal2 s 43884 0 43940 800 6 la_data_out[84]
port 353 nsew default output
rlabel metal2 s 44252 0 44308 800 6 la_data_out[85]
port 354 nsew default output
rlabel metal2 s 44620 0 44676 800 6 la_data_out[86]
port 355 nsew default output
rlabel metal2 s 44988 0 45044 800 6 la_data_out[87]
port 356 nsew default output
rlabel metal2 s 45356 0 45412 800 6 la_data_out[88]
port 357 nsew default output
rlabel metal2 s 45724 0 45780 800 6 la_data_out[89]
port 358 nsew default output
rlabel metal2 s 16008 0 16064 800 6 la_data_out[8]
port 359 nsew default output
rlabel metal2 s 46092 0 46148 800 6 la_data_out[90]
port 360 nsew default output
rlabel metal2 s 46460 0 46516 800 6 la_data_out[91]
port 361 nsew default output
rlabel metal2 s 46828 0 46884 800 6 la_data_out[92]
port 362 nsew default output
rlabel metal2 s 47196 0 47252 800 6 la_data_out[93]
port 363 nsew default output
rlabel metal2 s 47564 0 47620 800 6 la_data_out[94]
port 364 nsew default output
rlabel metal2 s 47932 0 47988 800 6 la_data_out[95]
port 365 nsew default output
rlabel metal2 s 48300 0 48356 800 6 la_data_out[96]
port 366 nsew default output
rlabel metal2 s 48668 0 48724 800 6 la_data_out[97]
port 367 nsew default output
rlabel metal2 s 49036 0 49092 800 6 la_data_out[98]
port 368 nsew default output
rlabel metal2 s 49404 0 49460 800 6 la_data_out[99]
port 369 nsew default output
rlabel metal2 s 16376 0 16432 800 6 la_data_out[9]
port 370 nsew default output
rlabel metal2 s 13156 0 13212 800 6 la_oen[0]
port 371 nsew default input
rlabel metal2 s 49864 0 49920 800 6 la_oen[100]
port 372 nsew default input
rlabel metal2 s 50232 0 50288 800 6 la_oen[101]
port 373 nsew default input
rlabel metal2 s 50600 0 50656 800 6 la_oen[102]
port 374 nsew default input
rlabel metal2 s 50968 0 51024 800 6 la_oen[103]
port 375 nsew default input
rlabel metal2 s 51336 0 51392 800 6 la_oen[104]
port 376 nsew default input
rlabel metal2 s 51704 0 51760 800 6 la_oen[105]
port 377 nsew default input
rlabel metal2 s 52072 0 52128 800 6 la_oen[106]
port 378 nsew default input
rlabel metal2 s 52440 0 52496 800 6 la_oen[107]
port 379 nsew default input
rlabel metal2 s 52808 0 52864 800 6 la_oen[108]
port 380 nsew default input
rlabel metal2 s 53176 0 53232 800 6 la_oen[109]
port 381 nsew default input
rlabel metal2 s 16836 0 16892 800 6 la_oen[10]
port 382 nsew default input
rlabel metal2 s 53544 0 53600 800 6 la_oen[110]
port 383 nsew default input
rlabel metal2 s 53912 0 53968 800 6 la_oen[111]
port 384 nsew default input
rlabel metal2 s 54280 0 54336 800 6 la_oen[112]
port 385 nsew default input
rlabel metal2 s 54648 0 54704 800 6 la_oen[113]
port 386 nsew default input
rlabel metal2 s 55016 0 55072 800 6 la_oen[114]
port 387 nsew default input
rlabel metal2 s 55384 0 55440 800 6 la_oen[115]
port 388 nsew default input
rlabel metal2 s 55752 0 55808 800 6 la_oen[116]
port 389 nsew default input
rlabel metal2 s 56120 0 56176 800 6 la_oen[117]
port 390 nsew default input
rlabel metal2 s 56488 0 56544 800 6 la_oen[118]
port 391 nsew default input
rlabel metal2 s 56856 0 56912 800 6 la_oen[119]
port 392 nsew default input
rlabel metal2 s 17204 0 17260 800 6 la_oen[11]
port 393 nsew default input
rlabel metal2 s 57224 0 57280 800 6 la_oen[120]
port 394 nsew default input
rlabel metal2 s 57592 0 57648 800 6 la_oen[121]
port 395 nsew default input
rlabel metal2 s 57960 0 58016 800 6 la_oen[122]
port 396 nsew default input
rlabel metal2 s 58328 0 58384 800 6 la_oen[123]
port 397 nsew default input
rlabel metal2 s 58696 0 58752 800 6 la_oen[124]
port 398 nsew default input
rlabel metal2 s 59064 0 59120 800 6 la_oen[125]
port 399 nsew default input
rlabel metal2 s 59432 0 59488 800 6 la_oen[126]
port 400 nsew default input
rlabel metal2 s 59800 0 59856 800 6 la_oen[127]
port 401 nsew default input
rlabel metal2 s 17572 0 17628 800 6 la_oen[12]
port 402 nsew default input
rlabel metal2 s 17940 0 17996 800 6 la_oen[13]
port 403 nsew default input
rlabel metal2 s 18308 0 18364 800 6 la_oen[14]
port 404 nsew default input
rlabel metal2 s 18676 0 18732 800 6 la_oen[15]
port 405 nsew default input
rlabel metal2 s 19044 0 19100 800 6 la_oen[16]
port 406 nsew default input
rlabel metal2 s 19412 0 19468 800 6 la_oen[17]
port 407 nsew default input
rlabel metal2 s 19780 0 19836 800 6 la_oen[18]
port 408 nsew default input
rlabel metal2 s 20148 0 20204 800 6 la_oen[19]
port 409 nsew default input
rlabel metal2 s 13524 0 13580 800 6 la_oen[1]
port 410 nsew default input
rlabel metal2 s 20516 0 20572 800 6 la_oen[20]
port 411 nsew default input
rlabel metal2 s 20884 0 20940 800 6 la_oen[21]
port 412 nsew default input
rlabel metal2 s 21252 0 21308 800 6 la_oen[22]
port 413 nsew default input
rlabel metal2 s 21620 0 21676 800 6 la_oen[23]
port 414 nsew default input
rlabel metal2 s 21988 0 22044 800 6 la_oen[24]
port 415 nsew default input
rlabel metal2 s 22356 0 22412 800 6 la_oen[25]
port 416 nsew default input
rlabel metal2 s 22724 0 22780 800 6 la_oen[26]
port 417 nsew default input
rlabel metal2 s 23092 0 23148 800 6 la_oen[27]
port 418 nsew default input
rlabel metal2 s 23460 0 23516 800 6 la_oen[28]
port 419 nsew default input
rlabel metal2 s 23828 0 23884 800 6 la_oen[29]
port 420 nsew default input
rlabel metal2 s 13892 0 13948 800 6 la_oen[2]
port 421 nsew default input
rlabel metal2 s 24196 0 24252 800 6 la_oen[30]
port 422 nsew default input
rlabel metal2 s 24564 0 24620 800 6 la_oen[31]
port 423 nsew default input
rlabel metal2 s 24932 0 24988 800 6 la_oen[32]
port 424 nsew default input
rlabel metal2 s 25300 0 25356 800 6 la_oen[33]
port 425 nsew default input
rlabel metal2 s 25668 0 25724 800 6 la_oen[34]
port 426 nsew default input
rlabel metal2 s 26036 0 26092 800 6 la_oen[35]
port 427 nsew default input
rlabel metal2 s 26404 0 26460 800 6 la_oen[36]
port 428 nsew default input
rlabel metal2 s 26772 0 26828 800 6 la_oen[37]
port 429 nsew default input
rlabel metal2 s 27140 0 27196 800 6 la_oen[38]
port 430 nsew default input
rlabel metal2 s 27508 0 27564 800 6 la_oen[39]
port 431 nsew default input
rlabel metal2 s 14260 0 14316 800 6 la_oen[3]
port 432 nsew default input
rlabel metal2 s 27876 0 27932 800 6 la_oen[40]
port 433 nsew default input
rlabel metal2 s 28244 0 28300 800 6 la_oen[41]
port 434 nsew default input
rlabel metal2 s 28612 0 28668 800 6 la_oen[42]
port 435 nsew default input
rlabel metal2 s 28980 0 29036 800 6 la_oen[43]
port 436 nsew default input
rlabel metal2 s 29348 0 29404 800 6 la_oen[44]
port 437 nsew default input
rlabel metal2 s 29716 0 29772 800 6 la_oen[45]
port 438 nsew default input
rlabel metal2 s 30084 0 30140 800 6 la_oen[46]
port 439 nsew default input
rlabel metal2 s 30452 0 30508 800 6 la_oen[47]
port 440 nsew default input
rlabel metal2 s 30820 0 30876 800 6 la_oen[48]
port 441 nsew default input
rlabel metal2 s 31188 0 31244 800 6 la_oen[49]
port 442 nsew default input
rlabel metal2 s 14628 0 14684 800 6 la_oen[4]
port 443 nsew default input
rlabel metal2 s 31556 0 31612 800 6 la_oen[50]
port 444 nsew default input
rlabel metal2 s 31924 0 31980 800 6 la_oen[51]
port 445 nsew default input
rlabel metal2 s 32292 0 32348 800 6 la_oen[52]
port 446 nsew default input
rlabel metal2 s 32660 0 32716 800 6 la_oen[53]
port 447 nsew default input
rlabel metal2 s 33028 0 33084 800 6 la_oen[54]
port 448 nsew default input
rlabel metal2 s 33396 0 33452 800 6 la_oen[55]
port 449 nsew default input
rlabel metal2 s 33764 0 33820 800 6 la_oen[56]
port 450 nsew default input
rlabel metal2 s 34132 0 34188 800 6 la_oen[57]
port 451 nsew default input
rlabel metal2 s 34500 0 34556 800 6 la_oen[58]
port 452 nsew default input
rlabel metal2 s 34868 0 34924 800 6 la_oen[59]
port 453 nsew default input
rlabel metal2 s 14996 0 15052 800 6 la_oen[5]
port 454 nsew default input
rlabel metal2 s 35236 0 35292 800 6 la_oen[60]
port 455 nsew default input
rlabel metal2 s 35604 0 35660 800 6 la_oen[61]
port 456 nsew default input
rlabel metal2 s 35972 0 36028 800 6 la_oen[62]
port 457 nsew default input
rlabel metal2 s 36340 0 36396 800 6 la_oen[63]
port 458 nsew default input
rlabel metal2 s 36708 0 36764 800 6 la_oen[64]
port 459 nsew default input
rlabel metal2 s 37076 0 37132 800 6 la_oen[65]
port 460 nsew default input
rlabel metal2 s 37444 0 37500 800 6 la_oen[66]
port 461 nsew default input
rlabel metal2 s 37812 0 37868 800 6 la_oen[67]
port 462 nsew default input
rlabel metal2 s 38180 0 38236 800 6 la_oen[68]
port 463 nsew default input
rlabel metal2 s 38548 0 38604 800 6 la_oen[69]
port 464 nsew default input
rlabel metal2 s 15364 0 15420 800 6 la_oen[6]
port 465 nsew default input
rlabel metal2 s 38916 0 38972 800 6 la_oen[70]
port 466 nsew default input
rlabel metal2 s 39284 0 39340 800 6 la_oen[71]
port 467 nsew default input
rlabel metal2 s 39652 0 39708 800 6 la_oen[72]
port 468 nsew default input
rlabel metal2 s 40020 0 40076 800 6 la_oen[73]
port 469 nsew default input
rlabel metal2 s 40388 0 40444 800 6 la_oen[74]
port 470 nsew default input
rlabel metal2 s 40756 0 40812 800 6 la_oen[75]
port 471 nsew default input
rlabel metal2 s 41124 0 41180 800 6 la_oen[76]
port 472 nsew default input
rlabel metal2 s 41492 0 41548 800 6 la_oen[77]
port 473 nsew default input
rlabel metal2 s 41860 0 41916 800 6 la_oen[78]
port 474 nsew default input
rlabel metal2 s 42228 0 42284 800 6 la_oen[79]
port 475 nsew default input
rlabel metal2 s 15732 0 15788 800 6 la_oen[7]
port 476 nsew default input
rlabel metal2 s 42596 0 42652 800 6 la_oen[80]
port 477 nsew default input
rlabel metal2 s 42964 0 43020 800 6 la_oen[81]
port 478 nsew default input
rlabel metal2 s 43332 0 43388 800 6 la_oen[82]
port 479 nsew default input
rlabel metal2 s 43700 0 43756 800 6 la_oen[83]
port 480 nsew default input
rlabel metal2 s 44068 0 44124 800 6 la_oen[84]
port 481 nsew default input
rlabel metal2 s 44436 0 44492 800 6 la_oen[85]
port 482 nsew default input
rlabel metal2 s 44804 0 44860 800 6 la_oen[86]
port 483 nsew default input
rlabel metal2 s 45080 0 45136 800 6 la_oen[87]
port 484 nsew default input
rlabel metal2 s 45448 0 45504 800 6 la_oen[88]
port 485 nsew default input
rlabel metal2 s 45816 0 45872 800 6 la_oen[89]
port 486 nsew default input
rlabel metal2 s 16100 0 16156 800 6 la_oen[8]
port 487 nsew default input
rlabel metal2 s 46184 0 46240 800 6 la_oen[90]
port 488 nsew default input
rlabel metal2 s 46552 0 46608 800 6 la_oen[91]
port 489 nsew default input
rlabel metal2 s 46920 0 46976 800 6 la_oen[92]
port 490 nsew default input
rlabel metal2 s 47288 0 47344 800 6 la_oen[93]
port 491 nsew default input
rlabel metal2 s 47656 0 47712 800 6 la_oen[94]
port 492 nsew default input
rlabel metal2 s 48024 0 48080 800 6 la_oen[95]
port 493 nsew default input
rlabel metal2 s 48392 0 48448 800 6 la_oen[96]
port 494 nsew default input
rlabel metal2 s 48760 0 48816 800 6 la_oen[97]
port 495 nsew default input
rlabel metal2 s 49128 0 49184 800 6 la_oen[98]
port 496 nsew default input
rlabel metal2 s 49496 0 49552 800 6 la_oen[99]
port 497 nsew default input
rlabel metal2 s 16468 0 16524 800 6 la_oen[9]
port 498 nsew default input
rlabel metal2 s 0 0 56 800 6 wb_clk_i
port 499 nsew default input
rlabel metal2 s 92 0 148 800 6 wb_rst_i
port 500 nsew default input
rlabel metal2 s 184 0 240 800 6 wbs_ack_o
port 501 nsew default output
rlabel metal2 s 644 0 700 800 6 wbs_adr_i[0]
port 502 nsew default input
rlabel metal2 s 4876 0 4932 800 6 wbs_adr_i[10]
port 503 nsew default input
rlabel metal2 s 5244 0 5300 800 6 wbs_adr_i[11]
port 504 nsew default input
rlabel metal2 s 5612 0 5668 800 6 wbs_adr_i[12]
port 505 nsew default input
rlabel metal2 s 5980 0 6036 800 6 wbs_adr_i[13]
port 506 nsew default input
rlabel metal2 s 6348 0 6404 800 6 wbs_adr_i[14]
port 507 nsew default input
rlabel metal2 s 6716 0 6772 800 6 wbs_adr_i[15]
port 508 nsew default input
rlabel metal2 s 7084 0 7140 800 6 wbs_adr_i[16]
port 509 nsew default input
rlabel metal2 s 7452 0 7508 800 6 wbs_adr_i[17]
port 510 nsew default input
rlabel metal2 s 7820 0 7876 800 6 wbs_adr_i[18]
port 511 nsew default input
rlabel metal2 s 8188 0 8244 800 6 wbs_adr_i[19]
port 512 nsew default input
rlabel metal2 s 1196 0 1252 800 6 wbs_adr_i[1]
port 513 nsew default input
rlabel metal2 s 8556 0 8612 800 6 wbs_adr_i[20]
port 514 nsew default input
rlabel metal2 s 8924 0 8980 800 6 wbs_adr_i[21]
port 515 nsew default input
rlabel metal2 s 9292 0 9348 800 6 wbs_adr_i[22]
port 516 nsew default input
rlabel metal2 s 9660 0 9716 800 6 wbs_adr_i[23]
port 517 nsew default input
rlabel metal2 s 10028 0 10084 800 6 wbs_adr_i[24]
port 518 nsew default input
rlabel metal2 s 10396 0 10452 800 6 wbs_adr_i[25]
port 519 nsew default input
rlabel metal2 s 10764 0 10820 800 6 wbs_adr_i[26]
port 520 nsew default input
rlabel metal2 s 11132 0 11188 800 6 wbs_adr_i[27]
port 521 nsew default input
rlabel metal2 s 11500 0 11556 800 6 wbs_adr_i[28]
port 522 nsew default input
rlabel metal2 s 11868 0 11924 800 6 wbs_adr_i[29]
port 523 nsew default input
rlabel metal2 s 1656 0 1712 800 6 wbs_adr_i[2]
port 524 nsew default input
rlabel metal2 s 12236 0 12292 800 6 wbs_adr_i[30]
port 525 nsew default input
rlabel metal2 s 12604 0 12660 800 6 wbs_adr_i[31]
port 526 nsew default input
rlabel metal2 s 2116 0 2172 800 6 wbs_adr_i[3]
port 527 nsew default input
rlabel metal2 s 2668 0 2724 800 6 wbs_adr_i[4]
port 528 nsew default input
rlabel metal2 s 3036 0 3092 800 6 wbs_adr_i[5]
port 529 nsew default input
rlabel metal2 s 3404 0 3460 800 6 wbs_adr_i[6]
port 530 nsew default input
rlabel metal2 s 3772 0 3828 800 6 wbs_adr_i[7]
port 531 nsew default input
rlabel metal2 s 4140 0 4196 800 6 wbs_adr_i[8]
port 532 nsew default input
rlabel metal2 s 4508 0 4564 800 6 wbs_adr_i[9]
port 533 nsew default input
rlabel metal2 s 276 0 332 800 6 wbs_cyc_i
port 534 nsew default input
rlabel metal2 s 828 0 884 800 6 wbs_dat_i[0]
port 535 nsew default input
rlabel metal2 s 4968 0 5024 800 6 wbs_dat_i[10]
port 536 nsew default input
rlabel metal2 s 5336 0 5392 800 6 wbs_dat_i[11]
port 537 nsew default input
rlabel metal2 s 5704 0 5760 800 6 wbs_dat_i[12]
port 538 nsew default input
rlabel metal2 s 6072 0 6128 800 6 wbs_dat_i[13]
port 539 nsew default input
rlabel metal2 s 6440 0 6496 800 6 wbs_dat_i[14]
port 540 nsew default input
rlabel metal2 s 6808 0 6864 800 6 wbs_dat_i[15]
port 541 nsew default input
rlabel metal2 s 7176 0 7232 800 6 wbs_dat_i[16]
port 542 nsew default input
rlabel metal2 s 7544 0 7600 800 6 wbs_dat_i[17]
port 543 nsew default input
rlabel metal2 s 7912 0 7968 800 6 wbs_dat_i[18]
port 544 nsew default input
rlabel metal2 s 8280 0 8336 800 6 wbs_dat_i[19]
port 545 nsew default input
rlabel metal2 s 1288 0 1344 800 6 wbs_dat_i[1]
port 546 nsew default input
rlabel metal2 s 8648 0 8704 800 6 wbs_dat_i[20]
port 547 nsew default input
rlabel metal2 s 9016 0 9072 800 6 wbs_dat_i[21]
port 548 nsew default input
rlabel metal2 s 9384 0 9440 800 6 wbs_dat_i[22]
port 549 nsew default input
rlabel metal2 s 9752 0 9808 800 6 wbs_dat_i[23]
port 550 nsew default input
rlabel metal2 s 10120 0 10176 800 6 wbs_dat_i[24]
port 551 nsew default input
rlabel metal2 s 10488 0 10544 800 6 wbs_dat_i[25]
port 552 nsew default input
rlabel metal2 s 10856 0 10912 800 6 wbs_dat_i[26]
port 553 nsew default input
rlabel metal2 s 11224 0 11280 800 6 wbs_dat_i[27]
port 554 nsew default input
rlabel metal2 s 11592 0 11648 800 6 wbs_dat_i[28]
port 555 nsew default input
rlabel metal2 s 11960 0 12016 800 6 wbs_dat_i[29]
port 556 nsew default input
rlabel metal2 s 1748 0 1804 800 6 wbs_dat_i[2]
port 557 nsew default input
rlabel metal2 s 12328 0 12384 800 6 wbs_dat_i[30]
port 558 nsew default input
rlabel metal2 s 12696 0 12752 800 6 wbs_dat_i[31]
port 559 nsew default input
rlabel metal2 s 2300 0 2356 800 6 wbs_dat_i[3]
port 560 nsew default input
rlabel metal2 s 2760 0 2816 800 6 wbs_dat_i[4]
port 561 nsew default input
rlabel metal2 s 3128 0 3184 800 6 wbs_dat_i[5]
port 562 nsew default input
rlabel metal2 s 3496 0 3552 800 6 wbs_dat_i[6]
port 563 nsew default input
rlabel metal2 s 3864 0 3920 800 6 wbs_dat_i[7]
port 564 nsew default input
rlabel metal2 s 4232 0 4288 800 6 wbs_dat_i[8]
port 565 nsew default input
rlabel metal2 s 4600 0 4656 800 6 wbs_dat_i[9]
port 566 nsew default input
rlabel metal2 s 920 0 976 800 6 wbs_dat_o[0]
port 567 nsew default output
rlabel metal2 s 5060 0 5116 800 6 wbs_dat_o[10]
port 568 nsew default output
rlabel metal2 s 5428 0 5484 800 6 wbs_dat_o[11]
port 569 nsew default output
rlabel metal2 s 5796 0 5852 800 6 wbs_dat_o[12]
port 570 nsew default output
rlabel metal2 s 6164 0 6220 800 6 wbs_dat_o[13]
port 571 nsew default output
rlabel metal2 s 6532 0 6588 800 6 wbs_dat_o[14]
port 572 nsew default output
rlabel metal2 s 6900 0 6956 800 6 wbs_dat_o[15]
port 573 nsew default output
rlabel metal2 s 7268 0 7324 800 6 wbs_dat_o[16]
port 574 nsew default output
rlabel metal2 s 7636 0 7692 800 6 wbs_dat_o[17]
port 575 nsew default output
rlabel metal2 s 8004 0 8060 800 6 wbs_dat_o[18]
port 576 nsew default output
rlabel metal2 s 8372 0 8428 800 6 wbs_dat_o[19]
port 577 nsew default output
rlabel metal2 s 1380 0 1436 800 6 wbs_dat_o[1]
port 578 nsew default output
rlabel metal2 s 8740 0 8796 800 6 wbs_dat_o[20]
port 579 nsew default output
rlabel metal2 s 9108 0 9164 800 6 wbs_dat_o[21]
port 580 nsew default output
rlabel metal2 s 9476 0 9532 800 6 wbs_dat_o[22]
port 581 nsew default output
rlabel metal2 s 9844 0 9900 800 6 wbs_dat_o[23]
port 582 nsew default output
rlabel metal2 s 10212 0 10268 800 6 wbs_dat_o[24]
port 583 nsew default output
rlabel metal2 s 10580 0 10636 800 6 wbs_dat_o[25]
port 584 nsew default output
rlabel metal2 s 10948 0 11004 800 6 wbs_dat_o[26]
port 585 nsew default output
rlabel metal2 s 11316 0 11372 800 6 wbs_dat_o[27]
port 586 nsew default output
rlabel metal2 s 11684 0 11740 800 6 wbs_dat_o[28]
port 587 nsew default output
rlabel metal2 s 12052 0 12108 800 6 wbs_dat_o[29]
port 588 nsew default output
rlabel metal2 s 1932 0 1988 800 6 wbs_dat_o[2]
port 589 nsew default output
rlabel metal2 s 12420 0 12476 800 6 wbs_dat_o[30]
port 590 nsew default output
rlabel metal2 s 12788 0 12844 800 6 wbs_dat_o[31]
port 591 nsew default output
rlabel metal2 s 2392 0 2448 800 6 wbs_dat_o[3]
port 592 nsew default output
rlabel metal2 s 2852 0 2908 800 6 wbs_dat_o[4]
port 593 nsew default output
rlabel metal2 s 3220 0 3276 800 6 wbs_dat_o[5]
port 594 nsew default output
rlabel metal2 s 3588 0 3644 800 6 wbs_dat_o[6]
port 595 nsew default output
rlabel metal2 s 3956 0 4012 800 6 wbs_dat_o[7]
port 596 nsew default output
rlabel metal2 s 4324 0 4380 800 6 wbs_dat_o[8]
port 597 nsew default output
rlabel metal2 s 4692 0 4748 800 6 wbs_dat_o[9]
port 598 nsew default output
rlabel metal2 s 1012 0 1068 800 6 wbs_sel_i[0]
port 599 nsew default input
rlabel metal2 s 1564 0 1620 800 6 wbs_sel_i[1]
port 600 nsew default input
rlabel metal2 s 2024 0 2080 800 6 wbs_sel_i[2]
port 601 nsew default input
rlabel metal2 s 2484 0 2540 800 6 wbs_sel_i[3]
port 602 nsew default input
rlabel metal2 s 460 0 516 800 6 wbs_stb_i
port 603 nsew default input
rlabel metal2 s 552 0 608 800 6 wbs_we_i
port 604 nsew default input
rlabel metal4 s 4190 2128 4510 57712 6 VPWR
port 605 nsew power input
rlabel metal4 s 19550 2128 19870 57712 6 VGND
port 606 nsew ground input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 59856 60000
string LEFview TRUE
<< end >>
