MACRO INVX1
 CLASS CORE ;
 ORIGIN 0.0 0.0 ;
 FOREIGN INVX1 0.0 0.0 ;
 SIZE 1.84 BY 2.72 ;
 SYMMETRY X Y R90 ;
 SITE unithd ;
  PIN vdd
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 0.00000000 2.52500000 1.84000000 2.91500000 ;
    END
  END vdd

  PIN gnd
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        RECT 0.00000000 -0.19500000 1.84000000 0.19500000 ;
    END
  END gnd

  PIN Y
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        POLYGON 1.26500000 0.60000000 1.26500000 0.83000000 1.31000000 0.83000000 1.31000000 1.90000000 1.26500000 1.90000000 1.26500000 2.13000000 1.49500000 2.13000000 1.49500000 1.90000000 1.45000000 1.90000000 1.45000000 0.83000000 1.49500000 0.83000000 1.49500000 0.60000000 ;
    END
  END Y

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER met2 ;
        POLYGON 0.80500000 0.99000000 0.80500000 1.22000000 0.85000000 1.22000000 0.85000000 1.51000000 0.80500000 1.51000000 0.80500000 1.74000000 1.03500000 1.74000000 1.03500000 1.51000000 0.99000000 1.51000000 0.99000000 1.22000000 1.03500000 1.22000000 1.03500000 0.99000000 ;
    END
  END A


END INVX1
