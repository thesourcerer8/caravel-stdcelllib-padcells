VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO OAI22X1
  CLASS CORE ;
  FOREIGN OAI22X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 4.600 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 4.600 2.960 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 4.600 0.240 ;
    END
  END gnd
  PIN Y
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.320 2.230 0.610 2.310 ;
        RECT 0.320 2.090 1.450 2.230 ;
        RECT 0.320 2.020 0.610 2.090 ;
        RECT 1.310 2.050 1.450 2.090 ;
        RECT 4.000 2.050 4.290 2.310 ;
        RECT 1.310 2.020 4.290 2.050 ;
        RECT 1.310 1.910 4.210 2.020 ;
        RECT 1.310 1.410 1.450 1.910 ;
        RECT 1.240 1.120 1.530 1.410 ;
    END
  END Y
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 3.540 1.480 3.830 1.770 ;
        RECT 3.610 1.230 3.750 1.480 ;
        RECT 3.540 0.940 3.830 1.230 ;
    END
  END B
  PIN C
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 1.700 1.120 1.990 1.770 ;
    END
  END C
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.780 1.480 1.070 1.770 ;
    END
  END D
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 2.620 1.480 2.910 1.770 ;
        RECT 2.690 1.230 2.830 1.480 ;
        RECT 2.620 0.940 2.910 1.230 ;
    END
  END A
END OAI22X1
END LIBRARY

