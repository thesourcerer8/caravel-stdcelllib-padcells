MACRO LATCH
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN LATCH 0 0 ;
 SITE CORE ;
 SYMMETRY X Y R90 ;
  PIN VDD
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.00000000 2.52500000 6.44000000 2.91500000 ;
    END
  END VDD

  PIN GND
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.00000000 -0.19500000 6.44000000 0.19500000 ;
    END
  END GND

  PIN Q
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        POLYGON 5.86500000 0.60000000 5.86500000 0.83000000 5.91000000 0.83000000 5.91000000 1.90000000 5.86500000 1.90000000 5.86500000 2.13000000 6.09500000 2.13000000 6.09500000 1.90000000 6.05000000 1.90000000 6.05000000 0.83000000 6.09500000 0.83000000 6.09500000 0.60000000 ;
       LAYER metal2 ;
        RECT 4.48500000 1.51000000 4.71500000 1.74000000 ;
       LAYER metal2 ;
        RECT 4.48500000 0.99000000 4.71500000 1.22000000 ;
    END
  END Q

  PIN D
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 1.72500000 0.99000000 1.95500000 1.35000000 ;
    END
  END D

  PIN CLK
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 3.56500000 1.51000000 3.79500000 1.74000000 ;
       LAYER metal2 ;
        RECT 0.80500000 0.99000000 1.03500000 1.22000000 ;
       LAYER metal2 ;
        RECT 3.10500000 1.51000000 3.33500000 1.74000000 ;
    END
  END CLK


END LATCH
