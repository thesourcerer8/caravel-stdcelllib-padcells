VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO XNOR2X1
  CLASS CORE ;
  FOREIGN XNOR2X1 ;
  ORIGIN 0.000 0.200 ;
  SIZE 6.440 BY 3.120 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
        RECT 0.000 2.530 6.440 2.920 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
        RECT 0.000 -0.200 6.440 0.200 ;
    END
  END gnd
  PIN Y
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
        RECT 3.110 0.860 3.340 1.090 ;
    END
  END Y
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
        RECT 0.810 1.180 1.040 1.220 ;
        RECT 1.730 1.180 1.960 1.350 ;
        RECT 0.810 1.040 1.960 1.180 ;
        RECT 0.810 0.990 1.040 1.040 ;
        RECT 1.730 0.990 1.960 1.040 ;
    END
  END B
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
        RECT 2.650 1.900 2.880 2.130 ;
    END
    PORT
      LAYER met2 ;
        RECT 3.570 0.990 3.800 1.220 ;
    END
    PORT
      LAYER met2 ;
        RECT 5.410 1.510 5.640 1.740 ;
        RECT 5.450 1.220 5.590 1.510 ;
        RECT 5.410 0.990 5.640 1.220 ;
    END
  END A
END XNOR2X1
END LIBRARY

