magic
tech sky130A
timestamp 1607784737
<< end >>
