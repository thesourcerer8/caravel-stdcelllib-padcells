VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO CLKBUF1
  CLASS CORE ;
  FOREIGN CLKBUF1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 8.280 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 8.280 2.960 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 8.280 0.240 ;
    END
  END gnd
  PIN Y
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 6.760 1.960 7.050 2.030 ;
        RECT 6.760 1.820 7.890 1.960 ;
        RECT 6.760 1.740 7.050 1.820 ;
        RECT 7.750 0.920 7.890 1.820 ;
        RECT 6.830 0.860 7.890 0.920 ;
        RECT 6.760 0.780 7.890 0.860 ;
        RECT 6.760 0.570 7.050 0.780 ;
    END
  END Y
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.780 1.570 1.070 1.640 ;
        RECT 1.700 1.570 1.990 1.640 ;
        RECT 0.780 1.430 1.990 1.570 ;
        RECT 0.780 1.090 1.070 1.430 ;
        RECT 1.700 1.090 1.990 1.430 ;
    END
  END A
END CLKBUF1
END LIBRARY

