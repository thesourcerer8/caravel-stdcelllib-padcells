VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO NAND2X1
  CLASS CORE ;
  FOREIGN NAND2X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 2.760 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 2.760 2.960 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 2.760 0.240 ;
    END
  END gnd
  PIN Y
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.320 2.230 0.610 2.310 ;
        RECT 2.160 2.230 2.450 2.310 ;
        RECT 0.320 2.090 2.450 2.230 ;
        RECT 0.320 2.020 0.610 2.090 ;
        RECT 2.160 2.020 2.450 2.090 ;
        RECT 2.230 0.690 2.370 2.020 ;
        RECT 2.160 0.400 2.450 0.690 ;
    END
  END Y
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.780 1.480 1.070 1.770 ;
        RECT 0.850 1.230 0.990 1.480 ;
        RECT 0.780 0.940 1.070 1.230 ;
    END
  END A
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 1.700 1.480 1.990 1.770 ;
        RECT 1.770 1.230 1.910 1.480 ;
        RECT 1.700 0.940 1.990 1.230 ;
    END
  END B
END NAND2X1
END LIBRARY

