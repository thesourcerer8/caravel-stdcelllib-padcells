MACRO TBUFX2
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN TBUFX2 0 0 ;
 SITE CORE ;
 SYMMETRY X Y R90 ;
  PIN VDD
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.00000000 2.52500000 5.52000000 2.91500000 ;
    END
  END VDD

  PIN GND
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.00000000 -0.19500000 5.52000000 0.19500000 ;
    END
  END GND

  PIN Y
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 3.10500000 0.60000000 3.33500000 0.83000000 ;
       LAYER metal2 ;
        RECT 3.10500000 1.90000000 3.33500000 2.13000000 ;
    END
  END Y

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        POLYGON 4.48500000 0.99000000 4.48500000 1.22000000 4.53000000 1.22000000 4.53000000 1.51000000 4.48500000 1.51000000 4.48500000 1.55500000 1.95500000 1.55500000 1.95500000 1.51000000 1.72500000 1.51000000 1.72500000 1.74000000 1.95500000 1.74000000 1.95500000 1.69500000 4.48500000 1.69500000 4.48500000 1.74000000 4.71500000 1.74000000 4.71500000 1.51000000 4.67000000 1.51000000 4.67000000 1.22000000 4.71500000 1.22000000 4.71500000 0.99000000 ;
    END
  END A

  PIN EN
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        POLYGON 0.80500000 0.99000000 0.80500000 1.22000000 0.85000000 1.22000000 0.85000000 1.51000000 0.80500000 1.51000000 0.80500000 1.74000000 1.03500000 1.74000000 1.03500000 1.51000000 0.99000000 1.51000000 0.99000000 1.22000000 1.03500000 1.22000000 1.03500000 1.17500000 2.64500000 1.17500000 2.64500000 1.22000000 2.87500000 1.22000000 2.87500000 1.17500000 3.56500000 1.17500000 3.56500000 1.22000000 3.79500000 1.22000000 3.79500000 0.99000000 3.56500000 0.99000000 3.56500000 1.03500000 2.87500000 1.03500000 2.87500000 0.99000000 2.64500000 0.99000000 2.64500000 1.03500000 1.03500000 1.03500000 1.03500000 0.99000000 ;
    END
  END EN


END TBUFX2
