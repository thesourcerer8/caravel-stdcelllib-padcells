MACRO NOR2X1
 CLASS CORE ;
 ORIGIN 0.0 0.0 ;
 FOREIGN NOR2X1 0.0 0.0 ;
 SITE CORE ;
 SYMMETRY X Y R90 ;
  PIN VDD
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.00000000 3.96500000 3.12000000 4.35500000 ;
    END
  END VDD

  PIN GND
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.00000000 -0.19500000 3.12000000 0.19500000 ;
    END
  END GND

  PIN Y
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        POLYGON 0.40500000 0.73000000 0.40500000 0.96000000 0.63500000 0.96000000 0.63500000 0.91500000 2.48500000 0.91500000 2.48500000 0.96000000 2.53000000 0.96000000 2.53000000 3.20000000 2.48500000 3.20000000 2.48500000 3.43000000 2.71500000 3.43000000 2.71500000 3.20000000 2.67000000 3.20000000 2.67000000 0.96000000 2.71500000 0.96000000 2.71500000 0.73000000 2.48500000 0.73000000 2.48500000 0.77500000 0.63500000 0.77500000 0.63500000 0.73000000 ;
    END
  END Y

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        POLYGON 1.96500000 1.12000000 1.96500000 1.35000000 2.01000000 1.35000000 2.01000000 2.81000000 1.96500000 2.81000000 1.96500000 3.04000000 2.19500000 3.04000000 2.19500000 2.81000000 2.15000000 2.81000000 2.15000000 1.35000000 2.19500000 1.35000000 2.19500000 1.12000000 ;
    END
  END B

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        POLYGON 0.92500000 1.12000000 0.92500000 1.35000000 0.97000000 1.35000000 0.97000000 2.81000000 0.92500000 2.81000000 0.92500000 3.04000000 1.15500000 3.04000000 1.15500000 2.81000000 1.11000000 2.81000000 1.11000000 1.35000000 1.15500000 1.35000000 1.15500000 1.12000000 ;
    END
  END A


END NOR2X1
