VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO HAX1
  CLASS CORE ;
  FOREIGN HAX1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.200 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 2.480 9.200 2.960 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.000 -0.240 9.200 0.240 ;
    END
  END gnd
  PIN YC
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 0.320 1.740 0.610 2.030 ;
        RECT 0.390 0.860 0.530 1.740 ;
        RECT 0.320 0.570 0.610 0.860 ;
    END
  END YC
  PIN YS
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 7.680 0.570 7.970 0.860 ;
    END
  END YS
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 2.620 1.180 2.910 1.640 ;
        RECT 5.380 1.180 5.670 1.640 ;
        RECT 2.620 1.090 5.670 1.180 ;
        RECT 2.690 1.040 5.590 1.090 ;
    END
  END B
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met1 ;
        RECT 6.300 1.090 6.590 1.640 ;
    END
    PORT
      LAYER met1 ;
        RECT 3.540 1.350 3.830 1.640 ;
    END
  END A
END HAX1
END LIBRARY

