VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO NAND3X1
  CLASS CORE ;
  FOREIGN NAND3X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.680 BY 2.720 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
        RECT 0.000 2.480 3.680 2.960 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
        RECT 0.000 -0.240 3.680 0.240 ;
    END
  END gnd
  PIN Y
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
        RECT 0.320 1.960 0.610 2.030 ;
        RECT 2.160 1.960 2.450 2.030 ;
        RECT 0.320 1.820 2.450 1.960 ;
        RECT 0.320 1.740 0.610 1.820 ;
        RECT 2.160 1.740 2.450 1.820 ;
        RECT 0.390 0.860 0.530 1.740 ;
        RECT 0.320 0.570 0.610 0.860 ;
    END
  END Y
  PIN C
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
        RECT 0.780 1.090 1.070 1.640 ;
    END
  END C
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
        RECT 1.700 1.090 1.990 1.640 ;
    END
  END B
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    SHAPE ABUTMENT ;
    PORT
      LAYER met2 ;
        RECT 2.620 1.090 2.910 1.640 ;
    END
  END A
END NAND3X1
END LIBRARY

