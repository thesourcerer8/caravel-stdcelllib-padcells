MACRO INVX8
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN INVX8 0 0 ;
 SITE CORE ;
 SYMMETRY X Y R90 ;
  PIN VDD
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.00000000 2.48000000 4.60000000 2.96000000 ;
    END
  END VDD

  PIN GND
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.00000000 -0.24000000 4.60000000 0.24000000 ;
    END
  END GND

  PIN Y
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.31500000 0.57000000 0.60500000 0.64500000 ;
        RECT 2.15500000 0.57000000 2.44500000 0.64500000 ;
        RECT 0.31500000 0.64500000 2.44500000 0.78500000 ;
        RECT 0.31500000 0.78500000 0.60500000 0.86000000 ;
        RECT 2.15500000 0.78500000 2.44500000 0.86000000 ;
        RECT 3.99500000 0.57000000 4.28500000 0.86000000 ;
        RECT 0.39000000 0.86000000 0.53000000 1.74000000 ;
        RECT 4.07000000 0.86000000 4.21000000 1.74000000 ;
        RECT 0.31500000 1.74000000 0.60500000 1.81500000 ;
        RECT 2.15500000 1.74000000 2.44500000 1.81500000 ;
        RECT 3.99500000 1.74000000 4.28500000 1.81500000 ;
        RECT 0.31500000 1.81500000 4.28500000 1.95500000 ;
        RECT 0.31500000 1.95500000 0.60500000 2.03000000 ;
        RECT 2.15500000 1.95500000 2.44500000 2.03000000 ;
        RECT 3.99500000 1.95500000 4.28500000 2.03000000 ;
    END
  END Y

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.77500000 1.09000000 1.06500000 1.16500000 ;
        RECT 1.69500000 1.09000000 1.98500000 1.16500000 ;
        RECT 2.61500000 1.09000000 2.90500000 1.16500000 ;
        RECT 3.53500000 1.09000000 3.82500000 1.16500000 ;
        RECT 0.77500000 1.16500000 3.82500000 1.30500000 ;
        RECT 0.77500000 1.30500000 1.06500000 1.64000000 ;
        RECT 1.69500000 1.30500000 1.98500000 1.64000000 ;
        RECT 2.61500000 1.30500000 2.90500000 1.64000000 ;
        RECT 3.53500000 1.30500000 3.82500000 1.64000000 ;
    END
  END A


END INVX8
