MACRO MUX2X1
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN MUX2X1 0 0 ;
 SITE CORE ;
 SYMMETRY X Y R90 ;
  PIN VDD
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.00000000 2.52500000 5.52000000 2.91500000 ;
    END
  END VDD

  PIN GND
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.00000000 -0.19500000 5.52000000 0.19500000 ;
    END
  END GND

  PIN Y
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        POLYGON 3.10500000 0.60000000 3.10500000 0.83000000 3.33500000 0.83000000 3.33500000 0.78500000 4.07000000 0.78500000 4.07000000 1.94500000 3.33500000 1.94500000 3.33500000 1.90000000 3.10500000 1.90000000 3.10500000 2.13000000 3.33500000 2.13000000 3.33500000 2.08500000 4.21000000 2.08500000 4.21000000 0.64500000 3.33500000 0.64500000 3.33500000 0.60000000 ;
    END
  END Y

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 1.72500000 0.99000000 1.95500000 1.35000000 ;
    END
  END A

  PIN S
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.80500000 0.99000000 1.03500000 1.35000000 ;
       LAYER metal2 ;
        RECT 3.56500000 1.51000000 3.79500000 1.74000000 ;
       LAYER metal2 ;
        RECT 3.10500000 1.51000000 3.33500000 1.74000000 ;
    END
  END S

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        POLYGON 4.48500000 0.99000000 4.48500000 1.22000000 4.53000000 1.22000000 4.53000000 1.51000000 4.48500000 1.51000000 4.48500000 1.74000000 4.71500000 1.74000000 4.71500000 1.51000000 4.67000000 1.51000000 4.67000000 1.22000000 4.71500000 1.22000000 4.71500000 0.99000000 ;
    END
  END B


END MUX2X1
