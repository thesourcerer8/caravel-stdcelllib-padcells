* NGSPICE file created from user_proj_example.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for NAND2X1 abstract view
.subckt NAND2X1 vdd gnd Y A B
.ends

* Black-box entry subcircuit for XNOR2X1 abstract view
.subckt XNOR2X1 vdd gnd Y A B
.ends

* Black-box entry subcircuit for AOI21X1 abstract view
.subckt AOI21X1 vdd gnd Y C B A
.ends

* Black-box entry subcircuit for XOR2X1 abstract view
.subckt XOR2X1 vdd gnd Y A B
.ends

* Black-box entry subcircuit for LATCH abstract view
.subckt LATCH vdd gnd Q CLK D
.ends

* Black-box entry subcircuit for INVX1 abstract view
.subckt INVX1 vdd gnd Y A
.ends

* Black-box entry subcircuit for INVX2 abstract view
.subckt INVX2 vdd gnd Y A
.ends

* Black-box entry subcircuit for NOR2X1 abstract view
.subckt NOR2X1 vdd gnd Y B A
.ends

* Black-box entry subcircuit for INVX4 abstract view
.subckt INVX4 vdd gnd Y A
.ends

* Black-box entry subcircuit for OR2X1 abstract view
.subckt OR2X1 vdd gnd Y B A
.ends

* Black-box entry subcircuit for OR2X2 abstract view
.subckt OR2X2 vdd gnd Y B A
.ends

* Black-box entry subcircuit for INVX8 abstract view
.subckt INVX8 vdd gnd Y A
.ends

* Black-box entry subcircuit for OAI22X1 abstract view
.subckt OAI22X1 vdd gnd Y B C D A
.ends

* Black-box entry subcircuit for BUFX2 abstract view
.subckt BUFX2 vdd gnd Y A
.ends

* Black-box entry subcircuit for NAND3X1 abstract view
.subckt NAND3X1 vdd gnd Y B A C
.ends

* Black-box entry subcircuit for INV abstract view
.subckt INV vdd gnd Y A
.ends

* Black-box entry subcircuit for TBUFX1 abstract view
.subckt TBUFX1 vdd gnd Y A EN
.ends

* Black-box entry subcircuit for BUFX4 abstract view
.subckt BUFX4 vdd gnd Y A
.ends

* Black-box entry subcircuit for TBUFX2 abstract view
.subckt TBUFX2 vdd gnd Y A EN
.ends

* Black-box entry subcircuit for AOI22X1 abstract view
.subckt AOI22X1 vdd gnd Y B A D C
.ends

* Black-box entry subcircuit for NOR3X1 abstract view
.subckt NOR3X1 vdd gnd Y B C A
.ends

* Black-box entry subcircuit for CLKBUF1 abstract view
.subckt CLKBUF1 vdd gnd Y A
.ends

* Black-box entry subcircuit for MUX2X1 abstract view
.subckt MUX2X1 vdd gnd Y A S B
.ends

* Black-box entry subcircuit for AND2X1 abstract view
.subckt AND2X1 vdd gnd Y B A
.ends

* Black-box entry subcircuit for AND2X2 abstract view
.subckt AND2X2 vdd gnd Y B A
.ends

* Black-box entry subcircuit for OAI21X1 abstract view
.subckt OAI21X1 vdd gnd Y C B A
.ends

* Black-box entry subcircuit for HAX1 abstract view
.subckt HAX1 vdd gnd YC YS A B
.ends

.subckt user_proj_example io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ la_data_in[0] la_data_in[100] la_data_in[101] la_data_in[102] la_data_in[103] la_data_in[104]
+ la_data_in[105] la_data_in[106] la_data_in[107] la_data_in[108] la_data_in[109]
+ la_data_in[10] la_data_in[110] la_data_in[111] la_data_in[112] la_data_in[113] la_data_in[114]
+ la_data_in[115] la_data_in[116] la_data_in[117] la_data_in[118] la_data_in[119]
+ la_data_in[11] la_data_in[120] la_data_in[121] la_data_in[122] la_data_in[123] la_data_in[124]
+ la_data_in[125] la_data_in[126] la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14]
+ la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1]
+ la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25]
+ la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30]
+ la_data_in[31] la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36]
+ la_data_in[37] la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41]
+ la_data_in[42] la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47]
+ la_data_in[48] la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52]
+ la_data_in[53] la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58]
+ la_data_in[59] la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63]
+ la_data_in[64] la_data_in[65] la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69]
+ la_data_in[6] la_data_in[70] la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74]
+ la_data_in[75] la_data_in[76] la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7]
+ la_data_in[80] la_data_in[81] la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85]
+ la_data_in[86] la_data_in[87] la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90]
+ la_data_in[91] la_data_in[92] la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96]
+ la_data_in[97] la_data_in[98] la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100]
+ la_data_out[101] la_data_out[102] la_data_out[103] la_data_out[104] la_data_out[105]
+ la_data_out[106] la_data_out[107] la_data_out[108] la_data_out[109] la_data_out[10]
+ la_data_out[110] la_data_out[111] la_data_out[112] la_data_out[113] la_data_out[114]
+ la_data_out[115] la_data_out[116] la_data_out[117] la_data_out[118] la_data_out[119]
+ la_data_out[11] la_data_out[120] la_data_out[121] la_data_out[122] la_data_out[123]
+ la_data_out[124] la_data_out[125] la_data_out[126] la_data_out[127] la_data_out[12]
+ la_data_out[13] la_data_out[14] la_data_out[15] la_data_out[16] la_data_out[17]
+ la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22]
+ la_data_out[23] la_data_out[24] la_data_out[25] la_data_out[26] la_data_out[27]
+ la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32]
+ la_data_out[33] la_data_out[34] la_data_out[35] la_data_out[36] la_data_out[37]
+ la_data_out[38] la_data_out[39] la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42]
+ la_data_out[43] la_data_out[44] la_data_out[45] la_data_out[46] la_data_out[47]
+ la_data_out[48] la_data_out[49] la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52]
+ la_data_out[53] la_data_out[54] la_data_out[55] la_data_out[56] la_data_out[57]
+ la_data_out[58] la_data_out[59] la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62]
+ la_data_out[63] la_data_out[64] la_data_out[65] la_data_out[66] la_data_out[67]
+ la_data_out[68] la_data_out[69] la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72]
+ la_data_out[73] la_data_out[74] la_data_out[75] la_data_out[76] la_data_out[77]
+ la_data_out[78] la_data_out[79] la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82]
+ la_data_out[83] la_data_out[84] la_data_out[85] la_data_out[86] la_data_out[87]
+ la_data_out[88] la_data_out[89] la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92]
+ la_data_out[93] la_data_out[94] la_data_out[95] la_data_out[96] la_data_out[97]
+ la_data_out[98] la_data_out[99] la_data_out[9] la_oen[0] la_oen[100] la_oen[101]
+ la_oen[102] la_oen[103] la_oen[104] la_oen[105] la_oen[106] la_oen[107] la_oen[108]
+ la_oen[109] la_oen[10] la_oen[110] la_oen[111] la_oen[112] la_oen[113] la_oen[114]
+ la_oen[115] la_oen[116] la_oen[117] la_oen[118] la_oen[119] la_oen[11] la_oen[120]
+ la_oen[121] la_oen[122] la_oen[123] la_oen[124] la_oen[125] la_oen[126] la_oen[127]
+ la_oen[12] la_oen[13] la_oen[14] la_oen[15] la_oen[16] la_oen[17] la_oen[18] la_oen[19]
+ la_oen[1] la_oen[20] la_oen[21] la_oen[22] la_oen[23] la_oen[24] la_oen[25] la_oen[26]
+ la_oen[27] la_oen[28] la_oen[29] la_oen[2] la_oen[30] la_oen[31] la_oen[32] la_oen[33]
+ la_oen[34] la_oen[35] la_oen[36] la_oen[37] la_oen[38] la_oen[39] la_oen[3] la_oen[40]
+ la_oen[41] la_oen[42] la_oen[43] la_oen[44] la_oen[45] la_oen[46] la_oen[47] la_oen[48]
+ la_oen[49] la_oen[4] la_oen[50] la_oen[51] la_oen[52] la_oen[53] la_oen[54] la_oen[55]
+ la_oen[56] la_oen[57] la_oen[58] la_oen[59] la_oen[5] la_oen[60] la_oen[61] la_oen[62]
+ la_oen[63] la_oen[64] la_oen[65] la_oen[66] la_oen[67] la_oen[68] la_oen[69] la_oen[6]
+ la_oen[70] la_oen[71] la_oen[72] la_oen[73] la_oen[74] la_oen[75] la_oen[76] la_oen[77]
+ la_oen[78] la_oen[79] la_oen[7] la_oen[80] la_oen[81] la_oen[82] la_oen[83] la_oen[84]
+ la_oen[85] la_oen[86] la_oen[87] la_oen[88] la_oen[89] la_oen[8] la_oen[90] la_oen[91]
+ la_oen[92] la_oen[93] la_oen[94] la_oen[95] la_oen[96] la_oen[97] la_oen[98] la_oen[99]
+ la_oen[9] wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12]
+ wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18]
+ wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23]
+ wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29]
+ wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5]
+ wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10]
+ wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15] wbs_dat_i[16]
+ wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20] wbs_dat_i[21]
+ wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26] wbs_dat_i[27]
+ wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31] wbs_dat_i[3]
+ wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9] wbs_dat_o[0]
+ wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14] wbs_dat_o[15]
+ wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1] wbs_dat_o[20]
+ wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25] wbs_dat_o[26]
+ wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30] wbs_dat_o[31]
+ wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9]
+ wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i VPWR VGND
XFILLER_79_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_12_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_37_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_200_ VGND VGND VPWR VPWR _200_/HI wbs_dat_o[26] sky130_fd_sc_hd__conb_1
XPHY_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_131_ VGND VGND VPWR VPWR _131_/HI la_data_out[86] sky130_fd_sc_hd__conb_1
XPHY_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_062_ VGND VGND VPWR VPWR _062_/HI la_data_out[5] sky130_fd_sc_hd__conb_1
XFILLER_3_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_2_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_69_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_114_ VGND VGND VPWR VPWR _114_/HI la_data_out[69] sky130_fd_sc_hd__conb_1
X_045_ VGND VGND VPWR VPWR _045_/HI io_out[13] sky130_fd_sc_hd__conb_1
XFILLER_98_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_40_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_028_ VGND VGND VPWR VPWR _028_/HI io_oeb[24] sky130_fd_sc_hd__conb_1
XFILLER_98_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_15_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_32_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_55_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_46_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_14_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XNAND2X1 VPWR VGND la_data_out[6] la_data_in[5] la_data_in[4] NAND2X1
XFILLER_73_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_1_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_130_ VGND VGND VPWR VPWR _130_/HI la_data_out[85] sky130_fd_sc_hd__conb_1
XFILLER_7_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_061_ VGND VGND VPWR VPWR _061_/HI la_data_out[4] sky130_fd_sc_hd__conb_1
XFILLER_23_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_113_ VGND VGND VPWR VPWR _113_/HI la_data_out[68] sky130_fd_sc_hd__conb_1
XFILLER_7_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_044_ VGND VGND VPWR VPWR _044_/HI io_out[12] sky130_fd_sc_hd__conb_1
XFILLER_3_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_78_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_61_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_71_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_027_ VGND VGND VPWR VPWR _027_/HI io_oeb[23] sky130_fd_sc_hd__conb_1
XFILLER_3_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_4_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_50_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_99_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_060_ VGND VGND VPWR VPWR _060_/HI la_data_out[2] sky130_fd_sc_hd__conb_1
XFILLER_99_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_189_ VGND VGND VPWR VPWR _189_/HI wbs_dat_o[15] sky130_fd_sc_hd__conb_1
XFILLER_6_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_33_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_55_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_112_ VGND VGND VPWR VPWR _112_/HI la_data_out[67] sky130_fd_sc_hd__conb_1
X_043_ VGND VGND VPWR VPWR _043_/HI io_out[11] sky130_fd_sc_hd__conb_1
XFILLER_3_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_59_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_21_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_026_ VGND VGND VPWR VPWR _026_/HI io_oeb[20] sky130_fd_sc_hd__conb_1
XFILLER_3_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_44_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_16_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_009_ VGND VGND VPWR VPWR io_oeb[29] _009_/LO sky130_fd_sc_hd__conb_1
XFILLER_4_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_99_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_70_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_94_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_46_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_34_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_188_ VGND VGND VPWR VPWR _188_/HI wbs_dat_o[14] sky130_fd_sc_hd__conb_1
XFILLER_69_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_92_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_111_ VGND VGND VPWR VPWR _111_/HI la_data_out[66] sky130_fd_sc_hd__conb_1
XPHY_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_042_ VGND VGND VPWR VPWR _042_/HI io_out[10] sky130_fd_sc_hd__conb_1
XFILLER_59_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_025_ VGND VGND VPWR VPWR _025_/HI io_oeb[18] sky130_fd_sc_hd__conb_1
XFILLER_3_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_008_ VGND VGND VPWR VPWR io_oeb[27] _008_/LO sky130_fd_sc_hd__conb_1
XFILLER_67_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_29_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XXNOR2X1 VPWR VGND la_data_out[41] la_data_in[40] la_data_in[39] XNOR2X1
XFILLER_83_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_99_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_187_ VGND VGND VPWR VPWR _187_/HI wbs_dat_o[13] sky130_fd_sc_hd__conb_1
XFILLER_96_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_49_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_110_ VGND VGND VPWR VPWR _110_/HI la_data_out[65] sky130_fd_sc_hd__conb_1
XPHY_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_041_ VGND VGND VPWR VPWR _041_/HI io_out[8] sky130_fd_sc_hd__conb_1
XFILLER_3_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_29_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_024_ VGND VGND VPWR VPWR _024_/HI io_oeb[16] sky130_fd_sc_hd__conb_1
XFILLER_3_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_33_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_5_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_24_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_007_ VGND VGND VPWR VPWR io_oeb[25] _007_/LO sky130_fd_sc_hd__conb_1
XFILLER_98_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_3_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XAOI21X1 VPWR VGND io_out[9] io_in[6] io_in[7] io_in[8] AOI21X1
XFILLER_12_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_68_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_186_ VGND VGND VPWR VPWR _186_/HI wbs_dat_o[12] sky130_fd_sc_hd__conb_1
XFILLER_10_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_49_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_040_ VGND VGND VPWR VPWR _040_/HI io_out[7] sky130_fd_sc_hd__conb_1
XFILLER_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_169_ VGND VGND VPWR VPWR _169_/HI la_data_out[124] sky130_fd_sc_hd__conb_1
XFILLER_6_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_97_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_023_ VGND VGND VPWR VPWR _023_/HI io_oeb[14] sky130_fd_sc_hd__conb_1
XFILLER_3_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XXOR2X1 VPWR VGND la_data_out[44] la_data_in[43] la_data_in[42] XOR2X1
XFILLER_66_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_25_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_006_ VGND VGND VPWR VPWR io_oeb[22] _006_/LO sky130_fd_sc_hd__conb_1
XFILLER_98_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_16_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_23_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XLATCH VPWR VGND io_out[37] io_in[36] io_in[35] LATCH
XFILLER_80_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_185_ VGND VGND VPWR VPWR _185_/HI wbs_dat_o[11] sky130_fd_sc_hd__conb_1
XFILLER_89_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_43_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_30_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_168_ VGND VGND VPWR VPWR _168_/HI la_data_out[123] sky130_fd_sc_hd__conb_1
XFILLER_6_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_099_ VGND VGND VPWR VPWR _099_/HI la_data_out[54] sky130_fd_sc_hd__conb_1
XFILLER_97_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_1_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_88_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_022_ VGND VGND VPWR VPWR io_oeb[11] _022_/LO sky130_fd_sc_hd__conb_1
XFILLER_79_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_005_ VGND VGND VPWR VPWR io_oeb[21] _005_/LO sky130_fd_sc_hd__conb_1
XFILLER_98_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_13_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_67_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_40_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XINVX1 VPWR VGND io_out[28] io_in[27] INVX1
XFILLER_100_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_80_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_184_ VGND VGND VPWR VPWR _184_/HI wbs_dat_o[10] sky130_fd_sc_hd__conb_1
XFILLER_6_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_77_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_55_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_54_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_91_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_167_ VGND VGND VPWR VPWR _167_/HI la_data_out[122] sky130_fd_sc_hd__conb_1
XFILLER_40_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_098_ VGND VGND VPWR VPWR _098_/HI la_data_out[53] sky130_fd_sc_hd__conb_1
XFILLER_97_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_37_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_021_ VGND VGND VPWR VPWR io_oeb[10] _021_/LO sky130_fd_sc_hd__conb_1
XFILLER_79_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_59_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_004_ VGND VGND VPWR VPWR io_oeb[19] _004_/LO sky130_fd_sc_hd__conb_1
XFILLER_4_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_23_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_15_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_97_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_38_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_90_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_37_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_94_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XINVX2 VPWR VGND io_out[30] io_in[29] INVX2
XFILLER_58_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_183_ VGND VGND VPWR VPWR _183_/HI wbs_dat_o[9] sky130_fd_sc_hd__conb_1
XFILLER_10_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_13_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_166_ VGND VGND VPWR VPWR _166_/HI la_data_out[121] sky130_fd_sc_hd__conb_1
XFILLER_6_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_097_ VGND VGND VPWR VPWR _097_/HI la_data_out[52] sky130_fd_sc_hd__conb_1
XFILLER_97_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_37_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_020_ VGND VGND VPWR VPWR io_oeb[8] _020_/LO sky130_fd_sc_hd__conb_1
XFILLER_79_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_149_ VGND VGND VPWR VPWR _149_/HI la_data_out[104] sky130_fd_sc_hd__conb_1
XFILLER_7_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XNOR2X1 VPWR VGND la_data_out[13] la_data_in[11] la_data_in[12] NOR2X1
XFILLER_21_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_16_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_003_ VGND VGND VPWR VPWR io_oeb[17] _003_/LO sky130_fd_sc_hd__conb_1
XFILLER_4_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_46_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_7_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_38_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_57_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_39_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_10_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_22_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_182_ VGND VGND VPWR VPWR _182_/HI wbs_dat_o[8] sky130_fd_sc_hd__conb_1
XFILLER_80_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_70_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_165_ VGND VGND VPWR VPWR _165_/HI la_data_out[120] sky130_fd_sc_hd__conb_1
X_096_ VGND VGND VPWR VPWR _096_/HI la_data_out[51] sky130_fd_sc_hd__conb_1
XFILLER_6_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_92_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_148_ VGND VGND VPWR VPWR _148_/HI la_data_out[103] sky130_fd_sc_hd__conb_1
XFILLER_7_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_079_ VGND VGND VPWR VPWR _079_/HI la_data_out[28] sky130_fd_sc_hd__conb_1
XFILLER_97_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_21_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_52_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_002_ VGND VGND VPWR VPWR io_oeb[15] _002_/LO sky130_fd_sc_hd__conb_1
XFILLER_21_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_94_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_17_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XINVX4 VPWR VGND io_out[32] io_in[31] INVX4
XFILLER_86_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_181_ VGND VGND VPWR VPWR _181_/HI wbs_dat_o[7] sky130_fd_sc_hd__conb_1
XFILLER_13_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_64_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_70_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_27_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_164_ VGND VGND VPWR VPWR _164_/HI la_data_out[119] sky130_fd_sc_hd__conb_1
X_095_ VGND VGND VPWR VPWR _095_/HI la_data_out[50] sky130_fd_sc_hd__conb_1
XFILLER_69_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_101_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_147_ VGND VGND VPWR VPWR _147_/HI la_data_out[102] sky130_fd_sc_hd__conb_1
XFILLER_7_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_078_ VGND VGND VPWR VPWR _078_/HI la_data_out[27] sky130_fd_sc_hd__conb_1
XFILLER_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_93_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_001_ VGND VGND VPWR VPWR io_oeb[13] _001_/LO sky130_fd_sc_hd__conb_1
XFILLER_21_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_15_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_30_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_12_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XOR2X1 VPWR VGND la_data_out[29] la_data_in[27] la_data_in[28] OR2X1
XFILLER_13_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_36_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_180_ VGND VGND VPWR VPWR _180_/HI wbs_dat_o[6] sky130_fd_sc_hd__conb_1
XFILLER_50_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_49_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_18_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_54_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_163_ VGND VGND VPWR VPWR _163_/HI la_data_out[118] sky130_fd_sc_hd__conb_1
XFILLER_6_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_094_ VGND VGND VPWR VPWR _094_/HI la_data_out[49] sky130_fd_sc_hd__conb_1
XFILLER_77_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_61_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_146_ VGND VGND VPWR VPWR _146_/HI la_data_out[101] sky130_fd_sc_hd__conb_1
X_077_ VGND VGND VPWR VPWR _077_/HI la_data_out[25] sky130_fd_sc_hd__conb_1
XFILLER_38_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_61_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_000_ VGND VGND VPWR VPWR io_oeb[12] _000_/LO sky130_fd_sc_hd__conb_1
XFILLER_101_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_47_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_129_ VGND VGND VPWR VPWR _129_/HI la_data_out[84] sky130_fd_sc_hd__conb_1
XFILLER_97_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_78_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_7_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_72_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XOR2X2 VPWR VGND la_data_out[32] la_data_in[30] la_data_in[31] OR2X2
XFILLER_9_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_36_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_162_ VGND VGND VPWR VPWR _162_/HI la_data_out[117] sky130_fd_sc_hd__conb_1
XFILLER_10_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_093_ VGND VGND VPWR VPWR _093_/HI la_data_out[48] sky130_fd_sc_hd__conb_1
XFILLER_40_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_101_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_42_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_145_ VGND VGND VPWR VPWR _145_/HI la_data_out[100] sky130_fd_sc_hd__conb_1
X_076_ VGND VGND VPWR VPWR _076_/HI la_data_out[24] sky130_fd_sc_hd__conb_1
XFILLER_78_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_128_ VGND VGND VPWR VPWR _128_/HI la_data_out[83] sky130_fd_sc_hd__conb_1
X_059_ VGND VGND VPWR VPWR _059_/HI la_data_out[1] sky130_fd_sc_hd__conb_1
XFILLER_97_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_81_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_26_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_2_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_41_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_86_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_161_ VGND VGND VPWR VPWR _161_/HI la_data_out[116] sky130_fd_sc_hd__conb_1
XFILLER_6_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_10_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_092_ VGND VGND VPWR VPWR _092_/HI la_data_out[47] sky130_fd_sc_hd__conb_1
XFILLER_2_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_60_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_20_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_144_ VGND VGND VPWR VPWR _144_/HI la_data_out[99] sky130_fd_sc_hd__conb_1
X_075_ VGND VGND VPWR VPWR _075_/HI la_data_out[23] sky130_fd_sc_hd__conb_1
XFILLER_97_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_64_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_127_ VGND VGND VPWR VPWR _127_/HI la_data_out[82] sky130_fd_sc_hd__conb_1
X_058_ VGND VGND VPWR VPWR _058_/HI la_data_out[0] sky130_fd_sc_hd__conb_1
XFILLER_97_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_5_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XINVX8 VPWR VGND io_out[34] io_in[33] INVX8
XFILLER_58_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_10_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_160_ VGND VGND VPWR VPWR _160_/HI la_data_out[115] sky130_fd_sc_hd__conb_1
X_091_ VGND VGND VPWR VPWR _091_/HI la_data_out[46] sky130_fd_sc_hd__conb_1
XFILLER_40_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_65_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_24_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_20_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_74_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_143_ VGND VGND VPWR VPWR _143_/HI la_data_out[98] sky130_fd_sc_hd__conb_1
X_074_ VGND VGND VPWR VPWR _074_/HI la_data_out[22] sky130_fd_sc_hd__conb_1
XFILLER_97_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_96_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_24_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_20_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_28_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_126_ VGND VGND VPWR VPWR _126_/HI la_data_out[81] sky130_fd_sc_hd__conb_1
XFILLER_98_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_057_ VGND VGND VPWR VPWR _057_/HI io_out[36] sky130_fd_sc_hd__conb_1
XFILLER_3_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XOAI22X1 VPWR VGND la_data_out[26] la_data_in[24] la_data_in[23] la_data_in[22] la_data_in[25]
+ OAI22X1
XPHY_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_109_ VGND VGND VPWR VPWR _109_/HI la_data_out[64] sky130_fd_sc_hd__conb_1
XFILLER_98_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_93_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_76_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_51_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_090_ VGND VGND VPWR VPWR _090_/HI la_data_out[45] sky130_fd_sc_hd__conb_1
XFILLER_40_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_142_ VGND VGND VPWR VPWR _142_/HI la_data_out[97] sky130_fd_sc_hd__conb_1
XFILLER_50_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_073_ VGND VGND VPWR VPWR _073_/HI la_data_out[20] sky130_fd_sc_hd__conb_1
XFILLER_78_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_125_ VGND VGND VPWR VPWR _125_/HI la_data_out[80] sky130_fd_sc_hd__conb_1
XFILLER_7_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_056_ VGND VGND VPWR VPWR _056_/HI io_out[35] sky130_fd_sc_hd__conb_1
XFILLER_98_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_78_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_21_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_21_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_31_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_108_ VGND VGND VPWR VPWR _108_/HI la_data_out[63] sky130_fd_sc_hd__conb_1
X_039_ VGND VGND VPWR VPWR _039_/HI io_out[6] sky130_fd_sc_hd__conb_1
XFILLER_98_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_13_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_4_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_66_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_79_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_32_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_36_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBUFX2 VPWR VGND io_out[16] io_in[15] BUFX2
XFILLER_87_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_141_ VGND VGND VPWR VPWR _141_/HI la_data_out[96] sky130_fd_sc_hd__conb_1
X_072_ VGND VGND VPWR VPWR _072_/HI la_data_out[19] sky130_fd_sc_hd__conb_1
XFILLER_2_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_93_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_18_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_2_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_124_ VGND VGND VPWR VPWR _124_/HI la_data_out[79] sky130_fd_sc_hd__conb_1
X_055_ VGND VGND VPWR VPWR _055_/HI io_out[33] sky130_fd_sc_hd__conb_1
XFILLER_3_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_87_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_12_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_107_ VGND VGND VPWR VPWR _107_/HI la_data_out[62] sky130_fd_sc_hd__conb_1
X_038_ VGND VGND VPWR VPWR _038_/HI io_out[4] sky130_fd_sc_hd__conb_1
XFILLER_98_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_90_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_100_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_89_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_54_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_72_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_81_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_50_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XNAND3X1 VPWR VGND la_data_out[10] la_data_in[8] la_data_in[9] la_data_in[7] NAND3X1
XFILLER_81_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_32_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_101_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_140_ VGND VGND VPWR VPWR _140_/HI la_data_out[95] sky130_fd_sc_hd__conb_1
X_071_ VGND VGND VPWR VPWR _071_/HI la_data_out[18] sky130_fd_sc_hd__conb_1
XFILLER_2_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XINV VPWR VGND io_out[26] io_in[25] INV
XFILLER_21_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_87_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_123_ VGND VGND VPWR VPWR _123_/HI la_data_out[78] sky130_fd_sc_hd__conb_1
XFILLER_7_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_054_ VGND VGND VPWR VPWR _054_/HI io_out[31] sky130_fd_sc_hd__conb_1
XFILLER_3_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_106_ VGND VGND VPWR VPWR _106_/HI la_data_out[61] sky130_fd_sc_hd__conb_1
XPHY_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_037_ VGND VGND VPWR VPWR _037_/HI io_out[3] sky130_fd_sc_hd__conb_1
XFILLER_93_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_75_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_79_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_24_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_81_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTBUFX1 VPWR VGND la_data_out[35] la_data_in[34] la_data_in[33] TBUFX1
XFILLER_5_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_68_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_64_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XBUFX4 VPWR VGND io_out[18] io_in[17] BUFX4
XFILLER_99_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_070_ VGND VGND VPWR VPWR _070_/HI la_data_out[16] sky130_fd_sc_hd__conb_1
XFILLER_4_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_34_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_73_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_61_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_199_ VGND VGND VPWR VPWR _199_/HI wbs_dat_o[25] sky130_fd_sc_hd__conb_1
XFILLER_96_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_43_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_122_ VGND VGND VPWR VPWR _122_/HI la_data_out[77] sky130_fd_sc_hd__conb_1
X_053_ VGND VGND VPWR VPWR _053_/HI io_out[29] sky130_fd_sc_hd__conb_1
XFILLER_78_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_19_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_57_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_52_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_80_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_105_ VGND VGND VPWR VPWR _105_/HI la_data_out[60] sky130_fd_sc_hd__conb_1
XFILLER_11_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_036_ VGND VGND VPWR VPWR _036_/HI io_out[1] sky130_fd_sc_hd__conb_1
XFILLER_78_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_53_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_019_ VGND VGND VPWR VPWR io_oeb[7] _019_/LO sky130_fd_sc_hd__conb_1
XFILLER_67_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_85_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_26_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XTBUFX2 VPWR VGND la_data_out[38] la_data_in[37] la_data_in[36] TBUFX2
XFILLER_5_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_27_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_27_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_23_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_198_ VGND VGND VPWR VPWR _198_/HI wbs_dat_o[24] sky130_fd_sc_hd__conb_1
XFILLER_96_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_121_ VGND VGND VPWR VPWR _121_/HI la_data_out[76] sky130_fd_sc_hd__conb_1
XPHY_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_052_ VGND VGND VPWR VPWR _052_/HI io_out[27] sky130_fd_sc_hd__conb_1
XFILLER_78_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_104_ VGND VGND VPWR VPWR _104_/HI la_data_out[59] sky130_fd_sc_hd__conb_1
XPHY_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_035_ VGND VGND VPWR VPWR _035_/HI io_out[0] sky130_fd_sc_hd__conb_1
XFILLER_22_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_48_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_018_ VGND VGND VPWR VPWR io_oeb[6] _018_/LO sky130_fd_sc_hd__conb_1
XFILLER_98_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_76_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_44_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_8_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_58_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_58_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_197_ VGND VGND VPWR VPWR _197_/HI wbs_dat_o[23] sky130_fd_sc_hd__conb_1
XFILLER_96_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_120_ VGND VGND VPWR VPWR _120_/HI la_data_out[75] sky130_fd_sc_hd__conb_1
XFILLER_23_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_051_ VGND VGND VPWR VPWR _051_/HI io_out[25] sky130_fd_sc_hd__conb_1
XFILLER_11_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_42_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_103_ VGND VGND VPWR VPWR _103_/HI la_data_out[58] sky130_fd_sc_hd__conb_1
XPHY_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_034_ VGND VGND VPWR VPWR _034_/HI io_oeb[37] sky130_fd_sc_hd__conb_1
XFILLER_98_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_017_ VGND VGND VPWR VPWR io_oeb[4] _017_/LO sky130_fd_sc_hd__conb_1
XFILLER_98_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_97_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XAOI22X1 VPWR VGND io_out[14] io_in[12] io_in[13] io_in[10] io_in[11] AOI22X1
XFILLER_49_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_1_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_95_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_196_ VGND VGND VPWR VPWR _196_/HI wbs_dat_o[22] sky130_fd_sc_hd__conb_1
XFILLER_1_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_17_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_62_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_050_ VGND VGND VPWR VPWR _050_/HI io_out[22] sky130_fd_sc_hd__conb_1
XFILLER_11_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_3_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_59_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_179_ VGND VGND VPWR VPWR _179_/HI wbs_dat_o[5] sky130_fd_sc_hd__conb_1
XFILLER_6_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_97_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_80_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_20_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_102_ VGND VGND VPWR VPWR _102_/HI la_data_out[57] sky130_fd_sc_hd__conb_1
XPHY_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_033_ VGND VGND VPWR VPWR _033_/HI io_oeb[34] sky130_fd_sc_hd__conb_1
XFILLER_98_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_78_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_4_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_75_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_016_ VGND VGND VPWR VPWR io_oeb[3] _016_/LO sky130_fd_sc_hd__conb_1
XFILLER_98_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_41_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_65_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_17_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_95_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_73_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_195_ VGND VGND VPWR VPWR _195_/HI wbs_dat_o[21] sky130_fd_sc_hd__conb_1
XFILLER_6_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_178_ VGND VGND VPWR VPWR _178_/HI wbs_dat_o[4] sky130_fd_sc_hd__conb_1
XFILLER_69_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_101_ VGND VGND VPWR VPWR _101_/HI la_data_out[56] sky130_fd_sc_hd__conb_1
XPHY_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_032_ VGND VGND VPWR VPWR _032_/HI io_oeb[32] sky130_fd_sc_hd__conb_1
XFILLER_98_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_15_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_62_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_69_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_75_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_71_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_015_ VGND VGND VPWR VPWR io_oeb[1] _015_/LO sky130_fd_sc_hd__conb_1
XFILLER_3_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_26_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_71_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_12_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_49_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_41_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_194_ VGND VGND VPWR VPWR _194_/HI wbs_dat_o[20] sky130_fd_sc_hd__conb_1
XFILLER_41_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_78_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_177_ VGND VGND VPWR VPWR _177_/HI wbs_dat_o[3] sky130_fd_sc_hd__conb_1
XFILLER_2_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_37_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_87_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_100_ VGND VGND VPWR VPWR _100_/HI la_data_out[55] sky130_fd_sc_hd__conb_1
XFILLER_11_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_031_ VGND VGND VPWR VPWR _031_/HI io_oeb[30] sky130_fd_sc_hd__conb_1
XFILLER_98_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_101_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_19_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_88_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_76_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_8_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_014_ VGND VGND VPWR VPWR io_oeb[0] _014_/LO sky130_fd_sc_hd__conb_1
XFILLER_3_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_85_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_88_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_91_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_4_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_89_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_49_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_13_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_35_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_193_ VGND VGND VPWR VPWR _193_/HI wbs_dat_o[19] sky130_fd_sc_hd__conb_1
XFILLER_41_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_6_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_2_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_32_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_83_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_14_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_176_ VGND VGND VPWR VPWR _176_/HI wbs_dat_o[2] sky130_fd_sc_hd__conb_1
XFILLER_6_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_37_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_73_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_030_ VGND VGND VPWR VPWR _030_/HI io_oeb[28] sky130_fd_sc_hd__conb_1
XFILLER_0_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_47_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_159_ VGND VGND VPWR VPWR _159_/HI la_data_out[114] sky130_fd_sc_hd__conb_1
XFILLER_6_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_53_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XNOR3X1 VPWR VGND la_data_out[17] la_data_in[15] la_data_in[14] la_data_in[16] NOR3X1
XFILLER_88_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_83_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_71_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_013_ VGND VGND VPWR VPWR io_oeb[36] _013_/LO sky130_fd_sc_hd__conb_1
XFILLER_79_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_97_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_76_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_14_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_39_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_55_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_67_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_50_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_192_ VGND VGND VPWR VPWR _192_/HI wbs_dat_o[18] sky130_fd_sc_hd__conb_1
XFILLER_41_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_175_ VGND VGND VPWR VPWR _175_/HI wbs_dat_o[1] sky130_fd_sc_hd__conb_1
XFILLER_6_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_65_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_45_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_33_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_60_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XCLKBUF1 VPWR VGND io_out[20] io_in[19] CLKBUF1
XFILLER_88_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_42_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_158_ VGND VGND VPWR VPWR _158_/HI la_data_out[113] sky130_fd_sc_hd__conb_1
X_089_ VGND VGND VPWR VPWR _089_/HI la_data_out[43] sky130_fd_sc_hd__conb_1
XFILLER_69_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_012_ VGND VGND VPWR VPWR io_oeb[35] _012_/LO sky130_fd_sc_hd__conb_1
XFILLER_79_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_97_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_50_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_71_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_14_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_81_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_10_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_191_ VGND VGND VPWR VPWR _191_/HI wbs_dat_o[17] sky130_fd_sc_hd__conb_1
XFILLER_41_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_95_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_63_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_87_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_46_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_22_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_174_ VGND VGND VPWR VPWR _174_/HI wbs_dat_o[0] sky130_fd_sc_hd__conb_1
XFILLER_6_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XMUX2X1 VPWR VGND la_data_out[3] la_data_in[2] la_data_in[0] la_data_in[1] MUX2X1
XFILLER_96_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_45_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_3_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_78_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_27_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_157_ VGND VGND VPWR VPWR _157_/HI la_data_out[112] sky130_fd_sc_hd__conb_1
X_088_ VGND VGND VPWR VPWR _088_/HI la_data_out[42] sky130_fd_sc_hd__conb_1
XFILLER_97_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_83_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_83_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_011_ VGND VGND VPWR VPWR io_oeb[33] _011_/LO sky130_fd_sc_hd__conb_1
XFILLER_3_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_38_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_65_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_84_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_40_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_12_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_69_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_47_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_55_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_44_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_63_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_100_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_190_ VGND VGND VPWR VPWR _190_/HI wbs_dat_o[16] sky130_fd_sc_hd__conb_1
XFILLER_10_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_99_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_51_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_173_ VGND VGND VPWR VPWR _173_/HI wbs_ack_o sky130_fd_sc_hd__conb_1
XFILLER_6_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_77_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_156_ VGND VGND VPWR VPWR _156_/HI la_data_out[111] sky130_fd_sc_hd__conb_1
XFILLER_6_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_087_ VGND VGND VPWR VPWR _087_/HI la_data_out[40] sky130_fd_sc_hd__conb_1
XFILLER_97_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_010_ VGND VGND VPWR VPWR io_oeb[31] _010_/LO sky130_fd_sc_hd__conb_1
XFILLER_3_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_208_ VGND VGND VPWR VPWR _208_/HI io_oeb[9] sky130_fd_sc_hd__conb_1
X_139_ VGND VGND VPWR VPWR _139_/HI la_data_out[94] sky130_fd_sc_hd__conb_1
XFILLER_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_85_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_79_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_57_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_9_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_63_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_98_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_41_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_5_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_59_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_86_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_172_ VGND VGND VPWR VPWR _172_/HI la_data_out[127] sky130_fd_sc_hd__conb_1
XFILLER_10_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_64_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XAND2X1 VPWR VGND io_out[2] io_in[0] io_in[1] AND2X1
XPHY_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_155_ VGND VGND VPWR VPWR _155_/HI la_data_out[110] sky130_fd_sc_hd__conb_1
XFILLER_12_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_086_ VGND VGND VPWR VPWR _086_/HI la_data_out[39] sky130_fd_sc_hd__conb_1
XFILLER_2_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_20_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_43_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_207_ VGND VGND VPWR VPWR _207_/HI io_oeb[5] sky130_fd_sc_hd__conb_1
X_138_ VGND VGND VPWR VPWR _138_/HI la_data_out[93] sky130_fd_sc_hd__conb_1
X_069_ VGND VGND VPWR VPWR _069_/HI la_data_out[15] sky130_fd_sc_hd__conb_1
XFILLER_97_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_38_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_52_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_40_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_35_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_100_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_39_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_42_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_34_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_9_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_55_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_51_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_11_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_171_ VGND VGND VPWR VPWR _171_/HI la_data_out[126] sky130_fd_sc_hd__conb_1
XFILLER_52_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_6_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_91_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XAND2X2 VPWR VGND io_out[5] io_in[3] io_in[4] AND2X2
XFILLER_55_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_15_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_154_ VGND VGND VPWR VPWR _154_/HI la_data_out[109] sky130_fd_sc_hd__conb_1
X_085_ VGND VGND VPWR VPWR _085_/HI la_data_out[37] sky130_fd_sc_hd__conb_1
XFILLER_6_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_93_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_77_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_21_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_96_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_52_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_58_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_74_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_206_ VGND VGND VPWR VPWR _206_/HI io_oeb[2] sky130_fd_sc_hd__conb_1
XFILLER_7_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_137_ VGND VGND VPWR VPWR _137_/HI la_data_out[92] sky130_fd_sc_hd__conb_1
XFILLER_99_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_068_ VGND VGND VPWR VPWR _068_/HI la_data_out[14] sky130_fd_sc_hd__conb_1
XFILLER_97_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_57_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_56_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_25_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_79_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_98_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_22_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_89_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_29_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_13_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_4_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_89_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_5_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_86_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_14_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_170_ VGND VGND VPWR VPWR _170_/HI la_data_out[125] sky130_fd_sc_hd__conb_1
XFILLER_6_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_3_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_59_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_74_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_153_ VGND VGND VPWR VPWR _153_/HI la_data_out[108] sky130_fd_sc_hd__conb_1
X_084_ VGND VGND VPWR VPWR _084_/HI la_data_out[36] sky130_fd_sc_hd__conb_1
XFILLER_12_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_56_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_58_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_205_ VGND VGND VPWR VPWR _205_/HI wbs_dat_o[31] sky130_fd_sc_hd__conb_1
X_136_ VGND VGND VPWR VPWR _136_/HI la_data_out[91] sky130_fd_sc_hd__conb_1
XFILLER_99_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_067_ VGND VGND VPWR VPWR _067_/HI la_data_out[12] sky130_fd_sc_hd__conb_1
XFILLER_38_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_19_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_69_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_87_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_85_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_119_ VGND VGND VPWR VPWR _119_/HI la_data_out[74] sky130_fd_sc_hd__conb_1
XFILLER_100_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_1_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_57_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_90_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_77_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_66_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_25_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_1_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_76_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_50_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_45_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_95_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_152_ VGND VGND VPWR VPWR _152_/HI la_data_out[107] sky130_fd_sc_hd__conb_1
XPHY_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_083_ VGND VGND VPWR VPWR _083_/HI la_data_out[34] sky130_fd_sc_hd__conb_1
XFILLER_88_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_53_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_33_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_59_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_90_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_74_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_204_ VGND VGND VPWR VPWR _204_/HI wbs_dat_o[30] sky130_fd_sc_hd__conb_1
XFILLER_11_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_135_ VGND VGND VPWR VPWR _135_/HI la_data_out[90] sky130_fd_sc_hd__conb_1
X_066_ VGND VGND VPWR VPWR _066_/HI la_data_out[11] sky130_fd_sc_hd__conb_1
XFILLER_7_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_34_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_88_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_84_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_44_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_47_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_118_ VGND VGND VPWR VPWR _118_/HI la_data_out[73] sky130_fd_sc_hd__conb_1
XFILLER_50_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_049_ VGND VGND VPWR VPWR _049_/HI io_out[21] sky130_fd_sc_hd__conb_1
XFILLER_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_85_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_81_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_29_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_48_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_22_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_17_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_72_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_40_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_31_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_98_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_54_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_51_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_101_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_86_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_67_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_82_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_151_ VGND VGND VPWR VPWR _151_/HI la_data_out[106] sky130_fd_sc_hd__conb_1
XFILLER_50_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_082_ VGND VGND VPWR VPWR _082_/HI la_data_out[33] sky130_fd_sc_hd__conb_1
XFILLER_88_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_18_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_68_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_68_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_52_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_87_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_43_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_203_ VGND VGND VPWR VPWR _203_/HI wbs_dat_o[29] sky130_fd_sc_hd__conb_1
XFILLER_11_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_134_ VGND VGND VPWR VPWR _134_/HI la_data_out[89] sky130_fd_sc_hd__conb_1
X_065_ VGND VGND VPWR VPWR _065_/HI la_data_out[9] sky130_fd_sc_hd__conb_1
XFILLER_99_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_80_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_88_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_100_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_12_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_31_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_117_ VGND VGND VPWR VPWR _117_/HI la_data_out[72] sky130_fd_sc_hd__conb_1
X_048_ VGND VGND VPWR VPWR _048_/HI io_out[19] sky130_fd_sc_hd__conb_1
XFILLER_93_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_72_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_96_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_54_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_13_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_31_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_82_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_67_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_54_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_54_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_82_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_10_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_83_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_32_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_27_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_82_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_150_ VGND VGND VPWR VPWR _150_/HI la_data_out[105] sky130_fd_sc_hd__conb_1
X_081_ VGND VGND VPWR VPWR _081_/HI la_data_out[31] sky130_fd_sc_hd__conb_1
XFILLER_10_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_77_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_33_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_14_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_3_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_87_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_90_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_11_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_70_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_202_ VGND VGND VPWR VPWR _202_/HI wbs_dat_o[28] sky130_fd_sc_hd__conb_1
XFILLER_7_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_7_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_133_ VGND VGND VPWR VPWR _133_/HI la_data_out[88] sky130_fd_sc_hd__conb_1
X_064_ VGND VGND VPWR VPWR _064_/HI la_data_out[8] sky130_fd_sc_hd__conb_1
XFILLER_78_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_65_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_29_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_25_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_48_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_28_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_116_ VGND VGND VPWR VPWR _116_/HI la_data_out[71] sky130_fd_sc_hd__conb_1
XFILLER_50_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_047_ VGND VGND VPWR VPWR _047_/HI io_out[17] sky130_fd_sc_hd__conb_1
XFILLER_78_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_93_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_46_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_30_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_39_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_96_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_90_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_35_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_16_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XOAI21X1 VPWR VGND la_data_out[21] la_data_in[18] la_data_in[19] la_data_in[20] OAI21X1
XFILLER_12_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_98_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_26_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_62_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_41_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_15_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_9_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_31_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_72_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_75_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_8_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_86_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_67_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_23_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_22_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_10_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_89_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_26_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_60_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_9_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_5_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_95_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_49_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_36_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_101_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_47_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_27_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_42_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_23_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_080_ VGND VGND VPWR VPWR _080_/HI la_data_out[30] sky130_fd_sc_hd__conb_1
XFILLER_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_2_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_88_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_5_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_77_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_92_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_18_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_33_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_41_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_76_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_24_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_64_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_99_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_59_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_74_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_28_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_43_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_201_ VGND VGND VPWR VPWR _201_/HI wbs_dat_o[27] sky130_fd_sc_hd__conb_1
XPHY_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_132_ VGND VGND VPWR VPWR _132_/HI la_data_out[87] sky130_fd_sc_hd__conb_1
XFILLER_7_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_7_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_23_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_063_ VGND VGND VPWR VPWR _063_/HI la_data_out[7] sky130_fd_sc_hd__conb_1
XFILLER_97_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_78_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_66_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_93_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_48_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_58_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_46_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_73_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_56_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_25_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_100_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_79_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_48_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_75_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_75_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_28_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_55_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_70_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_115_ VGND VGND VPWR VPWR _115_/HI la_data_out[70] sky130_fd_sc_hd__conb_1
XFILLER_7_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
X_046_ VGND VGND VPWR VPWR _046_/HI io_out[15] sky130_fd_sc_hd__conb_1
XFILLER_3_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_38_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_34_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_46_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_61_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_97_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_57_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_69_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_45_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_55_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_84_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_37_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_13_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_52_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_71_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_80_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_4_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_96_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_29_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_29_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_63_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_8_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_6_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_6_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_029_ VGND VGND VPWR VPWR _029_/HI io_oeb[26] sky130_fd_sc_hd__conb_1
XFILLER_79_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_94_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_39_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_66_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_19_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_34_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_81_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XHAX1 VPWR VGND io_out[24] io_out[23] io_in[22] io_in[21] HAX1
XFILLER_97_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_85_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_45_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_82_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_41_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_25_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_9_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_40_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_21_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_31_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_31_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_95_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_0_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_76_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_91_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_56_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_63_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_44_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_8_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_68_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_99_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_100_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
XFILLER_98_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_12
.ends

