MACRO INVX8
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN INVX8 0 0 ;
 SITE CORE ;
 SYMMETRY X Y R90 ;
  PIN VDD
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.00000000 2.52500000 4.60000000 2.91500000 ;
    END
  END VDD

  PIN GND
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.00000000 -0.19500000 4.60000000 0.19500000 ;
    END
  END GND

  PIN Y
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        POLYGON 0.34500000 0.60000000 0.34500000 0.83000000 0.39000000 0.83000000 0.39000000 1.90000000 0.34500000 1.90000000 0.34500000 2.13000000 0.57500000 2.13000000 0.57500000 2.08500000 2.18500000 2.08500000 2.18500000 2.13000000 2.41500000 2.13000000 2.41500000 2.08500000 4.02500000 2.08500000 4.02500000 2.13000000 4.25500000 2.13000000 4.25500000 1.90000000 4.21000000 1.90000000 4.21000000 0.83000000 4.25500000 0.83000000 4.25500000 0.60000000 4.02500000 0.60000000 4.02500000 0.83000000 4.07000000 0.83000000 4.07000000 1.90000000 4.02500000 1.90000000 4.02500000 1.94500000 2.41500000 1.94500000 2.41500000 1.90000000 2.18500000 1.90000000 2.18500000 1.94500000 0.57500000 1.94500000 0.57500000 1.90000000 0.53000000 1.90000000 0.53000000 0.83000000 0.57500000 0.83000000 0.57500000 0.78500000 2.18500000 0.78500000 2.18500000 0.83000000 2.41500000 0.83000000 2.41500000 0.60000000 2.18500000 0.60000000 2.18500000 0.64500000 0.57500000 0.64500000 0.57500000 0.60000000 ;
    END
  END Y

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        POLYGON 0.80500000 0.99000000 0.80500000 1.22000000 0.85000000 1.22000000 0.85000000 1.51000000 0.80500000 1.51000000 0.80500000 1.74000000 1.03500000 1.74000000 1.03500000 1.69500000 1.72500000 1.69500000 1.72500000 1.74000000 1.95500000 1.74000000 1.95500000 1.69500000 2.64500000 1.69500000 2.64500000 1.74000000 2.87500000 1.74000000 2.87500000 1.69500000 3.56500000 1.69500000 3.56500000 1.74000000 3.79500000 1.74000000 3.79500000 1.51000000 3.75000000 1.51000000 3.75000000 1.22000000 3.79500000 1.22000000 3.79500000 0.99000000 3.56500000 0.99000000 3.56500000 1.22000000 3.61000000 1.22000000 3.61000000 1.51000000 3.56500000 1.51000000 3.56500000 1.55500000 2.87500000 1.55500000 2.87500000 1.51000000 2.83000000 1.51000000 2.83000000 1.22000000 2.87500000 1.22000000 2.87500000 0.99000000 2.64500000 0.99000000 2.64500000 1.22000000 2.69000000 1.22000000 2.69000000 1.51000000 2.64500000 1.51000000 2.64500000 1.55500000 1.95500000 1.55500000 1.95500000 1.51000000 1.91000000 1.51000000 1.91000000 1.22000000 1.95500000 1.22000000 1.95500000 0.99000000 1.72500000 0.99000000 1.72500000 1.22000000 1.77000000 1.22000000 1.77000000 1.51000000 1.72500000 1.51000000 1.72500000 1.55500000 1.03500000 1.55500000 1.03500000 1.51000000 0.99000000 1.51000000 0.99000000 1.22000000 1.03500000 1.22000000 1.03500000 0.99000000 ;
    END
  END A


END INVX8
