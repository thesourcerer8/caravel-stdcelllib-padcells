MACRO TBUFX1
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN TBUFX1 0 0 ;
 SITE CORE ;
 SYMMETRY X Y R90 ;
  PIN VDD
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.00000000 2.48000000 3.68000000 2.96000000 ;
    END
  END VDD

  PIN GND
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.00000000 -0.24000000 3.68000000 0.24000000 ;
    END
  END GND

  PIN Y
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 3.07500000 0.39500000 3.36500000 0.68500000 ;
        RECT 3.15000000 0.68500000 3.29000000 2.01500000 ;
        RECT 3.07500000 2.01500000 3.36500000 2.30500000 ;
    END
  END Y

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 1.69500000 1.29500000 1.98500000 1.58500000 ;
    END
  END A

  PIN EN
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.77500000 0.93500000 1.06500000 1.01000000 ;
        RECT 2.61500000 0.93500000 2.90500000 1.01000000 ;
        RECT 0.77500000 1.01000000 2.90500000 1.15000000 ;
        RECT 2.61500000 1.15000000 2.90500000 1.22500000 ;
        RECT 0.77500000 1.15000000 1.06500000 1.58500000 ;
    END
  END EN


END TBUFX1
