MACRO AND2X2
 CLASS CORE ;
 ORIGIN 0 0 ;
 FOREIGN AND2X2 0 0 ;
 SITE CORE ;
 SYMMETRY X Y R90 ;
  PIN VDD
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.00000000 3965.00000000 4160.00000000 4355.00000000 ;
    END
  END VDD

  PIN GND
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        RECT 0.00000000 -195.00000000 4160.00000000 195.00000000 ;
    END
  END GND

  PIN Y
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        POLYGON 3525.00000000 730.00000000 3525.00000000 960.00000000 3570.00000000 960.00000000 3570.00000000 3200.00000000 3525.00000000 3200.00000000 3525.00000000 3430.00000000 3755.00000000 3430.00000000 3755.00000000 3200.00000000 3710.00000000 3200.00000000 3710.00000000 960.00000000 3755.00000000 960.00000000 3755.00000000 730.00000000 ;
    END
  END Y

  PIN B
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        POLYGON 1965.00000000 1120.00000000 1965.00000000 1350.00000000 2010.00000000 1350.00000000 2010.00000000 2810.00000000 1965.00000000 2810.00000000 1965.00000000 3040.00000000 2195.00000000 3040.00000000 2195.00000000 2810.00000000 2150.00000000 2810.00000000 2150.00000000 1350.00000000 2195.00000000 1350.00000000 2195.00000000 1120.00000000 ;
    END
  END B

  PIN A
   DIRECTION INOUT ;
   USE SIGNAL ;
   SHAPE ABUTMENT ;
    PORT
     CLASS CORE ;
       LAYER metal2 ;
        POLYGON 925.00000000 1120.00000000 925.00000000 1350.00000000 970.00000000 1350.00000000 970.00000000 2810.00000000 925.00000000 2810.00000000 925.00000000 3040.00000000 1155.00000000 3040.00000000 1155.00000000 2810.00000000 1110.00000000 2810.00000000 1110.00000000 1350.00000000 1155.00000000 1350.00000000 1155.00000000 1120.00000000 ;
    END
  END A


END AND2X2
